magic
tech sky130A
magscale 1 2
timestamp 1757832390
<< metal3 >>
rect -3928 1292 -3156 1320
rect -3928 868 -3240 1292
rect -3176 868 -3156 1292
rect -3928 840 -3156 868
rect -2916 1292 -2144 1320
rect -2916 868 -2228 1292
rect -2164 868 -2144 1292
rect -2916 840 -2144 868
rect -1904 1292 -1132 1320
rect -1904 868 -1216 1292
rect -1152 868 -1132 1292
rect -1904 840 -1132 868
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect 1132 1292 1904 1320
rect 1132 868 1820 1292
rect 1884 868 1904 1292
rect 1132 840 1904 868
rect 2144 1292 2916 1320
rect 2144 868 2832 1292
rect 2896 868 2916 1292
rect 2144 840 2916 868
rect 3156 1292 3928 1320
rect 3156 868 3844 1292
rect 3908 868 3928 1292
rect 3156 840 3928 868
rect -3928 572 -3156 600
rect -3928 148 -3240 572
rect -3176 148 -3156 572
rect -3928 120 -3156 148
rect -2916 572 -2144 600
rect -2916 148 -2228 572
rect -2164 148 -2144 572
rect -2916 120 -2144 148
rect -1904 572 -1132 600
rect -1904 148 -1216 572
rect -1152 148 -1132 572
rect -1904 120 -1132 148
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect 1132 572 1904 600
rect 1132 148 1820 572
rect 1884 148 1904 572
rect 1132 120 1904 148
rect 2144 572 2916 600
rect 2144 148 2832 572
rect 2896 148 2916 572
rect 2144 120 2916 148
rect 3156 572 3928 600
rect 3156 148 3844 572
rect 3908 148 3928 572
rect 3156 120 3928 148
rect -3928 -148 -3156 -120
rect -3928 -572 -3240 -148
rect -3176 -572 -3156 -148
rect -3928 -600 -3156 -572
rect -2916 -148 -2144 -120
rect -2916 -572 -2228 -148
rect -2164 -572 -2144 -148
rect -2916 -600 -2144 -572
rect -1904 -148 -1132 -120
rect -1904 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -1904 -600 -1132 -572
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect 1132 -148 1904 -120
rect 1132 -572 1820 -148
rect 1884 -572 1904 -148
rect 1132 -600 1904 -572
rect 2144 -148 2916 -120
rect 2144 -572 2832 -148
rect 2896 -572 2916 -148
rect 2144 -600 2916 -572
rect 3156 -148 3928 -120
rect 3156 -572 3844 -148
rect 3908 -572 3928 -148
rect 3156 -600 3928 -572
rect -3928 -868 -3156 -840
rect -3928 -1292 -3240 -868
rect -3176 -1292 -3156 -868
rect -3928 -1320 -3156 -1292
rect -2916 -868 -2144 -840
rect -2916 -1292 -2228 -868
rect -2164 -1292 -2144 -868
rect -2916 -1320 -2144 -1292
rect -1904 -868 -1132 -840
rect -1904 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -1904 -1320 -1132 -1292
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect 1132 -868 1904 -840
rect 1132 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 1132 -1320 1904 -1292
rect 2144 -868 2916 -840
rect 2144 -1292 2832 -868
rect 2896 -1292 2916 -868
rect 2144 -1320 2916 -1292
rect 3156 -868 3928 -840
rect 3156 -1292 3844 -868
rect 3908 -1292 3928 -868
rect 3156 -1320 3928 -1292
<< via3 >>
rect -3240 868 -3176 1292
rect -2228 868 -2164 1292
rect -1216 868 -1152 1292
rect -204 868 -140 1292
rect 808 868 872 1292
rect 1820 868 1884 1292
rect 2832 868 2896 1292
rect 3844 868 3908 1292
rect -3240 148 -3176 572
rect -2228 148 -2164 572
rect -1216 148 -1152 572
rect -204 148 -140 572
rect 808 148 872 572
rect 1820 148 1884 572
rect 2832 148 2896 572
rect 3844 148 3908 572
rect -3240 -572 -3176 -148
rect -2228 -572 -2164 -148
rect -1216 -572 -1152 -148
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect 1820 -572 1884 -148
rect 2832 -572 2896 -148
rect 3844 -572 3908 -148
rect -3240 -1292 -3176 -868
rect -2228 -1292 -2164 -868
rect -1216 -1292 -1152 -868
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect 1820 -1292 1884 -868
rect 2832 -1292 2896 -868
rect 3844 -1292 3908 -868
<< mimcap >>
rect -3888 1240 -3488 1280
rect -3888 920 -3848 1240
rect -3528 920 -3488 1240
rect -3888 880 -3488 920
rect -2876 1240 -2476 1280
rect -2876 920 -2836 1240
rect -2516 920 -2476 1240
rect -2876 880 -2476 920
rect -1864 1240 -1464 1280
rect -1864 920 -1824 1240
rect -1504 920 -1464 1240
rect -1864 880 -1464 920
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect 1172 1240 1572 1280
rect 1172 920 1212 1240
rect 1532 920 1572 1240
rect 1172 880 1572 920
rect 2184 1240 2584 1280
rect 2184 920 2224 1240
rect 2544 920 2584 1240
rect 2184 880 2584 920
rect 3196 1240 3596 1280
rect 3196 920 3236 1240
rect 3556 920 3596 1240
rect 3196 880 3596 920
rect -3888 520 -3488 560
rect -3888 200 -3848 520
rect -3528 200 -3488 520
rect -3888 160 -3488 200
rect -2876 520 -2476 560
rect -2876 200 -2836 520
rect -2516 200 -2476 520
rect -2876 160 -2476 200
rect -1864 520 -1464 560
rect -1864 200 -1824 520
rect -1504 200 -1464 520
rect -1864 160 -1464 200
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect 1172 520 1572 560
rect 1172 200 1212 520
rect 1532 200 1572 520
rect 1172 160 1572 200
rect 2184 520 2584 560
rect 2184 200 2224 520
rect 2544 200 2584 520
rect 2184 160 2584 200
rect 3196 520 3596 560
rect 3196 200 3236 520
rect 3556 200 3596 520
rect 3196 160 3596 200
rect -3888 -200 -3488 -160
rect -3888 -520 -3848 -200
rect -3528 -520 -3488 -200
rect -3888 -560 -3488 -520
rect -2876 -200 -2476 -160
rect -2876 -520 -2836 -200
rect -2516 -520 -2476 -200
rect -2876 -560 -2476 -520
rect -1864 -200 -1464 -160
rect -1864 -520 -1824 -200
rect -1504 -520 -1464 -200
rect -1864 -560 -1464 -520
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect 1172 -200 1572 -160
rect 1172 -520 1212 -200
rect 1532 -520 1572 -200
rect 1172 -560 1572 -520
rect 2184 -200 2584 -160
rect 2184 -520 2224 -200
rect 2544 -520 2584 -200
rect 2184 -560 2584 -520
rect 3196 -200 3596 -160
rect 3196 -520 3236 -200
rect 3556 -520 3596 -200
rect 3196 -560 3596 -520
rect -3888 -920 -3488 -880
rect -3888 -1240 -3848 -920
rect -3528 -1240 -3488 -920
rect -3888 -1280 -3488 -1240
rect -2876 -920 -2476 -880
rect -2876 -1240 -2836 -920
rect -2516 -1240 -2476 -920
rect -2876 -1280 -2476 -1240
rect -1864 -920 -1464 -880
rect -1864 -1240 -1824 -920
rect -1504 -1240 -1464 -920
rect -1864 -1280 -1464 -1240
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect 1172 -920 1572 -880
rect 1172 -1240 1212 -920
rect 1532 -1240 1572 -920
rect 1172 -1280 1572 -1240
rect 2184 -920 2584 -880
rect 2184 -1240 2224 -920
rect 2544 -1240 2584 -920
rect 2184 -1280 2584 -1240
rect 3196 -920 3596 -880
rect 3196 -1240 3236 -920
rect 3556 -1240 3596 -920
rect 3196 -1280 3596 -1240
<< mimcapcontact >>
rect -3848 920 -3528 1240
rect -2836 920 -2516 1240
rect -1824 920 -1504 1240
rect -812 920 -492 1240
rect 200 920 520 1240
rect 1212 920 1532 1240
rect 2224 920 2544 1240
rect 3236 920 3556 1240
rect -3848 200 -3528 520
rect -2836 200 -2516 520
rect -1824 200 -1504 520
rect -812 200 -492 520
rect 200 200 520 520
rect 1212 200 1532 520
rect 2224 200 2544 520
rect 3236 200 3556 520
rect -3848 -520 -3528 -200
rect -2836 -520 -2516 -200
rect -1824 -520 -1504 -200
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect 1212 -520 1532 -200
rect 2224 -520 2544 -200
rect 3236 -520 3556 -200
rect -3848 -1240 -3528 -920
rect -2836 -1240 -2516 -920
rect -1824 -1240 -1504 -920
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect 1212 -1240 1532 -920
rect 2224 -1240 2544 -920
rect 3236 -1240 3556 -920
<< metal4 >>
rect -3740 1241 -3636 1440
rect -3260 1292 -3156 1440
rect -3849 1240 -3527 1241
rect -3849 920 -3848 1240
rect -3528 920 -3527 1240
rect -3849 919 -3527 920
rect -3740 521 -3636 919
rect -3260 868 -3240 1292
rect -3176 868 -3156 1292
rect -2728 1241 -2624 1440
rect -2248 1292 -2144 1440
rect -2837 1240 -2515 1241
rect -2837 920 -2836 1240
rect -2516 920 -2515 1240
rect -2837 919 -2515 920
rect -3260 572 -3156 868
rect -3849 520 -3527 521
rect -3849 200 -3848 520
rect -3528 200 -3527 520
rect -3849 199 -3527 200
rect -3740 -199 -3636 199
rect -3260 148 -3240 572
rect -3176 148 -3156 572
rect -2728 521 -2624 919
rect -2248 868 -2228 1292
rect -2164 868 -2144 1292
rect -1716 1241 -1612 1440
rect -1236 1292 -1132 1440
rect -1825 1240 -1503 1241
rect -1825 920 -1824 1240
rect -1504 920 -1503 1240
rect -1825 919 -1503 920
rect -2248 572 -2144 868
rect -2837 520 -2515 521
rect -2837 200 -2836 520
rect -2516 200 -2515 520
rect -2837 199 -2515 200
rect -3260 -148 -3156 148
rect -3849 -200 -3527 -199
rect -3849 -520 -3848 -200
rect -3528 -520 -3527 -200
rect -3849 -521 -3527 -520
rect -3740 -919 -3636 -521
rect -3260 -572 -3240 -148
rect -3176 -572 -3156 -148
rect -2728 -199 -2624 199
rect -2248 148 -2228 572
rect -2164 148 -2144 572
rect -1716 521 -1612 919
rect -1236 868 -1216 1292
rect -1152 868 -1132 1292
rect -704 1241 -600 1440
rect -224 1292 -120 1440
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -1236 572 -1132 868
rect -1825 520 -1503 521
rect -1825 200 -1824 520
rect -1504 200 -1503 520
rect -1825 199 -1503 200
rect -2248 -148 -2144 148
rect -2837 -200 -2515 -199
rect -2837 -520 -2836 -200
rect -2516 -520 -2515 -200
rect -2837 -521 -2515 -520
rect -3260 -868 -3156 -572
rect -3849 -920 -3527 -919
rect -3849 -1240 -3848 -920
rect -3528 -1240 -3527 -920
rect -3849 -1241 -3527 -1240
rect -3740 -1440 -3636 -1241
rect -3260 -1292 -3240 -868
rect -3176 -1292 -3156 -868
rect -2728 -919 -2624 -521
rect -2248 -572 -2228 -148
rect -2164 -572 -2144 -148
rect -1716 -199 -1612 199
rect -1236 148 -1216 572
rect -1152 148 -1132 572
rect -704 521 -600 919
rect -224 868 -204 1292
rect -140 868 -120 1292
rect 308 1241 412 1440
rect 788 1292 892 1440
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -224 572 -120 868
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -1236 -148 -1132 148
rect -1825 -200 -1503 -199
rect -1825 -520 -1824 -200
rect -1504 -520 -1503 -200
rect -1825 -521 -1503 -520
rect -2248 -868 -2144 -572
rect -2837 -920 -2515 -919
rect -2837 -1240 -2836 -920
rect -2516 -1240 -2515 -920
rect -2837 -1241 -2515 -1240
rect -3260 -1440 -3156 -1292
rect -2728 -1440 -2624 -1241
rect -2248 -1292 -2228 -868
rect -2164 -1292 -2144 -868
rect -1716 -919 -1612 -521
rect -1236 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -704 -199 -600 199
rect -224 148 -204 572
rect -140 148 -120 572
rect 308 521 412 919
rect 788 868 808 1292
rect 872 868 892 1292
rect 1320 1241 1424 1440
rect 1800 1292 1904 1440
rect 1211 1240 1533 1241
rect 1211 920 1212 1240
rect 1532 920 1533 1240
rect 1211 919 1533 920
rect 788 572 892 868
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -1236 -868 -1132 -572
rect -1825 -920 -1503 -919
rect -1825 -1240 -1824 -920
rect -1504 -1240 -1503 -920
rect -1825 -1241 -1503 -1240
rect -2248 -1440 -2144 -1292
rect -1716 -1440 -1612 -1241
rect -1236 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -704 -919 -600 -521
rect -224 -572 -204 -148
rect -140 -572 -120 -148
rect 308 -199 412 199
rect 788 148 808 572
rect 872 148 892 572
rect 1320 521 1424 919
rect 1800 868 1820 1292
rect 1884 868 1904 1292
rect 2332 1241 2436 1440
rect 2812 1292 2916 1440
rect 2223 1240 2545 1241
rect 2223 920 2224 1240
rect 2544 920 2545 1240
rect 2223 919 2545 920
rect 1800 572 1904 868
rect 1211 520 1533 521
rect 1211 200 1212 520
rect 1532 200 1533 520
rect 1211 199 1533 200
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -224 -868 -120 -572
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -1236 -1440 -1132 -1292
rect -704 -1440 -600 -1241
rect -224 -1292 -204 -868
rect -140 -1292 -120 -868
rect 308 -919 412 -521
rect 788 -572 808 -148
rect 872 -572 892 -148
rect 1320 -199 1424 199
rect 1800 148 1820 572
rect 1884 148 1904 572
rect 2332 521 2436 919
rect 2812 868 2832 1292
rect 2896 868 2916 1292
rect 3344 1241 3448 1440
rect 3824 1292 3928 1440
rect 3235 1240 3557 1241
rect 3235 920 3236 1240
rect 3556 920 3557 1240
rect 3235 919 3557 920
rect 2812 572 2916 868
rect 2223 520 2545 521
rect 2223 200 2224 520
rect 2544 200 2545 520
rect 2223 199 2545 200
rect 1800 -148 1904 148
rect 1211 -200 1533 -199
rect 1211 -520 1212 -200
rect 1532 -520 1533 -200
rect 1211 -521 1533 -520
rect 788 -868 892 -572
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -224 -1440 -120 -1292
rect 308 -1440 412 -1241
rect 788 -1292 808 -868
rect 872 -1292 892 -868
rect 1320 -919 1424 -521
rect 1800 -572 1820 -148
rect 1884 -572 1904 -148
rect 2332 -199 2436 199
rect 2812 148 2832 572
rect 2896 148 2916 572
rect 3344 521 3448 919
rect 3824 868 3844 1292
rect 3908 868 3928 1292
rect 3824 572 3928 868
rect 3235 520 3557 521
rect 3235 200 3236 520
rect 3556 200 3557 520
rect 3235 199 3557 200
rect 2812 -148 2916 148
rect 2223 -200 2545 -199
rect 2223 -520 2224 -200
rect 2544 -520 2545 -200
rect 2223 -521 2545 -520
rect 1800 -868 1904 -572
rect 1211 -920 1533 -919
rect 1211 -1240 1212 -920
rect 1532 -1240 1533 -920
rect 1211 -1241 1533 -1240
rect 788 -1440 892 -1292
rect 1320 -1440 1424 -1241
rect 1800 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 2332 -919 2436 -521
rect 2812 -572 2832 -148
rect 2896 -572 2916 -148
rect 3344 -199 3448 199
rect 3824 148 3844 572
rect 3908 148 3928 572
rect 3824 -148 3928 148
rect 3235 -200 3557 -199
rect 3235 -520 3236 -200
rect 3556 -520 3557 -200
rect 3235 -521 3557 -520
rect 2812 -868 2916 -572
rect 2223 -920 2545 -919
rect 2223 -1240 2224 -920
rect 2544 -1240 2545 -920
rect 2223 -1241 2545 -1240
rect 1800 -1440 1904 -1292
rect 2332 -1440 2436 -1241
rect 2812 -1292 2832 -868
rect 2896 -1292 2916 -868
rect 3344 -919 3448 -521
rect 3824 -572 3844 -148
rect 3908 -572 3928 -148
rect 3824 -868 3928 -572
rect 3235 -920 3557 -919
rect 3235 -1240 3236 -920
rect 3556 -1240 3557 -920
rect 3235 -1241 3557 -1240
rect 2812 -1440 2916 -1292
rect 3344 -1440 3448 -1241
rect 3824 -1292 3844 -868
rect 3908 -1292 3928 -868
rect 3824 -1440 3928 -1292
<< properties >>
string FIXED_BBOX 3156 840 3636 1320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 8 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
