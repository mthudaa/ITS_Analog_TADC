magic
tech sky130A
magscale 1 2
timestamp 1757383169
<< metal3 >>
rect -32264 2372 -31492 2400
rect -32264 1948 -31576 2372
rect -31512 1948 -31492 2372
rect -32264 1920 -31492 1948
rect -31252 2372 -30480 2400
rect -31252 1948 -30564 2372
rect -30500 1948 -30480 2372
rect -31252 1920 -30480 1948
rect -30240 2372 -29468 2400
rect -30240 1948 -29552 2372
rect -29488 1948 -29468 2372
rect -30240 1920 -29468 1948
rect -29228 2372 -28456 2400
rect -29228 1948 -28540 2372
rect -28476 1948 -28456 2372
rect -29228 1920 -28456 1948
rect -28216 2372 -27444 2400
rect -28216 1948 -27528 2372
rect -27464 1948 -27444 2372
rect -28216 1920 -27444 1948
rect -27204 2372 -26432 2400
rect -27204 1948 -26516 2372
rect -26452 1948 -26432 2372
rect -27204 1920 -26432 1948
rect -26192 2372 -25420 2400
rect -26192 1948 -25504 2372
rect -25440 1948 -25420 2372
rect -26192 1920 -25420 1948
rect -25180 2372 -24408 2400
rect -25180 1948 -24492 2372
rect -24428 1948 -24408 2372
rect -25180 1920 -24408 1948
rect -24168 2372 -23396 2400
rect -24168 1948 -23480 2372
rect -23416 1948 -23396 2372
rect -24168 1920 -23396 1948
rect -23156 2372 -22384 2400
rect -23156 1948 -22468 2372
rect -22404 1948 -22384 2372
rect -23156 1920 -22384 1948
rect -22144 2372 -21372 2400
rect -22144 1948 -21456 2372
rect -21392 1948 -21372 2372
rect -22144 1920 -21372 1948
rect -21132 2372 -20360 2400
rect -21132 1948 -20444 2372
rect -20380 1948 -20360 2372
rect -21132 1920 -20360 1948
rect -20120 2372 -19348 2400
rect -20120 1948 -19432 2372
rect -19368 1948 -19348 2372
rect -20120 1920 -19348 1948
rect -19108 2372 -18336 2400
rect -19108 1948 -18420 2372
rect -18356 1948 -18336 2372
rect -19108 1920 -18336 1948
rect -18096 2372 -17324 2400
rect -18096 1948 -17408 2372
rect -17344 1948 -17324 2372
rect -18096 1920 -17324 1948
rect -17084 2372 -16312 2400
rect -17084 1948 -16396 2372
rect -16332 1948 -16312 2372
rect -17084 1920 -16312 1948
rect -16072 2372 -15300 2400
rect -16072 1948 -15384 2372
rect -15320 1948 -15300 2372
rect -16072 1920 -15300 1948
rect -15060 2372 -14288 2400
rect -15060 1948 -14372 2372
rect -14308 1948 -14288 2372
rect -15060 1920 -14288 1948
rect -14048 2372 -13276 2400
rect -14048 1948 -13360 2372
rect -13296 1948 -13276 2372
rect -14048 1920 -13276 1948
rect -13036 2372 -12264 2400
rect -13036 1948 -12348 2372
rect -12284 1948 -12264 2372
rect -13036 1920 -12264 1948
rect -12024 2372 -11252 2400
rect -12024 1948 -11336 2372
rect -11272 1948 -11252 2372
rect -12024 1920 -11252 1948
rect -11012 2372 -10240 2400
rect -11012 1948 -10324 2372
rect -10260 1948 -10240 2372
rect -11012 1920 -10240 1948
rect -10000 2372 -9228 2400
rect -10000 1948 -9312 2372
rect -9248 1948 -9228 2372
rect -10000 1920 -9228 1948
rect -8988 2372 -8216 2400
rect -8988 1948 -8300 2372
rect -8236 1948 -8216 2372
rect -8988 1920 -8216 1948
rect -7976 2372 -7204 2400
rect -7976 1948 -7288 2372
rect -7224 1948 -7204 2372
rect -7976 1920 -7204 1948
rect -6964 2372 -6192 2400
rect -6964 1948 -6276 2372
rect -6212 1948 -6192 2372
rect -6964 1920 -6192 1948
rect -5952 2372 -5180 2400
rect -5952 1948 -5264 2372
rect -5200 1948 -5180 2372
rect -5952 1920 -5180 1948
rect -4940 2372 -4168 2400
rect -4940 1948 -4252 2372
rect -4188 1948 -4168 2372
rect -4940 1920 -4168 1948
rect -3928 2372 -3156 2400
rect -3928 1948 -3240 2372
rect -3176 1948 -3156 2372
rect -3928 1920 -3156 1948
rect -2916 2372 -2144 2400
rect -2916 1948 -2228 2372
rect -2164 1948 -2144 2372
rect -2916 1920 -2144 1948
rect -1904 2372 -1132 2400
rect -1904 1948 -1216 2372
rect -1152 1948 -1132 2372
rect -1904 1920 -1132 1948
rect -892 2372 -120 2400
rect -892 1948 -204 2372
rect -140 1948 -120 2372
rect -892 1920 -120 1948
rect 120 2372 892 2400
rect 120 1948 808 2372
rect 872 1948 892 2372
rect 120 1920 892 1948
rect 1132 2372 1904 2400
rect 1132 1948 1820 2372
rect 1884 1948 1904 2372
rect 1132 1920 1904 1948
rect 2144 2372 2916 2400
rect 2144 1948 2832 2372
rect 2896 1948 2916 2372
rect 2144 1920 2916 1948
rect 3156 2372 3928 2400
rect 3156 1948 3844 2372
rect 3908 1948 3928 2372
rect 3156 1920 3928 1948
rect 4168 2372 4940 2400
rect 4168 1948 4856 2372
rect 4920 1948 4940 2372
rect 4168 1920 4940 1948
rect 5180 2372 5952 2400
rect 5180 1948 5868 2372
rect 5932 1948 5952 2372
rect 5180 1920 5952 1948
rect 6192 2372 6964 2400
rect 6192 1948 6880 2372
rect 6944 1948 6964 2372
rect 6192 1920 6964 1948
rect 7204 2372 7976 2400
rect 7204 1948 7892 2372
rect 7956 1948 7976 2372
rect 7204 1920 7976 1948
rect 8216 2372 8988 2400
rect 8216 1948 8904 2372
rect 8968 1948 8988 2372
rect 8216 1920 8988 1948
rect 9228 2372 10000 2400
rect 9228 1948 9916 2372
rect 9980 1948 10000 2372
rect 9228 1920 10000 1948
rect 10240 2372 11012 2400
rect 10240 1948 10928 2372
rect 10992 1948 11012 2372
rect 10240 1920 11012 1948
rect 11252 2372 12024 2400
rect 11252 1948 11940 2372
rect 12004 1948 12024 2372
rect 11252 1920 12024 1948
rect 12264 2372 13036 2400
rect 12264 1948 12952 2372
rect 13016 1948 13036 2372
rect 12264 1920 13036 1948
rect 13276 2372 14048 2400
rect 13276 1948 13964 2372
rect 14028 1948 14048 2372
rect 13276 1920 14048 1948
rect 14288 2372 15060 2400
rect 14288 1948 14976 2372
rect 15040 1948 15060 2372
rect 14288 1920 15060 1948
rect 15300 2372 16072 2400
rect 15300 1948 15988 2372
rect 16052 1948 16072 2372
rect 15300 1920 16072 1948
rect 16312 2372 17084 2400
rect 16312 1948 17000 2372
rect 17064 1948 17084 2372
rect 16312 1920 17084 1948
rect 17324 2372 18096 2400
rect 17324 1948 18012 2372
rect 18076 1948 18096 2372
rect 17324 1920 18096 1948
rect 18336 2372 19108 2400
rect 18336 1948 19024 2372
rect 19088 1948 19108 2372
rect 18336 1920 19108 1948
rect 19348 2372 20120 2400
rect 19348 1948 20036 2372
rect 20100 1948 20120 2372
rect 19348 1920 20120 1948
rect 20360 2372 21132 2400
rect 20360 1948 21048 2372
rect 21112 1948 21132 2372
rect 20360 1920 21132 1948
rect 21372 2372 22144 2400
rect 21372 1948 22060 2372
rect 22124 1948 22144 2372
rect 21372 1920 22144 1948
rect 22384 2372 23156 2400
rect 22384 1948 23072 2372
rect 23136 1948 23156 2372
rect 22384 1920 23156 1948
rect 23396 2372 24168 2400
rect 23396 1948 24084 2372
rect 24148 1948 24168 2372
rect 23396 1920 24168 1948
rect 24408 2372 25180 2400
rect 24408 1948 25096 2372
rect 25160 1948 25180 2372
rect 24408 1920 25180 1948
rect 25420 2372 26192 2400
rect 25420 1948 26108 2372
rect 26172 1948 26192 2372
rect 25420 1920 26192 1948
rect 26432 2372 27204 2400
rect 26432 1948 27120 2372
rect 27184 1948 27204 2372
rect 26432 1920 27204 1948
rect 27444 2372 28216 2400
rect 27444 1948 28132 2372
rect 28196 1948 28216 2372
rect 27444 1920 28216 1948
rect 28456 2372 29228 2400
rect 28456 1948 29144 2372
rect 29208 1948 29228 2372
rect 28456 1920 29228 1948
rect 29468 2372 30240 2400
rect 29468 1948 30156 2372
rect 30220 1948 30240 2372
rect 29468 1920 30240 1948
rect 30480 2372 31252 2400
rect 30480 1948 31168 2372
rect 31232 1948 31252 2372
rect 30480 1920 31252 1948
rect 31492 2372 32264 2400
rect 31492 1948 32180 2372
rect 32244 1948 32264 2372
rect 31492 1920 32264 1948
rect -32264 1652 -31492 1680
rect -32264 1228 -31576 1652
rect -31512 1228 -31492 1652
rect -32264 1200 -31492 1228
rect -31252 1652 -30480 1680
rect -31252 1228 -30564 1652
rect -30500 1228 -30480 1652
rect -31252 1200 -30480 1228
rect -30240 1652 -29468 1680
rect -30240 1228 -29552 1652
rect -29488 1228 -29468 1652
rect -30240 1200 -29468 1228
rect -29228 1652 -28456 1680
rect -29228 1228 -28540 1652
rect -28476 1228 -28456 1652
rect -29228 1200 -28456 1228
rect -28216 1652 -27444 1680
rect -28216 1228 -27528 1652
rect -27464 1228 -27444 1652
rect -28216 1200 -27444 1228
rect -27204 1652 -26432 1680
rect -27204 1228 -26516 1652
rect -26452 1228 -26432 1652
rect -27204 1200 -26432 1228
rect -26192 1652 -25420 1680
rect -26192 1228 -25504 1652
rect -25440 1228 -25420 1652
rect -26192 1200 -25420 1228
rect -25180 1652 -24408 1680
rect -25180 1228 -24492 1652
rect -24428 1228 -24408 1652
rect -25180 1200 -24408 1228
rect -24168 1652 -23396 1680
rect -24168 1228 -23480 1652
rect -23416 1228 -23396 1652
rect -24168 1200 -23396 1228
rect -23156 1652 -22384 1680
rect -23156 1228 -22468 1652
rect -22404 1228 -22384 1652
rect -23156 1200 -22384 1228
rect -22144 1652 -21372 1680
rect -22144 1228 -21456 1652
rect -21392 1228 -21372 1652
rect -22144 1200 -21372 1228
rect -21132 1652 -20360 1680
rect -21132 1228 -20444 1652
rect -20380 1228 -20360 1652
rect -21132 1200 -20360 1228
rect -20120 1652 -19348 1680
rect -20120 1228 -19432 1652
rect -19368 1228 -19348 1652
rect -20120 1200 -19348 1228
rect -19108 1652 -18336 1680
rect -19108 1228 -18420 1652
rect -18356 1228 -18336 1652
rect -19108 1200 -18336 1228
rect -18096 1652 -17324 1680
rect -18096 1228 -17408 1652
rect -17344 1228 -17324 1652
rect -18096 1200 -17324 1228
rect -17084 1652 -16312 1680
rect -17084 1228 -16396 1652
rect -16332 1228 -16312 1652
rect -17084 1200 -16312 1228
rect -16072 1652 -15300 1680
rect -16072 1228 -15384 1652
rect -15320 1228 -15300 1652
rect -16072 1200 -15300 1228
rect -15060 1652 -14288 1680
rect -15060 1228 -14372 1652
rect -14308 1228 -14288 1652
rect -15060 1200 -14288 1228
rect -14048 1652 -13276 1680
rect -14048 1228 -13360 1652
rect -13296 1228 -13276 1652
rect -14048 1200 -13276 1228
rect -13036 1652 -12264 1680
rect -13036 1228 -12348 1652
rect -12284 1228 -12264 1652
rect -13036 1200 -12264 1228
rect -12024 1652 -11252 1680
rect -12024 1228 -11336 1652
rect -11272 1228 -11252 1652
rect -12024 1200 -11252 1228
rect -11012 1652 -10240 1680
rect -11012 1228 -10324 1652
rect -10260 1228 -10240 1652
rect -11012 1200 -10240 1228
rect -10000 1652 -9228 1680
rect -10000 1228 -9312 1652
rect -9248 1228 -9228 1652
rect -10000 1200 -9228 1228
rect -8988 1652 -8216 1680
rect -8988 1228 -8300 1652
rect -8236 1228 -8216 1652
rect -8988 1200 -8216 1228
rect -7976 1652 -7204 1680
rect -7976 1228 -7288 1652
rect -7224 1228 -7204 1652
rect -7976 1200 -7204 1228
rect -6964 1652 -6192 1680
rect -6964 1228 -6276 1652
rect -6212 1228 -6192 1652
rect -6964 1200 -6192 1228
rect -5952 1652 -5180 1680
rect -5952 1228 -5264 1652
rect -5200 1228 -5180 1652
rect -5952 1200 -5180 1228
rect -4940 1652 -4168 1680
rect -4940 1228 -4252 1652
rect -4188 1228 -4168 1652
rect -4940 1200 -4168 1228
rect -3928 1652 -3156 1680
rect -3928 1228 -3240 1652
rect -3176 1228 -3156 1652
rect -3928 1200 -3156 1228
rect -2916 1652 -2144 1680
rect -2916 1228 -2228 1652
rect -2164 1228 -2144 1652
rect -2916 1200 -2144 1228
rect -1904 1652 -1132 1680
rect -1904 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -1904 1200 -1132 1228
rect -892 1652 -120 1680
rect -892 1228 -204 1652
rect -140 1228 -120 1652
rect -892 1200 -120 1228
rect 120 1652 892 1680
rect 120 1228 808 1652
rect 872 1228 892 1652
rect 120 1200 892 1228
rect 1132 1652 1904 1680
rect 1132 1228 1820 1652
rect 1884 1228 1904 1652
rect 1132 1200 1904 1228
rect 2144 1652 2916 1680
rect 2144 1228 2832 1652
rect 2896 1228 2916 1652
rect 2144 1200 2916 1228
rect 3156 1652 3928 1680
rect 3156 1228 3844 1652
rect 3908 1228 3928 1652
rect 3156 1200 3928 1228
rect 4168 1652 4940 1680
rect 4168 1228 4856 1652
rect 4920 1228 4940 1652
rect 4168 1200 4940 1228
rect 5180 1652 5952 1680
rect 5180 1228 5868 1652
rect 5932 1228 5952 1652
rect 5180 1200 5952 1228
rect 6192 1652 6964 1680
rect 6192 1228 6880 1652
rect 6944 1228 6964 1652
rect 6192 1200 6964 1228
rect 7204 1652 7976 1680
rect 7204 1228 7892 1652
rect 7956 1228 7976 1652
rect 7204 1200 7976 1228
rect 8216 1652 8988 1680
rect 8216 1228 8904 1652
rect 8968 1228 8988 1652
rect 8216 1200 8988 1228
rect 9228 1652 10000 1680
rect 9228 1228 9916 1652
rect 9980 1228 10000 1652
rect 9228 1200 10000 1228
rect 10240 1652 11012 1680
rect 10240 1228 10928 1652
rect 10992 1228 11012 1652
rect 10240 1200 11012 1228
rect 11252 1652 12024 1680
rect 11252 1228 11940 1652
rect 12004 1228 12024 1652
rect 11252 1200 12024 1228
rect 12264 1652 13036 1680
rect 12264 1228 12952 1652
rect 13016 1228 13036 1652
rect 12264 1200 13036 1228
rect 13276 1652 14048 1680
rect 13276 1228 13964 1652
rect 14028 1228 14048 1652
rect 13276 1200 14048 1228
rect 14288 1652 15060 1680
rect 14288 1228 14976 1652
rect 15040 1228 15060 1652
rect 14288 1200 15060 1228
rect 15300 1652 16072 1680
rect 15300 1228 15988 1652
rect 16052 1228 16072 1652
rect 15300 1200 16072 1228
rect 16312 1652 17084 1680
rect 16312 1228 17000 1652
rect 17064 1228 17084 1652
rect 16312 1200 17084 1228
rect 17324 1652 18096 1680
rect 17324 1228 18012 1652
rect 18076 1228 18096 1652
rect 17324 1200 18096 1228
rect 18336 1652 19108 1680
rect 18336 1228 19024 1652
rect 19088 1228 19108 1652
rect 18336 1200 19108 1228
rect 19348 1652 20120 1680
rect 19348 1228 20036 1652
rect 20100 1228 20120 1652
rect 19348 1200 20120 1228
rect 20360 1652 21132 1680
rect 20360 1228 21048 1652
rect 21112 1228 21132 1652
rect 20360 1200 21132 1228
rect 21372 1652 22144 1680
rect 21372 1228 22060 1652
rect 22124 1228 22144 1652
rect 21372 1200 22144 1228
rect 22384 1652 23156 1680
rect 22384 1228 23072 1652
rect 23136 1228 23156 1652
rect 22384 1200 23156 1228
rect 23396 1652 24168 1680
rect 23396 1228 24084 1652
rect 24148 1228 24168 1652
rect 23396 1200 24168 1228
rect 24408 1652 25180 1680
rect 24408 1228 25096 1652
rect 25160 1228 25180 1652
rect 24408 1200 25180 1228
rect 25420 1652 26192 1680
rect 25420 1228 26108 1652
rect 26172 1228 26192 1652
rect 25420 1200 26192 1228
rect 26432 1652 27204 1680
rect 26432 1228 27120 1652
rect 27184 1228 27204 1652
rect 26432 1200 27204 1228
rect 27444 1652 28216 1680
rect 27444 1228 28132 1652
rect 28196 1228 28216 1652
rect 27444 1200 28216 1228
rect 28456 1652 29228 1680
rect 28456 1228 29144 1652
rect 29208 1228 29228 1652
rect 28456 1200 29228 1228
rect 29468 1652 30240 1680
rect 29468 1228 30156 1652
rect 30220 1228 30240 1652
rect 29468 1200 30240 1228
rect 30480 1652 31252 1680
rect 30480 1228 31168 1652
rect 31232 1228 31252 1652
rect 30480 1200 31252 1228
rect 31492 1652 32264 1680
rect 31492 1228 32180 1652
rect 32244 1228 32264 1652
rect 31492 1200 32264 1228
rect -32264 932 -31492 960
rect -32264 508 -31576 932
rect -31512 508 -31492 932
rect -32264 480 -31492 508
rect -31252 932 -30480 960
rect -31252 508 -30564 932
rect -30500 508 -30480 932
rect -31252 480 -30480 508
rect -30240 932 -29468 960
rect -30240 508 -29552 932
rect -29488 508 -29468 932
rect -30240 480 -29468 508
rect -29228 932 -28456 960
rect -29228 508 -28540 932
rect -28476 508 -28456 932
rect -29228 480 -28456 508
rect -28216 932 -27444 960
rect -28216 508 -27528 932
rect -27464 508 -27444 932
rect -28216 480 -27444 508
rect -27204 932 -26432 960
rect -27204 508 -26516 932
rect -26452 508 -26432 932
rect -27204 480 -26432 508
rect -26192 932 -25420 960
rect -26192 508 -25504 932
rect -25440 508 -25420 932
rect -26192 480 -25420 508
rect -25180 932 -24408 960
rect -25180 508 -24492 932
rect -24428 508 -24408 932
rect -25180 480 -24408 508
rect -24168 932 -23396 960
rect -24168 508 -23480 932
rect -23416 508 -23396 932
rect -24168 480 -23396 508
rect -23156 932 -22384 960
rect -23156 508 -22468 932
rect -22404 508 -22384 932
rect -23156 480 -22384 508
rect -22144 932 -21372 960
rect -22144 508 -21456 932
rect -21392 508 -21372 932
rect -22144 480 -21372 508
rect -21132 932 -20360 960
rect -21132 508 -20444 932
rect -20380 508 -20360 932
rect -21132 480 -20360 508
rect -20120 932 -19348 960
rect -20120 508 -19432 932
rect -19368 508 -19348 932
rect -20120 480 -19348 508
rect -19108 932 -18336 960
rect -19108 508 -18420 932
rect -18356 508 -18336 932
rect -19108 480 -18336 508
rect -18096 932 -17324 960
rect -18096 508 -17408 932
rect -17344 508 -17324 932
rect -18096 480 -17324 508
rect -17084 932 -16312 960
rect -17084 508 -16396 932
rect -16332 508 -16312 932
rect -17084 480 -16312 508
rect -16072 932 -15300 960
rect -16072 508 -15384 932
rect -15320 508 -15300 932
rect -16072 480 -15300 508
rect -15060 932 -14288 960
rect -15060 508 -14372 932
rect -14308 508 -14288 932
rect -15060 480 -14288 508
rect -14048 932 -13276 960
rect -14048 508 -13360 932
rect -13296 508 -13276 932
rect -14048 480 -13276 508
rect -13036 932 -12264 960
rect -13036 508 -12348 932
rect -12284 508 -12264 932
rect -13036 480 -12264 508
rect -12024 932 -11252 960
rect -12024 508 -11336 932
rect -11272 508 -11252 932
rect -12024 480 -11252 508
rect -11012 932 -10240 960
rect -11012 508 -10324 932
rect -10260 508 -10240 932
rect -11012 480 -10240 508
rect -10000 932 -9228 960
rect -10000 508 -9312 932
rect -9248 508 -9228 932
rect -10000 480 -9228 508
rect -8988 932 -8216 960
rect -8988 508 -8300 932
rect -8236 508 -8216 932
rect -8988 480 -8216 508
rect -7976 932 -7204 960
rect -7976 508 -7288 932
rect -7224 508 -7204 932
rect -7976 480 -7204 508
rect -6964 932 -6192 960
rect -6964 508 -6276 932
rect -6212 508 -6192 932
rect -6964 480 -6192 508
rect -5952 932 -5180 960
rect -5952 508 -5264 932
rect -5200 508 -5180 932
rect -5952 480 -5180 508
rect -4940 932 -4168 960
rect -4940 508 -4252 932
rect -4188 508 -4168 932
rect -4940 480 -4168 508
rect -3928 932 -3156 960
rect -3928 508 -3240 932
rect -3176 508 -3156 932
rect -3928 480 -3156 508
rect -2916 932 -2144 960
rect -2916 508 -2228 932
rect -2164 508 -2144 932
rect -2916 480 -2144 508
rect -1904 932 -1132 960
rect -1904 508 -1216 932
rect -1152 508 -1132 932
rect -1904 480 -1132 508
rect -892 932 -120 960
rect -892 508 -204 932
rect -140 508 -120 932
rect -892 480 -120 508
rect 120 932 892 960
rect 120 508 808 932
rect 872 508 892 932
rect 120 480 892 508
rect 1132 932 1904 960
rect 1132 508 1820 932
rect 1884 508 1904 932
rect 1132 480 1904 508
rect 2144 932 2916 960
rect 2144 508 2832 932
rect 2896 508 2916 932
rect 2144 480 2916 508
rect 3156 932 3928 960
rect 3156 508 3844 932
rect 3908 508 3928 932
rect 3156 480 3928 508
rect 4168 932 4940 960
rect 4168 508 4856 932
rect 4920 508 4940 932
rect 4168 480 4940 508
rect 5180 932 5952 960
rect 5180 508 5868 932
rect 5932 508 5952 932
rect 5180 480 5952 508
rect 6192 932 6964 960
rect 6192 508 6880 932
rect 6944 508 6964 932
rect 6192 480 6964 508
rect 7204 932 7976 960
rect 7204 508 7892 932
rect 7956 508 7976 932
rect 7204 480 7976 508
rect 8216 932 8988 960
rect 8216 508 8904 932
rect 8968 508 8988 932
rect 8216 480 8988 508
rect 9228 932 10000 960
rect 9228 508 9916 932
rect 9980 508 10000 932
rect 9228 480 10000 508
rect 10240 932 11012 960
rect 10240 508 10928 932
rect 10992 508 11012 932
rect 10240 480 11012 508
rect 11252 932 12024 960
rect 11252 508 11940 932
rect 12004 508 12024 932
rect 11252 480 12024 508
rect 12264 932 13036 960
rect 12264 508 12952 932
rect 13016 508 13036 932
rect 12264 480 13036 508
rect 13276 932 14048 960
rect 13276 508 13964 932
rect 14028 508 14048 932
rect 13276 480 14048 508
rect 14288 932 15060 960
rect 14288 508 14976 932
rect 15040 508 15060 932
rect 14288 480 15060 508
rect 15300 932 16072 960
rect 15300 508 15988 932
rect 16052 508 16072 932
rect 15300 480 16072 508
rect 16312 932 17084 960
rect 16312 508 17000 932
rect 17064 508 17084 932
rect 16312 480 17084 508
rect 17324 932 18096 960
rect 17324 508 18012 932
rect 18076 508 18096 932
rect 17324 480 18096 508
rect 18336 932 19108 960
rect 18336 508 19024 932
rect 19088 508 19108 932
rect 18336 480 19108 508
rect 19348 932 20120 960
rect 19348 508 20036 932
rect 20100 508 20120 932
rect 19348 480 20120 508
rect 20360 932 21132 960
rect 20360 508 21048 932
rect 21112 508 21132 932
rect 20360 480 21132 508
rect 21372 932 22144 960
rect 21372 508 22060 932
rect 22124 508 22144 932
rect 21372 480 22144 508
rect 22384 932 23156 960
rect 22384 508 23072 932
rect 23136 508 23156 932
rect 22384 480 23156 508
rect 23396 932 24168 960
rect 23396 508 24084 932
rect 24148 508 24168 932
rect 23396 480 24168 508
rect 24408 932 25180 960
rect 24408 508 25096 932
rect 25160 508 25180 932
rect 24408 480 25180 508
rect 25420 932 26192 960
rect 25420 508 26108 932
rect 26172 508 26192 932
rect 25420 480 26192 508
rect 26432 932 27204 960
rect 26432 508 27120 932
rect 27184 508 27204 932
rect 26432 480 27204 508
rect 27444 932 28216 960
rect 27444 508 28132 932
rect 28196 508 28216 932
rect 27444 480 28216 508
rect 28456 932 29228 960
rect 28456 508 29144 932
rect 29208 508 29228 932
rect 28456 480 29228 508
rect 29468 932 30240 960
rect 29468 508 30156 932
rect 30220 508 30240 932
rect 29468 480 30240 508
rect 30480 932 31252 960
rect 30480 508 31168 932
rect 31232 508 31252 932
rect 30480 480 31252 508
rect 31492 932 32264 960
rect 31492 508 32180 932
rect 32244 508 32264 932
rect 31492 480 32264 508
rect -32264 212 -31492 240
rect -32264 -212 -31576 212
rect -31512 -212 -31492 212
rect -32264 -240 -31492 -212
rect -31252 212 -30480 240
rect -31252 -212 -30564 212
rect -30500 -212 -30480 212
rect -31252 -240 -30480 -212
rect -30240 212 -29468 240
rect -30240 -212 -29552 212
rect -29488 -212 -29468 212
rect -30240 -240 -29468 -212
rect -29228 212 -28456 240
rect -29228 -212 -28540 212
rect -28476 -212 -28456 212
rect -29228 -240 -28456 -212
rect -28216 212 -27444 240
rect -28216 -212 -27528 212
rect -27464 -212 -27444 212
rect -28216 -240 -27444 -212
rect -27204 212 -26432 240
rect -27204 -212 -26516 212
rect -26452 -212 -26432 212
rect -27204 -240 -26432 -212
rect -26192 212 -25420 240
rect -26192 -212 -25504 212
rect -25440 -212 -25420 212
rect -26192 -240 -25420 -212
rect -25180 212 -24408 240
rect -25180 -212 -24492 212
rect -24428 -212 -24408 212
rect -25180 -240 -24408 -212
rect -24168 212 -23396 240
rect -24168 -212 -23480 212
rect -23416 -212 -23396 212
rect -24168 -240 -23396 -212
rect -23156 212 -22384 240
rect -23156 -212 -22468 212
rect -22404 -212 -22384 212
rect -23156 -240 -22384 -212
rect -22144 212 -21372 240
rect -22144 -212 -21456 212
rect -21392 -212 -21372 212
rect -22144 -240 -21372 -212
rect -21132 212 -20360 240
rect -21132 -212 -20444 212
rect -20380 -212 -20360 212
rect -21132 -240 -20360 -212
rect -20120 212 -19348 240
rect -20120 -212 -19432 212
rect -19368 -212 -19348 212
rect -20120 -240 -19348 -212
rect -19108 212 -18336 240
rect -19108 -212 -18420 212
rect -18356 -212 -18336 212
rect -19108 -240 -18336 -212
rect -18096 212 -17324 240
rect -18096 -212 -17408 212
rect -17344 -212 -17324 212
rect -18096 -240 -17324 -212
rect -17084 212 -16312 240
rect -17084 -212 -16396 212
rect -16332 -212 -16312 212
rect -17084 -240 -16312 -212
rect -16072 212 -15300 240
rect -16072 -212 -15384 212
rect -15320 -212 -15300 212
rect -16072 -240 -15300 -212
rect -15060 212 -14288 240
rect -15060 -212 -14372 212
rect -14308 -212 -14288 212
rect -15060 -240 -14288 -212
rect -14048 212 -13276 240
rect -14048 -212 -13360 212
rect -13296 -212 -13276 212
rect -14048 -240 -13276 -212
rect -13036 212 -12264 240
rect -13036 -212 -12348 212
rect -12284 -212 -12264 212
rect -13036 -240 -12264 -212
rect -12024 212 -11252 240
rect -12024 -212 -11336 212
rect -11272 -212 -11252 212
rect -12024 -240 -11252 -212
rect -11012 212 -10240 240
rect -11012 -212 -10324 212
rect -10260 -212 -10240 212
rect -11012 -240 -10240 -212
rect -10000 212 -9228 240
rect -10000 -212 -9312 212
rect -9248 -212 -9228 212
rect -10000 -240 -9228 -212
rect -8988 212 -8216 240
rect -8988 -212 -8300 212
rect -8236 -212 -8216 212
rect -8988 -240 -8216 -212
rect -7976 212 -7204 240
rect -7976 -212 -7288 212
rect -7224 -212 -7204 212
rect -7976 -240 -7204 -212
rect -6964 212 -6192 240
rect -6964 -212 -6276 212
rect -6212 -212 -6192 212
rect -6964 -240 -6192 -212
rect -5952 212 -5180 240
rect -5952 -212 -5264 212
rect -5200 -212 -5180 212
rect -5952 -240 -5180 -212
rect -4940 212 -4168 240
rect -4940 -212 -4252 212
rect -4188 -212 -4168 212
rect -4940 -240 -4168 -212
rect -3928 212 -3156 240
rect -3928 -212 -3240 212
rect -3176 -212 -3156 212
rect -3928 -240 -3156 -212
rect -2916 212 -2144 240
rect -2916 -212 -2228 212
rect -2164 -212 -2144 212
rect -2916 -240 -2144 -212
rect -1904 212 -1132 240
rect -1904 -212 -1216 212
rect -1152 -212 -1132 212
rect -1904 -240 -1132 -212
rect -892 212 -120 240
rect -892 -212 -204 212
rect -140 -212 -120 212
rect -892 -240 -120 -212
rect 120 212 892 240
rect 120 -212 808 212
rect 872 -212 892 212
rect 120 -240 892 -212
rect 1132 212 1904 240
rect 1132 -212 1820 212
rect 1884 -212 1904 212
rect 1132 -240 1904 -212
rect 2144 212 2916 240
rect 2144 -212 2832 212
rect 2896 -212 2916 212
rect 2144 -240 2916 -212
rect 3156 212 3928 240
rect 3156 -212 3844 212
rect 3908 -212 3928 212
rect 3156 -240 3928 -212
rect 4168 212 4940 240
rect 4168 -212 4856 212
rect 4920 -212 4940 212
rect 4168 -240 4940 -212
rect 5180 212 5952 240
rect 5180 -212 5868 212
rect 5932 -212 5952 212
rect 5180 -240 5952 -212
rect 6192 212 6964 240
rect 6192 -212 6880 212
rect 6944 -212 6964 212
rect 6192 -240 6964 -212
rect 7204 212 7976 240
rect 7204 -212 7892 212
rect 7956 -212 7976 212
rect 7204 -240 7976 -212
rect 8216 212 8988 240
rect 8216 -212 8904 212
rect 8968 -212 8988 212
rect 8216 -240 8988 -212
rect 9228 212 10000 240
rect 9228 -212 9916 212
rect 9980 -212 10000 212
rect 9228 -240 10000 -212
rect 10240 212 11012 240
rect 10240 -212 10928 212
rect 10992 -212 11012 212
rect 10240 -240 11012 -212
rect 11252 212 12024 240
rect 11252 -212 11940 212
rect 12004 -212 12024 212
rect 11252 -240 12024 -212
rect 12264 212 13036 240
rect 12264 -212 12952 212
rect 13016 -212 13036 212
rect 12264 -240 13036 -212
rect 13276 212 14048 240
rect 13276 -212 13964 212
rect 14028 -212 14048 212
rect 13276 -240 14048 -212
rect 14288 212 15060 240
rect 14288 -212 14976 212
rect 15040 -212 15060 212
rect 14288 -240 15060 -212
rect 15300 212 16072 240
rect 15300 -212 15988 212
rect 16052 -212 16072 212
rect 15300 -240 16072 -212
rect 16312 212 17084 240
rect 16312 -212 17000 212
rect 17064 -212 17084 212
rect 16312 -240 17084 -212
rect 17324 212 18096 240
rect 17324 -212 18012 212
rect 18076 -212 18096 212
rect 17324 -240 18096 -212
rect 18336 212 19108 240
rect 18336 -212 19024 212
rect 19088 -212 19108 212
rect 18336 -240 19108 -212
rect 19348 212 20120 240
rect 19348 -212 20036 212
rect 20100 -212 20120 212
rect 19348 -240 20120 -212
rect 20360 212 21132 240
rect 20360 -212 21048 212
rect 21112 -212 21132 212
rect 20360 -240 21132 -212
rect 21372 212 22144 240
rect 21372 -212 22060 212
rect 22124 -212 22144 212
rect 21372 -240 22144 -212
rect 22384 212 23156 240
rect 22384 -212 23072 212
rect 23136 -212 23156 212
rect 22384 -240 23156 -212
rect 23396 212 24168 240
rect 23396 -212 24084 212
rect 24148 -212 24168 212
rect 23396 -240 24168 -212
rect 24408 212 25180 240
rect 24408 -212 25096 212
rect 25160 -212 25180 212
rect 24408 -240 25180 -212
rect 25420 212 26192 240
rect 25420 -212 26108 212
rect 26172 -212 26192 212
rect 25420 -240 26192 -212
rect 26432 212 27204 240
rect 26432 -212 27120 212
rect 27184 -212 27204 212
rect 26432 -240 27204 -212
rect 27444 212 28216 240
rect 27444 -212 28132 212
rect 28196 -212 28216 212
rect 27444 -240 28216 -212
rect 28456 212 29228 240
rect 28456 -212 29144 212
rect 29208 -212 29228 212
rect 28456 -240 29228 -212
rect 29468 212 30240 240
rect 29468 -212 30156 212
rect 30220 -212 30240 212
rect 29468 -240 30240 -212
rect 30480 212 31252 240
rect 30480 -212 31168 212
rect 31232 -212 31252 212
rect 30480 -240 31252 -212
rect 31492 212 32264 240
rect 31492 -212 32180 212
rect 32244 -212 32264 212
rect 31492 -240 32264 -212
rect -32264 -508 -31492 -480
rect -32264 -932 -31576 -508
rect -31512 -932 -31492 -508
rect -32264 -960 -31492 -932
rect -31252 -508 -30480 -480
rect -31252 -932 -30564 -508
rect -30500 -932 -30480 -508
rect -31252 -960 -30480 -932
rect -30240 -508 -29468 -480
rect -30240 -932 -29552 -508
rect -29488 -932 -29468 -508
rect -30240 -960 -29468 -932
rect -29228 -508 -28456 -480
rect -29228 -932 -28540 -508
rect -28476 -932 -28456 -508
rect -29228 -960 -28456 -932
rect -28216 -508 -27444 -480
rect -28216 -932 -27528 -508
rect -27464 -932 -27444 -508
rect -28216 -960 -27444 -932
rect -27204 -508 -26432 -480
rect -27204 -932 -26516 -508
rect -26452 -932 -26432 -508
rect -27204 -960 -26432 -932
rect -26192 -508 -25420 -480
rect -26192 -932 -25504 -508
rect -25440 -932 -25420 -508
rect -26192 -960 -25420 -932
rect -25180 -508 -24408 -480
rect -25180 -932 -24492 -508
rect -24428 -932 -24408 -508
rect -25180 -960 -24408 -932
rect -24168 -508 -23396 -480
rect -24168 -932 -23480 -508
rect -23416 -932 -23396 -508
rect -24168 -960 -23396 -932
rect -23156 -508 -22384 -480
rect -23156 -932 -22468 -508
rect -22404 -932 -22384 -508
rect -23156 -960 -22384 -932
rect -22144 -508 -21372 -480
rect -22144 -932 -21456 -508
rect -21392 -932 -21372 -508
rect -22144 -960 -21372 -932
rect -21132 -508 -20360 -480
rect -21132 -932 -20444 -508
rect -20380 -932 -20360 -508
rect -21132 -960 -20360 -932
rect -20120 -508 -19348 -480
rect -20120 -932 -19432 -508
rect -19368 -932 -19348 -508
rect -20120 -960 -19348 -932
rect -19108 -508 -18336 -480
rect -19108 -932 -18420 -508
rect -18356 -932 -18336 -508
rect -19108 -960 -18336 -932
rect -18096 -508 -17324 -480
rect -18096 -932 -17408 -508
rect -17344 -932 -17324 -508
rect -18096 -960 -17324 -932
rect -17084 -508 -16312 -480
rect -17084 -932 -16396 -508
rect -16332 -932 -16312 -508
rect -17084 -960 -16312 -932
rect -16072 -508 -15300 -480
rect -16072 -932 -15384 -508
rect -15320 -932 -15300 -508
rect -16072 -960 -15300 -932
rect -15060 -508 -14288 -480
rect -15060 -932 -14372 -508
rect -14308 -932 -14288 -508
rect -15060 -960 -14288 -932
rect -14048 -508 -13276 -480
rect -14048 -932 -13360 -508
rect -13296 -932 -13276 -508
rect -14048 -960 -13276 -932
rect -13036 -508 -12264 -480
rect -13036 -932 -12348 -508
rect -12284 -932 -12264 -508
rect -13036 -960 -12264 -932
rect -12024 -508 -11252 -480
rect -12024 -932 -11336 -508
rect -11272 -932 -11252 -508
rect -12024 -960 -11252 -932
rect -11012 -508 -10240 -480
rect -11012 -932 -10324 -508
rect -10260 -932 -10240 -508
rect -11012 -960 -10240 -932
rect -10000 -508 -9228 -480
rect -10000 -932 -9312 -508
rect -9248 -932 -9228 -508
rect -10000 -960 -9228 -932
rect -8988 -508 -8216 -480
rect -8988 -932 -8300 -508
rect -8236 -932 -8216 -508
rect -8988 -960 -8216 -932
rect -7976 -508 -7204 -480
rect -7976 -932 -7288 -508
rect -7224 -932 -7204 -508
rect -7976 -960 -7204 -932
rect -6964 -508 -6192 -480
rect -6964 -932 -6276 -508
rect -6212 -932 -6192 -508
rect -6964 -960 -6192 -932
rect -5952 -508 -5180 -480
rect -5952 -932 -5264 -508
rect -5200 -932 -5180 -508
rect -5952 -960 -5180 -932
rect -4940 -508 -4168 -480
rect -4940 -932 -4252 -508
rect -4188 -932 -4168 -508
rect -4940 -960 -4168 -932
rect -3928 -508 -3156 -480
rect -3928 -932 -3240 -508
rect -3176 -932 -3156 -508
rect -3928 -960 -3156 -932
rect -2916 -508 -2144 -480
rect -2916 -932 -2228 -508
rect -2164 -932 -2144 -508
rect -2916 -960 -2144 -932
rect -1904 -508 -1132 -480
rect -1904 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -1904 -960 -1132 -932
rect -892 -508 -120 -480
rect -892 -932 -204 -508
rect -140 -932 -120 -508
rect -892 -960 -120 -932
rect 120 -508 892 -480
rect 120 -932 808 -508
rect 872 -932 892 -508
rect 120 -960 892 -932
rect 1132 -508 1904 -480
rect 1132 -932 1820 -508
rect 1884 -932 1904 -508
rect 1132 -960 1904 -932
rect 2144 -508 2916 -480
rect 2144 -932 2832 -508
rect 2896 -932 2916 -508
rect 2144 -960 2916 -932
rect 3156 -508 3928 -480
rect 3156 -932 3844 -508
rect 3908 -932 3928 -508
rect 3156 -960 3928 -932
rect 4168 -508 4940 -480
rect 4168 -932 4856 -508
rect 4920 -932 4940 -508
rect 4168 -960 4940 -932
rect 5180 -508 5952 -480
rect 5180 -932 5868 -508
rect 5932 -932 5952 -508
rect 5180 -960 5952 -932
rect 6192 -508 6964 -480
rect 6192 -932 6880 -508
rect 6944 -932 6964 -508
rect 6192 -960 6964 -932
rect 7204 -508 7976 -480
rect 7204 -932 7892 -508
rect 7956 -932 7976 -508
rect 7204 -960 7976 -932
rect 8216 -508 8988 -480
rect 8216 -932 8904 -508
rect 8968 -932 8988 -508
rect 8216 -960 8988 -932
rect 9228 -508 10000 -480
rect 9228 -932 9916 -508
rect 9980 -932 10000 -508
rect 9228 -960 10000 -932
rect 10240 -508 11012 -480
rect 10240 -932 10928 -508
rect 10992 -932 11012 -508
rect 10240 -960 11012 -932
rect 11252 -508 12024 -480
rect 11252 -932 11940 -508
rect 12004 -932 12024 -508
rect 11252 -960 12024 -932
rect 12264 -508 13036 -480
rect 12264 -932 12952 -508
rect 13016 -932 13036 -508
rect 12264 -960 13036 -932
rect 13276 -508 14048 -480
rect 13276 -932 13964 -508
rect 14028 -932 14048 -508
rect 13276 -960 14048 -932
rect 14288 -508 15060 -480
rect 14288 -932 14976 -508
rect 15040 -932 15060 -508
rect 14288 -960 15060 -932
rect 15300 -508 16072 -480
rect 15300 -932 15988 -508
rect 16052 -932 16072 -508
rect 15300 -960 16072 -932
rect 16312 -508 17084 -480
rect 16312 -932 17000 -508
rect 17064 -932 17084 -508
rect 16312 -960 17084 -932
rect 17324 -508 18096 -480
rect 17324 -932 18012 -508
rect 18076 -932 18096 -508
rect 17324 -960 18096 -932
rect 18336 -508 19108 -480
rect 18336 -932 19024 -508
rect 19088 -932 19108 -508
rect 18336 -960 19108 -932
rect 19348 -508 20120 -480
rect 19348 -932 20036 -508
rect 20100 -932 20120 -508
rect 19348 -960 20120 -932
rect 20360 -508 21132 -480
rect 20360 -932 21048 -508
rect 21112 -932 21132 -508
rect 20360 -960 21132 -932
rect 21372 -508 22144 -480
rect 21372 -932 22060 -508
rect 22124 -932 22144 -508
rect 21372 -960 22144 -932
rect 22384 -508 23156 -480
rect 22384 -932 23072 -508
rect 23136 -932 23156 -508
rect 22384 -960 23156 -932
rect 23396 -508 24168 -480
rect 23396 -932 24084 -508
rect 24148 -932 24168 -508
rect 23396 -960 24168 -932
rect 24408 -508 25180 -480
rect 24408 -932 25096 -508
rect 25160 -932 25180 -508
rect 24408 -960 25180 -932
rect 25420 -508 26192 -480
rect 25420 -932 26108 -508
rect 26172 -932 26192 -508
rect 25420 -960 26192 -932
rect 26432 -508 27204 -480
rect 26432 -932 27120 -508
rect 27184 -932 27204 -508
rect 26432 -960 27204 -932
rect 27444 -508 28216 -480
rect 27444 -932 28132 -508
rect 28196 -932 28216 -508
rect 27444 -960 28216 -932
rect 28456 -508 29228 -480
rect 28456 -932 29144 -508
rect 29208 -932 29228 -508
rect 28456 -960 29228 -932
rect 29468 -508 30240 -480
rect 29468 -932 30156 -508
rect 30220 -932 30240 -508
rect 29468 -960 30240 -932
rect 30480 -508 31252 -480
rect 30480 -932 31168 -508
rect 31232 -932 31252 -508
rect 30480 -960 31252 -932
rect 31492 -508 32264 -480
rect 31492 -932 32180 -508
rect 32244 -932 32264 -508
rect 31492 -960 32264 -932
rect -32264 -1228 -31492 -1200
rect -32264 -1652 -31576 -1228
rect -31512 -1652 -31492 -1228
rect -32264 -1680 -31492 -1652
rect -31252 -1228 -30480 -1200
rect -31252 -1652 -30564 -1228
rect -30500 -1652 -30480 -1228
rect -31252 -1680 -30480 -1652
rect -30240 -1228 -29468 -1200
rect -30240 -1652 -29552 -1228
rect -29488 -1652 -29468 -1228
rect -30240 -1680 -29468 -1652
rect -29228 -1228 -28456 -1200
rect -29228 -1652 -28540 -1228
rect -28476 -1652 -28456 -1228
rect -29228 -1680 -28456 -1652
rect -28216 -1228 -27444 -1200
rect -28216 -1652 -27528 -1228
rect -27464 -1652 -27444 -1228
rect -28216 -1680 -27444 -1652
rect -27204 -1228 -26432 -1200
rect -27204 -1652 -26516 -1228
rect -26452 -1652 -26432 -1228
rect -27204 -1680 -26432 -1652
rect -26192 -1228 -25420 -1200
rect -26192 -1652 -25504 -1228
rect -25440 -1652 -25420 -1228
rect -26192 -1680 -25420 -1652
rect -25180 -1228 -24408 -1200
rect -25180 -1652 -24492 -1228
rect -24428 -1652 -24408 -1228
rect -25180 -1680 -24408 -1652
rect -24168 -1228 -23396 -1200
rect -24168 -1652 -23480 -1228
rect -23416 -1652 -23396 -1228
rect -24168 -1680 -23396 -1652
rect -23156 -1228 -22384 -1200
rect -23156 -1652 -22468 -1228
rect -22404 -1652 -22384 -1228
rect -23156 -1680 -22384 -1652
rect -22144 -1228 -21372 -1200
rect -22144 -1652 -21456 -1228
rect -21392 -1652 -21372 -1228
rect -22144 -1680 -21372 -1652
rect -21132 -1228 -20360 -1200
rect -21132 -1652 -20444 -1228
rect -20380 -1652 -20360 -1228
rect -21132 -1680 -20360 -1652
rect -20120 -1228 -19348 -1200
rect -20120 -1652 -19432 -1228
rect -19368 -1652 -19348 -1228
rect -20120 -1680 -19348 -1652
rect -19108 -1228 -18336 -1200
rect -19108 -1652 -18420 -1228
rect -18356 -1652 -18336 -1228
rect -19108 -1680 -18336 -1652
rect -18096 -1228 -17324 -1200
rect -18096 -1652 -17408 -1228
rect -17344 -1652 -17324 -1228
rect -18096 -1680 -17324 -1652
rect -17084 -1228 -16312 -1200
rect -17084 -1652 -16396 -1228
rect -16332 -1652 -16312 -1228
rect -17084 -1680 -16312 -1652
rect -16072 -1228 -15300 -1200
rect -16072 -1652 -15384 -1228
rect -15320 -1652 -15300 -1228
rect -16072 -1680 -15300 -1652
rect -15060 -1228 -14288 -1200
rect -15060 -1652 -14372 -1228
rect -14308 -1652 -14288 -1228
rect -15060 -1680 -14288 -1652
rect -14048 -1228 -13276 -1200
rect -14048 -1652 -13360 -1228
rect -13296 -1652 -13276 -1228
rect -14048 -1680 -13276 -1652
rect -13036 -1228 -12264 -1200
rect -13036 -1652 -12348 -1228
rect -12284 -1652 -12264 -1228
rect -13036 -1680 -12264 -1652
rect -12024 -1228 -11252 -1200
rect -12024 -1652 -11336 -1228
rect -11272 -1652 -11252 -1228
rect -12024 -1680 -11252 -1652
rect -11012 -1228 -10240 -1200
rect -11012 -1652 -10324 -1228
rect -10260 -1652 -10240 -1228
rect -11012 -1680 -10240 -1652
rect -10000 -1228 -9228 -1200
rect -10000 -1652 -9312 -1228
rect -9248 -1652 -9228 -1228
rect -10000 -1680 -9228 -1652
rect -8988 -1228 -8216 -1200
rect -8988 -1652 -8300 -1228
rect -8236 -1652 -8216 -1228
rect -8988 -1680 -8216 -1652
rect -7976 -1228 -7204 -1200
rect -7976 -1652 -7288 -1228
rect -7224 -1652 -7204 -1228
rect -7976 -1680 -7204 -1652
rect -6964 -1228 -6192 -1200
rect -6964 -1652 -6276 -1228
rect -6212 -1652 -6192 -1228
rect -6964 -1680 -6192 -1652
rect -5952 -1228 -5180 -1200
rect -5952 -1652 -5264 -1228
rect -5200 -1652 -5180 -1228
rect -5952 -1680 -5180 -1652
rect -4940 -1228 -4168 -1200
rect -4940 -1652 -4252 -1228
rect -4188 -1652 -4168 -1228
rect -4940 -1680 -4168 -1652
rect -3928 -1228 -3156 -1200
rect -3928 -1652 -3240 -1228
rect -3176 -1652 -3156 -1228
rect -3928 -1680 -3156 -1652
rect -2916 -1228 -2144 -1200
rect -2916 -1652 -2228 -1228
rect -2164 -1652 -2144 -1228
rect -2916 -1680 -2144 -1652
rect -1904 -1228 -1132 -1200
rect -1904 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -1904 -1680 -1132 -1652
rect -892 -1228 -120 -1200
rect -892 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect -892 -1680 -120 -1652
rect 120 -1228 892 -1200
rect 120 -1652 808 -1228
rect 872 -1652 892 -1228
rect 120 -1680 892 -1652
rect 1132 -1228 1904 -1200
rect 1132 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 1132 -1680 1904 -1652
rect 2144 -1228 2916 -1200
rect 2144 -1652 2832 -1228
rect 2896 -1652 2916 -1228
rect 2144 -1680 2916 -1652
rect 3156 -1228 3928 -1200
rect 3156 -1652 3844 -1228
rect 3908 -1652 3928 -1228
rect 3156 -1680 3928 -1652
rect 4168 -1228 4940 -1200
rect 4168 -1652 4856 -1228
rect 4920 -1652 4940 -1228
rect 4168 -1680 4940 -1652
rect 5180 -1228 5952 -1200
rect 5180 -1652 5868 -1228
rect 5932 -1652 5952 -1228
rect 5180 -1680 5952 -1652
rect 6192 -1228 6964 -1200
rect 6192 -1652 6880 -1228
rect 6944 -1652 6964 -1228
rect 6192 -1680 6964 -1652
rect 7204 -1228 7976 -1200
rect 7204 -1652 7892 -1228
rect 7956 -1652 7976 -1228
rect 7204 -1680 7976 -1652
rect 8216 -1228 8988 -1200
rect 8216 -1652 8904 -1228
rect 8968 -1652 8988 -1228
rect 8216 -1680 8988 -1652
rect 9228 -1228 10000 -1200
rect 9228 -1652 9916 -1228
rect 9980 -1652 10000 -1228
rect 9228 -1680 10000 -1652
rect 10240 -1228 11012 -1200
rect 10240 -1652 10928 -1228
rect 10992 -1652 11012 -1228
rect 10240 -1680 11012 -1652
rect 11252 -1228 12024 -1200
rect 11252 -1652 11940 -1228
rect 12004 -1652 12024 -1228
rect 11252 -1680 12024 -1652
rect 12264 -1228 13036 -1200
rect 12264 -1652 12952 -1228
rect 13016 -1652 13036 -1228
rect 12264 -1680 13036 -1652
rect 13276 -1228 14048 -1200
rect 13276 -1652 13964 -1228
rect 14028 -1652 14048 -1228
rect 13276 -1680 14048 -1652
rect 14288 -1228 15060 -1200
rect 14288 -1652 14976 -1228
rect 15040 -1652 15060 -1228
rect 14288 -1680 15060 -1652
rect 15300 -1228 16072 -1200
rect 15300 -1652 15988 -1228
rect 16052 -1652 16072 -1228
rect 15300 -1680 16072 -1652
rect 16312 -1228 17084 -1200
rect 16312 -1652 17000 -1228
rect 17064 -1652 17084 -1228
rect 16312 -1680 17084 -1652
rect 17324 -1228 18096 -1200
rect 17324 -1652 18012 -1228
rect 18076 -1652 18096 -1228
rect 17324 -1680 18096 -1652
rect 18336 -1228 19108 -1200
rect 18336 -1652 19024 -1228
rect 19088 -1652 19108 -1228
rect 18336 -1680 19108 -1652
rect 19348 -1228 20120 -1200
rect 19348 -1652 20036 -1228
rect 20100 -1652 20120 -1228
rect 19348 -1680 20120 -1652
rect 20360 -1228 21132 -1200
rect 20360 -1652 21048 -1228
rect 21112 -1652 21132 -1228
rect 20360 -1680 21132 -1652
rect 21372 -1228 22144 -1200
rect 21372 -1652 22060 -1228
rect 22124 -1652 22144 -1228
rect 21372 -1680 22144 -1652
rect 22384 -1228 23156 -1200
rect 22384 -1652 23072 -1228
rect 23136 -1652 23156 -1228
rect 22384 -1680 23156 -1652
rect 23396 -1228 24168 -1200
rect 23396 -1652 24084 -1228
rect 24148 -1652 24168 -1228
rect 23396 -1680 24168 -1652
rect 24408 -1228 25180 -1200
rect 24408 -1652 25096 -1228
rect 25160 -1652 25180 -1228
rect 24408 -1680 25180 -1652
rect 25420 -1228 26192 -1200
rect 25420 -1652 26108 -1228
rect 26172 -1652 26192 -1228
rect 25420 -1680 26192 -1652
rect 26432 -1228 27204 -1200
rect 26432 -1652 27120 -1228
rect 27184 -1652 27204 -1228
rect 26432 -1680 27204 -1652
rect 27444 -1228 28216 -1200
rect 27444 -1652 28132 -1228
rect 28196 -1652 28216 -1228
rect 27444 -1680 28216 -1652
rect 28456 -1228 29228 -1200
rect 28456 -1652 29144 -1228
rect 29208 -1652 29228 -1228
rect 28456 -1680 29228 -1652
rect 29468 -1228 30240 -1200
rect 29468 -1652 30156 -1228
rect 30220 -1652 30240 -1228
rect 29468 -1680 30240 -1652
rect 30480 -1228 31252 -1200
rect 30480 -1652 31168 -1228
rect 31232 -1652 31252 -1228
rect 30480 -1680 31252 -1652
rect 31492 -1228 32264 -1200
rect 31492 -1652 32180 -1228
rect 32244 -1652 32264 -1228
rect 31492 -1680 32264 -1652
rect -32264 -1948 -31492 -1920
rect -32264 -2372 -31576 -1948
rect -31512 -2372 -31492 -1948
rect -32264 -2400 -31492 -2372
rect -31252 -1948 -30480 -1920
rect -31252 -2372 -30564 -1948
rect -30500 -2372 -30480 -1948
rect -31252 -2400 -30480 -2372
rect -30240 -1948 -29468 -1920
rect -30240 -2372 -29552 -1948
rect -29488 -2372 -29468 -1948
rect -30240 -2400 -29468 -2372
rect -29228 -1948 -28456 -1920
rect -29228 -2372 -28540 -1948
rect -28476 -2372 -28456 -1948
rect -29228 -2400 -28456 -2372
rect -28216 -1948 -27444 -1920
rect -28216 -2372 -27528 -1948
rect -27464 -2372 -27444 -1948
rect -28216 -2400 -27444 -2372
rect -27204 -1948 -26432 -1920
rect -27204 -2372 -26516 -1948
rect -26452 -2372 -26432 -1948
rect -27204 -2400 -26432 -2372
rect -26192 -1948 -25420 -1920
rect -26192 -2372 -25504 -1948
rect -25440 -2372 -25420 -1948
rect -26192 -2400 -25420 -2372
rect -25180 -1948 -24408 -1920
rect -25180 -2372 -24492 -1948
rect -24428 -2372 -24408 -1948
rect -25180 -2400 -24408 -2372
rect -24168 -1948 -23396 -1920
rect -24168 -2372 -23480 -1948
rect -23416 -2372 -23396 -1948
rect -24168 -2400 -23396 -2372
rect -23156 -1948 -22384 -1920
rect -23156 -2372 -22468 -1948
rect -22404 -2372 -22384 -1948
rect -23156 -2400 -22384 -2372
rect -22144 -1948 -21372 -1920
rect -22144 -2372 -21456 -1948
rect -21392 -2372 -21372 -1948
rect -22144 -2400 -21372 -2372
rect -21132 -1948 -20360 -1920
rect -21132 -2372 -20444 -1948
rect -20380 -2372 -20360 -1948
rect -21132 -2400 -20360 -2372
rect -20120 -1948 -19348 -1920
rect -20120 -2372 -19432 -1948
rect -19368 -2372 -19348 -1948
rect -20120 -2400 -19348 -2372
rect -19108 -1948 -18336 -1920
rect -19108 -2372 -18420 -1948
rect -18356 -2372 -18336 -1948
rect -19108 -2400 -18336 -2372
rect -18096 -1948 -17324 -1920
rect -18096 -2372 -17408 -1948
rect -17344 -2372 -17324 -1948
rect -18096 -2400 -17324 -2372
rect -17084 -1948 -16312 -1920
rect -17084 -2372 -16396 -1948
rect -16332 -2372 -16312 -1948
rect -17084 -2400 -16312 -2372
rect -16072 -1948 -15300 -1920
rect -16072 -2372 -15384 -1948
rect -15320 -2372 -15300 -1948
rect -16072 -2400 -15300 -2372
rect -15060 -1948 -14288 -1920
rect -15060 -2372 -14372 -1948
rect -14308 -2372 -14288 -1948
rect -15060 -2400 -14288 -2372
rect -14048 -1948 -13276 -1920
rect -14048 -2372 -13360 -1948
rect -13296 -2372 -13276 -1948
rect -14048 -2400 -13276 -2372
rect -13036 -1948 -12264 -1920
rect -13036 -2372 -12348 -1948
rect -12284 -2372 -12264 -1948
rect -13036 -2400 -12264 -2372
rect -12024 -1948 -11252 -1920
rect -12024 -2372 -11336 -1948
rect -11272 -2372 -11252 -1948
rect -12024 -2400 -11252 -2372
rect -11012 -1948 -10240 -1920
rect -11012 -2372 -10324 -1948
rect -10260 -2372 -10240 -1948
rect -11012 -2400 -10240 -2372
rect -10000 -1948 -9228 -1920
rect -10000 -2372 -9312 -1948
rect -9248 -2372 -9228 -1948
rect -10000 -2400 -9228 -2372
rect -8988 -1948 -8216 -1920
rect -8988 -2372 -8300 -1948
rect -8236 -2372 -8216 -1948
rect -8988 -2400 -8216 -2372
rect -7976 -1948 -7204 -1920
rect -7976 -2372 -7288 -1948
rect -7224 -2372 -7204 -1948
rect -7976 -2400 -7204 -2372
rect -6964 -1948 -6192 -1920
rect -6964 -2372 -6276 -1948
rect -6212 -2372 -6192 -1948
rect -6964 -2400 -6192 -2372
rect -5952 -1948 -5180 -1920
rect -5952 -2372 -5264 -1948
rect -5200 -2372 -5180 -1948
rect -5952 -2400 -5180 -2372
rect -4940 -1948 -4168 -1920
rect -4940 -2372 -4252 -1948
rect -4188 -2372 -4168 -1948
rect -4940 -2400 -4168 -2372
rect -3928 -1948 -3156 -1920
rect -3928 -2372 -3240 -1948
rect -3176 -2372 -3156 -1948
rect -3928 -2400 -3156 -2372
rect -2916 -1948 -2144 -1920
rect -2916 -2372 -2228 -1948
rect -2164 -2372 -2144 -1948
rect -2916 -2400 -2144 -2372
rect -1904 -1948 -1132 -1920
rect -1904 -2372 -1216 -1948
rect -1152 -2372 -1132 -1948
rect -1904 -2400 -1132 -2372
rect -892 -1948 -120 -1920
rect -892 -2372 -204 -1948
rect -140 -2372 -120 -1948
rect -892 -2400 -120 -2372
rect 120 -1948 892 -1920
rect 120 -2372 808 -1948
rect 872 -2372 892 -1948
rect 120 -2400 892 -2372
rect 1132 -1948 1904 -1920
rect 1132 -2372 1820 -1948
rect 1884 -2372 1904 -1948
rect 1132 -2400 1904 -2372
rect 2144 -1948 2916 -1920
rect 2144 -2372 2832 -1948
rect 2896 -2372 2916 -1948
rect 2144 -2400 2916 -2372
rect 3156 -1948 3928 -1920
rect 3156 -2372 3844 -1948
rect 3908 -2372 3928 -1948
rect 3156 -2400 3928 -2372
rect 4168 -1948 4940 -1920
rect 4168 -2372 4856 -1948
rect 4920 -2372 4940 -1948
rect 4168 -2400 4940 -2372
rect 5180 -1948 5952 -1920
rect 5180 -2372 5868 -1948
rect 5932 -2372 5952 -1948
rect 5180 -2400 5952 -2372
rect 6192 -1948 6964 -1920
rect 6192 -2372 6880 -1948
rect 6944 -2372 6964 -1948
rect 6192 -2400 6964 -2372
rect 7204 -1948 7976 -1920
rect 7204 -2372 7892 -1948
rect 7956 -2372 7976 -1948
rect 7204 -2400 7976 -2372
rect 8216 -1948 8988 -1920
rect 8216 -2372 8904 -1948
rect 8968 -2372 8988 -1948
rect 8216 -2400 8988 -2372
rect 9228 -1948 10000 -1920
rect 9228 -2372 9916 -1948
rect 9980 -2372 10000 -1948
rect 9228 -2400 10000 -2372
rect 10240 -1948 11012 -1920
rect 10240 -2372 10928 -1948
rect 10992 -2372 11012 -1948
rect 10240 -2400 11012 -2372
rect 11252 -1948 12024 -1920
rect 11252 -2372 11940 -1948
rect 12004 -2372 12024 -1948
rect 11252 -2400 12024 -2372
rect 12264 -1948 13036 -1920
rect 12264 -2372 12952 -1948
rect 13016 -2372 13036 -1948
rect 12264 -2400 13036 -2372
rect 13276 -1948 14048 -1920
rect 13276 -2372 13964 -1948
rect 14028 -2372 14048 -1948
rect 13276 -2400 14048 -2372
rect 14288 -1948 15060 -1920
rect 14288 -2372 14976 -1948
rect 15040 -2372 15060 -1948
rect 14288 -2400 15060 -2372
rect 15300 -1948 16072 -1920
rect 15300 -2372 15988 -1948
rect 16052 -2372 16072 -1948
rect 15300 -2400 16072 -2372
rect 16312 -1948 17084 -1920
rect 16312 -2372 17000 -1948
rect 17064 -2372 17084 -1948
rect 16312 -2400 17084 -2372
rect 17324 -1948 18096 -1920
rect 17324 -2372 18012 -1948
rect 18076 -2372 18096 -1948
rect 17324 -2400 18096 -2372
rect 18336 -1948 19108 -1920
rect 18336 -2372 19024 -1948
rect 19088 -2372 19108 -1948
rect 18336 -2400 19108 -2372
rect 19348 -1948 20120 -1920
rect 19348 -2372 20036 -1948
rect 20100 -2372 20120 -1948
rect 19348 -2400 20120 -2372
rect 20360 -1948 21132 -1920
rect 20360 -2372 21048 -1948
rect 21112 -2372 21132 -1948
rect 20360 -2400 21132 -2372
rect 21372 -1948 22144 -1920
rect 21372 -2372 22060 -1948
rect 22124 -2372 22144 -1948
rect 21372 -2400 22144 -2372
rect 22384 -1948 23156 -1920
rect 22384 -2372 23072 -1948
rect 23136 -2372 23156 -1948
rect 22384 -2400 23156 -2372
rect 23396 -1948 24168 -1920
rect 23396 -2372 24084 -1948
rect 24148 -2372 24168 -1948
rect 23396 -2400 24168 -2372
rect 24408 -1948 25180 -1920
rect 24408 -2372 25096 -1948
rect 25160 -2372 25180 -1948
rect 24408 -2400 25180 -2372
rect 25420 -1948 26192 -1920
rect 25420 -2372 26108 -1948
rect 26172 -2372 26192 -1948
rect 25420 -2400 26192 -2372
rect 26432 -1948 27204 -1920
rect 26432 -2372 27120 -1948
rect 27184 -2372 27204 -1948
rect 26432 -2400 27204 -2372
rect 27444 -1948 28216 -1920
rect 27444 -2372 28132 -1948
rect 28196 -2372 28216 -1948
rect 27444 -2400 28216 -2372
rect 28456 -1948 29228 -1920
rect 28456 -2372 29144 -1948
rect 29208 -2372 29228 -1948
rect 28456 -2400 29228 -2372
rect 29468 -1948 30240 -1920
rect 29468 -2372 30156 -1948
rect 30220 -2372 30240 -1948
rect 29468 -2400 30240 -2372
rect 30480 -1948 31252 -1920
rect 30480 -2372 31168 -1948
rect 31232 -2372 31252 -1948
rect 30480 -2400 31252 -2372
rect 31492 -1948 32264 -1920
rect 31492 -2372 32180 -1948
rect 32244 -2372 32264 -1948
rect 31492 -2400 32264 -2372
<< via3 >>
rect -31576 1948 -31512 2372
rect -30564 1948 -30500 2372
rect -29552 1948 -29488 2372
rect -28540 1948 -28476 2372
rect -27528 1948 -27464 2372
rect -26516 1948 -26452 2372
rect -25504 1948 -25440 2372
rect -24492 1948 -24428 2372
rect -23480 1948 -23416 2372
rect -22468 1948 -22404 2372
rect -21456 1948 -21392 2372
rect -20444 1948 -20380 2372
rect -19432 1948 -19368 2372
rect -18420 1948 -18356 2372
rect -17408 1948 -17344 2372
rect -16396 1948 -16332 2372
rect -15384 1948 -15320 2372
rect -14372 1948 -14308 2372
rect -13360 1948 -13296 2372
rect -12348 1948 -12284 2372
rect -11336 1948 -11272 2372
rect -10324 1948 -10260 2372
rect -9312 1948 -9248 2372
rect -8300 1948 -8236 2372
rect -7288 1948 -7224 2372
rect -6276 1948 -6212 2372
rect -5264 1948 -5200 2372
rect -4252 1948 -4188 2372
rect -3240 1948 -3176 2372
rect -2228 1948 -2164 2372
rect -1216 1948 -1152 2372
rect -204 1948 -140 2372
rect 808 1948 872 2372
rect 1820 1948 1884 2372
rect 2832 1948 2896 2372
rect 3844 1948 3908 2372
rect 4856 1948 4920 2372
rect 5868 1948 5932 2372
rect 6880 1948 6944 2372
rect 7892 1948 7956 2372
rect 8904 1948 8968 2372
rect 9916 1948 9980 2372
rect 10928 1948 10992 2372
rect 11940 1948 12004 2372
rect 12952 1948 13016 2372
rect 13964 1948 14028 2372
rect 14976 1948 15040 2372
rect 15988 1948 16052 2372
rect 17000 1948 17064 2372
rect 18012 1948 18076 2372
rect 19024 1948 19088 2372
rect 20036 1948 20100 2372
rect 21048 1948 21112 2372
rect 22060 1948 22124 2372
rect 23072 1948 23136 2372
rect 24084 1948 24148 2372
rect 25096 1948 25160 2372
rect 26108 1948 26172 2372
rect 27120 1948 27184 2372
rect 28132 1948 28196 2372
rect 29144 1948 29208 2372
rect 30156 1948 30220 2372
rect 31168 1948 31232 2372
rect 32180 1948 32244 2372
rect -31576 1228 -31512 1652
rect -30564 1228 -30500 1652
rect -29552 1228 -29488 1652
rect -28540 1228 -28476 1652
rect -27528 1228 -27464 1652
rect -26516 1228 -26452 1652
rect -25504 1228 -25440 1652
rect -24492 1228 -24428 1652
rect -23480 1228 -23416 1652
rect -22468 1228 -22404 1652
rect -21456 1228 -21392 1652
rect -20444 1228 -20380 1652
rect -19432 1228 -19368 1652
rect -18420 1228 -18356 1652
rect -17408 1228 -17344 1652
rect -16396 1228 -16332 1652
rect -15384 1228 -15320 1652
rect -14372 1228 -14308 1652
rect -13360 1228 -13296 1652
rect -12348 1228 -12284 1652
rect -11336 1228 -11272 1652
rect -10324 1228 -10260 1652
rect -9312 1228 -9248 1652
rect -8300 1228 -8236 1652
rect -7288 1228 -7224 1652
rect -6276 1228 -6212 1652
rect -5264 1228 -5200 1652
rect -4252 1228 -4188 1652
rect -3240 1228 -3176 1652
rect -2228 1228 -2164 1652
rect -1216 1228 -1152 1652
rect -204 1228 -140 1652
rect 808 1228 872 1652
rect 1820 1228 1884 1652
rect 2832 1228 2896 1652
rect 3844 1228 3908 1652
rect 4856 1228 4920 1652
rect 5868 1228 5932 1652
rect 6880 1228 6944 1652
rect 7892 1228 7956 1652
rect 8904 1228 8968 1652
rect 9916 1228 9980 1652
rect 10928 1228 10992 1652
rect 11940 1228 12004 1652
rect 12952 1228 13016 1652
rect 13964 1228 14028 1652
rect 14976 1228 15040 1652
rect 15988 1228 16052 1652
rect 17000 1228 17064 1652
rect 18012 1228 18076 1652
rect 19024 1228 19088 1652
rect 20036 1228 20100 1652
rect 21048 1228 21112 1652
rect 22060 1228 22124 1652
rect 23072 1228 23136 1652
rect 24084 1228 24148 1652
rect 25096 1228 25160 1652
rect 26108 1228 26172 1652
rect 27120 1228 27184 1652
rect 28132 1228 28196 1652
rect 29144 1228 29208 1652
rect 30156 1228 30220 1652
rect 31168 1228 31232 1652
rect 32180 1228 32244 1652
rect -31576 508 -31512 932
rect -30564 508 -30500 932
rect -29552 508 -29488 932
rect -28540 508 -28476 932
rect -27528 508 -27464 932
rect -26516 508 -26452 932
rect -25504 508 -25440 932
rect -24492 508 -24428 932
rect -23480 508 -23416 932
rect -22468 508 -22404 932
rect -21456 508 -21392 932
rect -20444 508 -20380 932
rect -19432 508 -19368 932
rect -18420 508 -18356 932
rect -17408 508 -17344 932
rect -16396 508 -16332 932
rect -15384 508 -15320 932
rect -14372 508 -14308 932
rect -13360 508 -13296 932
rect -12348 508 -12284 932
rect -11336 508 -11272 932
rect -10324 508 -10260 932
rect -9312 508 -9248 932
rect -8300 508 -8236 932
rect -7288 508 -7224 932
rect -6276 508 -6212 932
rect -5264 508 -5200 932
rect -4252 508 -4188 932
rect -3240 508 -3176 932
rect -2228 508 -2164 932
rect -1216 508 -1152 932
rect -204 508 -140 932
rect 808 508 872 932
rect 1820 508 1884 932
rect 2832 508 2896 932
rect 3844 508 3908 932
rect 4856 508 4920 932
rect 5868 508 5932 932
rect 6880 508 6944 932
rect 7892 508 7956 932
rect 8904 508 8968 932
rect 9916 508 9980 932
rect 10928 508 10992 932
rect 11940 508 12004 932
rect 12952 508 13016 932
rect 13964 508 14028 932
rect 14976 508 15040 932
rect 15988 508 16052 932
rect 17000 508 17064 932
rect 18012 508 18076 932
rect 19024 508 19088 932
rect 20036 508 20100 932
rect 21048 508 21112 932
rect 22060 508 22124 932
rect 23072 508 23136 932
rect 24084 508 24148 932
rect 25096 508 25160 932
rect 26108 508 26172 932
rect 27120 508 27184 932
rect 28132 508 28196 932
rect 29144 508 29208 932
rect 30156 508 30220 932
rect 31168 508 31232 932
rect 32180 508 32244 932
rect -31576 -212 -31512 212
rect -30564 -212 -30500 212
rect -29552 -212 -29488 212
rect -28540 -212 -28476 212
rect -27528 -212 -27464 212
rect -26516 -212 -26452 212
rect -25504 -212 -25440 212
rect -24492 -212 -24428 212
rect -23480 -212 -23416 212
rect -22468 -212 -22404 212
rect -21456 -212 -21392 212
rect -20444 -212 -20380 212
rect -19432 -212 -19368 212
rect -18420 -212 -18356 212
rect -17408 -212 -17344 212
rect -16396 -212 -16332 212
rect -15384 -212 -15320 212
rect -14372 -212 -14308 212
rect -13360 -212 -13296 212
rect -12348 -212 -12284 212
rect -11336 -212 -11272 212
rect -10324 -212 -10260 212
rect -9312 -212 -9248 212
rect -8300 -212 -8236 212
rect -7288 -212 -7224 212
rect -6276 -212 -6212 212
rect -5264 -212 -5200 212
rect -4252 -212 -4188 212
rect -3240 -212 -3176 212
rect -2228 -212 -2164 212
rect -1216 -212 -1152 212
rect -204 -212 -140 212
rect 808 -212 872 212
rect 1820 -212 1884 212
rect 2832 -212 2896 212
rect 3844 -212 3908 212
rect 4856 -212 4920 212
rect 5868 -212 5932 212
rect 6880 -212 6944 212
rect 7892 -212 7956 212
rect 8904 -212 8968 212
rect 9916 -212 9980 212
rect 10928 -212 10992 212
rect 11940 -212 12004 212
rect 12952 -212 13016 212
rect 13964 -212 14028 212
rect 14976 -212 15040 212
rect 15988 -212 16052 212
rect 17000 -212 17064 212
rect 18012 -212 18076 212
rect 19024 -212 19088 212
rect 20036 -212 20100 212
rect 21048 -212 21112 212
rect 22060 -212 22124 212
rect 23072 -212 23136 212
rect 24084 -212 24148 212
rect 25096 -212 25160 212
rect 26108 -212 26172 212
rect 27120 -212 27184 212
rect 28132 -212 28196 212
rect 29144 -212 29208 212
rect 30156 -212 30220 212
rect 31168 -212 31232 212
rect 32180 -212 32244 212
rect -31576 -932 -31512 -508
rect -30564 -932 -30500 -508
rect -29552 -932 -29488 -508
rect -28540 -932 -28476 -508
rect -27528 -932 -27464 -508
rect -26516 -932 -26452 -508
rect -25504 -932 -25440 -508
rect -24492 -932 -24428 -508
rect -23480 -932 -23416 -508
rect -22468 -932 -22404 -508
rect -21456 -932 -21392 -508
rect -20444 -932 -20380 -508
rect -19432 -932 -19368 -508
rect -18420 -932 -18356 -508
rect -17408 -932 -17344 -508
rect -16396 -932 -16332 -508
rect -15384 -932 -15320 -508
rect -14372 -932 -14308 -508
rect -13360 -932 -13296 -508
rect -12348 -932 -12284 -508
rect -11336 -932 -11272 -508
rect -10324 -932 -10260 -508
rect -9312 -932 -9248 -508
rect -8300 -932 -8236 -508
rect -7288 -932 -7224 -508
rect -6276 -932 -6212 -508
rect -5264 -932 -5200 -508
rect -4252 -932 -4188 -508
rect -3240 -932 -3176 -508
rect -2228 -932 -2164 -508
rect -1216 -932 -1152 -508
rect -204 -932 -140 -508
rect 808 -932 872 -508
rect 1820 -932 1884 -508
rect 2832 -932 2896 -508
rect 3844 -932 3908 -508
rect 4856 -932 4920 -508
rect 5868 -932 5932 -508
rect 6880 -932 6944 -508
rect 7892 -932 7956 -508
rect 8904 -932 8968 -508
rect 9916 -932 9980 -508
rect 10928 -932 10992 -508
rect 11940 -932 12004 -508
rect 12952 -932 13016 -508
rect 13964 -932 14028 -508
rect 14976 -932 15040 -508
rect 15988 -932 16052 -508
rect 17000 -932 17064 -508
rect 18012 -932 18076 -508
rect 19024 -932 19088 -508
rect 20036 -932 20100 -508
rect 21048 -932 21112 -508
rect 22060 -932 22124 -508
rect 23072 -932 23136 -508
rect 24084 -932 24148 -508
rect 25096 -932 25160 -508
rect 26108 -932 26172 -508
rect 27120 -932 27184 -508
rect 28132 -932 28196 -508
rect 29144 -932 29208 -508
rect 30156 -932 30220 -508
rect 31168 -932 31232 -508
rect 32180 -932 32244 -508
rect -31576 -1652 -31512 -1228
rect -30564 -1652 -30500 -1228
rect -29552 -1652 -29488 -1228
rect -28540 -1652 -28476 -1228
rect -27528 -1652 -27464 -1228
rect -26516 -1652 -26452 -1228
rect -25504 -1652 -25440 -1228
rect -24492 -1652 -24428 -1228
rect -23480 -1652 -23416 -1228
rect -22468 -1652 -22404 -1228
rect -21456 -1652 -21392 -1228
rect -20444 -1652 -20380 -1228
rect -19432 -1652 -19368 -1228
rect -18420 -1652 -18356 -1228
rect -17408 -1652 -17344 -1228
rect -16396 -1652 -16332 -1228
rect -15384 -1652 -15320 -1228
rect -14372 -1652 -14308 -1228
rect -13360 -1652 -13296 -1228
rect -12348 -1652 -12284 -1228
rect -11336 -1652 -11272 -1228
rect -10324 -1652 -10260 -1228
rect -9312 -1652 -9248 -1228
rect -8300 -1652 -8236 -1228
rect -7288 -1652 -7224 -1228
rect -6276 -1652 -6212 -1228
rect -5264 -1652 -5200 -1228
rect -4252 -1652 -4188 -1228
rect -3240 -1652 -3176 -1228
rect -2228 -1652 -2164 -1228
rect -1216 -1652 -1152 -1228
rect -204 -1652 -140 -1228
rect 808 -1652 872 -1228
rect 1820 -1652 1884 -1228
rect 2832 -1652 2896 -1228
rect 3844 -1652 3908 -1228
rect 4856 -1652 4920 -1228
rect 5868 -1652 5932 -1228
rect 6880 -1652 6944 -1228
rect 7892 -1652 7956 -1228
rect 8904 -1652 8968 -1228
rect 9916 -1652 9980 -1228
rect 10928 -1652 10992 -1228
rect 11940 -1652 12004 -1228
rect 12952 -1652 13016 -1228
rect 13964 -1652 14028 -1228
rect 14976 -1652 15040 -1228
rect 15988 -1652 16052 -1228
rect 17000 -1652 17064 -1228
rect 18012 -1652 18076 -1228
rect 19024 -1652 19088 -1228
rect 20036 -1652 20100 -1228
rect 21048 -1652 21112 -1228
rect 22060 -1652 22124 -1228
rect 23072 -1652 23136 -1228
rect 24084 -1652 24148 -1228
rect 25096 -1652 25160 -1228
rect 26108 -1652 26172 -1228
rect 27120 -1652 27184 -1228
rect 28132 -1652 28196 -1228
rect 29144 -1652 29208 -1228
rect 30156 -1652 30220 -1228
rect 31168 -1652 31232 -1228
rect 32180 -1652 32244 -1228
rect -31576 -2372 -31512 -1948
rect -30564 -2372 -30500 -1948
rect -29552 -2372 -29488 -1948
rect -28540 -2372 -28476 -1948
rect -27528 -2372 -27464 -1948
rect -26516 -2372 -26452 -1948
rect -25504 -2372 -25440 -1948
rect -24492 -2372 -24428 -1948
rect -23480 -2372 -23416 -1948
rect -22468 -2372 -22404 -1948
rect -21456 -2372 -21392 -1948
rect -20444 -2372 -20380 -1948
rect -19432 -2372 -19368 -1948
rect -18420 -2372 -18356 -1948
rect -17408 -2372 -17344 -1948
rect -16396 -2372 -16332 -1948
rect -15384 -2372 -15320 -1948
rect -14372 -2372 -14308 -1948
rect -13360 -2372 -13296 -1948
rect -12348 -2372 -12284 -1948
rect -11336 -2372 -11272 -1948
rect -10324 -2372 -10260 -1948
rect -9312 -2372 -9248 -1948
rect -8300 -2372 -8236 -1948
rect -7288 -2372 -7224 -1948
rect -6276 -2372 -6212 -1948
rect -5264 -2372 -5200 -1948
rect -4252 -2372 -4188 -1948
rect -3240 -2372 -3176 -1948
rect -2228 -2372 -2164 -1948
rect -1216 -2372 -1152 -1948
rect -204 -2372 -140 -1948
rect 808 -2372 872 -1948
rect 1820 -2372 1884 -1948
rect 2832 -2372 2896 -1948
rect 3844 -2372 3908 -1948
rect 4856 -2372 4920 -1948
rect 5868 -2372 5932 -1948
rect 6880 -2372 6944 -1948
rect 7892 -2372 7956 -1948
rect 8904 -2372 8968 -1948
rect 9916 -2372 9980 -1948
rect 10928 -2372 10992 -1948
rect 11940 -2372 12004 -1948
rect 12952 -2372 13016 -1948
rect 13964 -2372 14028 -1948
rect 14976 -2372 15040 -1948
rect 15988 -2372 16052 -1948
rect 17000 -2372 17064 -1948
rect 18012 -2372 18076 -1948
rect 19024 -2372 19088 -1948
rect 20036 -2372 20100 -1948
rect 21048 -2372 21112 -1948
rect 22060 -2372 22124 -1948
rect 23072 -2372 23136 -1948
rect 24084 -2372 24148 -1948
rect 25096 -2372 25160 -1948
rect 26108 -2372 26172 -1948
rect 27120 -2372 27184 -1948
rect 28132 -2372 28196 -1948
rect 29144 -2372 29208 -1948
rect 30156 -2372 30220 -1948
rect 31168 -2372 31232 -1948
rect 32180 -2372 32244 -1948
<< mimcap >>
rect -32224 2320 -31824 2360
rect -32224 2000 -32184 2320
rect -31864 2000 -31824 2320
rect -32224 1960 -31824 2000
rect -31212 2320 -30812 2360
rect -31212 2000 -31172 2320
rect -30852 2000 -30812 2320
rect -31212 1960 -30812 2000
rect -30200 2320 -29800 2360
rect -30200 2000 -30160 2320
rect -29840 2000 -29800 2320
rect -30200 1960 -29800 2000
rect -29188 2320 -28788 2360
rect -29188 2000 -29148 2320
rect -28828 2000 -28788 2320
rect -29188 1960 -28788 2000
rect -28176 2320 -27776 2360
rect -28176 2000 -28136 2320
rect -27816 2000 -27776 2320
rect -28176 1960 -27776 2000
rect -27164 2320 -26764 2360
rect -27164 2000 -27124 2320
rect -26804 2000 -26764 2320
rect -27164 1960 -26764 2000
rect -26152 2320 -25752 2360
rect -26152 2000 -26112 2320
rect -25792 2000 -25752 2320
rect -26152 1960 -25752 2000
rect -25140 2320 -24740 2360
rect -25140 2000 -25100 2320
rect -24780 2000 -24740 2320
rect -25140 1960 -24740 2000
rect -24128 2320 -23728 2360
rect -24128 2000 -24088 2320
rect -23768 2000 -23728 2320
rect -24128 1960 -23728 2000
rect -23116 2320 -22716 2360
rect -23116 2000 -23076 2320
rect -22756 2000 -22716 2320
rect -23116 1960 -22716 2000
rect -22104 2320 -21704 2360
rect -22104 2000 -22064 2320
rect -21744 2000 -21704 2320
rect -22104 1960 -21704 2000
rect -21092 2320 -20692 2360
rect -21092 2000 -21052 2320
rect -20732 2000 -20692 2320
rect -21092 1960 -20692 2000
rect -20080 2320 -19680 2360
rect -20080 2000 -20040 2320
rect -19720 2000 -19680 2320
rect -20080 1960 -19680 2000
rect -19068 2320 -18668 2360
rect -19068 2000 -19028 2320
rect -18708 2000 -18668 2320
rect -19068 1960 -18668 2000
rect -18056 2320 -17656 2360
rect -18056 2000 -18016 2320
rect -17696 2000 -17656 2320
rect -18056 1960 -17656 2000
rect -17044 2320 -16644 2360
rect -17044 2000 -17004 2320
rect -16684 2000 -16644 2320
rect -17044 1960 -16644 2000
rect -16032 2320 -15632 2360
rect -16032 2000 -15992 2320
rect -15672 2000 -15632 2320
rect -16032 1960 -15632 2000
rect -15020 2320 -14620 2360
rect -15020 2000 -14980 2320
rect -14660 2000 -14620 2320
rect -15020 1960 -14620 2000
rect -14008 2320 -13608 2360
rect -14008 2000 -13968 2320
rect -13648 2000 -13608 2320
rect -14008 1960 -13608 2000
rect -12996 2320 -12596 2360
rect -12996 2000 -12956 2320
rect -12636 2000 -12596 2320
rect -12996 1960 -12596 2000
rect -11984 2320 -11584 2360
rect -11984 2000 -11944 2320
rect -11624 2000 -11584 2320
rect -11984 1960 -11584 2000
rect -10972 2320 -10572 2360
rect -10972 2000 -10932 2320
rect -10612 2000 -10572 2320
rect -10972 1960 -10572 2000
rect -9960 2320 -9560 2360
rect -9960 2000 -9920 2320
rect -9600 2000 -9560 2320
rect -9960 1960 -9560 2000
rect -8948 2320 -8548 2360
rect -8948 2000 -8908 2320
rect -8588 2000 -8548 2320
rect -8948 1960 -8548 2000
rect -7936 2320 -7536 2360
rect -7936 2000 -7896 2320
rect -7576 2000 -7536 2320
rect -7936 1960 -7536 2000
rect -6924 2320 -6524 2360
rect -6924 2000 -6884 2320
rect -6564 2000 -6524 2320
rect -6924 1960 -6524 2000
rect -5912 2320 -5512 2360
rect -5912 2000 -5872 2320
rect -5552 2000 -5512 2320
rect -5912 1960 -5512 2000
rect -4900 2320 -4500 2360
rect -4900 2000 -4860 2320
rect -4540 2000 -4500 2320
rect -4900 1960 -4500 2000
rect -3888 2320 -3488 2360
rect -3888 2000 -3848 2320
rect -3528 2000 -3488 2320
rect -3888 1960 -3488 2000
rect -2876 2320 -2476 2360
rect -2876 2000 -2836 2320
rect -2516 2000 -2476 2320
rect -2876 1960 -2476 2000
rect -1864 2320 -1464 2360
rect -1864 2000 -1824 2320
rect -1504 2000 -1464 2320
rect -1864 1960 -1464 2000
rect -852 2320 -452 2360
rect -852 2000 -812 2320
rect -492 2000 -452 2320
rect -852 1960 -452 2000
rect 160 2320 560 2360
rect 160 2000 200 2320
rect 520 2000 560 2320
rect 160 1960 560 2000
rect 1172 2320 1572 2360
rect 1172 2000 1212 2320
rect 1532 2000 1572 2320
rect 1172 1960 1572 2000
rect 2184 2320 2584 2360
rect 2184 2000 2224 2320
rect 2544 2000 2584 2320
rect 2184 1960 2584 2000
rect 3196 2320 3596 2360
rect 3196 2000 3236 2320
rect 3556 2000 3596 2320
rect 3196 1960 3596 2000
rect 4208 2320 4608 2360
rect 4208 2000 4248 2320
rect 4568 2000 4608 2320
rect 4208 1960 4608 2000
rect 5220 2320 5620 2360
rect 5220 2000 5260 2320
rect 5580 2000 5620 2320
rect 5220 1960 5620 2000
rect 6232 2320 6632 2360
rect 6232 2000 6272 2320
rect 6592 2000 6632 2320
rect 6232 1960 6632 2000
rect 7244 2320 7644 2360
rect 7244 2000 7284 2320
rect 7604 2000 7644 2320
rect 7244 1960 7644 2000
rect 8256 2320 8656 2360
rect 8256 2000 8296 2320
rect 8616 2000 8656 2320
rect 8256 1960 8656 2000
rect 9268 2320 9668 2360
rect 9268 2000 9308 2320
rect 9628 2000 9668 2320
rect 9268 1960 9668 2000
rect 10280 2320 10680 2360
rect 10280 2000 10320 2320
rect 10640 2000 10680 2320
rect 10280 1960 10680 2000
rect 11292 2320 11692 2360
rect 11292 2000 11332 2320
rect 11652 2000 11692 2320
rect 11292 1960 11692 2000
rect 12304 2320 12704 2360
rect 12304 2000 12344 2320
rect 12664 2000 12704 2320
rect 12304 1960 12704 2000
rect 13316 2320 13716 2360
rect 13316 2000 13356 2320
rect 13676 2000 13716 2320
rect 13316 1960 13716 2000
rect 14328 2320 14728 2360
rect 14328 2000 14368 2320
rect 14688 2000 14728 2320
rect 14328 1960 14728 2000
rect 15340 2320 15740 2360
rect 15340 2000 15380 2320
rect 15700 2000 15740 2320
rect 15340 1960 15740 2000
rect 16352 2320 16752 2360
rect 16352 2000 16392 2320
rect 16712 2000 16752 2320
rect 16352 1960 16752 2000
rect 17364 2320 17764 2360
rect 17364 2000 17404 2320
rect 17724 2000 17764 2320
rect 17364 1960 17764 2000
rect 18376 2320 18776 2360
rect 18376 2000 18416 2320
rect 18736 2000 18776 2320
rect 18376 1960 18776 2000
rect 19388 2320 19788 2360
rect 19388 2000 19428 2320
rect 19748 2000 19788 2320
rect 19388 1960 19788 2000
rect 20400 2320 20800 2360
rect 20400 2000 20440 2320
rect 20760 2000 20800 2320
rect 20400 1960 20800 2000
rect 21412 2320 21812 2360
rect 21412 2000 21452 2320
rect 21772 2000 21812 2320
rect 21412 1960 21812 2000
rect 22424 2320 22824 2360
rect 22424 2000 22464 2320
rect 22784 2000 22824 2320
rect 22424 1960 22824 2000
rect 23436 2320 23836 2360
rect 23436 2000 23476 2320
rect 23796 2000 23836 2320
rect 23436 1960 23836 2000
rect 24448 2320 24848 2360
rect 24448 2000 24488 2320
rect 24808 2000 24848 2320
rect 24448 1960 24848 2000
rect 25460 2320 25860 2360
rect 25460 2000 25500 2320
rect 25820 2000 25860 2320
rect 25460 1960 25860 2000
rect 26472 2320 26872 2360
rect 26472 2000 26512 2320
rect 26832 2000 26872 2320
rect 26472 1960 26872 2000
rect 27484 2320 27884 2360
rect 27484 2000 27524 2320
rect 27844 2000 27884 2320
rect 27484 1960 27884 2000
rect 28496 2320 28896 2360
rect 28496 2000 28536 2320
rect 28856 2000 28896 2320
rect 28496 1960 28896 2000
rect 29508 2320 29908 2360
rect 29508 2000 29548 2320
rect 29868 2000 29908 2320
rect 29508 1960 29908 2000
rect 30520 2320 30920 2360
rect 30520 2000 30560 2320
rect 30880 2000 30920 2320
rect 30520 1960 30920 2000
rect 31532 2320 31932 2360
rect 31532 2000 31572 2320
rect 31892 2000 31932 2320
rect 31532 1960 31932 2000
rect -32224 1600 -31824 1640
rect -32224 1280 -32184 1600
rect -31864 1280 -31824 1600
rect -32224 1240 -31824 1280
rect -31212 1600 -30812 1640
rect -31212 1280 -31172 1600
rect -30852 1280 -30812 1600
rect -31212 1240 -30812 1280
rect -30200 1600 -29800 1640
rect -30200 1280 -30160 1600
rect -29840 1280 -29800 1600
rect -30200 1240 -29800 1280
rect -29188 1600 -28788 1640
rect -29188 1280 -29148 1600
rect -28828 1280 -28788 1600
rect -29188 1240 -28788 1280
rect -28176 1600 -27776 1640
rect -28176 1280 -28136 1600
rect -27816 1280 -27776 1600
rect -28176 1240 -27776 1280
rect -27164 1600 -26764 1640
rect -27164 1280 -27124 1600
rect -26804 1280 -26764 1600
rect -27164 1240 -26764 1280
rect -26152 1600 -25752 1640
rect -26152 1280 -26112 1600
rect -25792 1280 -25752 1600
rect -26152 1240 -25752 1280
rect -25140 1600 -24740 1640
rect -25140 1280 -25100 1600
rect -24780 1280 -24740 1600
rect -25140 1240 -24740 1280
rect -24128 1600 -23728 1640
rect -24128 1280 -24088 1600
rect -23768 1280 -23728 1600
rect -24128 1240 -23728 1280
rect -23116 1600 -22716 1640
rect -23116 1280 -23076 1600
rect -22756 1280 -22716 1600
rect -23116 1240 -22716 1280
rect -22104 1600 -21704 1640
rect -22104 1280 -22064 1600
rect -21744 1280 -21704 1600
rect -22104 1240 -21704 1280
rect -21092 1600 -20692 1640
rect -21092 1280 -21052 1600
rect -20732 1280 -20692 1600
rect -21092 1240 -20692 1280
rect -20080 1600 -19680 1640
rect -20080 1280 -20040 1600
rect -19720 1280 -19680 1600
rect -20080 1240 -19680 1280
rect -19068 1600 -18668 1640
rect -19068 1280 -19028 1600
rect -18708 1280 -18668 1600
rect -19068 1240 -18668 1280
rect -18056 1600 -17656 1640
rect -18056 1280 -18016 1600
rect -17696 1280 -17656 1600
rect -18056 1240 -17656 1280
rect -17044 1600 -16644 1640
rect -17044 1280 -17004 1600
rect -16684 1280 -16644 1600
rect -17044 1240 -16644 1280
rect -16032 1600 -15632 1640
rect -16032 1280 -15992 1600
rect -15672 1280 -15632 1600
rect -16032 1240 -15632 1280
rect -15020 1600 -14620 1640
rect -15020 1280 -14980 1600
rect -14660 1280 -14620 1600
rect -15020 1240 -14620 1280
rect -14008 1600 -13608 1640
rect -14008 1280 -13968 1600
rect -13648 1280 -13608 1600
rect -14008 1240 -13608 1280
rect -12996 1600 -12596 1640
rect -12996 1280 -12956 1600
rect -12636 1280 -12596 1600
rect -12996 1240 -12596 1280
rect -11984 1600 -11584 1640
rect -11984 1280 -11944 1600
rect -11624 1280 -11584 1600
rect -11984 1240 -11584 1280
rect -10972 1600 -10572 1640
rect -10972 1280 -10932 1600
rect -10612 1280 -10572 1600
rect -10972 1240 -10572 1280
rect -9960 1600 -9560 1640
rect -9960 1280 -9920 1600
rect -9600 1280 -9560 1600
rect -9960 1240 -9560 1280
rect -8948 1600 -8548 1640
rect -8948 1280 -8908 1600
rect -8588 1280 -8548 1600
rect -8948 1240 -8548 1280
rect -7936 1600 -7536 1640
rect -7936 1280 -7896 1600
rect -7576 1280 -7536 1600
rect -7936 1240 -7536 1280
rect -6924 1600 -6524 1640
rect -6924 1280 -6884 1600
rect -6564 1280 -6524 1600
rect -6924 1240 -6524 1280
rect -5912 1600 -5512 1640
rect -5912 1280 -5872 1600
rect -5552 1280 -5512 1600
rect -5912 1240 -5512 1280
rect -4900 1600 -4500 1640
rect -4900 1280 -4860 1600
rect -4540 1280 -4500 1600
rect -4900 1240 -4500 1280
rect -3888 1600 -3488 1640
rect -3888 1280 -3848 1600
rect -3528 1280 -3488 1600
rect -3888 1240 -3488 1280
rect -2876 1600 -2476 1640
rect -2876 1280 -2836 1600
rect -2516 1280 -2476 1600
rect -2876 1240 -2476 1280
rect -1864 1600 -1464 1640
rect -1864 1280 -1824 1600
rect -1504 1280 -1464 1600
rect -1864 1240 -1464 1280
rect -852 1600 -452 1640
rect -852 1280 -812 1600
rect -492 1280 -452 1600
rect -852 1240 -452 1280
rect 160 1600 560 1640
rect 160 1280 200 1600
rect 520 1280 560 1600
rect 160 1240 560 1280
rect 1172 1600 1572 1640
rect 1172 1280 1212 1600
rect 1532 1280 1572 1600
rect 1172 1240 1572 1280
rect 2184 1600 2584 1640
rect 2184 1280 2224 1600
rect 2544 1280 2584 1600
rect 2184 1240 2584 1280
rect 3196 1600 3596 1640
rect 3196 1280 3236 1600
rect 3556 1280 3596 1600
rect 3196 1240 3596 1280
rect 4208 1600 4608 1640
rect 4208 1280 4248 1600
rect 4568 1280 4608 1600
rect 4208 1240 4608 1280
rect 5220 1600 5620 1640
rect 5220 1280 5260 1600
rect 5580 1280 5620 1600
rect 5220 1240 5620 1280
rect 6232 1600 6632 1640
rect 6232 1280 6272 1600
rect 6592 1280 6632 1600
rect 6232 1240 6632 1280
rect 7244 1600 7644 1640
rect 7244 1280 7284 1600
rect 7604 1280 7644 1600
rect 7244 1240 7644 1280
rect 8256 1600 8656 1640
rect 8256 1280 8296 1600
rect 8616 1280 8656 1600
rect 8256 1240 8656 1280
rect 9268 1600 9668 1640
rect 9268 1280 9308 1600
rect 9628 1280 9668 1600
rect 9268 1240 9668 1280
rect 10280 1600 10680 1640
rect 10280 1280 10320 1600
rect 10640 1280 10680 1600
rect 10280 1240 10680 1280
rect 11292 1600 11692 1640
rect 11292 1280 11332 1600
rect 11652 1280 11692 1600
rect 11292 1240 11692 1280
rect 12304 1600 12704 1640
rect 12304 1280 12344 1600
rect 12664 1280 12704 1600
rect 12304 1240 12704 1280
rect 13316 1600 13716 1640
rect 13316 1280 13356 1600
rect 13676 1280 13716 1600
rect 13316 1240 13716 1280
rect 14328 1600 14728 1640
rect 14328 1280 14368 1600
rect 14688 1280 14728 1600
rect 14328 1240 14728 1280
rect 15340 1600 15740 1640
rect 15340 1280 15380 1600
rect 15700 1280 15740 1600
rect 15340 1240 15740 1280
rect 16352 1600 16752 1640
rect 16352 1280 16392 1600
rect 16712 1280 16752 1600
rect 16352 1240 16752 1280
rect 17364 1600 17764 1640
rect 17364 1280 17404 1600
rect 17724 1280 17764 1600
rect 17364 1240 17764 1280
rect 18376 1600 18776 1640
rect 18376 1280 18416 1600
rect 18736 1280 18776 1600
rect 18376 1240 18776 1280
rect 19388 1600 19788 1640
rect 19388 1280 19428 1600
rect 19748 1280 19788 1600
rect 19388 1240 19788 1280
rect 20400 1600 20800 1640
rect 20400 1280 20440 1600
rect 20760 1280 20800 1600
rect 20400 1240 20800 1280
rect 21412 1600 21812 1640
rect 21412 1280 21452 1600
rect 21772 1280 21812 1600
rect 21412 1240 21812 1280
rect 22424 1600 22824 1640
rect 22424 1280 22464 1600
rect 22784 1280 22824 1600
rect 22424 1240 22824 1280
rect 23436 1600 23836 1640
rect 23436 1280 23476 1600
rect 23796 1280 23836 1600
rect 23436 1240 23836 1280
rect 24448 1600 24848 1640
rect 24448 1280 24488 1600
rect 24808 1280 24848 1600
rect 24448 1240 24848 1280
rect 25460 1600 25860 1640
rect 25460 1280 25500 1600
rect 25820 1280 25860 1600
rect 25460 1240 25860 1280
rect 26472 1600 26872 1640
rect 26472 1280 26512 1600
rect 26832 1280 26872 1600
rect 26472 1240 26872 1280
rect 27484 1600 27884 1640
rect 27484 1280 27524 1600
rect 27844 1280 27884 1600
rect 27484 1240 27884 1280
rect 28496 1600 28896 1640
rect 28496 1280 28536 1600
rect 28856 1280 28896 1600
rect 28496 1240 28896 1280
rect 29508 1600 29908 1640
rect 29508 1280 29548 1600
rect 29868 1280 29908 1600
rect 29508 1240 29908 1280
rect 30520 1600 30920 1640
rect 30520 1280 30560 1600
rect 30880 1280 30920 1600
rect 30520 1240 30920 1280
rect 31532 1600 31932 1640
rect 31532 1280 31572 1600
rect 31892 1280 31932 1600
rect 31532 1240 31932 1280
rect -32224 880 -31824 920
rect -32224 560 -32184 880
rect -31864 560 -31824 880
rect -32224 520 -31824 560
rect -31212 880 -30812 920
rect -31212 560 -31172 880
rect -30852 560 -30812 880
rect -31212 520 -30812 560
rect -30200 880 -29800 920
rect -30200 560 -30160 880
rect -29840 560 -29800 880
rect -30200 520 -29800 560
rect -29188 880 -28788 920
rect -29188 560 -29148 880
rect -28828 560 -28788 880
rect -29188 520 -28788 560
rect -28176 880 -27776 920
rect -28176 560 -28136 880
rect -27816 560 -27776 880
rect -28176 520 -27776 560
rect -27164 880 -26764 920
rect -27164 560 -27124 880
rect -26804 560 -26764 880
rect -27164 520 -26764 560
rect -26152 880 -25752 920
rect -26152 560 -26112 880
rect -25792 560 -25752 880
rect -26152 520 -25752 560
rect -25140 880 -24740 920
rect -25140 560 -25100 880
rect -24780 560 -24740 880
rect -25140 520 -24740 560
rect -24128 880 -23728 920
rect -24128 560 -24088 880
rect -23768 560 -23728 880
rect -24128 520 -23728 560
rect -23116 880 -22716 920
rect -23116 560 -23076 880
rect -22756 560 -22716 880
rect -23116 520 -22716 560
rect -22104 880 -21704 920
rect -22104 560 -22064 880
rect -21744 560 -21704 880
rect -22104 520 -21704 560
rect -21092 880 -20692 920
rect -21092 560 -21052 880
rect -20732 560 -20692 880
rect -21092 520 -20692 560
rect -20080 880 -19680 920
rect -20080 560 -20040 880
rect -19720 560 -19680 880
rect -20080 520 -19680 560
rect -19068 880 -18668 920
rect -19068 560 -19028 880
rect -18708 560 -18668 880
rect -19068 520 -18668 560
rect -18056 880 -17656 920
rect -18056 560 -18016 880
rect -17696 560 -17656 880
rect -18056 520 -17656 560
rect -17044 880 -16644 920
rect -17044 560 -17004 880
rect -16684 560 -16644 880
rect -17044 520 -16644 560
rect -16032 880 -15632 920
rect -16032 560 -15992 880
rect -15672 560 -15632 880
rect -16032 520 -15632 560
rect -15020 880 -14620 920
rect -15020 560 -14980 880
rect -14660 560 -14620 880
rect -15020 520 -14620 560
rect -14008 880 -13608 920
rect -14008 560 -13968 880
rect -13648 560 -13608 880
rect -14008 520 -13608 560
rect -12996 880 -12596 920
rect -12996 560 -12956 880
rect -12636 560 -12596 880
rect -12996 520 -12596 560
rect -11984 880 -11584 920
rect -11984 560 -11944 880
rect -11624 560 -11584 880
rect -11984 520 -11584 560
rect -10972 880 -10572 920
rect -10972 560 -10932 880
rect -10612 560 -10572 880
rect -10972 520 -10572 560
rect -9960 880 -9560 920
rect -9960 560 -9920 880
rect -9600 560 -9560 880
rect -9960 520 -9560 560
rect -8948 880 -8548 920
rect -8948 560 -8908 880
rect -8588 560 -8548 880
rect -8948 520 -8548 560
rect -7936 880 -7536 920
rect -7936 560 -7896 880
rect -7576 560 -7536 880
rect -7936 520 -7536 560
rect -6924 880 -6524 920
rect -6924 560 -6884 880
rect -6564 560 -6524 880
rect -6924 520 -6524 560
rect -5912 880 -5512 920
rect -5912 560 -5872 880
rect -5552 560 -5512 880
rect -5912 520 -5512 560
rect -4900 880 -4500 920
rect -4900 560 -4860 880
rect -4540 560 -4500 880
rect -4900 520 -4500 560
rect -3888 880 -3488 920
rect -3888 560 -3848 880
rect -3528 560 -3488 880
rect -3888 520 -3488 560
rect -2876 880 -2476 920
rect -2876 560 -2836 880
rect -2516 560 -2476 880
rect -2876 520 -2476 560
rect -1864 880 -1464 920
rect -1864 560 -1824 880
rect -1504 560 -1464 880
rect -1864 520 -1464 560
rect -852 880 -452 920
rect -852 560 -812 880
rect -492 560 -452 880
rect -852 520 -452 560
rect 160 880 560 920
rect 160 560 200 880
rect 520 560 560 880
rect 160 520 560 560
rect 1172 880 1572 920
rect 1172 560 1212 880
rect 1532 560 1572 880
rect 1172 520 1572 560
rect 2184 880 2584 920
rect 2184 560 2224 880
rect 2544 560 2584 880
rect 2184 520 2584 560
rect 3196 880 3596 920
rect 3196 560 3236 880
rect 3556 560 3596 880
rect 3196 520 3596 560
rect 4208 880 4608 920
rect 4208 560 4248 880
rect 4568 560 4608 880
rect 4208 520 4608 560
rect 5220 880 5620 920
rect 5220 560 5260 880
rect 5580 560 5620 880
rect 5220 520 5620 560
rect 6232 880 6632 920
rect 6232 560 6272 880
rect 6592 560 6632 880
rect 6232 520 6632 560
rect 7244 880 7644 920
rect 7244 560 7284 880
rect 7604 560 7644 880
rect 7244 520 7644 560
rect 8256 880 8656 920
rect 8256 560 8296 880
rect 8616 560 8656 880
rect 8256 520 8656 560
rect 9268 880 9668 920
rect 9268 560 9308 880
rect 9628 560 9668 880
rect 9268 520 9668 560
rect 10280 880 10680 920
rect 10280 560 10320 880
rect 10640 560 10680 880
rect 10280 520 10680 560
rect 11292 880 11692 920
rect 11292 560 11332 880
rect 11652 560 11692 880
rect 11292 520 11692 560
rect 12304 880 12704 920
rect 12304 560 12344 880
rect 12664 560 12704 880
rect 12304 520 12704 560
rect 13316 880 13716 920
rect 13316 560 13356 880
rect 13676 560 13716 880
rect 13316 520 13716 560
rect 14328 880 14728 920
rect 14328 560 14368 880
rect 14688 560 14728 880
rect 14328 520 14728 560
rect 15340 880 15740 920
rect 15340 560 15380 880
rect 15700 560 15740 880
rect 15340 520 15740 560
rect 16352 880 16752 920
rect 16352 560 16392 880
rect 16712 560 16752 880
rect 16352 520 16752 560
rect 17364 880 17764 920
rect 17364 560 17404 880
rect 17724 560 17764 880
rect 17364 520 17764 560
rect 18376 880 18776 920
rect 18376 560 18416 880
rect 18736 560 18776 880
rect 18376 520 18776 560
rect 19388 880 19788 920
rect 19388 560 19428 880
rect 19748 560 19788 880
rect 19388 520 19788 560
rect 20400 880 20800 920
rect 20400 560 20440 880
rect 20760 560 20800 880
rect 20400 520 20800 560
rect 21412 880 21812 920
rect 21412 560 21452 880
rect 21772 560 21812 880
rect 21412 520 21812 560
rect 22424 880 22824 920
rect 22424 560 22464 880
rect 22784 560 22824 880
rect 22424 520 22824 560
rect 23436 880 23836 920
rect 23436 560 23476 880
rect 23796 560 23836 880
rect 23436 520 23836 560
rect 24448 880 24848 920
rect 24448 560 24488 880
rect 24808 560 24848 880
rect 24448 520 24848 560
rect 25460 880 25860 920
rect 25460 560 25500 880
rect 25820 560 25860 880
rect 25460 520 25860 560
rect 26472 880 26872 920
rect 26472 560 26512 880
rect 26832 560 26872 880
rect 26472 520 26872 560
rect 27484 880 27884 920
rect 27484 560 27524 880
rect 27844 560 27884 880
rect 27484 520 27884 560
rect 28496 880 28896 920
rect 28496 560 28536 880
rect 28856 560 28896 880
rect 28496 520 28896 560
rect 29508 880 29908 920
rect 29508 560 29548 880
rect 29868 560 29908 880
rect 29508 520 29908 560
rect 30520 880 30920 920
rect 30520 560 30560 880
rect 30880 560 30920 880
rect 30520 520 30920 560
rect 31532 880 31932 920
rect 31532 560 31572 880
rect 31892 560 31932 880
rect 31532 520 31932 560
rect -32224 160 -31824 200
rect -32224 -160 -32184 160
rect -31864 -160 -31824 160
rect -32224 -200 -31824 -160
rect -31212 160 -30812 200
rect -31212 -160 -31172 160
rect -30852 -160 -30812 160
rect -31212 -200 -30812 -160
rect -30200 160 -29800 200
rect -30200 -160 -30160 160
rect -29840 -160 -29800 160
rect -30200 -200 -29800 -160
rect -29188 160 -28788 200
rect -29188 -160 -29148 160
rect -28828 -160 -28788 160
rect -29188 -200 -28788 -160
rect -28176 160 -27776 200
rect -28176 -160 -28136 160
rect -27816 -160 -27776 160
rect -28176 -200 -27776 -160
rect -27164 160 -26764 200
rect -27164 -160 -27124 160
rect -26804 -160 -26764 160
rect -27164 -200 -26764 -160
rect -26152 160 -25752 200
rect -26152 -160 -26112 160
rect -25792 -160 -25752 160
rect -26152 -200 -25752 -160
rect -25140 160 -24740 200
rect -25140 -160 -25100 160
rect -24780 -160 -24740 160
rect -25140 -200 -24740 -160
rect -24128 160 -23728 200
rect -24128 -160 -24088 160
rect -23768 -160 -23728 160
rect -24128 -200 -23728 -160
rect -23116 160 -22716 200
rect -23116 -160 -23076 160
rect -22756 -160 -22716 160
rect -23116 -200 -22716 -160
rect -22104 160 -21704 200
rect -22104 -160 -22064 160
rect -21744 -160 -21704 160
rect -22104 -200 -21704 -160
rect -21092 160 -20692 200
rect -21092 -160 -21052 160
rect -20732 -160 -20692 160
rect -21092 -200 -20692 -160
rect -20080 160 -19680 200
rect -20080 -160 -20040 160
rect -19720 -160 -19680 160
rect -20080 -200 -19680 -160
rect -19068 160 -18668 200
rect -19068 -160 -19028 160
rect -18708 -160 -18668 160
rect -19068 -200 -18668 -160
rect -18056 160 -17656 200
rect -18056 -160 -18016 160
rect -17696 -160 -17656 160
rect -18056 -200 -17656 -160
rect -17044 160 -16644 200
rect -17044 -160 -17004 160
rect -16684 -160 -16644 160
rect -17044 -200 -16644 -160
rect -16032 160 -15632 200
rect -16032 -160 -15992 160
rect -15672 -160 -15632 160
rect -16032 -200 -15632 -160
rect -15020 160 -14620 200
rect -15020 -160 -14980 160
rect -14660 -160 -14620 160
rect -15020 -200 -14620 -160
rect -14008 160 -13608 200
rect -14008 -160 -13968 160
rect -13648 -160 -13608 160
rect -14008 -200 -13608 -160
rect -12996 160 -12596 200
rect -12996 -160 -12956 160
rect -12636 -160 -12596 160
rect -12996 -200 -12596 -160
rect -11984 160 -11584 200
rect -11984 -160 -11944 160
rect -11624 -160 -11584 160
rect -11984 -200 -11584 -160
rect -10972 160 -10572 200
rect -10972 -160 -10932 160
rect -10612 -160 -10572 160
rect -10972 -200 -10572 -160
rect -9960 160 -9560 200
rect -9960 -160 -9920 160
rect -9600 -160 -9560 160
rect -9960 -200 -9560 -160
rect -8948 160 -8548 200
rect -8948 -160 -8908 160
rect -8588 -160 -8548 160
rect -8948 -200 -8548 -160
rect -7936 160 -7536 200
rect -7936 -160 -7896 160
rect -7576 -160 -7536 160
rect -7936 -200 -7536 -160
rect -6924 160 -6524 200
rect -6924 -160 -6884 160
rect -6564 -160 -6524 160
rect -6924 -200 -6524 -160
rect -5912 160 -5512 200
rect -5912 -160 -5872 160
rect -5552 -160 -5512 160
rect -5912 -200 -5512 -160
rect -4900 160 -4500 200
rect -4900 -160 -4860 160
rect -4540 -160 -4500 160
rect -4900 -200 -4500 -160
rect -3888 160 -3488 200
rect -3888 -160 -3848 160
rect -3528 -160 -3488 160
rect -3888 -200 -3488 -160
rect -2876 160 -2476 200
rect -2876 -160 -2836 160
rect -2516 -160 -2476 160
rect -2876 -200 -2476 -160
rect -1864 160 -1464 200
rect -1864 -160 -1824 160
rect -1504 -160 -1464 160
rect -1864 -200 -1464 -160
rect -852 160 -452 200
rect -852 -160 -812 160
rect -492 -160 -452 160
rect -852 -200 -452 -160
rect 160 160 560 200
rect 160 -160 200 160
rect 520 -160 560 160
rect 160 -200 560 -160
rect 1172 160 1572 200
rect 1172 -160 1212 160
rect 1532 -160 1572 160
rect 1172 -200 1572 -160
rect 2184 160 2584 200
rect 2184 -160 2224 160
rect 2544 -160 2584 160
rect 2184 -200 2584 -160
rect 3196 160 3596 200
rect 3196 -160 3236 160
rect 3556 -160 3596 160
rect 3196 -200 3596 -160
rect 4208 160 4608 200
rect 4208 -160 4248 160
rect 4568 -160 4608 160
rect 4208 -200 4608 -160
rect 5220 160 5620 200
rect 5220 -160 5260 160
rect 5580 -160 5620 160
rect 5220 -200 5620 -160
rect 6232 160 6632 200
rect 6232 -160 6272 160
rect 6592 -160 6632 160
rect 6232 -200 6632 -160
rect 7244 160 7644 200
rect 7244 -160 7284 160
rect 7604 -160 7644 160
rect 7244 -200 7644 -160
rect 8256 160 8656 200
rect 8256 -160 8296 160
rect 8616 -160 8656 160
rect 8256 -200 8656 -160
rect 9268 160 9668 200
rect 9268 -160 9308 160
rect 9628 -160 9668 160
rect 9268 -200 9668 -160
rect 10280 160 10680 200
rect 10280 -160 10320 160
rect 10640 -160 10680 160
rect 10280 -200 10680 -160
rect 11292 160 11692 200
rect 11292 -160 11332 160
rect 11652 -160 11692 160
rect 11292 -200 11692 -160
rect 12304 160 12704 200
rect 12304 -160 12344 160
rect 12664 -160 12704 160
rect 12304 -200 12704 -160
rect 13316 160 13716 200
rect 13316 -160 13356 160
rect 13676 -160 13716 160
rect 13316 -200 13716 -160
rect 14328 160 14728 200
rect 14328 -160 14368 160
rect 14688 -160 14728 160
rect 14328 -200 14728 -160
rect 15340 160 15740 200
rect 15340 -160 15380 160
rect 15700 -160 15740 160
rect 15340 -200 15740 -160
rect 16352 160 16752 200
rect 16352 -160 16392 160
rect 16712 -160 16752 160
rect 16352 -200 16752 -160
rect 17364 160 17764 200
rect 17364 -160 17404 160
rect 17724 -160 17764 160
rect 17364 -200 17764 -160
rect 18376 160 18776 200
rect 18376 -160 18416 160
rect 18736 -160 18776 160
rect 18376 -200 18776 -160
rect 19388 160 19788 200
rect 19388 -160 19428 160
rect 19748 -160 19788 160
rect 19388 -200 19788 -160
rect 20400 160 20800 200
rect 20400 -160 20440 160
rect 20760 -160 20800 160
rect 20400 -200 20800 -160
rect 21412 160 21812 200
rect 21412 -160 21452 160
rect 21772 -160 21812 160
rect 21412 -200 21812 -160
rect 22424 160 22824 200
rect 22424 -160 22464 160
rect 22784 -160 22824 160
rect 22424 -200 22824 -160
rect 23436 160 23836 200
rect 23436 -160 23476 160
rect 23796 -160 23836 160
rect 23436 -200 23836 -160
rect 24448 160 24848 200
rect 24448 -160 24488 160
rect 24808 -160 24848 160
rect 24448 -200 24848 -160
rect 25460 160 25860 200
rect 25460 -160 25500 160
rect 25820 -160 25860 160
rect 25460 -200 25860 -160
rect 26472 160 26872 200
rect 26472 -160 26512 160
rect 26832 -160 26872 160
rect 26472 -200 26872 -160
rect 27484 160 27884 200
rect 27484 -160 27524 160
rect 27844 -160 27884 160
rect 27484 -200 27884 -160
rect 28496 160 28896 200
rect 28496 -160 28536 160
rect 28856 -160 28896 160
rect 28496 -200 28896 -160
rect 29508 160 29908 200
rect 29508 -160 29548 160
rect 29868 -160 29908 160
rect 29508 -200 29908 -160
rect 30520 160 30920 200
rect 30520 -160 30560 160
rect 30880 -160 30920 160
rect 30520 -200 30920 -160
rect 31532 160 31932 200
rect 31532 -160 31572 160
rect 31892 -160 31932 160
rect 31532 -200 31932 -160
rect -32224 -560 -31824 -520
rect -32224 -880 -32184 -560
rect -31864 -880 -31824 -560
rect -32224 -920 -31824 -880
rect -31212 -560 -30812 -520
rect -31212 -880 -31172 -560
rect -30852 -880 -30812 -560
rect -31212 -920 -30812 -880
rect -30200 -560 -29800 -520
rect -30200 -880 -30160 -560
rect -29840 -880 -29800 -560
rect -30200 -920 -29800 -880
rect -29188 -560 -28788 -520
rect -29188 -880 -29148 -560
rect -28828 -880 -28788 -560
rect -29188 -920 -28788 -880
rect -28176 -560 -27776 -520
rect -28176 -880 -28136 -560
rect -27816 -880 -27776 -560
rect -28176 -920 -27776 -880
rect -27164 -560 -26764 -520
rect -27164 -880 -27124 -560
rect -26804 -880 -26764 -560
rect -27164 -920 -26764 -880
rect -26152 -560 -25752 -520
rect -26152 -880 -26112 -560
rect -25792 -880 -25752 -560
rect -26152 -920 -25752 -880
rect -25140 -560 -24740 -520
rect -25140 -880 -25100 -560
rect -24780 -880 -24740 -560
rect -25140 -920 -24740 -880
rect -24128 -560 -23728 -520
rect -24128 -880 -24088 -560
rect -23768 -880 -23728 -560
rect -24128 -920 -23728 -880
rect -23116 -560 -22716 -520
rect -23116 -880 -23076 -560
rect -22756 -880 -22716 -560
rect -23116 -920 -22716 -880
rect -22104 -560 -21704 -520
rect -22104 -880 -22064 -560
rect -21744 -880 -21704 -560
rect -22104 -920 -21704 -880
rect -21092 -560 -20692 -520
rect -21092 -880 -21052 -560
rect -20732 -880 -20692 -560
rect -21092 -920 -20692 -880
rect -20080 -560 -19680 -520
rect -20080 -880 -20040 -560
rect -19720 -880 -19680 -560
rect -20080 -920 -19680 -880
rect -19068 -560 -18668 -520
rect -19068 -880 -19028 -560
rect -18708 -880 -18668 -560
rect -19068 -920 -18668 -880
rect -18056 -560 -17656 -520
rect -18056 -880 -18016 -560
rect -17696 -880 -17656 -560
rect -18056 -920 -17656 -880
rect -17044 -560 -16644 -520
rect -17044 -880 -17004 -560
rect -16684 -880 -16644 -560
rect -17044 -920 -16644 -880
rect -16032 -560 -15632 -520
rect -16032 -880 -15992 -560
rect -15672 -880 -15632 -560
rect -16032 -920 -15632 -880
rect -15020 -560 -14620 -520
rect -15020 -880 -14980 -560
rect -14660 -880 -14620 -560
rect -15020 -920 -14620 -880
rect -14008 -560 -13608 -520
rect -14008 -880 -13968 -560
rect -13648 -880 -13608 -560
rect -14008 -920 -13608 -880
rect -12996 -560 -12596 -520
rect -12996 -880 -12956 -560
rect -12636 -880 -12596 -560
rect -12996 -920 -12596 -880
rect -11984 -560 -11584 -520
rect -11984 -880 -11944 -560
rect -11624 -880 -11584 -560
rect -11984 -920 -11584 -880
rect -10972 -560 -10572 -520
rect -10972 -880 -10932 -560
rect -10612 -880 -10572 -560
rect -10972 -920 -10572 -880
rect -9960 -560 -9560 -520
rect -9960 -880 -9920 -560
rect -9600 -880 -9560 -560
rect -9960 -920 -9560 -880
rect -8948 -560 -8548 -520
rect -8948 -880 -8908 -560
rect -8588 -880 -8548 -560
rect -8948 -920 -8548 -880
rect -7936 -560 -7536 -520
rect -7936 -880 -7896 -560
rect -7576 -880 -7536 -560
rect -7936 -920 -7536 -880
rect -6924 -560 -6524 -520
rect -6924 -880 -6884 -560
rect -6564 -880 -6524 -560
rect -6924 -920 -6524 -880
rect -5912 -560 -5512 -520
rect -5912 -880 -5872 -560
rect -5552 -880 -5512 -560
rect -5912 -920 -5512 -880
rect -4900 -560 -4500 -520
rect -4900 -880 -4860 -560
rect -4540 -880 -4500 -560
rect -4900 -920 -4500 -880
rect -3888 -560 -3488 -520
rect -3888 -880 -3848 -560
rect -3528 -880 -3488 -560
rect -3888 -920 -3488 -880
rect -2876 -560 -2476 -520
rect -2876 -880 -2836 -560
rect -2516 -880 -2476 -560
rect -2876 -920 -2476 -880
rect -1864 -560 -1464 -520
rect -1864 -880 -1824 -560
rect -1504 -880 -1464 -560
rect -1864 -920 -1464 -880
rect -852 -560 -452 -520
rect -852 -880 -812 -560
rect -492 -880 -452 -560
rect -852 -920 -452 -880
rect 160 -560 560 -520
rect 160 -880 200 -560
rect 520 -880 560 -560
rect 160 -920 560 -880
rect 1172 -560 1572 -520
rect 1172 -880 1212 -560
rect 1532 -880 1572 -560
rect 1172 -920 1572 -880
rect 2184 -560 2584 -520
rect 2184 -880 2224 -560
rect 2544 -880 2584 -560
rect 2184 -920 2584 -880
rect 3196 -560 3596 -520
rect 3196 -880 3236 -560
rect 3556 -880 3596 -560
rect 3196 -920 3596 -880
rect 4208 -560 4608 -520
rect 4208 -880 4248 -560
rect 4568 -880 4608 -560
rect 4208 -920 4608 -880
rect 5220 -560 5620 -520
rect 5220 -880 5260 -560
rect 5580 -880 5620 -560
rect 5220 -920 5620 -880
rect 6232 -560 6632 -520
rect 6232 -880 6272 -560
rect 6592 -880 6632 -560
rect 6232 -920 6632 -880
rect 7244 -560 7644 -520
rect 7244 -880 7284 -560
rect 7604 -880 7644 -560
rect 7244 -920 7644 -880
rect 8256 -560 8656 -520
rect 8256 -880 8296 -560
rect 8616 -880 8656 -560
rect 8256 -920 8656 -880
rect 9268 -560 9668 -520
rect 9268 -880 9308 -560
rect 9628 -880 9668 -560
rect 9268 -920 9668 -880
rect 10280 -560 10680 -520
rect 10280 -880 10320 -560
rect 10640 -880 10680 -560
rect 10280 -920 10680 -880
rect 11292 -560 11692 -520
rect 11292 -880 11332 -560
rect 11652 -880 11692 -560
rect 11292 -920 11692 -880
rect 12304 -560 12704 -520
rect 12304 -880 12344 -560
rect 12664 -880 12704 -560
rect 12304 -920 12704 -880
rect 13316 -560 13716 -520
rect 13316 -880 13356 -560
rect 13676 -880 13716 -560
rect 13316 -920 13716 -880
rect 14328 -560 14728 -520
rect 14328 -880 14368 -560
rect 14688 -880 14728 -560
rect 14328 -920 14728 -880
rect 15340 -560 15740 -520
rect 15340 -880 15380 -560
rect 15700 -880 15740 -560
rect 15340 -920 15740 -880
rect 16352 -560 16752 -520
rect 16352 -880 16392 -560
rect 16712 -880 16752 -560
rect 16352 -920 16752 -880
rect 17364 -560 17764 -520
rect 17364 -880 17404 -560
rect 17724 -880 17764 -560
rect 17364 -920 17764 -880
rect 18376 -560 18776 -520
rect 18376 -880 18416 -560
rect 18736 -880 18776 -560
rect 18376 -920 18776 -880
rect 19388 -560 19788 -520
rect 19388 -880 19428 -560
rect 19748 -880 19788 -560
rect 19388 -920 19788 -880
rect 20400 -560 20800 -520
rect 20400 -880 20440 -560
rect 20760 -880 20800 -560
rect 20400 -920 20800 -880
rect 21412 -560 21812 -520
rect 21412 -880 21452 -560
rect 21772 -880 21812 -560
rect 21412 -920 21812 -880
rect 22424 -560 22824 -520
rect 22424 -880 22464 -560
rect 22784 -880 22824 -560
rect 22424 -920 22824 -880
rect 23436 -560 23836 -520
rect 23436 -880 23476 -560
rect 23796 -880 23836 -560
rect 23436 -920 23836 -880
rect 24448 -560 24848 -520
rect 24448 -880 24488 -560
rect 24808 -880 24848 -560
rect 24448 -920 24848 -880
rect 25460 -560 25860 -520
rect 25460 -880 25500 -560
rect 25820 -880 25860 -560
rect 25460 -920 25860 -880
rect 26472 -560 26872 -520
rect 26472 -880 26512 -560
rect 26832 -880 26872 -560
rect 26472 -920 26872 -880
rect 27484 -560 27884 -520
rect 27484 -880 27524 -560
rect 27844 -880 27884 -560
rect 27484 -920 27884 -880
rect 28496 -560 28896 -520
rect 28496 -880 28536 -560
rect 28856 -880 28896 -560
rect 28496 -920 28896 -880
rect 29508 -560 29908 -520
rect 29508 -880 29548 -560
rect 29868 -880 29908 -560
rect 29508 -920 29908 -880
rect 30520 -560 30920 -520
rect 30520 -880 30560 -560
rect 30880 -880 30920 -560
rect 30520 -920 30920 -880
rect 31532 -560 31932 -520
rect 31532 -880 31572 -560
rect 31892 -880 31932 -560
rect 31532 -920 31932 -880
rect -32224 -1280 -31824 -1240
rect -32224 -1600 -32184 -1280
rect -31864 -1600 -31824 -1280
rect -32224 -1640 -31824 -1600
rect -31212 -1280 -30812 -1240
rect -31212 -1600 -31172 -1280
rect -30852 -1600 -30812 -1280
rect -31212 -1640 -30812 -1600
rect -30200 -1280 -29800 -1240
rect -30200 -1600 -30160 -1280
rect -29840 -1600 -29800 -1280
rect -30200 -1640 -29800 -1600
rect -29188 -1280 -28788 -1240
rect -29188 -1600 -29148 -1280
rect -28828 -1600 -28788 -1280
rect -29188 -1640 -28788 -1600
rect -28176 -1280 -27776 -1240
rect -28176 -1600 -28136 -1280
rect -27816 -1600 -27776 -1280
rect -28176 -1640 -27776 -1600
rect -27164 -1280 -26764 -1240
rect -27164 -1600 -27124 -1280
rect -26804 -1600 -26764 -1280
rect -27164 -1640 -26764 -1600
rect -26152 -1280 -25752 -1240
rect -26152 -1600 -26112 -1280
rect -25792 -1600 -25752 -1280
rect -26152 -1640 -25752 -1600
rect -25140 -1280 -24740 -1240
rect -25140 -1600 -25100 -1280
rect -24780 -1600 -24740 -1280
rect -25140 -1640 -24740 -1600
rect -24128 -1280 -23728 -1240
rect -24128 -1600 -24088 -1280
rect -23768 -1600 -23728 -1280
rect -24128 -1640 -23728 -1600
rect -23116 -1280 -22716 -1240
rect -23116 -1600 -23076 -1280
rect -22756 -1600 -22716 -1280
rect -23116 -1640 -22716 -1600
rect -22104 -1280 -21704 -1240
rect -22104 -1600 -22064 -1280
rect -21744 -1600 -21704 -1280
rect -22104 -1640 -21704 -1600
rect -21092 -1280 -20692 -1240
rect -21092 -1600 -21052 -1280
rect -20732 -1600 -20692 -1280
rect -21092 -1640 -20692 -1600
rect -20080 -1280 -19680 -1240
rect -20080 -1600 -20040 -1280
rect -19720 -1600 -19680 -1280
rect -20080 -1640 -19680 -1600
rect -19068 -1280 -18668 -1240
rect -19068 -1600 -19028 -1280
rect -18708 -1600 -18668 -1280
rect -19068 -1640 -18668 -1600
rect -18056 -1280 -17656 -1240
rect -18056 -1600 -18016 -1280
rect -17696 -1600 -17656 -1280
rect -18056 -1640 -17656 -1600
rect -17044 -1280 -16644 -1240
rect -17044 -1600 -17004 -1280
rect -16684 -1600 -16644 -1280
rect -17044 -1640 -16644 -1600
rect -16032 -1280 -15632 -1240
rect -16032 -1600 -15992 -1280
rect -15672 -1600 -15632 -1280
rect -16032 -1640 -15632 -1600
rect -15020 -1280 -14620 -1240
rect -15020 -1600 -14980 -1280
rect -14660 -1600 -14620 -1280
rect -15020 -1640 -14620 -1600
rect -14008 -1280 -13608 -1240
rect -14008 -1600 -13968 -1280
rect -13648 -1600 -13608 -1280
rect -14008 -1640 -13608 -1600
rect -12996 -1280 -12596 -1240
rect -12996 -1600 -12956 -1280
rect -12636 -1600 -12596 -1280
rect -12996 -1640 -12596 -1600
rect -11984 -1280 -11584 -1240
rect -11984 -1600 -11944 -1280
rect -11624 -1600 -11584 -1280
rect -11984 -1640 -11584 -1600
rect -10972 -1280 -10572 -1240
rect -10972 -1600 -10932 -1280
rect -10612 -1600 -10572 -1280
rect -10972 -1640 -10572 -1600
rect -9960 -1280 -9560 -1240
rect -9960 -1600 -9920 -1280
rect -9600 -1600 -9560 -1280
rect -9960 -1640 -9560 -1600
rect -8948 -1280 -8548 -1240
rect -8948 -1600 -8908 -1280
rect -8588 -1600 -8548 -1280
rect -8948 -1640 -8548 -1600
rect -7936 -1280 -7536 -1240
rect -7936 -1600 -7896 -1280
rect -7576 -1600 -7536 -1280
rect -7936 -1640 -7536 -1600
rect -6924 -1280 -6524 -1240
rect -6924 -1600 -6884 -1280
rect -6564 -1600 -6524 -1280
rect -6924 -1640 -6524 -1600
rect -5912 -1280 -5512 -1240
rect -5912 -1600 -5872 -1280
rect -5552 -1600 -5512 -1280
rect -5912 -1640 -5512 -1600
rect -4900 -1280 -4500 -1240
rect -4900 -1600 -4860 -1280
rect -4540 -1600 -4500 -1280
rect -4900 -1640 -4500 -1600
rect -3888 -1280 -3488 -1240
rect -3888 -1600 -3848 -1280
rect -3528 -1600 -3488 -1280
rect -3888 -1640 -3488 -1600
rect -2876 -1280 -2476 -1240
rect -2876 -1600 -2836 -1280
rect -2516 -1600 -2476 -1280
rect -2876 -1640 -2476 -1600
rect -1864 -1280 -1464 -1240
rect -1864 -1600 -1824 -1280
rect -1504 -1600 -1464 -1280
rect -1864 -1640 -1464 -1600
rect -852 -1280 -452 -1240
rect -852 -1600 -812 -1280
rect -492 -1600 -452 -1280
rect -852 -1640 -452 -1600
rect 160 -1280 560 -1240
rect 160 -1600 200 -1280
rect 520 -1600 560 -1280
rect 160 -1640 560 -1600
rect 1172 -1280 1572 -1240
rect 1172 -1600 1212 -1280
rect 1532 -1600 1572 -1280
rect 1172 -1640 1572 -1600
rect 2184 -1280 2584 -1240
rect 2184 -1600 2224 -1280
rect 2544 -1600 2584 -1280
rect 2184 -1640 2584 -1600
rect 3196 -1280 3596 -1240
rect 3196 -1600 3236 -1280
rect 3556 -1600 3596 -1280
rect 3196 -1640 3596 -1600
rect 4208 -1280 4608 -1240
rect 4208 -1600 4248 -1280
rect 4568 -1600 4608 -1280
rect 4208 -1640 4608 -1600
rect 5220 -1280 5620 -1240
rect 5220 -1600 5260 -1280
rect 5580 -1600 5620 -1280
rect 5220 -1640 5620 -1600
rect 6232 -1280 6632 -1240
rect 6232 -1600 6272 -1280
rect 6592 -1600 6632 -1280
rect 6232 -1640 6632 -1600
rect 7244 -1280 7644 -1240
rect 7244 -1600 7284 -1280
rect 7604 -1600 7644 -1280
rect 7244 -1640 7644 -1600
rect 8256 -1280 8656 -1240
rect 8256 -1600 8296 -1280
rect 8616 -1600 8656 -1280
rect 8256 -1640 8656 -1600
rect 9268 -1280 9668 -1240
rect 9268 -1600 9308 -1280
rect 9628 -1600 9668 -1280
rect 9268 -1640 9668 -1600
rect 10280 -1280 10680 -1240
rect 10280 -1600 10320 -1280
rect 10640 -1600 10680 -1280
rect 10280 -1640 10680 -1600
rect 11292 -1280 11692 -1240
rect 11292 -1600 11332 -1280
rect 11652 -1600 11692 -1280
rect 11292 -1640 11692 -1600
rect 12304 -1280 12704 -1240
rect 12304 -1600 12344 -1280
rect 12664 -1600 12704 -1280
rect 12304 -1640 12704 -1600
rect 13316 -1280 13716 -1240
rect 13316 -1600 13356 -1280
rect 13676 -1600 13716 -1280
rect 13316 -1640 13716 -1600
rect 14328 -1280 14728 -1240
rect 14328 -1600 14368 -1280
rect 14688 -1600 14728 -1280
rect 14328 -1640 14728 -1600
rect 15340 -1280 15740 -1240
rect 15340 -1600 15380 -1280
rect 15700 -1600 15740 -1280
rect 15340 -1640 15740 -1600
rect 16352 -1280 16752 -1240
rect 16352 -1600 16392 -1280
rect 16712 -1600 16752 -1280
rect 16352 -1640 16752 -1600
rect 17364 -1280 17764 -1240
rect 17364 -1600 17404 -1280
rect 17724 -1600 17764 -1280
rect 17364 -1640 17764 -1600
rect 18376 -1280 18776 -1240
rect 18376 -1600 18416 -1280
rect 18736 -1600 18776 -1280
rect 18376 -1640 18776 -1600
rect 19388 -1280 19788 -1240
rect 19388 -1600 19428 -1280
rect 19748 -1600 19788 -1280
rect 19388 -1640 19788 -1600
rect 20400 -1280 20800 -1240
rect 20400 -1600 20440 -1280
rect 20760 -1600 20800 -1280
rect 20400 -1640 20800 -1600
rect 21412 -1280 21812 -1240
rect 21412 -1600 21452 -1280
rect 21772 -1600 21812 -1280
rect 21412 -1640 21812 -1600
rect 22424 -1280 22824 -1240
rect 22424 -1600 22464 -1280
rect 22784 -1600 22824 -1280
rect 22424 -1640 22824 -1600
rect 23436 -1280 23836 -1240
rect 23436 -1600 23476 -1280
rect 23796 -1600 23836 -1280
rect 23436 -1640 23836 -1600
rect 24448 -1280 24848 -1240
rect 24448 -1600 24488 -1280
rect 24808 -1600 24848 -1280
rect 24448 -1640 24848 -1600
rect 25460 -1280 25860 -1240
rect 25460 -1600 25500 -1280
rect 25820 -1600 25860 -1280
rect 25460 -1640 25860 -1600
rect 26472 -1280 26872 -1240
rect 26472 -1600 26512 -1280
rect 26832 -1600 26872 -1280
rect 26472 -1640 26872 -1600
rect 27484 -1280 27884 -1240
rect 27484 -1600 27524 -1280
rect 27844 -1600 27884 -1280
rect 27484 -1640 27884 -1600
rect 28496 -1280 28896 -1240
rect 28496 -1600 28536 -1280
rect 28856 -1600 28896 -1280
rect 28496 -1640 28896 -1600
rect 29508 -1280 29908 -1240
rect 29508 -1600 29548 -1280
rect 29868 -1600 29908 -1280
rect 29508 -1640 29908 -1600
rect 30520 -1280 30920 -1240
rect 30520 -1600 30560 -1280
rect 30880 -1600 30920 -1280
rect 30520 -1640 30920 -1600
rect 31532 -1280 31932 -1240
rect 31532 -1600 31572 -1280
rect 31892 -1600 31932 -1280
rect 31532 -1640 31932 -1600
rect -32224 -2000 -31824 -1960
rect -32224 -2320 -32184 -2000
rect -31864 -2320 -31824 -2000
rect -32224 -2360 -31824 -2320
rect -31212 -2000 -30812 -1960
rect -31212 -2320 -31172 -2000
rect -30852 -2320 -30812 -2000
rect -31212 -2360 -30812 -2320
rect -30200 -2000 -29800 -1960
rect -30200 -2320 -30160 -2000
rect -29840 -2320 -29800 -2000
rect -30200 -2360 -29800 -2320
rect -29188 -2000 -28788 -1960
rect -29188 -2320 -29148 -2000
rect -28828 -2320 -28788 -2000
rect -29188 -2360 -28788 -2320
rect -28176 -2000 -27776 -1960
rect -28176 -2320 -28136 -2000
rect -27816 -2320 -27776 -2000
rect -28176 -2360 -27776 -2320
rect -27164 -2000 -26764 -1960
rect -27164 -2320 -27124 -2000
rect -26804 -2320 -26764 -2000
rect -27164 -2360 -26764 -2320
rect -26152 -2000 -25752 -1960
rect -26152 -2320 -26112 -2000
rect -25792 -2320 -25752 -2000
rect -26152 -2360 -25752 -2320
rect -25140 -2000 -24740 -1960
rect -25140 -2320 -25100 -2000
rect -24780 -2320 -24740 -2000
rect -25140 -2360 -24740 -2320
rect -24128 -2000 -23728 -1960
rect -24128 -2320 -24088 -2000
rect -23768 -2320 -23728 -2000
rect -24128 -2360 -23728 -2320
rect -23116 -2000 -22716 -1960
rect -23116 -2320 -23076 -2000
rect -22756 -2320 -22716 -2000
rect -23116 -2360 -22716 -2320
rect -22104 -2000 -21704 -1960
rect -22104 -2320 -22064 -2000
rect -21744 -2320 -21704 -2000
rect -22104 -2360 -21704 -2320
rect -21092 -2000 -20692 -1960
rect -21092 -2320 -21052 -2000
rect -20732 -2320 -20692 -2000
rect -21092 -2360 -20692 -2320
rect -20080 -2000 -19680 -1960
rect -20080 -2320 -20040 -2000
rect -19720 -2320 -19680 -2000
rect -20080 -2360 -19680 -2320
rect -19068 -2000 -18668 -1960
rect -19068 -2320 -19028 -2000
rect -18708 -2320 -18668 -2000
rect -19068 -2360 -18668 -2320
rect -18056 -2000 -17656 -1960
rect -18056 -2320 -18016 -2000
rect -17696 -2320 -17656 -2000
rect -18056 -2360 -17656 -2320
rect -17044 -2000 -16644 -1960
rect -17044 -2320 -17004 -2000
rect -16684 -2320 -16644 -2000
rect -17044 -2360 -16644 -2320
rect -16032 -2000 -15632 -1960
rect -16032 -2320 -15992 -2000
rect -15672 -2320 -15632 -2000
rect -16032 -2360 -15632 -2320
rect -15020 -2000 -14620 -1960
rect -15020 -2320 -14980 -2000
rect -14660 -2320 -14620 -2000
rect -15020 -2360 -14620 -2320
rect -14008 -2000 -13608 -1960
rect -14008 -2320 -13968 -2000
rect -13648 -2320 -13608 -2000
rect -14008 -2360 -13608 -2320
rect -12996 -2000 -12596 -1960
rect -12996 -2320 -12956 -2000
rect -12636 -2320 -12596 -2000
rect -12996 -2360 -12596 -2320
rect -11984 -2000 -11584 -1960
rect -11984 -2320 -11944 -2000
rect -11624 -2320 -11584 -2000
rect -11984 -2360 -11584 -2320
rect -10972 -2000 -10572 -1960
rect -10972 -2320 -10932 -2000
rect -10612 -2320 -10572 -2000
rect -10972 -2360 -10572 -2320
rect -9960 -2000 -9560 -1960
rect -9960 -2320 -9920 -2000
rect -9600 -2320 -9560 -2000
rect -9960 -2360 -9560 -2320
rect -8948 -2000 -8548 -1960
rect -8948 -2320 -8908 -2000
rect -8588 -2320 -8548 -2000
rect -8948 -2360 -8548 -2320
rect -7936 -2000 -7536 -1960
rect -7936 -2320 -7896 -2000
rect -7576 -2320 -7536 -2000
rect -7936 -2360 -7536 -2320
rect -6924 -2000 -6524 -1960
rect -6924 -2320 -6884 -2000
rect -6564 -2320 -6524 -2000
rect -6924 -2360 -6524 -2320
rect -5912 -2000 -5512 -1960
rect -5912 -2320 -5872 -2000
rect -5552 -2320 -5512 -2000
rect -5912 -2360 -5512 -2320
rect -4900 -2000 -4500 -1960
rect -4900 -2320 -4860 -2000
rect -4540 -2320 -4500 -2000
rect -4900 -2360 -4500 -2320
rect -3888 -2000 -3488 -1960
rect -3888 -2320 -3848 -2000
rect -3528 -2320 -3488 -2000
rect -3888 -2360 -3488 -2320
rect -2876 -2000 -2476 -1960
rect -2876 -2320 -2836 -2000
rect -2516 -2320 -2476 -2000
rect -2876 -2360 -2476 -2320
rect -1864 -2000 -1464 -1960
rect -1864 -2320 -1824 -2000
rect -1504 -2320 -1464 -2000
rect -1864 -2360 -1464 -2320
rect -852 -2000 -452 -1960
rect -852 -2320 -812 -2000
rect -492 -2320 -452 -2000
rect -852 -2360 -452 -2320
rect 160 -2000 560 -1960
rect 160 -2320 200 -2000
rect 520 -2320 560 -2000
rect 160 -2360 560 -2320
rect 1172 -2000 1572 -1960
rect 1172 -2320 1212 -2000
rect 1532 -2320 1572 -2000
rect 1172 -2360 1572 -2320
rect 2184 -2000 2584 -1960
rect 2184 -2320 2224 -2000
rect 2544 -2320 2584 -2000
rect 2184 -2360 2584 -2320
rect 3196 -2000 3596 -1960
rect 3196 -2320 3236 -2000
rect 3556 -2320 3596 -2000
rect 3196 -2360 3596 -2320
rect 4208 -2000 4608 -1960
rect 4208 -2320 4248 -2000
rect 4568 -2320 4608 -2000
rect 4208 -2360 4608 -2320
rect 5220 -2000 5620 -1960
rect 5220 -2320 5260 -2000
rect 5580 -2320 5620 -2000
rect 5220 -2360 5620 -2320
rect 6232 -2000 6632 -1960
rect 6232 -2320 6272 -2000
rect 6592 -2320 6632 -2000
rect 6232 -2360 6632 -2320
rect 7244 -2000 7644 -1960
rect 7244 -2320 7284 -2000
rect 7604 -2320 7644 -2000
rect 7244 -2360 7644 -2320
rect 8256 -2000 8656 -1960
rect 8256 -2320 8296 -2000
rect 8616 -2320 8656 -2000
rect 8256 -2360 8656 -2320
rect 9268 -2000 9668 -1960
rect 9268 -2320 9308 -2000
rect 9628 -2320 9668 -2000
rect 9268 -2360 9668 -2320
rect 10280 -2000 10680 -1960
rect 10280 -2320 10320 -2000
rect 10640 -2320 10680 -2000
rect 10280 -2360 10680 -2320
rect 11292 -2000 11692 -1960
rect 11292 -2320 11332 -2000
rect 11652 -2320 11692 -2000
rect 11292 -2360 11692 -2320
rect 12304 -2000 12704 -1960
rect 12304 -2320 12344 -2000
rect 12664 -2320 12704 -2000
rect 12304 -2360 12704 -2320
rect 13316 -2000 13716 -1960
rect 13316 -2320 13356 -2000
rect 13676 -2320 13716 -2000
rect 13316 -2360 13716 -2320
rect 14328 -2000 14728 -1960
rect 14328 -2320 14368 -2000
rect 14688 -2320 14728 -2000
rect 14328 -2360 14728 -2320
rect 15340 -2000 15740 -1960
rect 15340 -2320 15380 -2000
rect 15700 -2320 15740 -2000
rect 15340 -2360 15740 -2320
rect 16352 -2000 16752 -1960
rect 16352 -2320 16392 -2000
rect 16712 -2320 16752 -2000
rect 16352 -2360 16752 -2320
rect 17364 -2000 17764 -1960
rect 17364 -2320 17404 -2000
rect 17724 -2320 17764 -2000
rect 17364 -2360 17764 -2320
rect 18376 -2000 18776 -1960
rect 18376 -2320 18416 -2000
rect 18736 -2320 18776 -2000
rect 18376 -2360 18776 -2320
rect 19388 -2000 19788 -1960
rect 19388 -2320 19428 -2000
rect 19748 -2320 19788 -2000
rect 19388 -2360 19788 -2320
rect 20400 -2000 20800 -1960
rect 20400 -2320 20440 -2000
rect 20760 -2320 20800 -2000
rect 20400 -2360 20800 -2320
rect 21412 -2000 21812 -1960
rect 21412 -2320 21452 -2000
rect 21772 -2320 21812 -2000
rect 21412 -2360 21812 -2320
rect 22424 -2000 22824 -1960
rect 22424 -2320 22464 -2000
rect 22784 -2320 22824 -2000
rect 22424 -2360 22824 -2320
rect 23436 -2000 23836 -1960
rect 23436 -2320 23476 -2000
rect 23796 -2320 23836 -2000
rect 23436 -2360 23836 -2320
rect 24448 -2000 24848 -1960
rect 24448 -2320 24488 -2000
rect 24808 -2320 24848 -2000
rect 24448 -2360 24848 -2320
rect 25460 -2000 25860 -1960
rect 25460 -2320 25500 -2000
rect 25820 -2320 25860 -2000
rect 25460 -2360 25860 -2320
rect 26472 -2000 26872 -1960
rect 26472 -2320 26512 -2000
rect 26832 -2320 26872 -2000
rect 26472 -2360 26872 -2320
rect 27484 -2000 27884 -1960
rect 27484 -2320 27524 -2000
rect 27844 -2320 27884 -2000
rect 27484 -2360 27884 -2320
rect 28496 -2000 28896 -1960
rect 28496 -2320 28536 -2000
rect 28856 -2320 28896 -2000
rect 28496 -2360 28896 -2320
rect 29508 -2000 29908 -1960
rect 29508 -2320 29548 -2000
rect 29868 -2320 29908 -2000
rect 29508 -2360 29908 -2320
rect 30520 -2000 30920 -1960
rect 30520 -2320 30560 -2000
rect 30880 -2320 30920 -2000
rect 30520 -2360 30920 -2320
rect 31532 -2000 31932 -1960
rect 31532 -2320 31572 -2000
rect 31892 -2320 31932 -2000
rect 31532 -2360 31932 -2320
<< mimcapcontact >>
rect -32184 2000 -31864 2320
rect -31172 2000 -30852 2320
rect -30160 2000 -29840 2320
rect -29148 2000 -28828 2320
rect -28136 2000 -27816 2320
rect -27124 2000 -26804 2320
rect -26112 2000 -25792 2320
rect -25100 2000 -24780 2320
rect -24088 2000 -23768 2320
rect -23076 2000 -22756 2320
rect -22064 2000 -21744 2320
rect -21052 2000 -20732 2320
rect -20040 2000 -19720 2320
rect -19028 2000 -18708 2320
rect -18016 2000 -17696 2320
rect -17004 2000 -16684 2320
rect -15992 2000 -15672 2320
rect -14980 2000 -14660 2320
rect -13968 2000 -13648 2320
rect -12956 2000 -12636 2320
rect -11944 2000 -11624 2320
rect -10932 2000 -10612 2320
rect -9920 2000 -9600 2320
rect -8908 2000 -8588 2320
rect -7896 2000 -7576 2320
rect -6884 2000 -6564 2320
rect -5872 2000 -5552 2320
rect -4860 2000 -4540 2320
rect -3848 2000 -3528 2320
rect -2836 2000 -2516 2320
rect -1824 2000 -1504 2320
rect -812 2000 -492 2320
rect 200 2000 520 2320
rect 1212 2000 1532 2320
rect 2224 2000 2544 2320
rect 3236 2000 3556 2320
rect 4248 2000 4568 2320
rect 5260 2000 5580 2320
rect 6272 2000 6592 2320
rect 7284 2000 7604 2320
rect 8296 2000 8616 2320
rect 9308 2000 9628 2320
rect 10320 2000 10640 2320
rect 11332 2000 11652 2320
rect 12344 2000 12664 2320
rect 13356 2000 13676 2320
rect 14368 2000 14688 2320
rect 15380 2000 15700 2320
rect 16392 2000 16712 2320
rect 17404 2000 17724 2320
rect 18416 2000 18736 2320
rect 19428 2000 19748 2320
rect 20440 2000 20760 2320
rect 21452 2000 21772 2320
rect 22464 2000 22784 2320
rect 23476 2000 23796 2320
rect 24488 2000 24808 2320
rect 25500 2000 25820 2320
rect 26512 2000 26832 2320
rect 27524 2000 27844 2320
rect 28536 2000 28856 2320
rect 29548 2000 29868 2320
rect 30560 2000 30880 2320
rect 31572 2000 31892 2320
rect -32184 1280 -31864 1600
rect -31172 1280 -30852 1600
rect -30160 1280 -29840 1600
rect -29148 1280 -28828 1600
rect -28136 1280 -27816 1600
rect -27124 1280 -26804 1600
rect -26112 1280 -25792 1600
rect -25100 1280 -24780 1600
rect -24088 1280 -23768 1600
rect -23076 1280 -22756 1600
rect -22064 1280 -21744 1600
rect -21052 1280 -20732 1600
rect -20040 1280 -19720 1600
rect -19028 1280 -18708 1600
rect -18016 1280 -17696 1600
rect -17004 1280 -16684 1600
rect -15992 1280 -15672 1600
rect -14980 1280 -14660 1600
rect -13968 1280 -13648 1600
rect -12956 1280 -12636 1600
rect -11944 1280 -11624 1600
rect -10932 1280 -10612 1600
rect -9920 1280 -9600 1600
rect -8908 1280 -8588 1600
rect -7896 1280 -7576 1600
rect -6884 1280 -6564 1600
rect -5872 1280 -5552 1600
rect -4860 1280 -4540 1600
rect -3848 1280 -3528 1600
rect -2836 1280 -2516 1600
rect -1824 1280 -1504 1600
rect -812 1280 -492 1600
rect 200 1280 520 1600
rect 1212 1280 1532 1600
rect 2224 1280 2544 1600
rect 3236 1280 3556 1600
rect 4248 1280 4568 1600
rect 5260 1280 5580 1600
rect 6272 1280 6592 1600
rect 7284 1280 7604 1600
rect 8296 1280 8616 1600
rect 9308 1280 9628 1600
rect 10320 1280 10640 1600
rect 11332 1280 11652 1600
rect 12344 1280 12664 1600
rect 13356 1280 13676 1600
rect 14368 1280 14688 1600
rect 15380 1280 15700 1600
rect 16392 1280 16712 1600
rect 17404 1280 17724 1600
rect 18416 1280 18736 1600
rect 19428 1280 19748 1600
rect 20440 1280 20760 1600
rect 21452 1280 21772 1600
rect 22464 1280 22784 1600
rect 23476 1280 23796 1600
rect 24488 1280 24808 1600
rect 25500 1280 25820 1600
rect 26512 1280 26832 1600
rect 27524 1280 27844 1600
rect 28536 1280 28856 1600
rect 29548 1280 29868 1600
rect 30560 1280 30880 1600
rect 31572 1280 31892 1600
rect -32184 560 -31864 880
rect -31172 560 -30852 880
rect -30160 560 -29840 880
rect -29148 560 -28828 880
rect -28136 560 -27816 880
rect -27124 560 -26804 880
rect -26112 560 -25792 880
rect -25100 560 -24780 880
rect -24088 560 -23768 880
rect -23076 560 -22756 880
rect -22064 560 -21744 880
rect -21052 560 -20732 880
rect -20040 560 -19720 880
rect -19028 560 -18708 880
rect -18016 560 -17696 880
rect -17004 560 -16684 880
rect -15992 560 -15672 880
rect -14980 560 -14660 880
rect -13968 560 -13648 880
rect -12956 560 -12636 880
rect -11944 560 -11624 880
rect -10932 560 -10612 880
rect -9920 560 -9600 880
rect -8908 560 -8588 880
rect -7896 560 -7576 880
rect -6884 560 -6564 880
rect -5872 560 -5552 880
rect -4860 560 -4540 880
rect -3848 560 -3528 880
rect -2836 560 -2516 880
rect -1824 560 -1504 880
rect -812 560 -492 880
rect 200 560 520 880
rect 1212 560 1532 880
rect 2224 560 2544 880
rect 3236 560 3556 880
rect 4248 560 4568 880
rect 5260 560 5580 880
rect 6272 560 6592 880
rect 7284 560 7604 880
rect 8296 560 8616 880
rect 9308 560 9628 880
rect 10320 560 10640 880
rect 11332 560 11652 880
rect 12344 560 12664 880
rect 13356 560 13676 880
rect 14368 560 14688 880
rect 15380 560 15700 880
rect 16392 560 16712 880
rect 17404 560 17724 880
rect 18416 560 18736 880
rect 19428 560 19748 880
rect 20440 560 20760 880
rect 21452 560 21772 880
rect 22464 560 22784 880
rect 23476 560 23796 880
rect 24488 560 24808 880
rect 25500 560 25820 880
rect 26512 560 26832 880
rect 27524 560 27844 880
rect 28536 560 28856 880
rect 29548 560 29868 880
rect 30560 560 30880 880
rect 31572 560 31892 880
rect -32184 -160 -31864 160
rect -31172 -160 -30852 160
rect -30160 -160 -29840 160
rect -29148 -160 -28828 160
rect -28136 -160 -27816 160
rect -27124 -160 -26804 160
rect -26112 -160 -25792 160
rect -25100 -160 -24780 160
rect -24088 -160 -23768 160
rect -23076 -160 -22756 160
rect -22064 -160 -21744 160
rect -21052 -160 -20732 160
rect -20040 -160 -19720 160
rect -19028 -160 -18708 160
rect -18016 -160 -17696 160
rect -17004 -160 -16684 160
rect -15992 -160 -15672 160
rect -14980 -160 -14660 160
rect -13968 -160 -13648 160
rect -12956 -160 -12636 160
rect -11944 -160 -11624 160
rect -10932 -160 -10612 160
rect -9920 -160 -9600 160
rect -8908 -160 -8588 160
rect -7896 -160 -7576 160
rect -6884 -160 -6564 160
rect -5872 -160 -5552 160
rect -4860 -160 -4540 160
rect -3848 -160 -3528 160
rect -2836 -160 -2516 160
rect -1824 -160 -1504 160
rect -812 -160 -492 160
rect 200 -160 520 160
rect 1212 -160 1532 160
rect 2224 -160 2544 160
rect 3236 -160 3556 160
rect 4248 -160 4568 160
rect 5260 -160 5580 160
rect 6272 -160 6592 160
rect 7284 -160 7604 160
rect 8296 -160 8616 160
rect 9308 -160 9628 160
rect 10320 -160 10640 160
rect 11332 -160 11652 160
rect 12344 -160 12664 160
rect 13356 -160 13676 160
rect 14368 -160 14688 160
rect 15380 -160 15700 160
rect 16392 -160 16712 160
rect 17404 -160 17724 160
rect 18416 -160 18736 160
rect 19428 -160 19748 160
rect 20440 -160 20760 160
rect 21452 -160 21772 160
rect 22464 -160 22784 160
rect 23476 -160 23796 160
rect 24488 -160 24808 160
rect 25500 -160 25820 160
rect 26512 -160 26832 160
rect 27524 -160 27844 160
rect 28536 -160 28856 160
rect 29548 -160 29868 160
rect 30560 -160 30880 160
rect 31572 -160 31892 160
rect -32184 -880 -31864 -560
rect -31172 -880 -30852 -560
rect -30160 -880 -29840 -560
rect -29148 -880 -28828 -560
rect -28136 -880 -27816 -560
rect -27124 -880 -26804 -560
rect -26112 -880 -25792 -560
rect -25100 -880 -24780 -560
rect -24088 -880 -23768 -560
rect -23076 -880 -22756 -560
rect -22064 -880 -21744 -560
rect -21052 -880 -20732 -560
rect -20040 -880 -19720 -560
rect -19028 -880 -18708 -560
rect -18016 -880 -17696 -560
rect -17004 -880 -16684 -560
rect -15992 -880 -15672 -560
rect -14980 -880 -14660 -560
rect -13968 -880 -13648 -560
rect -12956 -880 -12636 -560
rect -11944 -880 -11624 -560
rect -10932 -880 -10612 -560
rect -9920 -880 -9600 -560
rect -8908 -880 -8588 -560
rect -7896 -880 -7576 -560
rect -6884 -880 -6564 -560
rect -5872 -880 -5552 -560
rect -4860 -880 -4540 -560
rect -3848 -880 -3528 -560
rect -2836 -880 -2516 -560
rect -1824 -880 -1504 -560
rect -812 -880 -492 -560
rect 200 -880 520 -560
rect 1212 -880 1532 -560
rect 2224 -880 2544 -560
rect 3236 -880 3556 -560
rect 4248 -880 4568 -560
rect 5260 -880 5580 -560
rect 6272 -880 6592 -560
rect 7284 -880 7604 -560
rect 8296 -880 8616 -560
rect 9308 -880 9628 -560
rect 10320 -880 10640 -560
rect 11332 -880 11652 -560
rect 12344 -880 12664 -560
rect 13356 -880 13676 -560
rect 14368 -880 14688 -560
rect 15380 -880 15700 -560
rect 16392 -880 16712 -560
rect 17404 -880 17724 -560
rect 18416 -880 18736 -560
rect 19428 -880 19748 -560
rect 20440 -880 20760 -560
rect 21452 -880 21772 -560
rect 22464 -880 22784 -560
rect 23476 -880 23796 -560
rect 24488 -880 24808 -560
rect 25500 -880 25820 -560
rect 26512 -880 26832 -560
rect 27524 -880 27844 -560
rect 28536 -880 28856 -560
rect 29548 -880 29868 -560
rect 30560 -880 30880 -560
rect 31572 -880 31892 -560
rect -32184 -1600 -31864 -1280
rect -31172 -1600 -30852 -1280
rect -30160 -1600 -29840 -1280
rect -29148 -1600 -28828 -1280
rect -28136 -1600 -27816 -1280
rect -27124 -1600 -26804 -1280
rect -26112 -1600 -25792 -1280
rect -25100 -1600 -24780 -1280
rect -24088 -1600 -23768 -1280
rect -23076 -1600 -22756 -1280
rect -22064 -1600 -21744 -1280
rect -21052 -1600 -20732 -1280
rect -20040 -1600 -19720 -1280
rect -19028 -1600 -18708 -1280
rect -18016 -1600 -17696 -1280
rect -17004 -1600 -16684 -1280
rect -15992 -1600 -15672 -1280
rect -14980 -1600 -14660 -1280
rect -13968 -1600 -13648 -1280
rect -12956 -1600 -12636 -1280
rect -11944 -1600 -11624 -1280
rect -10932 -1600 -10612 -1280
rect -9920 -1600 -9600 -1280
rect -8908 -1600 -8588 -1280
rect -7896 -1600 -7576 -1280
rect -6884 -1600 -6564 -1280
rect -5872 -1600 -5552 -1280
rect -4860 -1600 -4540 -1280
rect -3848 -1600 -3528 -1280
rect -2836 -1600 -2516 -1280
rect -1824 -1600 -1504 -1280
rect -812 -1600 -492 -1280
rect 200 -1600 520 -1280
rect 1212 -1600 1532 -1280
rect 2224 -1600 2544 -1280
rect 3236 -1600 3556 -1280
rect 4248 -1600 4568 -1280
rect 5260 -1600 5580 -1280
rect 6272 -1600 6592 -1280
rect 7284 -1600 7604 -1280
rect 8296 -1600 8616 -1280
rect 9308 -1600 9628 -1280
rect 10320 -1600 10640 -1280
rect 11332 -1600 11652 -1280
rect 12344 -1600 12664 -1280
rect 13356 -1600 13676 -1280
rect 14368 -1600 14688 -1280
rect 15380 -1600 15700 -1280
rect 16392 -1600 16712 -1280
rect 17404 -1600 17724 -1280
rect 18416 -1600 18736 -1280
rect 19428 -1600 19748 -1280
rect 20440 -1600 20760 -1280
rect 21452 -1600 21772 -1280
rect 22464 -1600 22784 -1280
rect 23476 -1600 23796 -1280
rect 24488 -1600 24808 -1280
rect 25500 -1600 25820 -1280
rect 26512 -1600 26832 -1280
rect 27524 -1600 27844 -1280
rect 28536 -1600 28856 -1280
rect 29548 -1600 29868 -1280
rect 30560 -1600 30880 -1280
rect 31572 -1600 31892 -1280
rect -32184 -2320 -31864 -2000
rect -31172 -2320 -30852 -2000
rect -30160 -2320 -29840 -2000
rect -29148 -2320 -28828 -2000
rect -28136 -2320 -27816 -2000
rect -27124 -2320 -26804 -2000
rect -26112 -2320 -25792 -2000
rect -25100 -2320 -24780 -2000
rect -24088 -2320 -23768 -2000
rect -23076 -2320 -22756 -2000
rect -22064 -2320 -21744 -2000
rect -21052 -2320 -20732 -2000
rect -20040 -2320 -19720 -2000
rect -19028 -2320 -18708 -2000
rect -18016 -2320 -17696 -2000
rect -17004 -2320 -16684 -2000
rect -15992 -2320 -15672 -2000
rect -14980 -2320 -14660 -2000
rect -13968 -2320 -13648 -2000
rect -12956 -2320 -12636 -2000
rect -11944 -2320 -11624 -2000
rect -10932 -2320 -10612 -2000
rect -9920 -2320 -9600 -2000
rect -8908 -2320 -8588 -2000
rect -7896 -2320 -7576 -2000
rect -6884 -2320 -6564 -2000
rect -5872 -2320 -5552 -2000
rect -4860 -2320 -4540 -2000
rect -3848 -2320 -3528 -2000
rect -2836 -2320 -2516 -2000
rect -1824 -2320 -1504 -2000
rect -812 -2320 -492 -2000
rect 200 -2320 520 -2000
rect 1212 -2320 1532 -2000
rect 2224 -2320 2544 -2000
rect 3236 -2320 3556 -2000
rect 4248 -2320 4568 -2000
rect 5260 -2320 5580 -2000
rect 6272 -2320 6592 -2000
rect 7284 -2320 7604 -2000
rect 8296 -2320 8616 -2000
rect 9308 -2320 9628 -2000
rect 10320 -2320 10640 -2000
rect 11332 -2320 11652 -2000
rect 12344 -2320 12664 -2000
rect 13356 -2320 13676 -2000
rect 14368 -2320 14688 -2000
rect 15380 -2320 15700 -2000
rect 16392 -2320 16712 -2000
rect 17404 -2320 17724 -2000
rect 18416 -2320 18736 -2000
rect 19428 -2320 19748 -2000
rect 20440 -2320 20760 -2000
rect 21452 -2320 21772 -2000
rect 22464 -2320 22784 -2000
rect 23476 -2320 23796 -2000
rect 24488 -2320 24808 -2000
rect 25500 -2320 25820 -2000
rect 26512 -2320 26832 -2000
rect 27524 -2320 27844 -2000
rect 28536 -2320 28856 -2000
rect 29548 -2320 29868 -2000
rect 30560 -2320 30880 -2000
rect 31572 -2320 31892 -2000
<< metal4 >>
rect -32076 2321 -31972 2520
rect -31596 2372 -31492 2520
rect -32185 2320 -31863 2321
rect -32185 2000 -32184 2320
rect -31864 2000 -31863 2320
rect -32185 1999 -31863 2000
rect -32076 1601 -31972 1999
rect -31596 1948 -31576 2372
rect -31512 1948 -31492 2372
rect -31064 2321 -30960 2520
rect -30584 2372 -30480 2520
rect -31173 2320 -30851 2321
rect -31173 2000 -31172 2320
rect -30852 2000 -30851 2320
rect -31173 1999 -30851 2000
rect -31596 1652 -31492 1948
rect -32185 1600 -31863 1601
rect -32185 1280 -32184 1600
rect -31864 1280 -31863 1600
rect -32185 1279 -31863 1280
rect -32076 881 -31972 1279
rect -31596 1228 -31576 1652
rect -31512 1228 -31492 1652
rect -31064 1601 -30960 1999
rect -30584 1948 -30564 2372
rect -30500 1948 -30480 2372
rect -30052 2321 -29948 2520
rect -29572 2372 -29468 2520
rect -30161 2320 -29839 2321
rect -30161 2000 -30160 2320
rect -29840 2000 -29839 2320
rect -30161 1999 -29839 2000
rect -30584 1652 -30480 1948
rect -31173 1600 -30851 1601
rect -31173 1280 -31172 1600
rect -30852 1280 -30851 1600
rect -31173 1279 -30851 1280
rect -31596 932 -31492 1228
rect -32185 880 -31863 881
rect -32185 560 -32184 880
rect -31864 560 -31863 880
rect -32185 559 -31863 560
rect -32076 161 -31972 559
rect -31596 508 -31576 932
rect -31512 508 -31492 932
rect -31064 881 -30960 1279
rect -30584 1228 -30564 1652
rect -30500 1228 -30480 1652
rect -30052 1601 -29948 1999
rect -29572 1948 -29552 2372
rect -29488 1948 -29468 2372
rect -29040 2321 -28936 2520
rect -28560 2372 -28456 2520
rect -29149 2320 -28827 2321
rect -29149 2000 -29148 2320
rect -28828 2000 -28827 2320
rect -29149 1999 -28827 2000
rect -29572 1652 -29468 1948
rect -30161 1600 -29839 1601
rect -30161 1280 -30160 1600
rect -29840 1280 -29839 1600
rect -30161 1279 -29839 1280
rect -30584 932 -30480 1228
rect -31173 880 -30851 881
rect -31173 560 -31172 880
rect -30852 560 -30851 880
rect -31173 559 -30851 560
rect -31596 212 -31492 508
rect -32185 160 -31863 161
rect -32185 -160 -32184 160
rect -31864 -160 -31863 160
rect -32185 -161 -31863 -160
rect -32076 -559 -31972 -161
rect -31596 -212 -31576 212
rect -31512 -212 -31492 212
rect -31064 161 -30960 559
rect -30584 508 -30564 932
rect -30500 508 -30480 932
rect -30052 881 -29948 1279
rect -29572 1228 -29552 1652
rect -29488 1228 -29468 1652
rect -29040 1601 -28936 1999
rect -28560 1948 -28540 2372
rect -28476 1948 -28456 2372
rect -28028 2321 -27924 2520
rect -27548 2372 -27444 2520
rect -28137 2320 -27815 2321
rect -28137 2000 -28136 2320
rect -27816 2000 -27815 2320
rect -28137 1999 -27815 2000
rect -28560 1652 -28456 1948
rect -29149 1600 -28827 1601
rect -29149 1280 -29148 1600
rect -28828 1280 -28827 1600
rect -29149 1279 -28827 1280
rect -29572 932 -29468 1228
rect -30161 880 -29839 881
rect -30161 560 -30160 880
rect -29840 560 -29839 880
rect -30161 559 -29839 560
rect -30584 212 -30480 508
rect -31173 160 -30851 161
rect -31173 -160 -31172 160
rect -30852 -160 -30851 160
rect -31173 -161 -30851 -160
rect -31596 -508 -31492 -212
rect -32185 -560 -31863 -559
rect -32185 -880 -32184 -560
rect -31864 -880 -31863 -560
rect -32185 -881 -31863 -880
rect -32076 -1279 -31972 -881
rect -31596 -932 -31576 -508
rect -31512 -932 -31492 -508
rect -31064 -559 -30960 -161
rect -30584 -212 -30564 212
rect -30500 -212 -30480 212
rect -30052 161 -29948 559
rect -29572 508 -29552 932
rect -29488 508 -29468 932
rect -29040 881 -28936 1279
rect -28560 1228 -28540 1652
rect -28476 1228 -28456 1652
rect -28028 1601 -27924 1999
rect -27548 1948 -27528 2372
rect -27464 1948 -27444 2372
rect -27016 2321 -26912 2520
rect -26536 2372 -26432 2520
rect -27125 2320 -26803 2321
rect -27125 2000 -27124 2320
rect -26804 2000 -26803 2320
rect -27125 1999 -26803 2000
rect -27548 1652 -27444 1948
rect -28137 1600 -27815 1601
rect -28137 1280 -28136 1600
rect -27816 1280 -27815 1600
rect -28137 1279 -27815 1280
rect -28560 932 -28456 1228
rect -29149 880 -28827 881
rect -29149 560 -29148 880
rect -28828 560 -28827 880
rect -29149 559 -28827 560
rect -29572 212 -29468 508
rect -30161 160 -29839 161
rect -30161 -160 -30160 160
rect -29840 -160 -29839 160
rect -30161 -161 -29839 -160
rect -30584 -508 -30480 -212
rect -31173 -560 -30851 -559
rect -31173 -880 -31172 -560
rect -30852 -880 -30851 -560
rect -31173 -881 -30851 -880
rect -31596 -1228 -31492 -932
rect -32185 -1280 -31863 -1279
rect -32185 -1600 -32184 -1280
rect -31864 -1600 -31863 -1280
rect -32185 -1601 -31863 -1600
rect -32076 -1999 -31972 -1601
rect -31596 -1652 -31576 -1228
rect -31512 -1652 -31492 -1228
rect -31064 -1279 -30960 -881
rect -30584 -932 -30564 -508
rect -30500 -932 -30480 -508
rect -30052 -559 -29948 -161
rect -29572 -212 -29552 212
rect -29488 -212 -29468 212
rect -29040 161 -28936 559
rect -28560 508 -28540 932
rect -28476 508 -28456 932
rect -28028 881 -27924 1279
rect -27548 1228 -27528 1652
rect -27464 1228 -27444 1652
rect -27016 1601 -26912 1999
rect -26536 1948 -26516 2372
rect -26452 1948 -26432 2372
rect -26004 2321 -25900 2520
rect -25524 2372 -25420 2520
rect -26113 2320 -25791 2321
rect -26113 2000 -26112 2320
rect -25792 2000 -25791 2320
rect -26113 1999 -25791 2000
rect -26536 1652 -26432 1948
rect -27125 1600 -26803 1601
rect -27125 1280 -27124 1600
rect -26804 1280 -26803 1600
rect -27125 1279 -26803 1280
rect -27548 932 -27444 1228
rect -28137 880 -27815 881
rect -28137 560 -28136 880
rect -27816 560 -27815 880
rect -28137 559 -27815 560
rect -28560 212 -28456 508
rect -29149 160 -28827 161
rect -29149 -160 -29148 160
rect -28828 -160 -28827 160
rect -29149 -161 -28827 -160
rect -29572 -508 -29468 -212
rect -30161 -560 -29839 -559
rect -30161 -880 -30160 -560
rect -29840 -880 -29839 -560
rect -30161 -881 -29839 -880
rect -30584 -1228 -30480 -932
rect -31173 -1280 -30851 -1279
rect -31173 -1600 -31172 -1280
rect -30852 -1600 -30851 -1280
rect -31173 -1601 -30851 -1600
rect -31596 -1948 -31492 -1652
rect -32185 -2000 -31863 -1999
rect -32185 -2320 -32184 -2000
rect -31864 -2320 -31863 -2000
rect -32185 -2321 -31863 -2320
rect -32076 -2520 -31972 -2321
rect -31596 -2372 -31576 -1948
rect -31512 -2372 -31492 -1948
rect -31064 -1999 -30960 -1601
rect -30584 -1652 -30564 -1228
rect -30500 -1652 -30480 -1228
rect -30052 -1279 -29948 -881
rect -29572 -932 -29552 -508
rect -29488 -932 -29468 -508
rect -29040 -559 -28936 -161
rect -28560 -212 -28540 212
rect -28476 -212 -28456 212
rect -28028 161 -27924 559
rect -27548 508 -27528 932
rect -27464 508 -27444 932
rect -27016 881 -26912 1279
rect -26536 1228 -26516 1652
rect -26452 1228 -26432 1652
rect -26004 1601 -25900 1999
rect -25524 1948 -25504 2372
rect -25440 1948 -25420 2372
rect -24992 2321 -24888 2520
rect -24512 2372 -24408 2520
rect -25101 2320 -24779 2321
rect -25101 2000 -25100 2320
rect -24780 2000 -24779 2320
rect -25101 1999 -24779 2000
rect -25524 1652 -25420 1948
rect -26113 1600 -25791 1601
rect -26113 1280 -26112 1600
rect -25792 1280 -25791 1600
rect -26113 1279 -25791 1280
rect -26536 932 -26432 1228
rect -27125 880 -26803 881
rect -27125 560 -27124 880
rect -26804 560 -26803 880
rect -27125 559 -26803 560
rect -27548 212 -27444 508
rect -28137 160 -27815 161
rect -28137 -160 -28136 160
rect -27816 -160 -27815 160
rect -28137 -161 -27815 -160
rect -28560 -508 -28456 -212
rect -29149 -560 -28827 -559
rect -29149 -880 -29148 -560
rect -28828 -880 -28827 -560
rect -29149 -881 -28827 -880
rect -29572 -1228 -29468 -932
rect -30161 -1280 -29839 -1279
rect -30161 -1600 -30160 -1280
rect -29840 -1600 -29839 -1280
rect -30161 -1601 -29839 -1600
rect -30584 -1948 -30480 -1652
rect -31173 -2000 -30851 -1999
rect -31173 -2320 -31172 -2000
rect -30852 -2320 -30851 -2000
rect -31173 -2321 -30851 -2320
rect -31596 -2520 -31492 -2372
rect -31064 -2520 -30960 -2321
rect -30584 -2372 -30564 -1948
rect -30500 -2372 -30480 -1948
rect -30052 -1999 -29948 -1601
rect -29572 -1652 -29552 -1228
rect -29488 -1652 -29468 -1228
rect -29040 -1279 -28936 -881
rect -28560 -932 -28540 -508
rect -28476 -932 -28456 -508
rect -28028 -559 -27924 -161
rect -27548 -212 -27528 212
rect -27464 -212 -27444 212
rect -27016 161 -26912 559
rect -26536 508 -26516 932
rect -26452 508 -26432 932
rect -26004 881 -25900 1279
rect -25524 1228 -25504 1652
rect -25440 1228 -25420 1652
rect -24992 1601 -24888 1999
rect -24512 1948 -24492 2372
rect -24428 1948 -24408 2372
rect -23980 2321 -23876 2520
rect -23500 2372 -23396 2520
rect -24089 2320 -23767 2321
rect -24089 2000 -24088 2320
rect -23768 2000 -23767 2320
rect -24089 1999 -23767 2000
rect -24512 1652 -24408 1948
rect -25101 1600 -24779 1601
rect -25101 1280 -25100 1600
rect -24780 1280 -24779 1600
rect -25101 1279 -24779 1280
rect -25524 932 -25420 1228
rect -26113 880 -25791 881
rect -26113 560 -26112 880
rect -25792 560 -25791 880
rect -26113 559 -25791 560
rect -26536 212 -26432 508
rect -27125 160 -26803 161
rect -27125 -160 -27124 160
rect -26804 -160 -26803 160
rect -27125 -161 -26803 -160
rect -27548 -508 -27444 -212
rect -28137 -560 -27815 -559
rect -28137 -880 -28136 -560
rect -27816 -880 -27815 -560
rect -28137 -881 -27815 -880
rect -28560 -1228 -28456 -932
rect -29149 -1280 -28827 -1279
rect -29149 -1600 -29148 -1280
rect -28828 -1600 -28827 -1280
rect -29149 -1601 -28827 -1600
rect -29572 -1948 -29468 -1652
rect -30161 -2000 -29839 -1999
rect -30161 -2320 -30160 -2000
rect -29840 -2320 -29839 -2000
rect -30161 -2321 -29839 -2320
rect -30584 -2520 -30480 -2372
rect -30052 -2520 -29948 -2321
rect -29572 -2372 -29552 -1948
rect -29488 -2372 -29468 -1948
rect -29040 -1999 -28936 -1601
rect -28560 -1652 -28540 -1228
rect -28476 -1652 -28456 -1228
rect -28028 -1279 -27924 -881
rect -27548 -932 -27528 -508
rect -27464 -932 -27444 -508
rect -27016 -559 -26912 -161
rect -26536 -212 -26516 212
rect -26452 -212 -26432 212
rect -26004 161 -25900 559
rect -25524 508 -25504 932
rect -25440 508 -25420 932
rect -24992 881 -24888 1279
rect -24512 1228 -24492 1652
rect -24428 1228 -24408 1652
rect -23980 1601 -23876 1999
rect -23500 1948 -23480 2372
rect -23416 1948 -23396 2372
rect -22968 2321 -22864 2520
rect -22488 2372 -22384 2520
rect -23077 2320 -22755 2321
rect -23077 2000 -23076 2320
rect -22756 2000 -22755 2320
rect -23077 1999 -22755 2000
rect -23500 1652 -23396 1948
rect -24089 1600 -23767 1601
rect -24089 1280 -24088 1600
rect -23768 1280 -23767 1600
rect -24089 1279 -23767 1280
rect -24512 932 -24408 1228
rect -25101 880 -24779 881
rect -25101 560 -25100 880
rect -24780 560 -24779 880
rect -25101 559 -24779 560
rect -25524 212 -25420 508
rect -26113 160 -25791 161
rect -26113 -160 -26112 160
rect -25792 -160 -25791 160
rect -26113 -161 -25791 -160
rect -26536 -508 -26432 -212
rect -27125 -560 -26803 -559
rect -27125 -880 -27124 -560
rect -26804 -880 -26803 -560
rect -27125 -881 -26803 -880
rect -27548 -1228 -27444 -932
rect -28137 -1280 -27815 -1279
rect -28137 -1600 -28136 -1280
rect -27816 -1600 -27815 -1280
rect -28137 -1601 -27815 -1600
rect -28560 -1948 -28456 -1652
rect -29149 -2000 -28827 -1999
rect -29149 -2320 -29148 -2000
rect -28828 -2320 -28827 -2000
rect -29149 -2321 -28827 -2320
rect -29572 -2520 -29468 -2372
rect -29040 -2520 -28936 -2321
rect -28560 -2372 -28540 -1948
rect -28476 -2372 -28456 -1948
rect -28028 -1999 -27924 -1601
rect -27548 -1652 -27528 -1228
rect -27464 -1652 -27444 -1228
rect -27016 -1279 -26912 -881
rect -26536 -932 -26516 -508
rect -26452 -932 -26432 -508
rect -26004 -559 -25900 -161
rect -25524 -212 -25504 212
rect -25440 -212 -25420 212
rect -24992 161 -24888 559
rect -24512 508 -24492 932
rect -24428 508 -24408 932
rect -23980 881 -23876 1279
rect -23500 1228 -23480 1652
rect -23416 1228 -23396 1652
rect -22968 1601 -22864 1999
rect -22488 1948 -22468 2372
rect -22404 1948 -22384 2372
rect -21956 2321 -21852 2520
rect -21476 2372 -21372 2520
rect -22065 2320 -21743 2321
rect -22065 2000 -22064 2320
rect -21744 2000 -21743 2320
rect -22065 1999 -21743 2000
rect -22488 1652 -22384 1948
rect -23077 1600 -22755 1601
rect -23077 1280 -23076 1600
rect -22756 1280 -22755 1600
rect -23077 1279 -22755 1280
rect -23500 932 -23396 1228
rect -24089 880 -23767 881
rect -24089 560 -24088 880
rect -23768 560 -23767 880
rect -24089 559 -23767 560
rect -24512 212 -24408 508
rect -25101 160 -24779 161
rect -25101 -160 -25100 160
rect -24780 -160 -24779 160
rect -25101 -161 -24779 -160
rect -25524 -508 -25420 -212
rect -26113 -560 -25791 -559
rect -26113 -880 -26112 -560
rect -25792 -880 -25791 -560
rect -26113 -881 -25791 -880
rect -26536 -1228 -26432 -932
rect -27125 -1280 -26803 -1279
rect -27125 -1600 -27124 -1280
rect -26804 -1600 -26803 -1280
rect -27125 -1601 -26803 -1600
rect -27548 -1948 -27444 -1652
rect -28137 -2000 -27815 -1999
rect -28137 -2320 -28136 -2000
rect -27816 -2320 -27815 -2000
rect -28137 -2321 -27815 -2320
rect -28560 -2520 -28456 -2372
rect -28028 -2520 -27924 -2321
rect -27548 -2372 -27528 -1948
rect -27464 -2372 -27444 -1948
rect -27016 -1999 -26912 -1601
rect -26536 -1652 -26516 -1228
rect -26452 -1652 -26432 -1228
rect -26004 -1279 -25900 -881
rect -25524 -932 -25504 -508
rect -25440 -932 -25420 -508
rect -24992 -559 -24888 -161
rect -24512 -212 -24492 212
rect -24428 -212 -24408 212
rect -23980 161 -23876 559
rect -23500 508 -23480 932
rect -23416 508 -23396 932
rect -22968 881 -22864 1279
rect -22488 1228 -22468 1652
rect -22404 1228 -22384 1652
rect -21956 1601 -21852 1999
rect -21476 1948 -21456 2372
rect -21392 1948 -21372 2372
rect -20944 2321 -20840 2520
rect -20464 2372 -20360 2520
rect -21053 2320 -20731 2321
rect -21053 2000 -21052 2320
rect -20732 2000 -20731 2320
rect -21053 1999 -20731 2000
rect -21476 1652 -21372 1948
rect -22065 1600 -21743 1601
rect -22065 1280 -22064 1600
rect -21744 1280 -21743 1600
rect -22065 1279 -21743 1280
rect -22488 932 -22384 1228
rect -23077 880 -22755 881
rect -23077 560 -23076 880
rect -22756 560 -22755 880
rect -23077 559 -22755 560
rect -23500 212 -23396 508
rect -24089 160 -23767 161
rect -24089 -160 -24088 160
rect -23768 -160 -23767 160
rect -24089 -161 -23767 -160
rect -24512 -508 -24408 -212
rect -25101 -560 -24779 -559
rect -25101 -880 -25100 -560
rect -24780 -880 -24779 -560
rect -25101 -881 -24779 -880
rect -25524 -1228 -25420 -932
rect -26113 -1280 -25791 -1279
rect -26113 -1600 -26112 -1280
rect -25792 -1600 -25791 -1280
rect -26113 -1601 -25791 -1600
rect -26536 -1948 -26432 -1652
rect -27125 -2000 -26803 -1999
rect -27125 -2320 -27124 -2000
rect -26804 -2320 -26803 -2000
rect -27125 -2321 -26803 -2320
rect -27548 -2520 -27444 -2372
rect -27016 -2520 -26912 -2321
rect -26536 -2372 -26516 -1948
rect -26452 -2372 -26432 -1948
rect -26004 -1999 -25900 -1601
rect -25524 -1652 -25504 -1228
rect -25440 -1652 -25420 -1228
rect -24992 -1279 -24888 -881
rect -24512 -932 -24492 -508
rect -24428 -932 -24408 -508
rect -23980 -559 -23876 -161
rect -23500 -212 -23480 212
rect -23416 -212 -23396 212
rect -22968 161 -22864 559
rect -22488 508 -22468 932
rect -22404 508 -22384 932
rect -21956 881 -21852 1279
rect -21476 1228 -21456 1652
rect -21392 1228 -21372 1652
rect -20944 1601 -20840 1999
rect -20464 1948 -20444 2372
rect -20380 1948 -20360 2372
rect -19932 2321 -19828 2520
rect -19452 2372 -19348 2520
rect -20041 2320 -19719 2321
rect -20041 2000 -20040 2320
rect -19720 2000 -19719 2320
rect -20041 1999 -19719 2000
rect -20464 1652 -20360 1948
rect -21053 1600 -20731 1601
rect -21053 1280 -21052 1600
rect -20732 1280 -20731 1600
rect -21053 1279 -20731 1280
rect -21476 932 -21372 1228
rect -22065 880 -21743 881
rect -22065 560 -22064 880
rect -21744 560 -21743 880
rect -22065 559 -21743 560
rect -22488 212 -22384 508
rect -23077 160 -22755 161
rect -23077 -160 -23076 160
rect -22756 -160 -22755 160
rect -23077 -161 -22755 -160
rect -23500 -508 -23396 -212
rect -24089 -560 -23767 -559
rect -24089 -880 -24088 -560
rect -23768 -880 -23767 -560
rect -24089 -881 -23767 -880
rect -24512 -1228 -24408 -932
rect -25101 -1280 -24779 -1279
rect -25101 -1600 -25100 -1280
rect -24780 -1600 -24779 -1280
rect -25101 -1601 -24779 -1600
rect -25524 -1948 -25420 -1652
rect -26113 -2000 -25791 -1999
rect -26113 -2320 -26112 -2000
rect -25792 -2320 -25791 -2000
rect -26113 -2321 -25791 -2320
rect -26536 -2520 -26432 -2372
rect -26004 -2520 -25900 -2321
rect -25524 -2372 -25504 -1948
rect -25440 -2372 -25420 -1948
rect -24992 -1999 -24888 -1601
rect -24512 -1652 -24492 -1228
rect -24428 -1652 -24408 -1228
rect -23980 -1279 -23876 -881
rect -23500 -932 -23480 -508
rect -23416 -932 -23396 -508
rect -22968 -559 -22864 -161
rect -22488 -212 -22468 212
rect -22404 -212 -22384 212
rect -21956 161 -21852 559
rect -21476 508 -21456 932
rect -21392 508 -21372 932
rect -20944 881 -20840 1279
rect -20464 1228 -20444 1652
rect -20380 1228 -20360 1652
rect -19932 1601 -19828 1999
rect -19452 1948 -19432 2372
rect -19368 1948 -19348 2372
rect -18920 2321 -18816 2520
rect -18440 2372 -18336 2520
rect -19029 2320 -18707 2321
rect -19029 2000 -19028 2320
rect -18708 2000 -18707 2320
rect -19029 1999 -18707 2000
rect -19452 1652 -19348 1948
rect -20041 1600 -19719 1601
rect -20041 1280 -20040 1600
rect -19720 1280 -19719 1600
rect -20041 1279 -19719 1280
rect -20464 932 -20360 1228
rect -21053 880 -20731 881
rect -21053 560 -21052 880
rect -20732 560 -20731 880
rect -21053 559 -20731 560
rect -21476 212 -21372 508
rect -22065 160 -21743 161
rect -22065 -160 -22064 160
rect -21744 -160 -21743 160
rect -22065 -161 -21743 -160
rect -22488 -508 -22384 -212
rect -23077 -560 -22755 -559
rect -23077 -880 -23076 -560
rect -22756 -880 -22755 -560
rect -23077 -881 -22755 -880
rect -23500 -1228 -23396 -932
rect -24089 -1280 -23767 -1279
rect -24089 -1600 -24088 -1280
rect -23768 -1600 -23767 -1280
rect -24089 -1601 -23767 -1600
rect -24512 -1948 -24408 -1652
rect -25101 -2000 -24779 -1999
rect -25101 -2320 -25100 -2000
rect -24780 -2320 -24779 -2000
rect -25101 -2321 -24779 -2320
rect -25524 -2520 -25420 -2372
rect -24992 -2520 -24888 -2321
rect -24512 -2372 -24492 -1948
rect -24428 -2372 -24408 -1948
rect -23980 -1999 -23876 -1601
rect -23500 -1652 -23480 -1228
rect -23416 -1652 -23396 -1228
rect -22968 -1279 -22864 -881
rect -22488 -932 -22468 -508
rect -22404 -932 -22384 -508
rect -21956 -559 -21852 -161
rect -21476 -212 -21456 212
rect -21392 -212 -21372 212
rect -20944 161 -20840 559
rect -20464 508 -20444 932
rect -20380 508 -20360 932
rect -19932 881 -19828 1279
rect -19452 1228 -19432 1652
rect -19368 1228 -19348 1652
rect -18920 1601 -18816 1999
rect -18440 1948 -18420 2372
rect -18356 1948 -18336 2372
rect -17908 2321 -17804 2520
rect -17428 2372 -17324 2520
rect -18017 2320 -17695 2321
rect -18017 2000 -18016 2320
rect -17696 2000 -17695 2320
rect -18017 1999 -17695 2000
rect -18440 1652 -18336 1948
rect -19029 1600 -18707 1601
rect -19029 1280 -19028 1600
rect -18708 1280 -18707 1600
rect -19029 1279 -18707 1280
rect -19452 932 -19348 1228
rect -20041 880 -19719 881
rect -20041 560 -20040 880
rect -19720 560 -19719 880
rect -20041 559 -19719 560
rect -20464 212 -20360 508
rect -21053 160 -20731 161
rect -21053 -160 -21052 160
rect -20732 -160 -20731 160
rect -21053 -161 -20731 -160
rect -21476 -508 -21372 -212
rect -22065 -560 -21743 -559
rect -22065 -880 -22064 -560
rect -21744 -880 -21743 -560
rect -22065 -881 -21743 -880
rect -22488 -1228 -22384 -932
rect -23077 -1280 -22755 -1279
rect -23077 -1600 -23076 -1280
rect -22756 -1600 -22755 -1280
rect -23077 -1601 -22755 -1600
rect -23500 -1948 -23396 -1652
rect -24089 -2000 -23767 -1999
rect -24089 -2320 -24088 -2000
rect -23768 -2320 -23767 -2000
rect -24089 -2321 -23767 -2320
rect -24512 -2520 -24408 -2372
rect -23980 -2520 -23876 -2321
rect -23500 -2372 -23480 -1948
rect -23416 -2372 -23396 -1948
rect -22968 -1999 -22864 -1601
rect -22488 -1652 -22468 -1228
rect -22404 -1652 -22384 -1228
rect -21956 -1279 -21852 -881
rect -21476 -932 -21456 -508
rect -21392 -932 -21372 -508
rect -20944 -559 -20840 -161
rect -20464 -212 -20444 212
rect -20380 -212 -20360 212
rect -19932 161 -19828 559
rect -19452 508 -19432 932
rect -19368 508 -19348 932
rect -18920 881 -18816 1279
rect -18440 1228 -18420 1652
rect -18356 1228 -18336 1652
rect -17908 1601 -17804 1999
rect -17428 1948 -17408 2372
rect -17344 1948 -17324 2372
rect -16896 2321 -16792 2520
rect -16416 2372 -16312 2520
rect -17005 2320 -16683 2321
rect -17005 2000 -17004 2320
rect -16684 2000 -16683 2320
rect -17005 1999 -16683 2000
rect -17428 1652 -17324 1948
rect -18017 1600 -17695 1601
rect -18017 1280 -18016 1600
rect -17696 1280 -17695 1600
rect -18017 1279 -17695 1280
rect -18440 932 -18336 1228
rect -19029 880 -18707 881
rect -19029 560 -19028 880
rect -18708 560 -18707 880
rect -19029 559 -18707 560
rect -19452 212 -19348 508
rect -20041 160 -19719 161
rect -20041 -160 -20040 160
rect -19720 -160 -19719 160
rect -20041 -161 -19719 -160
rect -20464 -508 -20360 -212
rect -21053 -560 -20731 -559
rect -21053 -880 -21052 -560
rect -20732 -880 -20731 -560
rect -21053 -881 -20731 -880
rect -21476 -1228 -21372 -932
rect -22065 -1280 -21743 -1279
rect -22065 -1600 -22064 -1280
rect -21744 -1600 -21743 -1280
rect -22065 -1601 -21743 -1600
rect -22488 -1948 -22384 -1652
rect -23077 -2000 -22755 -1999
rect -23077 -2320 -23076 -2000
rect -22756 -2320 -22755 -2000
rect -23077 -2321 -22755 -2320
rect -23500 -2520 -23396 -2372
rect -22968 -2520 -22864 -2321
rect -22488 -2372 -22468 -1948
rect -22404 -2372 -22384 -1948
rect -21956 -1999 -21852 -1601
rect -21476 -1652 -21456 -1228
rect -21392 -1652 -21372 -1228
rect -20944 -1279 -20840 -881
rect -20464 -932 -20444 -508
rect -20380 -932 -20360 -508
rect -19932 -559 -19828 -161
rect -19452 -212 -19432 212
rect -19368 -212 -19348 212
rect -18920 161 -18816 559
rect -18440 508 -18420 932
rect -18356 508 -18336 932
rect -17908 881 -17804 1279
rect -17428 1228 -17408 1652
rect -17344 1228 -17324 1652
rect -16896 1601 -16792 1999
rect -16416 1948 -16396 2372
rect -16332 1948 -16312 2372
rect -15884 2321 -15780 2520
rect -15404 2372 -15300 2520
rect -15993 2320 -15671 2321
rect -15993 2000 -15992 2320
rect -15672 2000 -15671 2320
rect -15993 1999 -15671 2000
rect -16416 1652 -16312 1948
rect -17005 1600 -16683 1601
rect -17005 1280 -17004 1600
rect -16684 1280 -16683 1600
rect -17005 1279 -16683 1280
rect -17428 932 -17324 1228
rect -18017 880 -17695 881
rect -18017 560 -18016 880
rect -17696 560 -17695 880
rect -18017 559 -17695 560
rect -18440 212 -18336 508
rect -19029 160 -18707 161
rect -19029 -160 -19028 160
rect -18708 -160 -18707 160
rect -19029 -161 -18707 -160
rect -19452 -508 -19348 -212
rect -20041 -560 -19719 -559
rect -20041 -880 -20040 -560
rect -19720 -880 -19719 -560
rect -20041 -881 -19719 -880
rect -20464 -1228 -20360 -932
rect -21053 -1280 -20731 -1279
rect -21053 -1600 -21052 -1280
rect -20732 -1600 -20731 -1280
rect -21053 -1601 -20731 -1600
rect -21476 -1948 -21372 -1652
rect -22065 -2000 -21743 -1999
rect -22065 -2320 -22064 -2000
rect -21744 -2320 -21743 -2000
rect -22065 -2321 -21743 -2320
rect -22488 -2520 -22384 -2372
rect -21956 -2520 -21852 -2321
rect -21476 -2372 -21456 -1948
rect -21392 -2372 -21372 -1948
rect -20944 -1999 -20840 -1601
rect -20464 -1652 -20444 -1228
rect -20380 -1652 -20360 -1228
rect -19932 -1279 -19828 -881
rect -19452 -932 -19432 -508
rect -19368 -932 -19348 -508
rect -18920 -559 -18816 -161
rect -18440 -212 -18420 212
rect -18356 -212 -18336 212
rect -17908 161 -17804 559
rect -17428 508 -17408 932
rect -17344 508 -17324 932
rect -16896 881 -16792 1279
rect -16416 1228 -16396 1652
rect -16332 1228 -16312 1652
rect -15884 1601 -15780 1999
rect -15404 1948 -15384 2372
rect -15320 1948 -15300 2372
rect -14872 2321 -14768 2520
rect -14392 2372 -14288 2520
rect -14981 2320 -14659 2321
rect -14981 2000 -14980 2320
rect -14660 2000 -14659 2320
rect -14981 1999 -14659 2000
rect -15404 1652 -15300 1948
rect -15993 1600 -15671 1601
rect -15993 1280 -15992 1600
rect -15672 1280 -15671 1600
rect -15993 1279 -15671 1280
rect -16416 932 -16312 1228
rect -17005 880 -16683 881
rect -17005 560 -17004 880
rect -16684 560 -16683 880
rect -17005 559 -16683 560
rect -17428 212 -17324 508
rect -18017 160 -17695 161
rect -18017 -160 -18016 160
rect -17696 -160 -17695 160
rect -18017 -161 -17695 -160
rect -18440 -508 -18336 -212
rect -19029 -560 -18707 -559
rect -19029 -880 -19028 -560
rect -18708 -880 -18707 -560
rect -19029 -881 -18707 -880
rect -19452 -1228 -19348 -932
rect -20041 -1280 -19719 -1279
rect -20041 -1600 -20040 -1280
rect -19720 -1600 -19719 -1280
rect -20041 -1601 -19719 -1600
rect -20464 -1948 -20360 -1652
rect -21053 -2000 -20731 -1999
rect -21053 -2320 -21052 -2000
rect -20732 -2320 -20731 -2000
rect -21053 -2321 -20731 -2320
rect -21476 -2520 -21372 -2372
rect -20944 -2520 -20840 -2321
rect -20464 -2372 -20444 -1948
rect -20380 -2372 -20360 -1948
rect -19932 -1999 -19828 -1601
rect -19452 -1652 -19432 -1228
rect -19368 -1652 -19348 -1228
rect -18920 -1279 -18816 -881
rect -18440 -932 -18420 -508
rect -18356 -932 -18336 -508
rect -17908 -559 -17804 -161
rect -17428 -212 -17408 212
rect -17344 -212 -17324 212
rect -16896 161 -16792 559
rect -16416 508 -16396 932
rect -16332 508 -16312 932
rect -15884 881 -15780 1279
rect -15404 1228 -15384 1652
rect -15320 1228 -15300 1652
rect -14872 1601 -14768 1999
rect -14392 1948 -14372 2372
rect -14308 1948 -14288 2372
rect -13860 2321 -13756 2520
rect -13380 2372 -13276 2520
rect -13969 2320 -13647 2321
rect -13969 2000 -13968 2320
rect -13648 2000 -13647 2320
rect -13969 1999 -13647 2000
rect -14392 1652 -14288 1948
rect -14981 1600 -14659 1601
rect -14981 1280 -14980 1600
rect -14660 1280 -14659 1600
rect -14981 1279 -14659 1280
rect -15404 932 -15300 1228
rect -15993 880 -15671 881
rect -15993 560 -15992 880
rect -15672 560 -15671 880
rect -15993 559 -15671 560
rect -16416 212 -16312 508
rect -17005 160 -16683 161
rect -17005 -160 -17004 160
rect -16684 -160 -16683 160
rect -17005 -161 -16683 -160
rect -17428 -508 -17324 -212
rect -18017 -560 -17695 -559
rect -18017 -880 -18016 -560
rect -17696 -880 -17695 -560
rect -18017 -881 -17695 -880
rect -18440 -1228 -18336 -932
rect -19029 -1280 -18707 -1279
rect -19029 -1600 -19028 -1280
rect -18708 -1600 -18707 -1280
rect -19029 -1601 -18707 -1600
rect -19452 -1948 -19348 -1652
rect -20041 -2000 -19719 -1999
rect -20041 -2320 -20040 -2000
rect -19720 -2320 -19719 -2000
rect -20041 -2321 -19719 -2320
rect -20464 -2520 -20360 -2372
rect -19932 -2520 -19828 -2321
rect -19452 -2372 -19432 -1948
rect -19368 -2372 -19348 -1948
rect -18920 -1999 -18816 -1601
rect -18440 -1652 -18420 -1228
rect -18356 -1652 -18336 -1228
rect -17908 -1279 -17804 -881
rect -17428 -932 -17408 -508
rect -17344 -932 -17324 -508
rect -16896 -559 -16792 -161
rect -16416 -212 -16396 212
rect -16332 -212 -16312 212
rect -15884 161 -15780 559
rect -15404 508 -15384 932
rect -15320 508 -15300 932
rect -14872 881 -14768 1279
rect -14392 1228 -14372 1652
rect -14308 1228 -14288 1652
rect -13860 1601 -13756 1999
rect -13380 1948 -13360 2372
rect -13296 1948 -13276 2372
rect -12848 2321 -12744 2520
rect -12368 2372 -12264 2520
rect -12957 2320 -12635 2321
rect -12957 2000 -12956 2320
rect -12636 2000 -12635 2320
rect -12957 1999 -12635 2000
rect -13380 1652 -13276 1948
rect -13969 1600 -13647 1601
rect -13969 1280 -13968 1600
rect -13648 1280 -13647 1600
rect -13969 1279 -13647 1280
rect -14392 932 -14288 1228
rect -14981 880 -14659 881
rect -14981 560 -14980 880
rect -14660 560 -14659 880
rect -14981 559 -14659 560
rect -15404 212 -15300 508
rect -15993 160 -15671 161
rect -15993 -160 -15992 160
rect -15672 -160 -15671 160
rect -15993 -161 -15671 -160
rect -16416 -508 -16312 -212
rect -17005 -560 -16683 -559
rect -17005 -880 -17004 -560
rect -16684 -880 -16683 -560
rect -17005 -881 -16683 -880
rect -17428 -1228 -17324 -932
rect -18017 -1280 -17695 -1279
rect -18017 -1600 -18016 -1280
rect -17696 -1600 -17695 -1280
rect -18017 -1601 -17695 -1600
rect -18440 -1948 -18336 -1652
rect -19029 -2000 -18707 -1999
rect -19029 -2320 -19028 -2000
rect -18708 -2320 -18707 -2000
rect -19029 -2321 -18707 -2320
rect -19452 -2520 -19348 -2372
rect -18920 -2520 -18816 -2321
rect -18440 -2372 -18420 -1948
rect -18356 -2372 -18336 -1948
rect -17908 -1999 -17804 -1601
rect -17428 -1652 -17408 -1228
rect -17344 -1652 -17324 -1228
rect -16896 -1279 -16792 -881
rect -16416 -932 -16396 -508
rect -16332 -932 -16312 -508
rect -15884 -559 -15780 -161
rect -15404 -212 -15384 212
rect -15320 -212 -15300 212
rect -14872 161 -14768 559
rect -14392 508 -14372 932
rect -14308 508 -14288 932
rect -13860 881 -13756 1279
rect -13380 1228 -13360 1652
rect -13296 1228 -13276 1652
rect -12848 1601 -12744 1999
rect -12368 1948 -12348 2372
rect -12284 1948 -12264 2372
rect -11836 2321 -11732 2520
rect -11356 2372 -11252 2520
rect -11945 2320 -11623 2321
rect -11945 2000 -11944 2320
rect -11624 2000 -11623 2320
rect -11945 1999 -11623 2000
rect -12368 1652 -12264 1948
rect -12957 1600 -12635 1601
rect -12957 1280 -12956 1600
rect -12636 1280 -12635 1600
rect -12957 1279 -12635 1280
rect -13380 932 -13276 1228
rect -13969 880 -13647 881
rect -13969 560 -13968 880
rect -13648 560 -13647 880
rect -13969 559 -13647 560
rect -14392 212 -14288 508
rect -14981 160 -14659 161
rect -14981 -160 -14980 160
rect -14660 -160 -14659 160
rect -14981 -161 -14659 -160
rect -15404 -508 -15300 -212
rect -15993 -560 -15671 -559
rect -15993 -880 -15992 -560
rect -15672 -880 -15671 -560
rect -15993 -881 -15671 -880
rect -16416 -1228 -16312 -932
rect -17005 -1280 -16683 -1279
rect -17005 -1600 -17004 -1280
rect -16684 -1600 -16683 -1280
rect -17005 -1601 -16683 -1600
rect -17428 -1948 -17324 -1652
rect -18017 -2000 -17695 -1999
rect -18017 -2320 -18016 -2000
rect -17696 -2320 -17695 -2000
rect -18017 -2321 -17695 -2320
rect -18440 -2520 -18336 -2372
rect -17908 -2520 -17804 -2321
rect -17428 -2372 -17408 -1948
rect -17344 -2372 -17324 -1948
rect -16896 -1999 -16792 -1601
rect -16416 -1652 -16396 -1228
rect -16332 -1652 -16312 -1228
rect -15884 -1279 -15780 -881
rect -15404 -932 -15384 -508
rect -15320 -932 -15300 -508
rect -14872 -559 -14768 -161
rect -14392 -212 -14372 212
rect -14308 -212 -14288 212
rect -13860 161 -13756 559
rect -13380 508 -13360 932
rect -13296 508 -13276 932
rect -12848 881 -12744 1279
rect -12368 1228 -12348 1652
rect -12284 1228 -12264 1652
rect -11836 1601 -11732 1999
rect -11356 1948 -11336 2372
rect -11272 1948 -11252 2372
rect -10824 2321 -10720 2520
rect -10344 2372 -10240 2520
rect -10933 2320 -10611 2321
rect -10933 2000 -10932 2320
rect -10612 2000 -10611 2320
rect -10933 1999 -10611 2000
rect -11356 1652 -11252 1948
rect -11945 1600 -11623 1601
rect -11945 1280 -11944 1600
rect -11624 1280 -11623 1600
rect -11945 1279 -11623 1280
rect -12368 932 -12264 1228
rect -12957 880 -12635 881
rect -12957 560 -12956 880
rect -12636 560 -12635 880
rect -12957 559 -12635 560
rect -13380 212 -13276 508
rect -13969 160 -13647 161
rect -13969 -160 -13968 160
rect -13648 -160 -13647 160
rect -13969 -161 -13647 -160
rect -14392 -508 -14288 -212
rect -14981 -560 -14659 -559
rect -14981 -880 -14980 -560
rect -14660 -880 -14659 -560
rect -14981 -881 -14659 -880
rect -15404 -1228 -15300 -932
rect -15993 -1280 -15671 -1279
rect -15993 -1600 -15992 -1280
rect -15672 -1600 -15671 -1280
rect -15993 -1601 -15671 -1600
rect -16416 -1948 -16312 -1652
rect -17005 -2000 -16683 -1999
rect -17005 -2320 -17004 -2000
rect -16684 -2320 -16683 -2000
rect -17005 -2321 -16683 -2320
rect -17428 -2520 -17324 -2372
rect -16896 -2520 -16792 -2321
rect -16416 -2372 -16396 -1948
rect -16332 -2372 -16312 -1948
rect -15884 -1999 -15780 -1601
rect -15404 -1652 -15384 -1228
rect -15320 -1652 -15300 -1228
rect -14872 -1279 -14768 -881
rect -14392 -932 -14372 -508
rect -14308 -932 -14288 -508
rect -13860 -559 -13756 -161
rect -13380 -212 -13360 212
rect -13296 -212 -13276 212
rect -12848 161 -12744 559
rect -12368 508 -12348 932
rect -12284 508 -12264 932
rect -11836 881 -11732 1279
rect -11356 1228 -11336 1652
rect -11272 1228 -11252 1652
rect -10824 1601 -10720 1999
rect -10344 1948 -10324 2372
rect -10260 1948 -10240 2372
rect -9812 2321 -9708 2520
rect -9332 2372 -9228 2520
rect -9921 2320 -9599 2321
rect -9921 2000 -9920 2320
rect -9600 2000 -9599 2320
rect -9921 1999 -9599 2000
rect -10344 1652 -10240 1948
rect -10933 1600 -10611 1601
rect -10933 1280 -10932 1600
rect -10612 1280 -10611 1600
rect -10933 1279 -10611 1280
rect -11356 932 -11252 1228
rect -11945 880 -11623 881
rect -11945 560 -11944 880
rect -11624 560 -11623 880
rect -11945 559 -11623 560
rect -12368 212 -12264 508
rect -12957 160 -12635 161
rect -12957 -160 -12956 160
rect -12636 -160 -12635 160
rect -12957 -161 -12635 -160
rect -13380 -508 -13276 -212
rect -13969 -560 -13647 -559
rect -13969 -880 -13968 -560
rect -13648 -880 -13647 -560
rect -13969 -881 -13647 -880
rect -14392 -1228 -14288 -932
rect -14981 -1280 -14659 -1279
rect -14981 -1600 -14980 -1280
rect -14660 -1600 -14659 -1280
rect -14981 -1601 -14659 -1600
rect -15404 -1948 -15300 -1652
rect -15993 -2000 -15671 -1999
rect -15993 -2320 -15992 -2000
rect -15672 -2320 -15671 -2000
rect -15993 -2321 -15671 -2320
rect -16416 -2520 -16312 -2372
rect -15884 -2520 -15780 -2321
rect -15404 -2372 -15384 -1948
rect -15320 -2372 -15300 -1948
rect -14872 -1999 -14768 -1601
rect -14392 -1652 -14372 -1228
rect -14308 -1652 -14288 -1228
rect -13860 -1279 -13756 -881
rect -13380 -932 -13360 -508
rect -13296 -932 -13276 -508
rect -12848 -559 -12744 -161
rect -12368 -212 -12348 212
rect -12284 -212 -12264 212
rect -11836 161 -11732 559
rect -11356 508 -11336 932
rect -11272 508 -11252 932
rect -10824 881 -10720 1279
rect -10344 1228 -10324 1652
rect -10260 1228 -10240 1652
rect -9812 1601 -9708 1999
rect -9332 1948 -9312 2372
rect -9248 1948 -9228 2372
rect -8800 2321 -8696 2520
rect -8320 2372 -8216 2520
rect -8909 2320 -8587 2321
rect -8909 2000 -8908 2320
rect -8588 2000 -8587 2320
rect -8909 1999 -8587 2000
rect -9332 1652 -9228 1948
rect -9921 1600 -9599 1601
rect -9921 1280 -9920 1600
rect -9600 1280 -9599 1600
rect -9921 1279 -9599 1280
rect -10344 932 -10240 1228
rect -10933 880 -10611 881
rect -10933 560 -10932 880
rect -10612 560 -10611 880
rect -10933 559 -10611 560
rect -11356 212 -11252 508
rect -11945 160 -11623 161
rect -11945 -160 -11944 160
rect -11624 -160 -11623 160
rect -11945 -161 -11623 -160
rect -12368 -508 -12264 -212
rect -12957 -560 -12635 -559
rect -12957 -880 -12956 -560
rect -12636 -880 -12635 -560
rect -12957 -881 -12635 -880
rect -13380 -1228 -13276 -932
rect -13969 -1280 -13647 -1279
rect -13969 -1600 -13968 -1280
rect -13648 -1600 -13647 -1280
rect -13969 -1601 -13647 -1600
rect -14392 -1948 -14288 -1652
rect -14981 -2000 -14659 -1999
rect -14981 -2320 -14980 -2000
rect -14660 -2320 -14659 -2000
rect -14981 -2321 -14659 -2320
rect -15404 -2520 -15300 -2372
rect -14872 -2520 -14768 -2321
rect -14392 -2372 -14372 -1948
rect -14308 -2372 -14288 -1948
rect -13860 -1999 -13756 -1601
rect -13380 -1652 -13360 -1228
rect -13296 -1652 -13276 -1228
rect -12848 -1279 -12744 -881
rect -12368 -932 -12348 -508
rect -12284 -932 -12264 -508
rect -11836 -559 -11732 -161
rect -11356 -212 -11336 212
rect -11272 -212 -11252 212
rect -10824 161 -10720 559
rect -10344 508 -10324 932
rect -10260 508 -10240 932
rect -9812 881 -9708 1279
rect -9332 1228 -9312 1652
rect -9248 1228 -9228 1652
rect -8800 1601 -8696 1999
rect -8320 1948 -8300 2372
rect -8236 1948 -8216 2372
rect -7788 2321 -7684 2520
rect -7308 2372 -7204 2520
rect -7897 2320 -7575 2321
rect -7897 2000 -7896 2320
rect -7576 2000 -7575 2320
rect -7897 1999 -7575 2000
rect -8320 1652 -8216 1948
rect -8909 1600 -8587 1601
rect -8909 1280 -8908 1600
rect -8588 1280 -8587 1600
rect -8909 1279 -8587 1280
rect -9332 932 -9228 1228
rect -9921 880 -9599 881
rect -9921 560 -9920 880
rect -9600 560 -9599 880
rect -9921 559 -9599 560
rect -10344 212 -10240 508
rect -10933 160 -10611 161
rect -10933 -160 -10932 160
rect -10612 -160 -10611 160
rect -10933 -161 -10611 -160
rect -11356 -508 -11252 -212
rect -11945 -560 -11623 -559
rect -11945 -880 -11944 -560
rect -11624 -880 -11623 -560
rect -11945 -881 -11623 -880
rect -12368 -1228 -12264 -932
rect -12957 -1280 -12635 -1279
rect -12957 -1600 -12956 -1280
rect -12636 -1600 -12635 -1280
rect -12957 -1601 -12635 -1600
rect -13380 -1948 -13276 -1652
rect -13969 -2000 -13647 -1999
rect -13969 -2320 -13968 -2000
rect -13648 -2320 -13647 -2000
rect -13969 -2321 -13647 -2320
rect -14392 -2520 -14288 -2372
rect -13860 -2520 -13756 -2321
rect -13380 -2372 -13360 -1948
rect -13296 -2372 -13276 -1948
rect -12848 -1999 -12744 -1601
rect -12368 -1652 -12348 -1228
rect -12284 -1652 -12264 -1228
rect -11836 -1279 -11732 -881
rect -11356 -932 -11336 -508
rect -11272 -932 -11252 -508
rect -10824 -559 -10720 -161
rect -10344 -212 -10324 212
rect -10260 -212 -10240 212
rect -9812 161 -9708 559
rect -9332 508 -9312 932
rect -9248 508 -9228 932
rect -8800 881 -8696 1279
rect -8320 1228 -8300 1652
rect -8236 1228 -8216 1652
rect -7788 1601 -7684 1999
rect -7308 1948 -7288 2372
rect -7224 1948 -7204 2372
rect -6776 2321 -6672 2520
rect -6296 2372 -6192 2520
rect -6885 2320 -6563 2321
rect -6885 2000 -6884 2320
rect -6564 2000 -6563 2320
rect -6885 1999 -6563 2000
rect -7308 1652 -7204 1948
rect -7897 1600 -7575 1601
rect -7897 1280 -7896 1600
rect -7576 1280 -7575 1600
rect -7897 1279 -7575 1280
rect -8320 932 -8216 1228
rect -8909 880 -8587 881
rect -8909 560 -8908 880
rect -8588 560 -8587 880
rect -8909 559 -8587 560
rect -9332 212 -9228 508
rect -9921 160 -9599 161
rect -9921 -160 -9920 160
rect -9600 -160 -9599 160
rect -9921 -161 -9599 -160
rect -10344 -508 -10240 -212
rect -10933 -560 -10611 -559
rect -10933 -880 -10932 -560
rect -10612 -880 -10611 -560
rect -10933 -881 -10611 -880
rect -11356 -1228 -11252 -932
rect -11945 -1280 -11623 -1279
rect -11945 -1600 -11944 -1280
rect -11624 -1600 -11623 -1280
rect -11945 -1601 -11623 -1600
rect -12368 -1948 -12264 -1652
rect -12957 -2000 -12635 -1999
rect -12957 -2320 -12956 -2000
rect -12636 -2320 -12635 -2000
rect -12957 -2321 -12635 -2320
rect -13380 -2520 -13276 -2372
rect -12848 -2520 -12744 -2321
rect -12368 -2372 -12348 -1948
rect -12284 -2372 -12264 -1948
rect -11836 -1999 -11732 -1601
rect -11356 -1652 -11336 -1228
rect -11272 -1652 -11252 -1228
rect -10824 -1279 -10720 -881
rect -10344 -932 -10324 -508
rect -10260 -932 -10240 -508
rect -9812 -559 -9708 -161
rect -9332 -212 -9312 212
rect -9248 -212 -9228 212
rect -8800 161 -8696 559
rect -8320 508 -8300 932
rect -8236 508 -8216 932
rect -7788 881 -7684 1279
rect -7308 1228 -7288 1652
rect -7224 1228 -7204 1652
rect -6776 1601 -6672 1999
rect -6296 1948 -6276 2372
rect -6212 1948 -6192 2372
rect -5764 2321 -5660 2520
rect -5284 2372 -5180 2520
rect -5873 2320 -5551 2321
rect -5873 2000 -5872 2320
rect -5552 2000 -5551 2320
rect -5873 1999 -5551 2000
rect -6296 1652 -6192 1948
rect -6885 1600 -6563 1601
rect -6885 1280 -6884 1600
rect -6564 1280 -6563 1600
rect -6885 1279 -6563 1280
rect -7308 932 -7204 1228
rect -7897 880 -7575 881
rect -7897 560 -7896 880
rect -7576 560 -7575 880
rect -7897 559 -7575 560
rect -8320 212 -8216 508
rect -8909 160 -8587 161
rect -8909 -160 -8908 160
rect -8588 -160 -8587 160
rect -8909 -161 -8587 -160
rect -9332 -508 -9228 -212
rect -9921 -560 -9599 -559
rect -9921 -880 -9920 -560
rect -9600 -880 -9599 -560
rect -9921 -881 -9599 -880
rect -10344 -1228 -10240 -932
rect -10933 -1280 -10611 -1279
rect -10933 -1600 -10932 -1280
rect -10612 -1600 -10611 -1280
rect -10933 -1601 -10611 -1600
rect -11356 -1948 -11252 -1652
rect -11945 -2000 -11623 -1999
rect -11945 -2320 -11944 -2000
rect -11624 -2320 -11623 -2000
rect -11945 -2321 -11623 -2320
rect -12368 -2520 -12264 -2372
rect -11836 -2520 -11732 -2321
rect -11356 -2372 -11336 -1948
rect -11272 -2372 -11252 -1948
rect -10824 -1999 -10720 -1601
rect -10344 -1652 -10324 -1228
rect -10260 -1652 -10240 -1228
rect -9812 -1279 -9708 -881
rect -9332 -932 -9312 -508
rect -9248 -932 -9228 -508
rect -8800 -559 -8696 -161
rect -8320 -212 -8300 212
rect -8236 -212 -8216 212
rect -7788 161 -7684 559
rect -7308 508 -7288 932
rect -7224 508 -7204 932
rect -6776 881 -6672 1279
rect -6296 1228 -6276 1652
rect -6212 1228 -6192 1652
rect -5764 1601 -5660 1999
rect -5284 1948 -5264 2372
rect -5200 1948 -5180 2372
rect -4752 2321 -4648 2520
rect -4272 2372 -4168 2520
rect -4861 2320 -4539 2321
rect -4861 2000 -4860 2320
rect -4540 2000 -4539 2320
rect -4861 1999 -4539 2000
rect -5284 1652 -5180 1948
rect -5873 1600 -5551 1601
rect -5873 1280 -5872 1600
rect -5552 1280 -5551 1600
rect -5873 1279 -5551 1280
rect -6296 932 -6192 1228
rect -6885 880 -6563 881
rect -6885 560 -6884 880
rect -6564 560 -6563 880
rect -6885 559 -6563 560
rect -7308 212 -7204 508
rect -7897 160 -7575 161
rect -7897 -160 -7896 160
rect -7576 -160 -7575 160
rect -7897 -161 -7575 -160
rect -8320 -508 -8216 -212
rect -8909 -560 -8587 -559
rect -8909 -880 -8908 -560
rect -8588 -880 -8587 -560
rect -8909 -881 -8587 -880
rect -9332 -1228 -9228 -932
rect -9921 -1280 -9599 -1279
rect -9921 -1600 -9920 -1280
rect -9600 -1600 -9599 -1280
rect -9921 -1601 -9599 -1600
rect -10344 -1948 -10240 -1652
rect -10933 -2000 -10611 -1999
rect -10933 -2320 -10932 -2000
rect -10612 -2320 -10611 -2000
rect -10933 -2321 -10611 -2320
rect -11356 -2520 -11252 -2372
rect -10824 -2520 -10720 -2321
rect -10344 -2372 -10324 -1948
rect -10260 -2372 -10240 -1948
rect -9812 -1999 -9708 -1601
rect -9332 -1652 -9312 -1228
rect -9248 -1652 -9228 -1228
rect -8800 -1279 -8696 -881
rect -8320 -932 -8300 -508
rect -8236 -932 -8216 -508
rect -7788 -559 -7684 -161
rect -7308 -212 -7288 212
rect -7224 -212 -7204 212
rect -6776 161 -6672 559
rect -6296 508 -6276 932
rect -6212 508 -6192 932
rect -5764 881 -5660 1279
rect -5284 1228 -5264 1652
rect -5200 1228 -5180 1652
rect -4752 1601 -4648 1999
rect -4272 1948 -4252 2372
rect -4188 1948 -4168 2372
rect -3740 2321 -3636 2520
rect -3260 2372 -3156 2520
rect -3849 2320 -3527 2321
rect -3849 2000 -3848 2320
rect -3528 2000 -3527 2320
rect -3849 1999 -3527 2000
rect -4272 1652 -4168 1948
rect -4861 1600 -4539 1601
rect -4861 1280 -4860 1600
rect -4540 1280 -4539 1600
rect -4861 1279 -4539 1280
rect -5284 932 -5180 1228
rect -5873 880 -5551 881
rect -5873 560 -5872 880
rect -5552 560 -5551 880
rect -5873 559 -5551 560
rect -6296 212 -6192 508
rect -6885 160 -6563 161
rect -6885 -160 -6884 160
rect -6564 -160 -6563 160
rect -6885 -161 -6563 -160
rect -7308 -508 -7204 -212
rect -7897 -560 -7575 -559
rect -7897 -880 -7896 -560
rect -7576 -880 -7575 -560
rect -7897 -881 -7575 -880
rect -8320 -1228 -8216 -932
rect -8909 -1280 -8587 -1279
rect -8909 -1600 -8908 -1280
rect -8588 -1600 -8587 -1280
rect -8909 -1601 -8587 -1600
rect -9332 -1948 -9228 -1652
rect -9921 -2000 -9599 -1999
rect -9921 -2320 -9920 -2000
rect -9600 -2320 -9599 -2000
rect -9921 -2321 -9599 -2320
rect -10344 -2520 -10240 -2372
rect -9812 -2520 -9708 -2321
rect -9332 -2372 -9312 -1948
rect -9248 -2372 -9228 -1948
rect -8800 -1999 -8696 -1601
rect -8320 -1652 -8300 -1228
rect -8236 -1652 -8216 -1228
rect -7788 -1279 -7684 -881
rect -7308 -932 -7288 -508
rect -7224 -932 -7204 -508
rect -6776 -559 -6672 -161
rect -6296 -212 -6276 212
rect -6212 -212 -6192 212
rect -5764 161 -5660 559
rect -5284 508 -5264 932
rect -5200 508 -5180 932
rect -4752 881 -4648 1279
rect -4272 1228 -4252 1652
rect -4188 1228 -4168 1652
rect -3740 1601 -3636 1999
rect -3260 1948 -3240 2372
rect -3176 1948 -3156 2372
rect -2728 2321 -2624 2520
rect -2248 2372 -2144 2520
rect -2837 2320 -2515 2321
rect -2837 2000 -2836 2320
rect -2516 2000 -2515 2320
rect -2837 1999 -2515 2000
rect -3260 1652 -3156 1948
rect -3849 1600 -3527 1601
rect -3849 1280 -3848 1600
rect -3528 1280 -3527 1600
rect -3849 1279 -3527 1280
rect -4272 932 -4168 1228
rect -4861 880 -4539 881
rect -4861 560 -4860 880
rect -4540 560 -4539 880
rect -4861 559 -4539 560
rect -5284 212 -5180 508
rect -5873 160 -5551 161
rect -5873 -160 -5872 160
rect -5552 -160 -5551 160
rect -5873 -161 -5551 -160
rect -6296 -508 -6192 -212
rect -6885 -560 -6563 -559
rect -6885 -880 -6884 -560
rect -6564 -880 -6563 -560
rect -6885 -881 -6563 -880
rect -7308 -1228 -7204 -932
rect -7897 -1280 -7575 -1279
rect -7897 -1600 -7896 -1280
rect -7576 -1600 -7575 -1280
rect -7897 -1601 -7575 -1600
rect -8320 -1948 -8216 -1652
rect -8909 -2000 -8587 -1999
rect -8909 -2320 -8908 -2000
rect -8588 -2320 -8587 -2000
rect -8909 -2321 -8587 -2320
rect -9332 -2520 -9228 -2372
rect -8800 -2520 -8696 -2321
rect -8320 -2372 -8300 -1948
rect -8236 -2372 -8216 -1948
rect -7788 -1999 -7684 -1601
rect -7308 -1652 -7288 -1228
rect -7224 -1652 -7204 -1228
rect -6776 -1279 -6672 -881
rect -6296 -932 -6276 -508
rect -6212 -932 -6192 -508
rect -5764 -559 -5660 -161
rect -5284 -212 -5264 212
rect -5200 -212 -5180 212
rect -4752 161 -4648 559
rect -4272 508 -4252 932
rect -4188 508 -4168 932
rect -3740 881 -3636 1279
rect -3260 1228 -3240 1652
rect -3176 1228 -3156 1652
rect -2728 1601 -2624 1999
rect -2248 1948 -2228 2372
rect -2164 1948 -2144 2372
rect -1716 2321 -1612 2520
rect -1236 2372 -1132 2520
rect -1825 2320 -1503 2321
rect -1825 2000 -1824 2320
rect -1504 2000 -1503 2320
rect -1825 1999 -1503 2000
rect -2248 1652 -2144 1948
rect -2837 1600 -2515 1601
rect -2837 1280 -2836 1600
rect -2516 1280 -2515 1600
rect -2837 1279 -2515 1280
rect -3260 932 -3156 1228
rect -3849 880 -3527 881
rect -3849 560 -3848 880
rect -3528 560 -3527 880
rect -3849 559 -3527 560
rect -4272 212 -4168 508
rect -4861 160 -4539 161
rect -4861 -160 -4860 160
rect -4540 -160 -4539 160
rect -4861 -161 -4539 -160
rect -5284 -508 -5180 -212
rect -5873 -560 -5551 -559
rect -5873 -880 -5872 -560
rect -5552 -880 -5551 -560
rect -5873 -881 -5551 -880
rect -6296 -1228 -6192 -932
rect -6885 -1280 -6563 -1279
rect -6885 -1600 -6884 -1280
rect -6564 -1600 -6563 -1280
rect -6885 -1601 -6563 -1600
rect -7308 -1948 -7204 -1652
rect -7897 -2000 -7575 -1999
rect -7897 -2320 -7896 -2000
rect -7576 -2320 -7575 -2000
rect -7897 -2321 -7575 -2320
rect -8320 -2520 -8216 -2372
rect -7788 -2520 -7684 -2321
rect -7308 -2372 -7288 -1948
rect -7224 -2372 -7204 -1948
rect -6776 -1999 -6672 -1601
rect -6296 -1652 -6276 -1228
rect -6212 -1652 -6192 -1228
rect -5764 -1279 -5660 -881
rect -5284 -932 -5264 -508
rect -5200 -932 -5180 -508
rect -4752 -559 -4648 -161
rect -4272 -212 -4252 212
rect -4188 -212 -4168 212
rect -3740 161 -3636 559
rect -3260 508 -3240 932
rect -3176 508 -3156 932
rect -2728 881 -2624 1279
rect -2248 1228 -2228 1652
rect -2164 1228 -2144 1652
rect -1716 1601 -1612 1999
rect -1236 1948 -1216 2372
rect -1152 1948 -1132 2372
rect -704 2321 -600 2520
rect -224 2372 -120 2520
rect -813 2320 -491 2321
rect -813 2000 -812 2320
rect -492 2000 -491 2320
rect -813 1999 -491 2000
rect -1236 1652 -1132 1948
rect -1825 1600 -1503 1601
rect -1825 1280 -1824 1600
rect -1504 1280 -1503 1600
rect -1825 1279 -1503 1280
rect -2248 932 -2144 1228
rect -2837 880 -2515 881
rect -2837 560 -2836 880
rect -2516 560 -2515 880
rect -2837 559 -2515 560
rect -3260 212 -3156 508
rect -3849 160 -3527 161
rect -3849 -160 -3848 160
rect -3528 -160 -3527 160
rect -3849 -161 -3527 -160
rect -4272 -508 -4168 -212
rect -4861 -560 -4539 -559
rect -4861 -880 -4860 -560
rect -4540 -880 -4539 -560
rect -4861 -881 -4539 -880
rect -5284 -1228 -5180 -932
rect -5873 -1280 -5551 -1279
rect -5873 -1600 -5872 -1280
rect -5552 -1600 -5551 -1280
rect -5873 -1601 -5551 -1600
rect -6296 -1948 -6192 -1652
rect -6885 -2000 -6563 -1999
rect -6885 -2320 -6884 -2000
rect -6564 -2320 -6563 -2000
rect -6885 -2321 -6563 -2320
rect -7308 -2520 -7204 -2372
rect -6776 -2520 -6672 -2321
rect -6296 -2372 -6276 -1948
rect -6212 -2372 -6192 -1948
rect -5764 -1999 -5660 -1601
rect -5284 -1652 -5264 -1228
rect -5200 -1652 -5180 -1228
rect -4752 -1279 -4648 -881
rect -4272 -932 -4252 -508
rect -4188 -932 -4168 -508
rect -3740 -559 -3636 -161
rect -3260 -212 -3240 212
rect -3176 -212 -3156 212
rect -2728 161 -2624 559
rect -2248 508 -2228 932
rect -2164 508 -2144 932
rect -1716 881 -1612 1279
rect -1236 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -704 1601 -600 1999
rect -224 1948 -204 2372
rect -140 1948 -120 2372
rect 308 2321 412 2520
rect 788 2372 892 2520
rect 199 2320 521 2321
rect 199 2000 200 2320
rect 520 2000 521 2320
rect 199 1999 521 2000
rect -224 1652 -120 1948
rect -813 1600 -491 1601
rect -813 1280 -812 1600
rect -492 1280 -491 1600
rect -813 1279 -491 1280
rect -1236 932 -1132 1228
rect -1825 880 -1503 881
rect -1825 560 -1824 880
rect -1504 560 -1503 880
rect -1825 559 -1503 560
rect -2248 212 -2144 508
rect -2837 160 -2515 161
rect -2837 -160 -2836 160
rect -2516 -160 -2515 160
rect -2837 -161 -2515 -160
rect -3260 -508 -3156 -212
rect -3849 -560 -3527 -559
rect -3849 -880 -3848 -560
rect -3528 -880 -3527 -560
rect -3849 -881 -3527 -880
rect -4272 -1228 -4168 -932
rect -4861 -1280 -4539 -1279
rect -4861 -1600 -4860 -1280
rect -4540 -1600 -4539 -1280
rect -4861 -1601 -4539 -1600
rect -5284 -1948 -5180 -1652
rect -5873 -2000 -5551 -1999
rect -5873 -2320 -5872 -2000
rect -5552 -2320 -5551 -2000
rect -5873 -2321 -5551 -2320
rect -6296 -2520 -6192 -2372
rect -5764 -2520 -5660 -2321
rect -5284 -2372 -5264 -1948
rect -5200 -2372 -5180 -1948
rect -4752 -1999 -4648 -1601
rect -4272 -1652 -4252 -1228
rect -4188 -1652 -4168 -1228
rect -3740 -1279 -3636 -881
rect -3260 -932 -3240 -508
rect -3176 -932 -3156 -508
rect -2728 -559 -2624 -161
rect -2248 -212 -2228 212
rect -2164 -212 -2144 212
rect -1716 161 -1612 559
rect -1236 508 -1216 932
rect -1152 508 -1132 932
rect -704 881 -600 1279
rect -224 1228 -204 1652
rect -140 1228 -120 1652
rect 308 1601 412 1999
rect 788 1948 808 2372
rect 872 1948 892 2372
rect 1320 2321 1424 2520
rect 1800 2372 1904 2520
rect 1211 2320 1533 2321
rect 1211 2000 1212 2320
rect 1532 2000 1533 2320
rect 1211 1999 1533 2000
rect 788 1652 892 1948
rect 199 1600 521 1601
rect 199 1280 200 1600
rect 520 1280 521 1600
rect 199 1279 521 1280
rect -224 932 -120 1228
rect -813 880 -491 881
rect -813 560 -812 880
rect -492 560 -491 880
rect -813 559 -491 560
rect -1236 212 -1132 508
rect -1825 160 -1503 161
rect -1825 -160 -1824 160
rect -1504 -160 -1503 160
rect -1825 -161 -1503 -160
rect -2248 -508 -2144 -212
rect -2837 -560 -2515 -559
rect -2837 -880 -2836 -560
rect -2516 -880 -2515 -560
rect -2837 -881 -2515 -880
rect -3260 -1228 -3156 -932
rect -3849 -1280 -3527 -1279
rect -3849 -1600 -3848 -1280
rect -3528 -1600 -3527 -1280
rect -3849 -1601 -3527 -1600
rect -4272 -1948 -4168 -1652
rect -4861 -2000 -4539 -1999
rect -4861 -2320 -4860 -2000
rect -4540 -2320 -4539 -2000
rect -4861 -2321 -4539 -2320
rect -5284 -2520 -5180 -2372
rect -4752 -2520 -4648 -2321
rect -4272 -2372 -4252 -1948
rect -4188 -2372 -4168 -1948
rect -3740 -1999 -3636 -1601
rect -3260 -1652 -3240 -1228
rect -3176 -1652 -3156 -1228
rect -2728 -1279 -2624 -881
rect -2248 -932 -2228 -508
rect -2164 -932 -2144 -508
rect -1716 -559 -1612 -161
rect -1236 -212 -1216 212
rect -1152 -212 -1132 212
rect -704 161 -600 559
rect -224 508 -204 932
rect -140 508 -120 932
rect 308 881 412 1279
rect 788 1228 808 1652
rect 872 1228 892 1652
rect 1320 1601 1424 1999
rect 1800 1948 1820 2372
rect 1884 1948 1904 2372
rect 2332 2321 2436 2520
rect 2812 2372 2916 2520
rect 2223 2320 2545 2321
rect 2223 2000 2224 2320
rect 2544 2000 2545 2320
rect 2223 1999 2545 2000
rect 1800 1652 1904 1948
rect 1211 1600 1533 1601
rect 1211 1280 1212 1600
rect 1532 1280 1533 1600
rect 1211 1279 1533 1280
rect 788 932 892 1228
rect 199 880 521 881
rect 199 560 200 880
rect 520 560 521 880
rect 199 559 521 560
rect -224 212 -120 508
rect -813 160 -491 161
rect -813 -160 -812 160
rect -492 -160 -491 160
rect -813 -161 -491 -160
rect -1236 -508 -1132 -212
rect -1825 -560 -1503 -559
rect -1825 -880 -1824 -560
rect -1504 -880 -1503 -560
rect -1825 -881 -1503 -880
rect -2248 -1228 -2144 -932
rect -2837 -1280 -2515 -1279
rect -2837 -1600 -2836 -1280
rect -2516 -1600 -2515 -1280
rect -2837 -1601 -2515 -1600
rect -3260 -1948 -3156 -1652
rect -3849 -2000 -3527 -1999
rect -3849 -2320 -3848 -2000
rect -3528 -2320 -3527 -2000
rect -3849 -2321 -3527 -2320
rect -4272 -2520 -4168 -2372
rect -3740 -2520 -3636 -2321
rect -3260 -2372 -3240 -1948
rect -3176 -2372 -3156 -1948
rect -2728 -1999 -2624 -1601
rect -2248 -1652 -2228 -1228
rect -2164 -1652 -2144 -1228
rect -1716 -1279 -1612 -881
rect -1236 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -704 -559 -600 -161
rect -224 -212 -204 212
rect -140 -212 -120 212
rect 308 161 412 559
rect 788 508 808 932
rect 872 508 892 932
rect 1320 881 1424 1279
rect 1800 1228 1820 1652
rect 1884 1228 1904 1652
rect 2332 1601 2436 1999
rect 2812 1948 2832 2372
rect 2896 1948 2916 2372
rect 3344 2321 3448 2520
rect 3824 2372 3928 2520
rect 3235 2320 3557 2321
rect 3235 2000 3236 2320
rect 3556 2000 3557 2320
rect 3235 1999 3557 2000
rect 2812 1652 2916 1948
rect 2223 1600 2545 1601
rect 2223 1280 2224 1600
rect 2544 1280 2545 1600
rect 2223 1279 2545 1280
rect 1800 932 1904 1228
rect 1211 880 1533 881
rect 1211 560 1212 880
rect 1532 560 1533 880
rect 1211 559 1533 560
rect 788 212 892 508
rect 199 160 521 161
rect 199 -160 200 160
rect 520 -160 521 160
rect 199 -161 521 -160
rect -224 -508 -120 -212
rect -813 -560 -491 -559
rect -813 -880 -812 -560
rect -492 -880 -491 -560
rect -813 -881 -491 -880
rect -1236 -1228 -1132 -932
rect -1825 -1280 -1503 -1279
rect -1825 -1600 -1824 -1280
rect -1504 -1600 -1503 -1280
rect -1825 -1601 -1503 -1600
rect -2248 -1948 -2144 -1652
rect -2837 -2000 -2515 -1999
rect -2837 -2320 -2836 -2000
rect -2516 -2320 -2515 -2000
rect -2837 -2321 -2515 -2320
rect -3260 -2520 -3156 -2372
rect -2728 -2520 -2624 -2321
rect -2248 -2372 -2228 -1948
rect -2164 -2372 -2144 -1948
rect -1716 -1999 -1612 -1601
rect -1236 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -704 -1279 -600 -881
rect -224 -932 -204 -508
rect -140 -932 -120 -508
rect 308 -559 412 -161
rect 788 -212 808 212
rect 872 -212 892 212
rect 1320 161 1424 559
rect 1800 508 1820 932
rect 1884 508 1904 932
rect 2332 881 2436 1279
rect 2812 1228 2832 1652
rect 2896 1228 2916 1652
rect 3344 1601 3448 1999
rect 3824 1948 3844 2372
rect 3908 1948 3928 2372
rect 4356 2321 4460 2520
rect 4836 2372 4940 2520
rect 4247 2320 4569 2321
rect 4247 2000 4248 2320
rect 4568 2000 4569 2320
rect 4247 1999 4569 2000
rect 3824 1652 3928 1948
rect 3235 1600 3557 1601
rect 3235 1280 3236 1600
rect 3556 1280 3557 1600
rect 3235 1279 3557 1280
rect 2812 932 2916 1228
rect 2223 880 2545 881
rect 2223 560 2224 880
rect 2544 560 2545 880
rect 2223 559 2545 560
rect 1800 212 1904 508
rect 1211 160 1533 161
rect 1211 -160 1212 160
rect 1532 -160 1533 160
rect 1211 -161 1533 -160
rect 788 -508 892 -212
rect 199 -560 521 -559
rect 199 -880 200 -560
rect 520 -880 521 -560
rect 199 -881 521 -880
rect -224 -1228 -120 -932
rect -813 -1280 -491 -1279
rect -813 -1600 -812 -1280
rect -492 -1600 -491 -1280
rect -813 -1601 -491 -1600
rect -1236 -1948 -1132 -1652
rect -1825 -2000 -1503 -1999
rect -1825 -2320 -1824 -2000
rect -1504 -2320 -1503 -2000
rect -1825 -2321 -1503 -2320
rect -2248 -2520 -2144 -2372
rect -1716 -2520 -1612 -2321
rect -1236 -2372 -1216 -1948
rect -1152 -2372 -1132 -1948
rect -704 -1999 -600 -1601
rect -224 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect 308 -1279 412 -881
rect 788 -932 808 -508
rect 872 -932 892 -508
rect 1320 -559 1424 -161
rect 1800 -212 1820 212
rect 1884 -212 1904 212
rect 2332 161 2436 559
rect 2812 508 2832 932
rect 2896 508 2916 932
rect 3344 881 3448 1279
rect 3824 1228 3844 1652
rect 3908 1228 3928 1652
rect 4356 1601 4460 1999
rect 4836 1948 4856 2372
rect 4920 1948 4940 2372
rect 5368 2321 5472 2520
rect 5848 2372 5952 2520
rect 5259 2320 5581 2321
rect 5259 2000 5260 2320
rect 5580 2000 5581 2320
rect 5259 1999 5581 2000
rect 4836 1652 4940 1948
rect 4247 1600 4569 1601
rect 4247 1280 4248 1600
rect 4568 1280 4569 1600
rect 4247 1279 4569 1280
rect 3824 932 3928 1228
rect 3235 880 3557 881
rect 3235 560 3236 880
rect 3556 560 3557 880
rect 3235 559 3557 560
rect 2812 212 2916 508
rect 2223 160 2545 161
rect 2223 -160 2224 160
rect 2544 -160 2545 160
rect 2223 -161 2545 -160
rect 1800 -508 1904 -212
rect 1211 -560 1533 -559
rect 1211 -880 1212 -560
rect 1532 -880 1533 -560
rect 1211 -881 1533 -880
rect 788 -1228 892 -932
rect 199 -1280 521 -1279
rect 199 -1600 200 -1280
rect 520 -1600 521 -1280
rect 199 -1601 521 -1600
rect -224 -1948 -120 -1652
rect -813 -2000 -491 -1999
rect -813 -2320 -812 -2000
rect -492 -2320 -491 -2000
rect -813 -2321 -491 -2320
rect -1236 -2520 -1132 -2372
rect -704 -2520 -600 -2321
rect -224 -2372 -204 -1948
rect -140 -2372 -120 -1948
rect 308 -1999 412 -1601
rect 788 -1652 808 -1228
rect 872 -1652 892 -1228
rect 1320 -1279 1424 -881
rect 1800 -932 1820 -508
rect 1884 -932 1904 -508
rect 2332 -559 2436 -161
rect 2812 -212 2832 212
rect 2896 -212 2916 212
rect 3344 161 3448 559
rect 3824 508 3844 932
rect 3908 508 3928 932
rect 4356 881 4460 1279
rect 4836 1228 4856 1652
rect 4920 1228 4940 1652
rect 5368 1601 5472 1999
rect 5848 1948 5868 2372
rect 5932 1948 5952 2372
rect 6380 2321 6484 2520
rect 6860 2372 6964 2520
rect 6271 2320 6593 2321
rect 6271 2000 6272 2320
rect 6592 2000 6593 2320
rect 6271 1999 6593 2000
rect 5848 1652 5952 1948
rect 5259 1600 5581 1601
rect 5259 1280 5260 1600
rect 5580 1280 5581 1600
rect 5259 1279 5581 1280
rect 4836 932 4940 1228
rect 4247 880 4569 881
rect 4247 560 4248 880
rect 4568 560 4569 880
rect 4247 559 4569 560
rect 3824 212 3928 508
rect 3235 160 3557 161
rect 3235 -160 3236 160
rect 3556 -160 3557 160
rect 3235 -161 3557 -160
rect 2812 -508 2916 -212
rect 2223 -560 2545 -559
rect 2223 -880 2224 -560
rect 2544 -880 2545 -560
rect 2223 -881 2545 -880
rect 1800 -1228 1904 -932
rect 1211 -1280 1533 -1279
rect 1211 -1600 1212 -1280
rect 1532 -1600 1533 -1280
rect 1211 -1601 1533 -1600
rect 788 -1948 892 -1652
rect 199 -2000 521 -1999
rect 199 -2320 200 -2000
rect 520 -2320 521 -2000
rect 199 -2321 521 -2320
rect -224 -2520 -120 -2372
rect 308 -2520 412 -2321
rect 788 -2372 808 -1948
rect 872 -2372 892 -1948
rect 1320 -1999 1424 -1601
rect 1800 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 2332 -1279 2436 -881
rect 2812 -932 2832 -508
rect 2896 -932 2916 -508
rect 3344 -559 3448 -161
rect 3824 -212 3844 212
rect 3908 -212 3928 212
rect 4356 161 4460 559
rect 4836 508 4856 932
rect 4920 508 4940 932
rect 5368 881 5472 1279
rect 5848 1228 5868 1652
rect 5932 1228 5952 1652
rect 6380 1601 6484 1999
rect 6860 1948 6880 2372
rect 6944 1948 6964 2372
rect 7392 2321 7496 2520
rect 7872 2372 7976 2520
rect 7283 2320 7605 2321
rect 7283 2000 7284 2320
rect 7604 2000 7605 2320
rect 7283 1999 7605 2000
rect 6860 1652 6964 1948
rect 6271 1600 6593 1601
rect 6271 1280 6272 1600
rect 6592 1280 6593 1600
rect 6271 1279 6593 1280
rect 5848 932 5952 1228
rect 5259 880 5581 881
rect 5259 560 5260 880
rect 5580 560 5581 880
rect 5259 559 5581 560
rect 4836 212 4940 508
rect 4247 160 4569 161
rect 4247 -160 4248 160
rect 4568 -160 4569 160
rect 4247 -161 4569 -160
rect 3824 -508 3928 -212
rect 3235 -560 3557 -559
rect 3235 -880 3236 -560
rect 3556 -880 3557 -560
rect 3235 -881 3557 -880
rect 2812 -1228 2916 -932
rect 2223 -1280 2545 -1279
rect 2223 -1600 2224 -1280
rect 2544 -1600 2545 -1280
rect 2223 -1601 2545 -1600
rect 1800 -1948 1904 -1652
rect 1211 -2000 1533 -1999
rect 1211 -2320 1212 -2000
rect 1532 -2320 1533 -2000
rect 1211 -2321 1533 -2320
rect 788 -2520 892 -2372
rect 1320 -2520 1424 -2321
rect 1800 -2372 1820 -1948
rect 1884 -2372 1904 -1948
rect 2332 -1999 2436 -1601
rect 2812 -1652 2832 -1228
rect 2896 -1652 2916 -1228
rect 3344 -1279 3448 -881
rect 3824 -932 3844 -508
rect 3908 -932 3928 -508
rect 4356 -559 4460 -161
rect 4836 -212 4856 212
rect 4920 -212 4940 212
rect 5368 161 5472 559
rect 5848 508 5868 932
rect 5932 508 5952 932
rect 6380 881 6484 1279
rect 6860 1228 6880 1652
rect 6944 1228 6964 1652
rect 7392 1601 7496 1999
rect 7872 1948 7892 2372
rect 7956 1948 7976 2372
rect 8404 2321 8508 2520
rect 8884 2372 8988 2520
rect 8295 2320 8617 2321
rect 8295 2000 8296 2320
rect 8616 2000 8617 2320
rect 8295 1999 8617 2000
rect 7872 1652 7976 1948
rect 7283 1600 7605 1601
rect 7283 1280 7284 1600
rect 7604 1280 7605 1600
rect 7283 1279 7605 1280
rect 6860 932 6964 1228
rect 6271 880 6593 881
rect 6271 560 6272 880
rect 6592 560 6593 880
rect 6271 559 6593 560
rect 5848 212 5952 508
rect 5259 160 5581 161
rect 5259 -160 5260 160
rect 5580 -160 5581 160
rect 5259 -161 5581 -160
rect 4836 -508 4940 -212
rect 4247 -560 4569 -559
rect 4247 -880 4248 -560
rect 4568 -880 4569 -560
rect 4247 -881 4569 -880
rect 3824 -1228 3928 -932
rect 3235 -1280 3557 -1279
rect 3235 -1600 3236 -1280
rect 3556 -1600 3557 -1280
rect 3235 -1601 3557 -1600
rect 2812 -1948 2916 -1652
rect 2223 -2000 2545 -1999
rect 2223 -2320 2224 -2000
rect 2544 -2320 2545 -2000
rect 2223 -2321 2545 -2320
rect 1800 -2520 1904 -2372
rect 2332 -2520 2436 -2321
rect 2812 -2372 2832 -1948
rect 2896 -2372 2916 -1948
rect 3344 -1999 3448 -1601
rect 3824 -1652 3844 -1228
rect 3908 -1652 3928 -1228
rect 4356 -1279 4460 -881
rect 4836 -932 4856 -508
rect 4920 -932 4940 -508
rect 5368 -559 5472 -161
rect 5848 -212 5868 212
rect 5932 -212 5952 212
rect 6380 161 6484 559
rect 6860 508 6880 932
rect 6944 508 6964 932
rect 7392 881 7496 1279
rect 7872 1228 7892 1652
rect 7956 1228 7976 1652
rect 8404 1601 8508 1999
rect 8884 1948 8904 2372
rect 8968 1948 8988 2372
rect 9416 2321 9520 2520
rect 9896 2372 10000 2520
rect 9307 2320 9629 2321
rect 9307 2000 9308 2320
rect 9628 2000 9629 2320
rect 9307 1999 9629 2000
rect 8884 1652 8988 1948
rect 8295 1600 8617 1601
rect 8295 1280 8296 1600
rect 8616 1280 8617 1600
rect 8295 1279 8617 1280
rect 7872 932 7976 1228
rect 7283 880 7605 881
rect 7283 560 7284 880
rect 7604 560 7605 880
rect 7283 559 7605 560
rect 6860 212 6964 508
rect 6271 160 6593 161
rect 6271 -160 6272 160
rect 6592 -160 6593 160
rect 6271 -161 6593 -160
rect 5848 -508 5952 -212
rect 5259 -560 5581 -559
rect 5259 -880 5260 -560
rect 5580 -880 5581 -560
rect 5259 -881 5581 -880
rect 4836 -1228 4940 -932
rect 4247 -1280 4569 -1279
rect 4247 -1600 4248 -1280
rect 4568 -1600 4569 -1280
rect 4247 -1601 4569 -1600
rect 3824 -1948 3928 -1652
rect 3235 -2000 3557 -1999
rect 3235 -2320 3236 -2000
rect 3556 -2320 3557 -2000
rect 3235 -2321 3557 -2320
rect 2812 -2520 2916 -2372
rect 3344 -2520 3448 -2321
rect 3824 -2372 3844 -1948
rect 3908 -2372 3928 -1948
rect 4356 -1999 4460 -1601
rect 4836 -1652 4856 -1228
rect 4920 -1652 4940 -1228
rect 5368 -1279 5472 -881
rect 5848 -932 5868 -508
rect 5932 -932 5952 -508
rect 6380 -559 6484 -161
rect 6860 -212 6880 212
rect 6944 -212 6964 212
rect 7392 161 7496 559
rect 7872 508 7892 932
rect 7956 508 7976 932
rect 8404 881 8508 1279
rect 8884 1228 8904 1652
rect 8968 1228 8988 1652
rect 9416 1601 9520 1999
rect 9896 1948 9916 2372
rect 9980 1948 10000 2372
rect 10428 2321 10532 2520
rect 10908 2372 11012 2520
rect 10319 2320 10641 2321
rect 10319 2000 10320 2320
rect 10640 2000 10641 2320
rect 10319 1999 10641 2000
rect 9896 1652 10000 1948
rect 9307 1600 9629 1601
rect 9307 1280 9308 1600
rect 9628 1280 9629 1600
rect 9307 1279 9629 1280
rect 8884 932 8988 1228
rect 8295 880 8617 881
rect 8295 560 8296 880
rect 8616 560 8617 880
rect 8295 559 8617 560
rect 7872 212 7976 508
rect 7283 160 7605 161
rect 7283 -160 7284 160
rect 7604 -160 7605 160
rect 7283 -161 7605 -160
rect 6860 -508 6964 -212
rect 6271 -560 6593 -559
rect 6271 -880 6272 -560
rect 6592 -880 6593 -560
rect 6271 -881 6593 -880
rect 5848 -1228 5952 -932
rect 5259 -1280 5581 -1279
rect 5259 -1600 5260 -1280
rect 5580 -1600 5581 -1280
rect 5259 -1601 5581 -1600
rect 4836 -1948 4940 -1652
rect 4247 -2000 4569 -1999
rect 4247 -2320 4248 -2000
rect 4568 -2320 4569 -2000
rect 4247 -2321 4569 -2320
rect 3824 -2520 3928 -2372
rect 4356 -2520 4460 -2321
rect 4836 -2372 4856 -1948
rect 4920 -2372 4940 -1948
rect 5368 -1999 5472 -1601
rect 5848 -1652 5868 -1228
rect 5932 -1652 5952 -1228
rect 6380 -1279 6484 -881
rect 6860 -932 6880 -508
rect 6944 -932 6964 -508
rect 7392 -559 7496 -161
rect 7872 -212 7892 212
rect 7956 -212 7976 212
rect 8404 161 8508 559
rect 8884 508 8904 932
rect 8968 508 8988 932
rect 9416 881 9520 1279
rect 9896 1228 9916 1652
rect 9980 1228 10000 1652
rect 10428 1601 10532 1999
rect 10908 1948 10928 2372
rect 10992 1948 11012 2372
rect 11440 2321 11544 2520
rect 11920 2372 12024 2520
rect 11331 2320 11653 2321
rect 11331 2000 11332 2320
rect 11652 2000 11653 2320
rect 11331 1999 11653 2000
rect 10908 1652 11012 1948
rect 10319 1600 10641 1601
rect 10319 1280 10320 1600
rect 10640 1280 10641 1600
rect 10319 1279 10641 1280
rect 9896 932 10000 1228
rect 9307 880 9629 881
rect 9307 560 9308 880
rect 9628 560 9629 880
rect 9307 559 9629 560
rect 8884 212 8988 508
rect 8295 160 8617 161
rect 8295 -160 8296 160
rect 8616 -160 8617 160
rect 8295 -161 8617 -160
rect 7872 -508 7976 -212
rect 7283 -560 7605 -559
rect 7283 -880 7284 -560
rect 7604 -880 7605 -560
rect 7283 -881 7605 -880
rect 6860 -1228 6964 -932
rect 6271 -1280 6593 -1279
rect 6271 -1600 6272 -1280
rect 6592 -1600 6593 -1280
rect 6271 -1601 6593 -1600
rect 5848 -1948 5952 -1652
rect 5259 -2000 5581 -1999
rect 5259 -2320 5260 -2000
rect 5580 -2320 5581 -2000
rect 5259 -2321 5581 -2320
rect 4836 -2520 4940 -2372
rect 5368 -2520 5472 -2321
rect 5848 -2372 5868 -1948
rect 5932 -2372 5952 -1948
rect 6380 -1999 6484 -1601
rect 6860 -1652 6880 -1228
rect 6944 -1652 6964 -1228
rect 7392 -1279 7496 -881
rect 7872 -932 7892 -508
rect 7956 -932 7976 -508
rect 8404 -559 8508 -161
rect 8884 -212 8904 212
rect 8968 -212 8988 212
rect 9416 161 9520 559
rect 9896 508 9916 932
rect 9980 508 10000 932
rect 10428 881 10532 1279
rect 10908 1228 10928 1652
rect 10992 1228 11012 1652
rect 11440 1601 11544 1999
rect 11920 1948 11940 2372
rect 12004 1948 12024 2372
rect 12452 2321 12556 2520
rect 12932 2372 13036 2520
rect 12343 2320 12665 2321
rect 12343 2000 12344 2320
rect 12664 2000 12665 2320
rect 12343 1999 12665 2000
rect 11920 1652 12024 1948
rect 11331 1600 11653 1601
rect 11331 1280 11332 1600
rect 11652 1280 11653 1600
rect 11331 1279 11653 1280
rect 10908 932 11012 1228
rect 10319 880 10641 881
rect 10319 560 10320 880
rect 10640 560 10641 880
rect 10319 559 10641 560
rect 9896 212 10000 508
rect 9307 160 9629 161
rect 9307 -160 9308 160
rect 9628 -160 9629 160
rect 9307 -161 9629 -160
rect 8884 -508 8988 -212
rect 8295 -560 8617 -559
rect 8295 -880 8296 -560
rect 8616 -880 8617 -560
rect 8295 -881 8617 -880
rect 7872 -1228 7976 -932
rect 7283 -1280 7605 -1279
rect 7283 -1600 7284 -1280
rect 7604 -1600 7605 -1280
rect 7283 -1601 7605 -1600
rect 6860 -1948 6964 -1652
rect 6271 -2000 6593 -1999
rect 6271 -2320 6272 -2000
rect 6592 -2320 6593 -2000
rect 6271 -2321 6593 -2320
rect 5848 -2520 5952 -2372
rect 6380 -2520 6484 -2321
rect 6860 -2372 6880 -1948
rect 6944 -2372 6964 -1948
rect 7392 -1999 7496 -1601
rect 7872 -1652 7892 -1228
rect 7956 -1652 7976 -1228
rect 8404 -1279 8508 -881
rect 8884 -932 8904 -508
rect 8968 -932 8988 -508
rect 9416 -559 9520 -161
rect 9896 -212 9916 212
rect 9980 -212 10000 212
rect 10428 161 10532 559
rect 10908 508 10928 932
rect 10992 508 11012 932
rect 11440 881 11544 1279
rect 11920 1228 11940 1652
rect 12004 1228 12024 1652
rect 12452 1601 12556 1999
rect 12932 1948 12952 2372
rect 13016 1948 13036 2372
rect 13464 2321 13568 2520
rect 13944 2372 14048 2520
rect 13355 2320 13677 2321
rect 13355 2000 13356 2320
rect 13676 2000 13677 2320
rect 13355 1999 13677 2000
rect 12932 1652 13036 1948
rect 12343 1600 12665 1601
rect 12343 1280 12344 1600
rect 12664 1280 12665 1600
rect 12343 1279 12665 1280
rect 11920 932 12024 1228
rect 11331 880 11653 881
rect 11331 560 11332 880
rect 11652 560 11653 880
rect 11331 559 11653 560
rect 10908 212 11012 508
rect 10319 160 10641 161
rect 10319 -160 10320 160
rect 10640 -160 10641 160
rect 10319 -161 10641 -160
rect 9896 -508 10000 -212
rect 9307 -560 9629 -559
rect 9307 -880 9308 -560
rect 9628 -880 9629 -560
rect 9307 -881 9629 -880
rect 8884 -1228 8988 -932
rect 8295 -1280 8617 -1279
rect 8295 -1600 8296 -1280
rect 8616 -1600 8617 -1280
rect 8295 -1601 8617 -1600
rect 7872 -1948 7976 -1652
rect 7283 -2000 7605 -1999
rect 7283 -2320 7284 -2000
rect 7604 -2320 7605 -2000
rect 7283 -2321 7605 -2320
rect 6860 -2520 6964 -2372
rect 7392 -2520 7496 -2321
rect 7872 -2372 7892 -1948
rect 7956 -2372 7976 -1948
rect 8404 -1999 8508 -1601
rect 8884 -1652 8904 -1228
rect 8968 -1652 8988 -1228
rect 9416 -1279 9520 -881
rect 9896 -932 9916 -508
rect 9980 -932 10000 -508
rect 10428 -559 10532 -161
rect 10908 -212 10928 212
rect 10992 -212 11012 212
rect 11440 161 11544 559
rect 11920 508 11940 932
rect 12004 508 12024 932
rect 12452 881 12556 1279
rect 12932 1228 12952 1652
rect 13016 1228 13036 1652
rect 13464 1601 13568 1999
rect 13944 1948 13964 2372
rect 14028 1948 14048 2372
rect 14476 2321 14580 2520
rect 14956 2372 15060 2520
rect 14367 2320 14689 2321
rect 14367 2000 14368 2320
rect 14688 2000 14689 2320
rect 14367 1999 14689 2000
rect 13944 1652 14048 1948
rect 13355 1600 13677 1601
rect 13355 1280 13356 1600
rect 13676 1280 13677 1600
rect 13355 1279 13677 1280
rect 12932 932 13036 1228
rect 12343 880 12665 881
rect 12343 560 12344 880
rect 12664 560 12665 880
rect 12343 559 12665 560
rect 11920 212 12024 508
rect 11331 160 11653 161
rect 11331 -160 11332 160
rect 11652 -160 11653 160
rect 11331 -161 11653 -160
rect 10908 -508 11012 -212
rect 10319 -560 10641 -559
rect 10319 -880 10320 -560
rect 10640 -880 10641 -560
rect 10319 -881 10641 -880
rect 9896 -1228 10000 -932
rect 9307 -1280 9629 -1279
rect 9307 -1600 9308 -1280
rect 9628 -1600 9629 -1280
rect 9307 -1601 9629 -1600
rect 8884 -1948 8988 -1652
rect 8295 -2000 8617 -1999
rect 8295 -2320 8296 -2000
rect 8616 -2320 8617 -2000
rect 8295 -2321 8617 -2320
rect 7872 -2520 7976 -2372
rect 8404 -2520 8508 -2321
rect 8884 -2372 8904 -1948
rect 8968 -2372 8988 -1948
rect 9416 -1999 9520 -1601
rect 9896 -1652 9916 -1228
rect 9980 -1652 10000 -1228
rect 10428 -1279 10532 -881
rect 10908 -932 10928 -508
rect 10992 -932 11012 -508
rect 11440 -559 11544 -161
rect 11920 -212 11940 212
rect 12004 -212 12024 212
rect 12452 161 12556 559
rect 12932 508 12952 932
rect 13016 508 13036 932
rect 13464 881 13568 1279
rect 13944 1228 13964 1652
rect 14028 1228 14048 1652
rect 14476 1601 14580 1999
rect 14956 1948 14976 2372
rect 15040 1948 15060 2372
rect 15488 2321 15592 2520
rect 15968 2372 16072 2520
rect 15379 2320 15701 2321
rect 15379 2000 15380 2320
rect 15700 2000 15701 2320
rect 15379 1999 15701 2000
rect 14956 1652 15060 1948
rect 14367 1600 14689 1601
rect 14367 1280 14368 1600
rect 14688 1280 14689 1600
rect 14367 1279 14689 1280
rect 13944 932 14048 1228
rect 13355 880 13677 881
rect 13355 560 13356 880
rect 13676 560 13677 880
rect 13355 559 13677 560
rect 12932 212 13036 508
rect 12343 160 12665 161
rect 12343 -160 12344 160
rect 12664 -160 12665 160
rect 12343 -161 12665 -160
rect 11920 -508 12024 -212
rect 11331 -560 11653 -559
rect 11331 -880 11332 -560
rect 11652 -880 11653 -560
rect 11331 -881 11653 -880
rect 10908 -1228 11012 -932
rect 10319 -1280 10641 -1279
rect 10319 -1600 10320 -1280
rect 10640 -1600 10641 -1280
rect 10319 -1601 10641 -1600
rect 9896 -1948 10000 -1652
rect 9307 -2000 9629 -1999
rect 9307 -2320 9308 -2000
rect 9628 -2320 9629 -2000
rect 9307 -2321 9629 -2320
rect 8884 -2520 8988 -2372
rect 9416 -2520 9520 -2321
rect 9896 -2372 9916 -1948
rect 9980 -2372 10000 -1948
rect 10428 -1999 10532 -1601
rect 10908 -1652 10928 -1228
rect 10992 -1652 11012 -1228
rect 11440 -1279 11544 -881
rect 11920 -932 11940 -508
rect 12004 -932 12024 -508
rect 12452 -559 12556 -161
rect 12932 -212 12952 212
rect 13016 -212 13036 212
rect 13464 161 13568 559
rect 13944 508 13964 932
rect 14028 508 14048 932
rect 14476 881 14580 1279
rect 14956 1228 14976 1652
rect 15040 1228 15060 1652
rect 15488 1601 15592 1999
rect 15968 1948 15988 2372
rect 16052 1948 16072 2372
rect 16500 2321 16604 2520
rect 16980 2372 17084 2520
rect 16391 2320 16713 2321
rect 16391 2000 16392 2320
rect 16712 2000 16713 2320
rect 16391 1999 16713 2000
rect 15968 1652 16072 1948
rect 15379 1600 15701 1601
rect 15379 1280 15380 1600
rect 15700 1280 15701 1600
rect 15379 1279 15701 1280
rect 14956 932 15060 1228
rect 14367 880 14689 881
rect 14367 560 14368 880
rect 14688 560 14689 880
rect 14367 559 14689 560
rect 13944 212 14048 508
rect 13355 160 13677 161
rect 13355 -160 13356 160
rect 13676 -160 13677 160
rect 13355 -161 13677 -160
rect 12932 -508 13036 -212
rect 12343 -560 12665 -559
rect 12343 -880 12344 -560
rect 12664 -880 12665 -560
rect 12343 -881 12665 -880
rect 11920 -1228 12024 -932
rect 11331 -1280 11653 -1279
rect 11331 -1600 11332 -1280
rect 11652 -1600 11653 -1280
rect 11331 -1601 11653 -1600
rect 10908 -1948 11012 -1652
rect 10319 -2000 10641 -1999
rect 10319 -2320 10320 -2000
rect 10640 -2320 10641 -2000
rect 10319 -2321 10641 -2320
rect 9896 -2520 10000 -2372
rect 10428 -2520 10532 -2321
rect 10908 -2372 10928 -1948
rect 10992 -2372 11012 -1948
rect 11440 -1999 11544 -1601
rect 11920 -1652 11940 -1228
rect 12004 -1652 12024 -1228
rect 12452 -1279 12556 -881
rect 12932 -932 12952 -508
rect 13016 -932 13036 -508
rect 13464 -559 13568 -161
rect 13944 -212 13964 212
rect 14028 -212 14048 212
rect 14476 161 14580 559
rect 14956 508 14976 932
rect 15040 508 15060 932
rect 15488 881 15592 1279
rect 15968 1228 15988 1652
rect 16052 1228 16072 1652
rect 16500 1601 16604 1999
rect 16980 1948 17000 2372
rect 17064 1948 17084 2372
rect 17512 2321 17616 2520
rect 17992 2372 18096 2520
rect 17403 2320 17725 2321
rect 17403 2000 17404 2320
rect 17724 2000 17725 2320
rect 17403 1999 17725 2000
rect 16980 1652 17084 1948
rect 16391 1600 16713 1601
rect 16391 1280 16392 1600
rect 16712 1280 16713 1600
rect 16391 1279 16713 1280
rect 15968 932 16072 1228
rect 15379 880 15701 881
rect 15379 560 15380 880
rect 15700 560 15701 880
rect 15379 559 15701 560
rect 14956 212 15060 508
rect 14367 160 14689 161
rect 14367 -160 14368 160
rect 14688 -160 14689 160
rect 14367 -161 14689 -160
rect 13944 -508 14048 -212
rect 13355 -560 13677 -559
rect 13355 -880 13356 -560
rect 13676 -880 13677 -560
rect 13355 -881 13677 -880
rect 12932 -1228 13036 -932
rect 12343 -1280 12665 -1279
rect 12343 -1600 12344 -1280
rect 12664 -1600 12665 -1280
rect 12343 -1601 12665 -1600
rect 11920 -1948 12024 -1652
rect 11331 -2000 11653 -1999
rect 11331 -2320 11332 -2000
rect 11652 -2320 11653 -2000
rect 11331 -2321 11653 -2320
rect 10908 -2520 11012 -2372
rect 11440 -2520 11544 -2321
rect 11920 -2372 11940 -1948
rect 12004 -2372 12024 -1948
rect 12452 -1999 12556 -1601
rect 12932 -1652 12952 -1228
rect 13016 -1652 13036 -1228
rect 13464 -1279 13568 -881
rect 13944 -932 13964 -508
rect 14028 -932 14048 -508
rect 14476 -559 14580 -161
rect 14956 -212 14976 212
rect 15040 -212 15060 212
rect 15488 161 15592 559
rect 15968 508 15988 932
rect 16052 508 16072 932
rect 16500 881 16604 1279
rect 16980 1228 17000 1652
rect 17064 1228 17084 1652
rect 17512 1601 17616 1999
rect 17992 1948 18012 2372
rect 18076 1948 18096 2372
rect 18524 2321 18628 2520
rect 19004 2372 19108 2520
rect 18415 2320 18737 2321
rect 18415 2000 18416 2320
rect 18736 2000 18737 2320
rect 18415 1999 18737 2000
rect 17992 1652 18096 1948
rect 17403 1600 17725 1601
rect 17403 1280 17404 1600
rect 17724 1280 17725 1600
rect 17403 1279 17725 1280
rect 16980 932 17084 1228
rect 16391 880 16713 881
rect 16391 560 16392 880
rect 16712 560 16713 880
rect 16391 559 16713 560
rect 15968 212 16072 508
rect 15379 160 15701 161
rect 15379 -160 15380 160
rect 15700 -160 15701 160
rect 15379 -161 15701 -160
rect 14956 -508 15060 -212
rect 14367 -560 14689 -559
rect 14367 -880 14368 -560
rect 14688 -880 14689 -560
rect 14367 -881 14689 -880
rect 13944 -1228 14048 -932
rect 13355 -1280 13677 -1279
rect 13355 -1600 13356 -1280
rect 13676 -1600 13677 -1280
rect 13355 -1601 13677 -1600
rect 12932 -1948 13036 -1652
rect 12343 -2000 12665 -1999
rect 12343 -2320 12344 -2000
rect 12664 -2320 12665 -2000
rect 12343 -2321 12665 -2320
rect 11920 -2520 12024 -2372
rect 12452 -2520 12556 -2321
rect 12932 -2372 12952 -1948
rect 13016 -2372 13036 -1948
rect 13464 -1999 13568 -1601
rect 13944 -1652 13964 -1228
rect 14028 -1652 14048 -1228
rect 14476 -1279 14580 -881
rect 14956 -932 14976 -508
rect 15040 -932 15060 -508
rect 15488 -559 15592 -161
rect 15968 -212 15988 212
rect 16052 -212 16072 212
rect 16500 161 16604 559
rect 16980 508 17000 932
rect 17064 508 17084 932
rect 17512 881 17616 1279
rect 17992 1228 18012 1652
rect 18076 1228 18096 1652
rect 18524 1601 18628 1999
rect 19004 1948 19024 2372
rect 19088 1948 19108 2372
rect 19536 2321 19640 2520
rect 20016 2372 20120 2520
rect 19427 2320 19749 2321
rect 19427 2000 19428 2320
rect 19748 2000 19749 2320
rect 19427 1999 19749 2000
rect 19004 1652 19108 1948
rect 18415 1600 18737 1601
rect 18415 1280 18416 1600
rect 18736 1280 18737 1600
rect 18415 1279 18737 1280
rect 17992 932 18096 1228
rect 17403 880 17725 881
rect 17403 560 17404 880
rect 17724 560 17725 880
rect 17403 559 17725 560
rect 16980 212 17084 508
rect 16391 160 16713 161
rect 16391 -160 16392 160
rect 16712 -160 16713 160
rect 16391 -161 16713 -160
rect 15968 -508 16072 -212
rect 15379 -560 15701 -559
rect 15379 -880 15380 -560
rect 15700 -880 15701 -560
rect 15379 -881 15701 -880
rect 14956 -1228 15060 -932
rect 14367 -1280 14689 -1279
rect 14367 -1600 14368 -1280
rect 14688 -1600 14689 -1280
rect 14367 -1601 14689 -1600
rect 13944 -1948 14048 -1652
rect 13355 -2000 13677 -1999
rect 13355 -2320 13356 -2000
rect 13676 -2320 13677 -2000
rect 13355 -2321 13677 -2320
rect 12932 -2520 13036 -2372
rect 13464 -2520 13568 -2321
rect 13944 -2372 13964 -1948
rect 14028 -2372 14048 -1948
rect 14476 -1999 14580 -1601
rect 14956 -1652 14976 -1228
rect 15040 -1652 15060 -1228
rect 15488 -1279 15592 -881
rect 15968 -932 15988 -508
rect 16052 -932 16072 -508
rect 16500 -559 16604 -161
rect 16980 -212 17000 212
rect 17064 -212 17084 212
rect 17512 161 17616 559
rect 17992 508 18012 932
rect 18076 508 18096 932
rect 18524 881 18628 1279
rect 19004 1228 19024 1652
rect 19088 1228 19108 1652
rect 19536 1601 19640 1999
rect 20016 1948 20036 2372
rect 20100 1948 20120 2372
rect 20548 2321 20652 2520
rect 21028 2372 21132 2520
rect 20439 2320 20761 2321
rect 20439 2000 20440 2320
rect 20760 2000 20761 2320
rect 20439 1999 20761 2000
rect 20016 1652 20120 1948
rect 19427 1600 19749 1601
rect 19427 1280 19428 1600
rect 19748 1280 19749 1600
rect 19427 1279 19749 1280
rect 19004 932 19108 1228
rect 18415 880 18737 881
rect 18415 560 18416 880
rect 18736 560 18737 880
rect 18415 559 18737 560
rect 17992 212 18096 508
rect 17403 160 17725 161
rect 17403 -160 17404 160
rect 17724 -160 17725 160
rect 17403 -161 17725 -160
rect 16980 -508 17084 -212
rect 16391 -560 16713 -559
rect 16391 -880 16392 -560
rect 16712 -880 16713 -560
rect 16391 -881 16713 -880
rect 15968 -1228 16072 -932
rect 15379 -1280 15701 -1279
rect 15379 -1600 15380 -1280
rect 15700 -1600 15701 -1280
rect 15379 -1601 15701 -1600
rect 14956 -1948 15060 -1652
rect 14367 -2000 14689 -1999
rect 14367 -2320 14368 -2000
rect 14688 -2320 14689 -2000
rect 14367 -2321 14689 -2320
rect 13944 -2520 14048 -2372
rect 14476 -2520 14580 -2321
rect 14956 -2372 14976 -1948
rect 15040 -2372 15060 -1948
rect 15488 -1999 15592 -1601
rect 15968 -1652 15988 -1228
rect 16052 -1652 16072 -1228
rect 16500 -1279 16604 -881
rect 16980 -932 17000 -508
rect 17064 -932 17084 -508
rect 17512 -559 17616 -161
rect 17992 -212 18012 212
rect 18076 -212 18096 212
rect 18524 161 18628 559
rect 19004 508 19024 932
rect 19088 508 19108 932
rect 19536 881 19640 1279
rect 20016 1228 20036 1652
rect 20100 1228 20120 1652
rect 20548 1601 20652 1999
rect 21028 1948 21048 2372
rect 21112 1948 21132 2372
rect 21560 2321 21664 2520
rect 22040 2372 22144 2520
rect 21451 2320 21773 2321
rect 21451 2000 21452 2320
rect 21772 2000 21773 2320
rect 21451 1999 21773 2000
rect 21028 1652 21132 1948
rect 20439 1600 20761 1601
rect 20439 1280 20440 1600
rect 20760 1280 20761 1600
rect 20439 1279 20761 1280
rect 20016 932 20120 1228
rect 19427 880 19749 881
rect 19427 560 19428 880
rect 19748 560 19749 880
rect 19427 559 19749 560
rect 19004 212 19108 508
rect 18415 160 18737 161
rect 18415 -160 18416 160
rect 18736 -160 18737 160
rect 18415 -161 18737 -160
rect 17992 -508 18096 -212
rect 17403 -560 17725 -559
rect 17403 -880 17404 -560
rect 17724 -880 17725 -560
rect 17403 -881 17725 -880
rect 16980 -1228 17084 -932
rect 16391 -1280 16713 -1279
rect 16391 -1600 16392 -1280
rect 16712 -1600 16713 -1280
rect 16391 -1601 16713 -1600
rect 15968 -1948 16072 -1652
rect 15379 -2000 15701 -1999
rect 15379 -2320 15380 -2000
rect 15700 -2320 15701 -2000
rect 15379 -2321 15701 -2320
rect 14956 -2520 15060 -2372
rect 15488 -2520 15592 -2321
rect 15968 -2372 15988 -1948
rect 16052 -2372 16072 -1948
rect 16500 -1999 16604 -1601
rect 16980 -1652 17000 -1228
rect 17064 -1652 17084 -1228
rect 17512 -1279 17616 -881
rect 17992 -932 18012 -508
rect 18076 -932 18096 -508
rect 18524 -559 18628 -161
rect 19004 -212 19024 212
rect 19088 -212 19108 212
rect 19536 161 19640 559
rect 20016 508 20036 932
rect 20100 508 20120 932
rect 20548 881 20652 1279
rect 21028 1228 21048 1652
rect 21112 1228 21132 1652
rect 21560 1601 21664 1999
rect 22040 1948 22060 2372
rect 22124 1948 22144 2372
rect 22572 2321 22676 2520
rect 23052 2372 23156 2520
rect 22463 2320 22785 2321
rect 22463 2000 22464 2320
rect 22784 2000 22785 2320
rect 22463 1999 22785 2000
rect 22040 1652 22144 1948
rect 21451 1600 21773 1601
rect 21451 1280 21452 1600
rect 21772 1280 21773 1600
rect 21451 1279 21773 1280
rect 21028 932 21132 1228
rect 20439 880 20761 881
rect 20439 560 20440 880
rect 20760 560 20761 880
rect 20439 559 20761 560
rect 20016 212 20120 508
rect 19427 160 19749 161
rect 19427 -160 19428 160
rect 19748 -160 19749 160
rect 19427 -161 19749 -160
rect 19004 -508 19108 -212
rect 18415 -560 18737 -559
rect 18415 -880 18416 -560
rect 18736 -880 18737 -560
rect 18415 -881 18737 -880
rect 17992 -1228 18096 -932
rect 17403 -1280 17725 -1279
rect 17403 -1600 17404 -1280
rect 17724 -1600 17725 -1280
rect 17403 -1601 17725 -1600
rect 16980 -1948 17084 -1652
rect 16391 -2000 16713 -1999
rect 16391 -2320 16392 -2000
rect 16712 -2320 16713 -2000
rect 16391 -2321 16713 -2320
rect 15968 -2520 16072 -2372
rect 16500 -2520 16604 -2321
rect 16980 -2372 17000 -1948
rect 17064 -2372 17084 -1948
rect 17512 -1999 17616 -1601
rect 17992 -1652 18012 -1228
rect 18076 -1652 18096 -1228
rect 18524 -1279 18628 -881
rect 19004 -932 19024 -508
rect 19088 -932 19108 -508
rect 19536 -559 19640 -161
rect 20016 -212 20036 212
rect 20100 -212 20120 212
rect 20548 161 20652 559
rect 21028 508 21048 932
rect 21112 508 21132 932
rect 21560 881 21664 1279
rect 22040 1228 22060 1652
rect 22124 1228 22144 1652
rect 22572 1601 22676 1999
rect 23052 1948 23072 2372
rect 23136 1948 23156 2372
rect 23584 2321 23688 2520
rect 24064 2372 24168 2520
rect 23475 2320 23797 2321
rect 23475 2000 23476 2320
rect 23796 2000 23797 2320
rect 23475 1999 23797 2000
rect 23052 1652 23156 1948
rect 22463 1600 22785 1601
rect 22463 1280 22464 1600
rect 22784 1280 22785 1600
rect 22463 1279 22785 1280
rect 22040 932 22144 1228
rect 21451 880 21773 881
rect 21451 560 21452 880
rect 21772 560 21773 880
rect 21451 559 21773 560
rect 21028 212 21132 508
rect 20439 160 20761 161
rect 20439 -160 20440 160
rect 20760 -160 20761 160
rect 20439 -161 20761 -160
rect 20016 -508 20120 -212
rect 19427 -560 19749 -559
rect 19427 -880 19428 -560
rect 19748 -880 19749 -560
rect 19427 -881 19749 -880
rect 19004 -1228 19108 -932
rect 18415 -1280 18737 -1279
rect 18415 -1600 18416 -1280
rect 18736 -1600 18737 -1280
rect 18415 -1601 18737 -1600
rect 17992 -1948 18096 -1652
rect 17403 -2000 17725 -1999
rect 17403 -2320 17404 -2000
rect 17724 -2320 17725 -2000
rect 17403 -2321 17725 -2320
rect 16980 -2520 17084 -2372
rect 17512 -2520 17616 -2321
rect 17992 -2372 18012 -1948
rect 18076 -2372 18096 -1948
rect 18524 -1999 18628 -1601
rect 19004 -1652 19024 -1228
rect 19088 -1652 19108 -1228
rect 19536 -1279 19640 -881
rect 20016 -932 20036 -508
rect 20100 -932 20120 -508
rect 20548 -559 20652 -161
rect 21028 -212 21048 212
rect 21112 -212 21132 212
rect 21560 161 21664 559
rect 22040 508 22060 932
rect 22124 508 22144 932
rect 22572 881 22676 1279
rect 23052 1228 23072 1652
rect 23136 1228 23156 1652
rect 23584 1601 23688 1999
rect 24064 1948 24084 2372
rect 24148 1948 24168 2372
rect 24596 2321 24700 2520
rect 25076 2372 25180 2520
rect 24487 2320 24809 2321
rect 24487 2000 24488 2320
rect 24808 2000 24809 2320
rect 24487 1999 24809 2000
rect 24064 1652 24168 1948
rect 23475 1600 23797 1601
rect 23475 1280 23476 1600
rect 23796 1280 23797 1600
rect 23475 1279 23797 1280
rect 23052 932 23156 1228
rect 22463 880 22785 881
rect 22463 560 22464 880
rect 22784 560 22785 880
rect 22463 559 22785 560
rect 22040 212 22144 508
rect 21451 160 21773 161
rect 21451 -160 21452 160
rect 21772 -160 21773 160
rect 21451 -161 21773 -160
rect 21028 -508 21132 -212
rect 20439 -560 20761 -559
rect 20439 -880 20440 -560
rect 20760 -880 20761 -560
rect 20439 -881 20761 -880
rect 20016 -1228 20120 -932
rect 19427 -1280 19749 -1279
rect 19427 -1600 19428 -1280
rect 19748 -1600 19749 -1280
rect 19427 -1601 19749 -1600
rect 19004 -1948 19108 -1652
rect 18415 -2000 18737 -1999
rect 18415 -2320 18416 -2000
rect 18736 -2320 18737 -2000
rect 18415 -2321 18737 -2320
rect 17992 -2520 18096 -2372
rect 18524 -2520 18628 -2321
rect 19004 -2372 19024 -1948
rect 19088 -2372 19108 -1948
rect 19536 -1999 19640 -1601
rect 20016 -1652 20036 -1228
rect 20100 -1652 20120 -1228
rect 20548 -1279 20652 -881
rect 21028 -932 21048 -508
rect 21112 -932 21132 -508
rect 21560 -559 21664 -161
rect 22040 -212 22060 212
rect 22124 -212 22144 212
rect 22572 161 22676 559
rect 23052 508 23072 932
rect 23136 508 23156 932
rect 23584 881 23688 1279
rect 24064 1228 24084 1652
rect 24148 1228 24168 1652
rect 24596 1601 24700 1999
rect 25076 1948 25096 2372
rect 25160 1948 25180 2372
rect 25608 2321 25712 2520
rect 26088 2372 26192 2520
rect 25499 2320 25821 2321
rect 25499 2000 25500 2320
rect 25820 2000 25821 2320
rect 25499 1999 25821 2000
rect 25076 1652 25180 1948
rect 24487 1600 24809 1601
rect 24487 1280 24488 1600
rect 24808 1280 24809 1600
rect 24487 1279 24809 1280
rect 24064 932 24168 1228
rect 23475 880 23797 881
rect 23475 560 23476 880
rect 23796 560 23797 880
rect 23475 559 23797 560
rect 23052 212 23156 508
rect 22463 160 22785 161
rect 22463 -160 22464 160
rect 22784 -160 22785 160
rect 22463 -161 22785 -160
rect 22040 -508 22144 -212
rect 21451 -560 21773 -559
rect 21451 -880 21452 -560
rect 21772 -880 21773 -560
rect 21451 -881 21773 -880
rect 21028 -1228 21132 -932
rect 20439 -1280 20761 -1279
rect 20439 -1600 20440 -1280
rect 20760 -1600 20761 -1280
rect 20439 -1601 20761 -1600
rect 20016 -1948 20120 -1652
rect 19427 -2000 19749 -1999
rect 19427 -2320 19428 -2000
rect 19748 -2320 19749 -2000
rect 19427 -2321 19749 -2320
rect 19004 -2520 19108 -2372
rect 19536 -2520 19640 -2321
rect 20016 -2372 20036 -1948
rect 20100 -2372 20120 -1948
rect 20548 -1999 20652 -1601
rect 21028 -1652 21048 -1228
rect 21112 -1652 21132 -1228
rect 21560 -1279 21664 -881
rect 22040 -932 22060 -508
rect 22124 -932 22144 -508
rect 22572 -559 22676 -161
rect 23052 -212 23072 212
rect 23136 -212 23156 212
rect 23584 161 23688 559
rect 24064 508 24084 932
rect 24148 508 24168 932
rect 24596 881 24700 1279
rect 25076 1228 25096 1652
rect 25160 1228 25180 1652
rect 25608 1601 25712 1999
rect 26088 1948 26108 2372
rect 26172 1948 26192 2372
rect 26620 2321 26724 2520
rect 27100 2372 27204 2520
rect 26511 2320 26833 2321
rect 26511 2000 26512 2320
rect 26832 2000 26833 2320
rect 26511 1999 26833 2000
rect 26088 1652 26192 1948
rect 25499 1600 25821 1601
rect 25499 1280 25500 1600
rect 25820 1280 25821 1600
rect 25499 1279 25821 1280
rect 25076 932 25180 1228
rect 24487 880 24809 881
rect 24487 560 24488 880
rect 24808 560 24809 880
rect 24487 559 24809 560
rect 24064 212 24168 508
rect 23475 160 23797 161
rect 23475 -160 23476 160
rect 23796 -160 23797 160
rect 23475 -161 23797 -160
rect 23052 -508 23156 -212
rect 22463 -560 22785 -559
rect 22463 -880 22464 -560
rect 22784 -880 22785 -560
rect 22463 -881 22785 -880
rect 22040 -1228 22144 -932
rect 21451 -1280 21773 -1279
rect 21451 -1600 21452 -1280
rect 21772 -1600 21773 -1280
rect 21451 -1601 21773 -1600
rect 21028 -1948 21132 -1652
rect 20439 -2000 20761 -1999
rect 20439 -2320 20440 -2000
rect 20760 -2320 20761 -2000
rect 20439 -2321 20761 -2320
rect 20016 -2520 20120 -2372
rect 20548 -2520 20652 -2321
rect 21028 -2372 21048 -1948
rect 21112 -2372 21132 -1948
rect 21560 -1999 21664 -1601
rect 22040 -1652 22060 -1228
rect 22124 -1652 22144 -1228
rect 22572 -1279 22676 -881
rect 23052 -932 23072 -508
rect 23136 -932 23156 -508
rect 23584 -559 23688 -161
rect 24064 -212 24084 212
rect 24148 -212 24168 212
rect 24596 161 24700 559
rect 25076 508 25096 932
rect 25160 508 25180 932
rect 25608 881 25712 1279
rect 26088 1228 26108 1652
rect 26172 1228 26192 1652
rect 26620 1601 26724 1999
rect 27100 1948 27120 2372
rect 27184 1948 27204 2372
rect 27632 2321 27736 2520
rect 28112 2372 28216 2520
rect 27523 2320 27845 2321
rect 27523 2000 27524 2320
rect 27844 2000 27845 2320
rect 27523 1999 27845 2000
rect 27100 1652 27204 1948
rect 26511 1600 26833 1601
rect 26511 1280 26512 1600
rect 26832 1280 26833 1600
rect 26511 1279 26833 1280
rect 26088 932 26192 1228
rect 25499 880 25821 881
rect 25499 560 25500 880
rect 25820 560 25821 880
rect 25499 559 25821 560
rect 25076 212 25180 508
rect 24487 160 24809 161
rect 24487 -160 24488 160
rect 24808 -160 24809 160
rect 24487 -161 24809 -160
rect 24064 -508 24168 -212
rect 23475 -560 23797 -559
rect 23475 -880 23476 -560
rect 23796 -880 23797 -560
rect 23475 -881 23797 -880
rect 23052 -1228 23156 -932
rect 22463 -1280 22785 -1279
rect 22463 -1600 22464 -1280
rect 22784 -1600 22785 -1280
rect 22463 -1601 22785 -1600
rect 22040 -1948 22144 -1652
rect 21451 -2000 21773 -1999
rect 21451 -2320 21452 -2000
rect 21772 -2320 21773 -2000
rect 21451 -2321 21773 -2320
rect 21028 -2520 21132 -2372
rect 21560 -2520 21664 -2321
rect 22040 -2372 22060 -1948
rect 22124 -2372 22144 -1948
rect 22572 -1999 22676 -1601
rect 23052 -1652 23072 -1228
rect 23136 -1652 23156 -1228
rect 23584 -1279 23688 -881
rect 24064 -932 24084 -508
rect 24148 -932 24168 -508
rect 24596 -559 24700 -161
rect 25076 -212 25096 212
rect 25160 -212 25180 212
rect 25608 161 25712 559
rect 26088 508 26108 932
rect 26172 508 26192 932
rect 26620 881 26724 1279
rect 27100 1228 27120 1652
rect 27184 1228 27204 1652
rect 27632 1601 27736 1999
rect 28112 1948 28132 2372
rect 28196 1948 28216 2372
rect 28644 2321 28748 2520
rect 29124 2372 29228 2520
rect 28535 2320 28857 2321
rect 28535 2000 28536 2320
rect 28856 2000 28857 2320
rect 28535 1999 28857 2000
rect 28112 1652 28216 1948
rect 27523 1600 27845 1601
rect 27523 1280 27524 1600
rect 27844 1280 27845 1600
rect 27523 1279 27845 1280
rect 27100 932 27204 1228
rect 26511 880 26833 881
rect 26511 560 26512 880
rect 26832 560 26833 880
rect 26511 559 26833 560
rect 26088 212 26192 508
rect 25499 160 25821 161
rect 25499 -160 25500 160
rect 25820 -160 25821 160
rect 25499 -161 25821 -160
rect 25076 -508 25180 -212
rect 24487 -560 24809 -559
rect 24487 -880 24488 -560
rect 24808 -880 24809 -560
rect 24487 -881 24809 -880
rect 24064 -1228 24168 -932
rect 23475 -1280 23797 -1279
rect 23475 -1600 23476 -1280
rect 23796 -1600 23797 -1280
rect 23475 -1601 23797 -1600
rect 23052 -1948 23156 -1652
rect 22463 -2000 22785 -1999
rect 22463 -2320 22464 -2000
rect 22784 -2320 22785 -2000
rect 22463 -2321 22785 -2320
rect 22040 -2520 22144 -2372
rect 22572 -2520 22676 -2321
rect 23052 -2372 23072 -1948
rect 23136 -2372 23156 -1948
rect 23584 -1999 23688 -1601
rect 24064 -1652 24084 -1228
rect 24148 -1652 24168 -1228
rect 24596 -1279 24700 -881
rect 25076 -932 25096 -508
rect 25160 -932 25180 -508
rect 25608 -559 25712 -161
rect 26088 -212 26108 212
rect 26172 -212 26192 212
rect 26620 161 26724 559
rect 27100 508 27120 932
rect 27184 508 27204 932
rect 27632 881 27736 1279
rect 28112 1228 28132 1652
rect 28196 1228 28216 1652
rect 28644 1601 28748 1999
rect 29124 1948 29144 2372
rect 29208 1948 29228 2372
rect 29656 2321 29760 2520
rect 30136 2372 30240 2520
rect 29547 2320 29869 2321
rect 29547 2000 29548 2320
rect 29868 2000 29869 2320
rect 29547 1999 29869 2000
rect 29124 1652 29228 1948
rect 28535 1600 28857 1601
rect 28535 1280 28536 1600
rect 28856 1280 28857 1600
rect 28535 1279 28857 1280
rect 28112 932 28216 1228
rect 27523 880 27845 881
rect 27523 560 27524 880
rect 27844 560 27845 880
rect 27523 559 27845 560
rect 27100 212 27204 508
rect 26511 160 26833 161
rect 26511 -160 26512 160
rect 26832 -160 26833 160
rect 26511 -161 26833 -160
rect 26088 -508 26192 -212
rect 25499 -560 25821 -559
rect 25499 -880 25500 -560
rect 25820 -880 25821 -560
rect 25499 -881 25821 -880
rect 25076 -1228 25180 -932
rect 24487 -1280 24809 -1279
rect 24487 -1600 24488 -1280
rect 24808 -1600 24809 -1280
rect 24487 -1601 24809 -1600
rect 24064 -1948 24168 -1652
rect 23475 -2000 23797 -1999
rect 23475 -2320 23476 -2000
rect 23796 -2320 23797 -2000
rect 23475 -2321 23797 -2320
rect 23052 -2520 23156 -2372
rect 23584 -2520 23688 -2321
rect 24064 -2372 24084 -1948
rect 24148 -2372 24168 -1948
rect 24596 -1999 24700 -1601
rect 25076 -1652 25096 -1228
rect 25160 -1652 25180 -1228
rect 25608 -1279 25712 -881
rect 26088 -932 26108 -508
rect 26172 -932 26192 -508
rect 26620 -559 26724 -161
rect 27100 -212 27120 212
rect 27184 -212 27204 212
rect 27632 161 27736 559
rect 28112 508 28132 932
rect 28196 508 28216 932
rect 28644 881 28748 1279
rect 29124 1228 29144 1652
rect 29208 1228 29228 1652
rect 29656 1601 29760 1999
rect 30136 1948 30156 2372
rect 30220 1948 30240 2372
rect 30668 2321 30772 2520
rect 31148 2372 31252 2520
rect 30559 2320 30881 2321
rect 30559 2000 30560 2320
rect 30880 2000 30881 2320
rect 30559 1999 30881 2000
rect 30136 1652 30240 1948
rect 29547 1600 29869 1601
rect 29547 1280 29548 1600
rect 29868 1280 29869 1600
rect 29547 1279 29869 1280
rect 29124 932 29228 1228
rect 28535 880 28857 881
rect 28535 560 28536 880
rect 28856 560 28857 880
rect 28535 559 28857 560
rect 28112 212 28216 508
rect 27523 160 27845 161
rect 27523 -160 27524 160
rect 27844 -160 27845 160
rect 27523 -161 27845 -160
rect 27100 -508 27204 -212
rect 26511 -560 26833 -559
rect 26511 -880 26512 -560
rect 26832 -880 26833 -560
rect 26511 -881 26833 -880
rect 26088 -1228 26192 -932
rect 25499 -1280 25821 -1279
rect 25499 -1600 25500 -1280
rect 25820 -1600 25821 -1280
rect 25499 -1601 25821 -1600
rect 25076 -1948 25180 -1652
rect 24487 -2000 24809 -1999
rect 24487 -2320 24488 -2000
rect 24808 -2320 24809 -2000
rect 24487 -2321 24809 -2320
rect 24064 -2520 24168 -2372
rect 24596 -2520 24700 -2321
rect 25076 -2372 25096 -1948
rect 25160 -2372 25180 -1948
rect 25608 -1999 25712 -1601
rect 26088 -1652 26108 -1228
rect 26172 -1652 26192 -1228
rect 26620 -1279 26724 -881
rect 27100 -932 27120 -508
rect 27184 -932 27204 -508
rect 27632 -559 27736 -161
rect 28112 -212 28132 212
rect 28196 -212 28216 212
rect 28644 161 28748 559
rect 29124 508 29144 932
rect 29208 508 29228 932
rect 29656 881 29760 1279
rect 30136 1228 30156 1652
rect 30220 1228 30240 1652
rect 30668 1601 30772 1999
rect 31148 1948 31168 2372
rect 31232 1948 31252 2372
rect 31680 2321 31784 2520
rect 32160 2372 32264 2520
rect 31571 2320 31893 2321
rect 31571 2000 31572 2320
rect 31892 2000 31893 2320
rect 31571 1999 31893 2000
rect 31148 1652 31252 1948
rect 30559 1600 30881 1601
rect 30559 1280 30560 1600
rect 30880 1280 30881 1600
rect 30559 1279 30881 1280
rect 30136 932 30240 1228
rect 29547 880 29869 881
rect 29547 560 29548 880
rect 29868 560 29869 880
rect 29547 559 29869 560
rect 29124 212 29228 508
rect 28535 160 28857 161
rect 28535 -160 28536 160
rect 28856 -160 28857 160
rect 28535 -161 28857 -160
rect 28112 -508 28216 -212
rect 27523 -560 27845 -559
rect 27523 -880 27524 -560
rect 27844 -880 27845 -560
rect 27523 -881 27845 -880
rect 27100 -1228 27204 -932
rect 26511 -1280 26833 -1279
rect 26511 -1600 26512 -1280
rect 26832 -1600 26833 -1280
rect 26511 -1601 26833 -1600
rect 26088 -1948 26192 -1652
rect 25499 -2000 25821 -1999
rect 25499 -2320 25500 -2000
rect 25820 -2320 25821 -2000
rect 25499 -2321 25821 -2320
rect 25076 -2520 25180 -2372
rect 25608 -2520 25712 -2321
rect 26088 -2372 26108 -1948
rect 26172 -2372 26192 -1948
rect 26620 -1999 26724 -1601
rect 27100 -1652 27120 -1228
rect 27184 -1652 27204 -1228
rect 27632 -1279 27736 -881
rect 28112 -932 28132 -508
rect 28196 -932 28216 -508
rect 28644 -559 28748 -161
rect 29124 -212 29144 212
rect 29208 -212 29228 212
rect 29656 161 29760 559
rect 30136 508 30156 932
rect 30220 508 30240 932
rect 30668 881 30772 1279
rect 31148 1228 31168 1652
rect 31232 1228 31252 1652
rect 31680 1601 31784 1999
rect 32160 1948 32180 2372
rect 32244 1948 32264 2372
rect 32160 1652 32264 1948
rect 31571 1600 31893 1601
rect 31571 1280 31572 1600
rect 31892 1280 31893 1600
rect 31571 1279 31893 1280
rect 31148 932 31252 1228
rect 30559 880 30881 881
rect 30559 560 30560 880
rect 30880 560 30881 880
rect 30559 559 30881 560
rect 30136 212 30240 508
rect 29547 160 29869 161
rect 29547 -160 29548 160
rect 29868 -160 29869 160
rect 29547 -161 29869 -160
rect 29124 -508 29228 -212
rect 28535 -560 28857 -559
rect 28535 -880 28536 -560
rect 28856 -880 28857 -560
rect 28535 -881 28857 -880
rect 28112 -1228 28216 -932
rect 27523 -1280 27845 -1279
rect 27523 -1600 27524 -1280
rect 27844 -1600 27845 -1280
rect 27523 -1601 27845 -1600
rect 27100 -1948 27204 -1652
rect 26511 -2000 26833 -1999
rect 26511 -2320 26512 -2000
rect 26832 -2320 26833 -2000
rect 26511 -2321 26833 -2320
rect 26088 -2520 26192 -2372
rect 26620 -2520 26724 -2321
rect 27100 -2372 27120 -1948
rect 27184 -2372 27204 -1948
rect 27632 -1999 27736 -1601
rect 28112 -1652 28132 -1228
rect 28196 -1652 28216 -1228
rect 28644 -1279 28748 -881
rect 29124 -932 29144 -508
rect 29208 -932 29228 -508
rect 29656 -559 29760 -161
rect 30136 -212 30156 212
rect 30220 -212 30240 212
rect 30668 161 30772 559
rect 31148 508 31168 932
rect 31232 508 31252 932
rect 31680 881 31784 1279
rect 32160 1228 32180 1652
rect 32244 1228 32264 1652
rect 32160 932 32264 1228
rect 31571 880 31893 881
rect 31571 560 31572 880
rect 31892 560 31893 880
rect 31571 559 31893 560
rect 31148 212 31252 508
rect 30559 160 30881 161
rect 30559 -160 30560 160
rect 30880 -160 30881 160
rect 30559 -161 30881 -160
rect 30136 -508 30240 -212
rect 29547 -560 29869 -559
rect 29547 -880 29548 -560
rect 29868 -880 29869 -560
rect 29547 -881 29869 -880
rect 29124 -1228 29228 -932
rect 28535 -1280 28857 -1279
rect 28535 -1600 28536 -1280
rect 28856 -1600 28857 -1280
rect 28535 -1601 28857 -1600
rect 28112 -1948 28216 -1652
rect 27523 -2000 27845 -1999
rect 27523 -2320 27524 -2000
rect 27844 -2320 27845 -2000
rect 27523 -2321 27845 -2320
rect 27100 -2520 27204 -2372
rect 27632 -2520 27736 -2321
rect 28112 -2372 28132 -1948
rect 28196 -2372 28216 -1948
rect 28644 -1999 28748 -1601
rect 29124 -1652 29144 -1228
rect 29208 -1652 29228 -1228
rect 29656 -1279 29760 -881
rect 30136 -932 30156 -508
rect 30220 -932 30240 -508
rect 30668 -559 30772 -161
rect 31148 -212 31168 212
rect 31232 -212 31252 212
rect 31680 161 31784 559
rect 32160 508 32180 932
rect 32244 508 32264 932
rect 32160 212 32264 508
rect 31571 160 31893 161
rect 31571 -160 31572 160
rect 31892 -160 31893 160
rect 31571 -161 31893 -160
rect 31148 -508 31252 -212
rect 30559 -560 30881 -559
rect 30559 -880 30560 -560
rect 30880 -880 30881 -560
rect 30559 -881 30881 -880
rect 30136 -1228 30240 -932
rect 29547 -1280 29869 -1279
rect 29547 -1600 29548 -1280
rect 29868 -1600 29869 -1280
rect 29547 -1601 29869 -1600
rect 29124 -1948 29228 -1652
rect 28535 -2000 28857 -1999
rect 28535 -2320 28536 -2000
rect 28856 -2320 28857 -2000
rect 28535 -2321 28857 -2320
rect 28112 -2520 28216 -2372
rect 28644 -2520 28748 -2321
rect 29124 -2372 29144 -1948
rect 29208 -2372 29228 -1948
rect 29656 -1999 29760 -1601
rect 30136 -1652 30156 -1228
rect 30220 -1652 30240 -1228
rect 30668 -1279 30772 -881
rect 31148 -932 31168 -508
rect 31232 -932 31252 -508
rect 31680 -559 31784 -161
rect 32160 -212 32180 212
rect 32244 -212 32264 212
rect 32160 -508 32264 -212
rect 31571 -560 31893 -559
rect 31571 -880 31572 -560
rect 31892 -880 31893 -560
rect 31571 -881 31893 -880
rect 31148 -1228 31252 -932
rect 30559 -1280 30881 -1279
rect 30559 -1600 30560 -1280
rect 30880 -1600 30881 -1280
rect 30559 -1601 30881 -1600
rect 30136 -1948 30240 -1652
rect 29547 -2000 29869 -1999
rect 29547 -2320 29548 -2000
rect 29868 -2320 29869 -2000
rect 29547 -2321 29869 -2320
rect 29124 -2520 29228 -2372
rect 29656 -2520 29760 -2321
rect 30136 -2372 30156 -1948
rect 30220 -2372 30240 -1948
rect 30668 -1999 30772 -1601
rect 31148 -1652 31168 -1228
rect 31232 -1652 31252 -1228
rect 31680 -1279 31784 -881
rect 32160 -932 32180 -508
rect 32244 -932 32264 -508
rect 32160 -1228 32264 -932
rect 31571 -1280 31893 -1279
rect 31571 -1600 31572 -1280
rect 31892 -1600 31893 -1280
rect 31571 -1601 31893 -1600
rect 31148 -1948 31252 -1652
rect 30559 -2000 30881 -1999
rect 30559 -2320 30560 -2000
rect 30880 -2320 30881 -2000
rect 30559 -2321 30881 -2320
rect 30136 -2520 30240 -2372
rect 30668 -2520 30772 -2321
rect 31148 -2372 31168 -1948
rect 31232 -2372 31252 -1948
rect 31680 -1999 31784 -1601
rect 32160 -1652 32180 -1228
rect 32244 -1652 32264 -1228
rect 32160 -1948 32264 -1652
rect 31571 -2000 31893 -1999
rect 31571 -2320 31572 -2000
rect 31892 -2320 31893 -2000
rect 31571 -2321 31893 -2320
rect 31148 -2520 31252 -2372
rect 31680 -2520 31784 -2321
rect 32160 -2372 32180 -1948
rect 32244 -2372 32264 -1948
rect 32160 -2520 32264 -2372
<< properties >>
string FIXED_BBOX 31492 1920 31972 2400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 64 ny 7 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
