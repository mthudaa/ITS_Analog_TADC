magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -16 369 5 403
rect 39 369 77 403
rect 111 369 149 403
rect 183 369 221 403
rect 255 369 293 403
rect 327 369 365 403
rect 399 369 437 403
rect 471 369 509 403
rect 543 369 581 403
rect 615 369 653 403
rect 687 369 725 403
rect 759 369 797 403
rect 831 369 869 403
rect 903 369 941 403
rect 975 369 1013 403
rect 1047 369 1085 403
rect 1119 369 1157 403
rect 1191 369 1229 403
rect 1263 369 1301 403
rect 1335 369 1373 403
rect 1407 369 1445 403
rect 1479 369 1517 403
rect 1551 369 1589 403
rect 1623 369 1661 403
rect 1695 369 1733 403
rect 1767 369 1805 403
rect 1839 369 1877 403
rect 1911 369 1933 403
rect 2005 -17 2023 17
rect 2057 -17 2095 17
rect 2129 -17 2167 17
rect 2201 -17 2239 17
rect 2273 -17 2311 17
rect 2345 -17 2383 17
rect 2417 -17 2455 17
rect 2489 -17 2527 17
rect 2561 -17 2599 17
rect 2633 -17 2671 17
rect 2705 -17 2743 17
rect 2777 -17 2815 17
rect 2849 -17 2887 17
rect 2921 -17 2959 17
rect 2993 -17 3031 17
rect 3065 -17 3083 17
<< viali >>
rect 5 369 39 403
rect 77 369 111 403
rect 149 369 183 403
rect 221 369 255 403
rect 293 369 327 403
rect 365 369 399 403
rect 437 369 471 403
rect 509 369 543 403
rect 581 369 615 403
rect 653 369 687 403
rect 725 369 759 403
rect 797 369 831 403
rect 869 369 903 403
rect 941 369 975 403
rect 1013 369 1047 403
rect 1085 369 1119 403
rect 1157 369 1191 403
rect 1229 369 1263 403
rect 1301 369 1335 403
rect 1373 369 1407 403
rect 1445 369 1479 403
rect 1517 369 1551 403
rect 1589 369 1623 403
rect 1661 369 1695 403
rect 1733 369 1767 403
rect 1805 369 1839 403
rect 1877 369 1911 403
rect 2023 -17 2057 17
rect 2095 -17 2129 17
rect 2167 -17 2201 17
rect 2239 -17 2273 17
rect 2311 -17 2345 17
rect 2383 -17 2417 17
rect 2455 -17 2489 17
rect 2527 -17 2561 17
rect 2599 -17 2633 17
rect 2671 -17 2705 17
rect 2743 -17 2777 17
rect 2815 -17 2849 17
rect 2887 -17 2921 17
rect 2959 -17 2993 17
rect 3031 -17 3065 17
<< metal1 >>
rect -53 403 3119 439
rect -53 369 5 403
rect 39 369 77 403
rect 111 369 149 403
rect 183 369 221 403
rect 255 369 293 403
rect 327 369 365 403
rect 399 369 437 403
rect 471 369 509 403
rect 543 369 581 403
rect 615 369 653 403
rect 687 369 725 403
rect 759 369 797 403
rect 831 369 869 403
rect 903 369 941 403
rect 975 369 1013 403
rect 1047 369 1085 403
rect 1119 369 1157 403
rect 1191 369 1229 403
rect 1263 369 1301 403
rect 1335 369 1373 403
rect 1407 369 1445 403
rect 1479 369 1517 403
rect 1551 369 1589 403
rect 1623 369 1661 403
rect 1695 369 1733 403
rect 1767 369 1805 403
rect 1839 369 1877 403
rect 1911 369 3119 403
rect -53 363 3119 369
rect -53 289 3119 323
rect -53 143 125 243
rect 2941 143 3119 243
rect 166 63 3119 97
rect -53 17 3119 23
rect -53 -17 2023 17
rect 2057 -17 2095 17
rect 2129 -17 2167 17
rect 2201 -17 2239 17
rect 2273 -17 2311 17
rect 2345 -17 2383 17
rect 2417 -17 2455 17
rect 2489 -17 2527 17
rect 2561 -17 2599 17
rect 2633 -17 2671 17
rect 2705 -17 2743 17
rect 2777 -17 2815 17
rect 2849 -17 2887 17
rect 2921 -17 2959 17
rect 2993 -17 3031 17
rect 3065 -17 3119 17
rect -53 -53 3119 -17
use sky130_fd_pr__pfet_01v8_SEQ3W4  XM1
timestamp 1750100919
transform 0 1 958 -1 0 193
box -246 -1011 246 1011
use sky130_fd_pr__nfet_01v8_G4VVNX  XM2
timestamp 1750100919
transform 0 1 2544 -1 0 193
box -236 -565 236 565
<< labels >>
flabel metal1 s -40 400 -29 411 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -40 -18 -29 -7 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -43 302 -34 311 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -37 186 -28 195 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 3096 193 3106 202 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 3096 76 3106 85 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
