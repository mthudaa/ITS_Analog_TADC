magic
tech sky130A
magscale 1 2
timestamp 1757831936
<< metal1 >>
rect 1286 -29150 1296 -29050
rect 1396 -29150 1406 -29050
rect 6088 -29358 6098 -29258
rect 6198 -29358 6208 -29258
rect 10883 -29566 10893 -29466
rect 10993 -29566 11003 -29466
rect 15691 -29774 15701 -29674
rect 15801 -29774 15811 -29674
rect 20494 -29982 20504 -29882
rect 20604 -29982 20614 -29882
rect 25296 -30190 25306 -30090
rect 25406 -30190 25416 -30090
rect 30861 -30398 30871 -30298
rect 30971 -30398 30981 -30298
rect 34900 -30606 34910 -30506
rect 35010 -30606 35020 -30506
rect 39702 -30814 39712 -30714
rect 39812 -30814 39822 -30714
rect 44504 -31022 44514 -30922
rect 44614 -31022 44624 -30922
rect 46856 -36208 46956 -31199
rect 46846 -36308 46856 -36208
rect 46956 -36308 46966 -36208
rect 3228 -36848 3328 -36748
rect 3428 -36848 3528 -36748
rect 8030 -36848 8130 -36748
rect 8230 -36848 8330 -36748
rect 12832 -36848 12932 -36748
rect 13032 -36848 13132 -36748
rect 17634 -36848 17734 -36748
rect 17834 -36848 17934 -36748
rect 22436 -36848 22536 -36748
rect 22636 -36845 22736 -36745
rect 27238 -36848 27338 -36748
rect 27438 -36848 27538 -36748
rect 32040 -36848 32140 -36748
rect 32240 -36848 32340 -36748
rect 36842 -36848 36942 -36748
rect 37042 -36848 37142 -36748
rect 41644 -36848 41744 -36748
rect 41844 -36848 41944 -36748
rect 46446 -36848 46546 -36748
rect 46646 -36848 46746 -36748
<< via1 >>
rect 1296 -29150 1396 -29050
rect 6098 -29358 6198 -29258
rect 10893 -29566 10993 -29466
rect 15701 -29774 15801 -29674
rect 20504 -29982 20604 -29882
rect 25306 -30190 25406 -30090
rect 30871 -30398 30971 -30298
rect 34910 -30606 35010 -30506
rect 39712 -30814 39812 -30714
rect 44514 -31022 44614 -30922
rect 46856 -36308 46956 -36208
<< metal2 >>
rect 1296 -29050 1396 -29040
rect 1296 -31635 1396 -29150
rect 6098 -29258 6198 -29248
rect 6098 -31635 6198 -29358
rect 10893 -29466 10993 -29456
rect 10893 -31635 10993 -29566
rect 15701 -29674 15801 -29664
rect 15701 -31635 15801 -29774
rect 20504 -29882 20604 -29872
rect 20504 -31635 20604 -29982
rect 25306 -30090 25406 -30080
rect 25306 -31635 25406 -30190
rect 30871 -30298 30971 -30288
rect 30871 -31586 30971 -30398
rect 34910 -30506 35010 -30496
rect 34910 -31592 35010 -30606
rect 39712 -30714 39812 -30704
rect 39712 -31614 39812 -30814
rect 44514 -30922 44614 -30912
rect 44514 -31626 44614 -31022
rect 40630 -34722 40730 -33464
rect -748 -35108 -648 -35008
rect -745 -35308 -645 -35208
rect 46856 -36208 46956 -36198
rect -636 -36308 -536 -36208
rect 46756 -36308 46856 -36208
rect 46856 -36318 46956 -36308
<< metal4 >>
rect 895 -17114 999 -17010
use cap_array_10b  cap_array_10b_0
timestamp 1757830127
transform 1 0 63092 0 1 -17818
box -64236 -13426 292 808
use cdac_sw_10b  cdac_sw_10b_0
timestamp 1757827688
transform 0 -1 3588 1 0 -36329
box -519 -43168 5049 4732
<< labels >>
flabel metal1 46646 -36848 46746 -36748 0 FreeSans 320 0 0 0 CF[9]
port 0 nsew
flabel metal1 46446 -36848 46546 -36748 0 FreeSans 320 0 0 0 SW[9]
port 1 nsew
flabel metal1 41644 -36848 41744 -36748 0 FreeSans 320 0 0 0 SW[8]
port 2 nsew
flabel metal1 41844 -36848 41944 -36748 0 FreeSans 320 0 0 0 CF[8]
port 3 nsew
flabel metal1 37042 -36848 37142 -36748 0 FreeSans 320 0 0 0 CF[7]
port 4 nsew
flabel metal1 36842 -36848 36942 -36748 0 FreeSans 320 0 0 0 SW[7]
port 5 nsew
flabel metal1 32240 -36848 32340 -36748 0 FreeSans 320 0 0 0 CF[6]
port 6 nsew
flabel metal1 32040 -36848 32140 -36748 0 FreeSans 320 0 0 0 SW[6]
port 7 nsew
flabel metal1 27238 -36848 27338 -36748 0 FreeSans 320 0 0 0 SW[5]
port 8 nsew
flabel metal1 27438 -36848 27538 -36748 0 FreeSans 320 0 0 0 CF[5]
port 9 nsew
flabel metal1 22636 -36845 22736 -36745 0 FreeSans 320 0 0 0 CF[4]
port 10 nsew
flabel metal1 22436 -36848 22536 -36748 0 FreeSans 320 0 0 0 SW[4]
port 11 nsew
flabel metal1 17634 -36848 17734 -36748 0 FreeSans 320 0 0 0 SW[3]
port 12 nsew
flabel metal1 17834 -36848 17934 -36748 0 FreeSans 320 0 0 0 CF[3]
port 13 nsew
flabel metal1 13032 -36848 13132 -36748 0 FreeSans 320 0 0 0 CF[2]
port 14 nsew
flabel metal1 12832 -36848 12932 -36748 0 FreeSans 320 0 0 0 SW[2]
port 15 nsew
flabel metal1 8030 -36848 8130 -36748 0 FreeSans 320 0 0 0 SW[1]
port 16 nsew
flabel metal1 8230 -36848 8330 -36748 0 FreeSans 320 0 0 0 CF[1]
port 17 nsew
flabel metal1 3428 -36848 3528 -36748 0 FreeSans 320 0 0 0 CF[0]
port 18 nsew
flabel metal1 3228 -36848 3328 -36748 0 FreeSans 320 0 0 0 SW[0]
port 19 nsew
flabel metal2 -748 -35108 -648 -35008 0 FreeSans 320 0 0 0 VSS
port 20 nsew
flabel metal2 -745 -35308 -645 -35208 0 FreeSans 320 0 0 0 VDD
port 21 nsew
flabel metal4 895 -17114 999 -17010 0 FreeSans 320 0 0 0 VC
port 23 nsew
flabel metal2 -636 -36308 -536 -36208 0 FreeSans 320 0 0 0 VCM
port 25 nsew
<< end >>
