magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -109 -362 109 362
<< pmos >>
rect -15 -300 15 300
<< pdiff >>
rect -73 255 -15 300
rect -73 221 -61 255
rect -27 221 -15 255
rect -73 187 -15 221
rect -73 153 -61 187
rect -27 153 -15 187
rect -73 119 -15 153
rect -73 85 -61 119
rect -27 85 -15 119
rect -73 51 -15 85
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -85 -15 -51
rect -73 -119 -61 -85
rect -27 -119 -15 -85
rect -73 -153 -15 -119
rect -73 -187 -61 -153
rect -27 -187 -15 -153
rect -73 -221 -15 -187
rect -73 -255 -61 -221
rect -27 -255 -15 -221
rect -73 -300 -15 -255
rect 15 255 73 300
rect 15 221 27 255
rect 61 221 73 255
rect 15 187 73 221
rect 15 153 27 187
rect 61 153 73 187
rect 15 119 73 153
rect 15 85 27 119
rect 61 85 73 119
rect 15 51 73 85
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -85 73 -51
rect 15 -119 27 -85
rect 61 -119 73 -85
rect 15 -153 73 -119
rect 15 -187 27 -153
rect 61 -187 73 -153
rect 15 -221 73 -187
rect 15 -255 27 -221
rect 61 -255 73 -221
rect 15 -300 73 -255
<< pdiffc >>
rect -61 221 -27 255
rect -61 153 -27 187
rect -61 85 -27 119
rect -61 17 -27 51
rect -61 -51 -27 -17
rect -61 -119 -27 -85
rect -61 -187 -27 -153
rect -61 -255 -27 -221
rect 27 221 61 255
rect 27 153 61 187
rect 27 85 61 119
rect 27 17 61 51
rect 27 -51 61 -17
rect 27 -119 61 -85
rect 27 -187 61 -153
rect 27 -255 61 -221
<< poly >>
rect -15 300 15 326
rect -15 -326 15 -300
<< locali >>
rect -61 269 -27 304
rect -61 197 -27 221
rect -61 125 -27 153
rect -61 53 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -53
rect -61 -153 -27 -125
rect -61 -221 -27 -197
rect -61 -304 -27 -269
rect 27 269 61 304
rect 27 197 61 221
rect 27 125 61 153
rect 27 53 61 85
rect 27 -17 61 17
rect 27 -85 61 -53
rect 27 -153 61 -125
rect 27 -221 61 -197
rect 27 -304 61 -269
<< viali >>
rect -61 255 -27 269
rect -61 235 -27 255
rect -61 187 -27 197
rect -61 163 -27 187
rect -61 119 -27 125
rect -61 91 -27 119
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect -61 -119 -27 -91
rect -61 -125 -27 -119
rect -61 -187 -27 -163
rect -61 -197 -27 -187
rect -61 -255 -27 -235
rect -61 -269 -27 -255
rect 27 255 61 269
rect 27 235 61 255
rect 27 187 61 197
rect 27 163 61 187
rect 27 119 61 125
rect 27 91 61 119
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect 27 -119 61 -91
rect 27 -125 61 -119
rect 27 -187 61 -163
rect 27 -197 61 -187
rect 27 -255 61 -235
rect 27 -269 61 -255
<< metal1 >>
rect -67 269 -21 300
rect -67 235 -61 269
rect -27 235 -21 269
rect -67 197 -21 235
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -163 -21 -125
rect -67 -197 -61 -163
rect -27 -197 -21 -163
rect -67 -235 -21 -197
rect -67 -269 -61 -235
rect -27 -269 -21 -235
rect -67 -300 -21 -269
rect 21 269 67 300
rect 21 235 27 269
rect 61 235 67 269
rect 21 197 67 235
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -163 67 -125
rect 21 -197 27 -163
rect 61 -197 67 -163
rect 21 -235 67 -197
rect 21 -269 27 -235
rect 61 -269 67 -235
rect 21 -300 67 -269
<< end >>
