magic
tech sky130A
magscale 1 2
timestamp 1748279908
<< metal3 >>
rect -17084 11372 -16312 11400
rect -17084 10948 -16396 11372
rect -16332 10948 -16312 11372
rect -17084 10920 -16312 10948
rect -16072 11372 -15300 11400
rect -16072 10948 -15384 11372
rect -15320 10948 -15300 11372
rect -16072 10920 -15300 10948
rect -15060 11372 -14288 11400
rect -15060 10948 -14372 11372
rect -14308 10948 -14288 11372
rect -15060 10920 -14288 10948
rect -14048 11372 -13276 11400
rect -14048 10948 -13360 11372
rect -13296 10948 -13276 11372
rect -14048 10920 -13276 10948
rect -13036 11372 -12264 11400
rect -13036 10948 -12348 11372
rect -12284 10948 -12264 11372
rect -13036 10920 -12264 10948
rect -12024 11372 -11252 11400
rect -12024 10948 -11336 11372
rect -11272 10948 -11252 11372
rect -12024 10920 -11252 10948
rect -11012 11372 -10240 11400
rect -11012 10948 -10324 11372
rect -10260 10948 -10240 11372
rect -11012 10920 -10240 10948
rect -10000 11372 -9228 11400
rect -10000 10948 -9312 11372
rect -9248 10948 -9228 11372
rect -10000 10920 -9228 10948
rect -8988 11372 -8216 11400
rect -8988 10948 -8300 11372
rect -8236 10948 -8216 11372
rect -8988 10920 -8216 10948
rect -7976 11372 -7204 11400
rect -7976 10948 -7288 11372
rect -7224 10948 -7204 11372
rect -7976 10920 -7204 10948
rect -6964 11372 -6192 11400
rect -6964 10948 -6276 11372
rect -6212 10948 -6192 11372
rect -6964 10920 -6192 10948
rect -5952 11372 -5180 11400
rect -5952 10948 -5264 11372
rect -5200 10948 -5180 11372
rect -5952 10920 -5180 10948
rect -4940 11372 -4168 11400
rect -4940 10948 -4252 11372
rect -4188 10948 -4168 11372
rect -4940 10920 -4168 10948
rect -3928 11372 -3156 11400
rect -3928 10948 -3240 11372
rect -3176 10948 -3156 11372
rect -3928 10920 -3156 10948
rect -2916 11372 -2144 11400
rect -2916 10948 -2228 11372
rect -2164 10948 -2144 11372
rect -2916 10920 -2144 10948
rect -1904 11372 -1132 11400
rect -1904 10948 -1216 11372
rect -1152 10948 -1132 11372
rect -1904 10920 -1132 10948
rect -892 11372 -120 11400
rect -892 10948 -204 11372
rect -140 10948 -120 11372
rect -892 10920 -120 10948
rect 120 11372 892 11400
rect 120 10948 808 11372
rect 872 10948 892 11372
rect 120 10920 892 10948
rect 1132 11372 1904 11400
rect 1132 10948 1820 11372
rect 1884 10948 1904 11372
rect 1132 10920 1904 10948
rect 2144 11372 2916 11400
rect 2144 10948 2832 11372
rect 2896 10948 2916 11372
rect 2144 10920 2916 10948
rect 3156 11372 3928 11400
rect 3156 10948 3844 11372
rect 3908 10948 3928 11372
rect 3156 10920 3928 10948
rect 4168 11372 4940 11400
rect 4168 10948 4856 11372
rect 4920 10948 4940 11372
rect 4168 10920 4940 10948
rect 5180 11372 5952 11400
rect 5180 10948 5868 11372
rect 5932 10948 5952 11372
rect 5180 10920 5952 10948
rect 6192 11372 6964 11400
rect 6192 10948 6880 11372
rect 6944 10948 6964 11372
rect 6192 10920 6964 10948
rect 7204 11372 7976 11400
rect 7204 10948 7892 11372
rect 7956 10948 7976 11372
rect 7204 10920 7976 10948
rect 8216 11372 8988 11400
rect 8216 10948 8904 11372
rect 8968 10948 8988 11372
rect 8216 10920 8988 10948
rect 9228 11372 10000 11400
rect 9228 10948 9916 11372
rect 9980 10948 10000 11372
rect 9228 10920 10000 10948
rect 10240 11372 11012 11400
rect 10240 10948 10928 11372
rect 10992 10948 11012 11372
rect 10240 10920 11012 10948
rect 11252 11372 12024 11400
rect 11252 10948 11940 11372
rect 12004 10948 12024 11372
rect 11252 10920 12024 10948
rect 12264 11372 13036 11400
rect 12264 10948 12952 11372
rect 13016 10948 13036 11372
rect 12264 10920 13036 10948
rect 13276 11372 14048 11400
rect 13276 10948 13964 11372
rect 14028 10948 14048 11372
rect 13276 10920 14048 10948
rect 14288 11372 15060 11400
rect 14288 10948 14976 11372
rect 15040 10948 15060 11372
rect 14288 10920 15060 10948
rect 15300 11372 16072 11400
rect 15300 10948 15988 11372
rect 16052 10948 16072 11372
rect 15300 10920 16072 10948
rect 16312 11372 17084 11400
rect 16312 10948 17000 11372
rect 17064 10948 17084 11372
rect 16312 10920 17084 10948
rect -17084 10652 -16312 10680
rect -17084 10228 -16396 10652
rect -16332 10228 -16312 10652
rect -17084 10200 -16312 10228
rect -16072 10652 -15300 10680
rect -16072 10228 -15384 10652
rect -15320 10228 -15300 10652
rect -16072 10200 -15300 10228
rect -15060 10652 -14288 10680
rect -15060 10228 -14372 10652
rect -14308 10228 -14288 10652
rect -15060 10200 -14288 10228
rect -14048 10652 -13276 10680
rect -14048 10228 -13360 10652
rect -13296 10228 -13276 10652
rect -14048 10200 -13276 10228
rect -13036 10652 -12264 10680
rect -13036 10228 -12348 10652
rect -12284 10228 -12264 10652
rect -13036 10200 -12264 10228
rect -12024 10652 -11252 10680
rect -12024 10228 -11336 10652
rect -11272 10228 -11252 10652
rect -12024 10200 -11252 10228
rect -11012 10652 -10240 10680
rect -11012 10228 -10324 10652
rect -10260 10228 -10240 10652
rect -11012 10200 -10240 10228
rect -10000 10652 -9228 10680
rect -10000 10228 -9312 10652
rect -9248 10228 -9228 10652
rect -10000 10200 -9228 10228
rect -8988 10652 -8216 10680
rect -8988 10228 -8300 10652
rect -8236 10228 -8216 10652
rect -8988 10200 -8216 10228
rect -7976 10652 -7204 10680
rect -7976 10228 -7288 10652
rect -7224 10228 -7204 10652
rect -7976 10200 -7204 10228
rect -6964 10652 -6192 10680
rect -6964 10228 -6276 10652
rect -6212 10228 -6192 10652
rect -6964 10200 -6192 10228
rect -5952 10652 -5180 10680
rect -5952 10228 -5264 10652
rect -5200 10228 -5180 10652
rect -5952 10200 -5180 10228
rect -4940 10652 -4168 10680
rect -4940 10228 -4252 10652
rect -4188 10228 -4168 10652
rect -4940 10200 -4168 10228
rect -3928 10652 -3156 10680
rect -3928 10228 -3240 10652
rect -3176 10228 -3156 10652
rect -3928 10200 -3156 10228
rect -2916 10652 -2144 10680
rect -2916 10228 -2228 10652
rect -2164 10228 -2144 10652
rect -2916 10200 -2144 10228
rect -1904 10652 -1132 10680
rect -1904 10228 -1216 10652
rect -1152 10228 -1132 10652
rect -1904 10200 -1132 10228
rect -892 10652 -120 10680
rect -892 10228 -204 10652
rect -140 10228 -120 10652
rect -892 10200 -120 10228
rect 120 10652 892 10680
rect 120 10228 808 10652
rect 872 10228 892 10652
rect 120 10200 892 10228
rect 1132 10652 1904 10680
rect 1132 10228 1820 10652
rect 1884 10228 1904 10652
rect 1132 10200 1904 10228
rect 2144 10652 2916 10680
rect 2144 10228 2832 10652
rect 2896 10228 2916 10652
rect 2144 10200 2916 10228
rect 3156 10652 3928 10680
rect 3156 10228 3844 10652
rect 3908 10228 3928 10652
rect 3156 10200 3928 10228
rect 4168 10652 4940 10680
rect 4168 10228 4856 10652
rect 4920 10228 4940 10652
rect 4168 10200 4940 10228
rect 5180 10652 5952 10680
rect 5180 10228 5868 10652
rect 5932 10228 5952 10652
rect 5180 10200 5952 10228
rect 6192 10652 6964 10680
rect 6192 10228 6880 10652
rect 6944 10228 6964 10652
rect 6192 10200 6964 10228
rect 7204 10652 7976 10680
rect 7204 10228 7892 10652
rect 7956 10228 7976 10652
rect 7204 10200 7976 10228
rect 8216 10652 8988 10680
rect 8216 10228 8904 10652
rect 8968 10228 8988 10652
rect 8216 10200 8988 10228
rect 9228 10652 10000 10680
rect 9228 10228 9916 10652
rect 9980 10228 10000 10652
rect 9228 10200 10000 10228
rect 10240 10652 11012 10680
rect 10240 10228 10928 10652
rect 10992 10228 11012 10652
rect 10240 10200 11012 10228
rect 11252 10652 12024 10680
rect 11252 10228 11940 10652
rect 12004 10228 12024 10652
rect 11252 10200 12024 10228
rect 12264 10652 13036 10680
rect 12264 10228 12952 10652
rect 13016 10228 13036 10652
rect 12264 10200 13036 10228
rect 13276 10652 14048 10680
rect 13276 10228 13964 10652
rect 14028 10228 14048 10652
rect 13276 10200 14048 10228
rect 14288 10652 15060 10680
rect 14288 10228 14976 10652
rect 15040 10228 15060 10652
rect 14288 10200 15060 10228
rect 15300 10652 16072 10680
rect 15300 10228 15988 10652
rect 16052 10228 16072 10652
rect 15300 10200 16072 10228
rect 16312 10652 17084 10680
rect 16312 10228 17000 10652
rect 17064 10228 17084 10652
rect 16312 10200 17084 10228
rect -17084 9932 -16312 9960
rect -17084 9508 -16396 9932
rect -16332 9508 -16312 9932
rect -17084 9480 -16312 9508
rect -16072 9932 -15300 9960
rect -16072 9508 -15384 9932
rect -15320 9508 -15300 9932
rect -16072 9480 -15300 9508
rect -15060 9932 -14288 9960
rect -15060 9508 -14372 9932
rect -14308 9508 -14288 9932
rect -15060 9480 -14288 9508
rect -14048 9932 -13276 9960
rect -14048 9508 -13360 9932
rect -13296 9508 -13276 9932
rect -14048 9480 -13276 9508
rect -13036 9932 -12264 9960
rect -13036 9508 -12348 9932
rect -12284 9508 -12264 9932
rect -13036 9480 -12264 9508
rect -12024 9932 -11252 9960
rect -12024 9508 -11336 9932
rect -11272 9508 -11252 9932
rect -12024 9480 -11252 9508
rect -11012 9932 -10240 9960
rect -11012 9508 -10324 9932
rect -10260 9508 -10240 9932
rect -11012 9480 -10240 9508
rect -10000 9932 -9228 9960
rect -10000 9508 -9312 9932
rect -9248 9508 -9228 9932
rect -10000 9480 -9228 9508
rect -8988 9932 -8216 9960
rect -8988 9508 -8300 9932
rect -8236 9508 -8216 9932
rect -8988 9480 -8216 9508
rect -7976 9932 -7204 9960
rect -7976 9508 -7288 9932
rect -7224 9508 -7204 9932
rect -7976 9480 -7204 9508
rect -6964 9932 -6192 9960
rect -6964 9508 -6276 9932
rect -6212 9508 -6192 9932
rect -6964 9480 -6192 9508
rect -5952 9932 -5180 9960
rect -5952 9508 -5264 9932
rect -5200 9508 -5180 9932
rect -5952 9480 -5180 9508
rect -4940 9932 -4168 9960
rect -4940 9508 -4252 9932
rect -4188 9508 -4168 9932
rect -4940 9480 -4168 9508
rect -3928 9932 -3156 9960
rect -3928 9508 -3240 9932
rect -3176 9508 -3156 9932
rect -3928 9480 -3156 9508
rect -2916 9932 -2144 9960
rect -2916 9508 -2228 9932
rect -2164 9508 -2144 9932
rect -2916 9480 -2144 9508
rect -1904 9932 -1132 9960
rect -1904 9508 -1216 9932
rect -1152 9508 -1132 9932
rect -1904 9480 -1132 9508
rect -892 9932 -120 9960
rect -892 9508 -204 9932
rect -140 9508 -120 9932
rect -892 9480 -120 9508
rect 120 9932 892 9960
rect 120 9508 808 9932
rect 872 9508 892 9932
rect 120 9480 892 9508
rect 1132 9932 1904 9960
rect 1132 9508 1820 9932
rect 1884 9508 1904 9932
rect 1132 9480 1904 9508
rect 2144 9932 2916 9960
rect 2144 9508 2832 9932
rect 2896 9508 2916 9932
rect 2144 9480 2916 9508
rect 3156 9932 3928 9960
rect 3156 9508 3844 9932
rect 3908 9508 3928 9932
rect 3156 9480 3928 9508
rect 4168 9932 4940 9960
rect 4168 9508 4856 9932
rect 4920 9508 4940 9932
rect 4168 9480 4940 9508
rect 5180 9932 5952 9960
rect 5180 9508 5868 9932
rect 5932 9508 5952 9932
rect 5180 9480 5952 9508
rect 6192 9932 6964 9960
rect 6192 9508 6880 9932
rect 6944 9508 6964 9932
rect 6192 9480 6964 9508
rect 7204 9932 7976 9960
rect 7204 9508 7892 9932
rect 7956 9508 7976 9932
rect 7204 9480 7976 9508
rect 8216 9932 8988 9960
rect 8216 9508 8904 9932
rect 8968 9508 8988 9932
rect 8216 9480 8988 9508
rect 9228 9932 10000 9960
rect 9228 9508 9916 9932
rect 9980 9508 10000 9932
rect 9228 9480 10000 9508
rect 10240 9932 11012 9960
rect 10240 9508 10928 9932
rect 10992 9508 11012 9932
rect 10240 9480 11012 9508
rect 11252 9932 12024 9960
rect 11252 9508 11940 9932
rect 12004 9508 12024 9932
rect 11252 9480 12024 9508
rect 12264 9932 13036 9960
rect 12264 9508 12952 9932
rect 13016 9508 13036 9932
rect 12264 9480 13036 9508
rect 13276 9932 14048 9960
rect 13276 9508 13964 9932
rect 14028 9508 14048 9932
rect 13276 9480 14048 9508
rect 14288 9932 15060 9960
rect 14288 9508 14976 9932
rect 15040 9508 15060 9932
rect 14288 9480 15060 9508
rect 15300 9932 16072 9960
rect 15300 9508 15988 9932
rect 16052 9508 16072 9932
rect 15300 9480 16072 9508
rect 16312 9932 17084 9960
rect 16312 9508 17000 9932
rect 17064 9508 17084 9932
rect 16312 9480 17084 9508
rect -17084 9212 -16312 9240
rect -17084 8788 -16396 9212
rect -16332 8788 -16312 9212
rect -17084 8760 -16312 8788
rect -16072 9212 -15300 9240
rect -16072 8788 -15384 9212
rect -15320 8788 -15300 9212
rect -16072 8760 -15300 8788
rect -15060 9212 -14288 9240
rect -15060 8788 -14372 9212
rect -14308 8788 -14288 9212
rect -15060 8760 -14288 8788
rect -14048 9212 -13276 9240
rect -14048 8788 -13360 9212
rect -13296 8788 -13276 9212
rect -14048 8760 -13276 8788
rect -13036 9212 -12264 9240
rect -13036 8788 -12348 9212
rect -12284 8788 -12264 9212
rect -13036 8760 -12264 8788
rect -12024 9212 -11252 9240
rect -12024 8788 -11336 9212
rect -11272 8788 -11252 9212
rect -12024 8760 -11252 8788
rect -11012 9212 -10240 9240
rect -11012 8788 -10324 9212
rect -10260 8788 -10240 9212
rect -11012 8760 -10240 8788
rect -10000 9212 -9228 9240
rect -10000 8788 -9312 9212
rect -9248 8788 -9228 9212
rect -10000 8760 -9228 8788
rect -8988 9212 -8216 9240
rect -8988 8788 -8300 9212
rect -8236 8788 -8216 9212
rect -8988 8760 -8216 8788
rect -7976 9212 -7204 9240
rect -7976 8788 -7288 9212
rect -7224 8788 -7204 9212
rect -7976 8760 -7204 8788
rect -6964 9212 -6192 9240
rect -6964 8788 -6276 9212
rect -6212 8788 -6192 9212
rect -6964 8760 -6192 8788
rect -5952 9212 -5180 9240
rect -5952 8788 -5264 9212
rect -5200 8788 -5180 9212
rect -5952 8760 -5180 8788
rect -4940 9212 -4168 9240
rect -4940 8788 -4252 9212
rect -4188 8788 -4168 9212
rect -4940 8760 -4168 8788
rect -3928 9212 -3156 9240
rect -3928 8788 -3240 9212
rect -3176 8788 -3156 9212
rect -3928 8760 -3156 8788
rect -2916 9212 -2144 9240
rect -2916 8788 -2228 9212
rect -2164 8788 -2144 9212
rect -2916 8760 -2144 8788
rect -1904 9212 -1132 9240
rect -1904 8788 -1216 9212
rect -1152 8788 -1132 9212
rect -1904 8760 -1132 8788
rect -892 9212 -120 9240
rect -892 8788 -204 9212
rect -140 8788 -120 9212
rect -892 8760 -120 8788
rect 120 9212 892 9240
rect 120 8788 808 9212
rect 872 8788 892 9212
rect 120 8760 892 8788
rect 1132 9212 1904 9240
rect 1132 8788 1820 9212
rect 1884 8788 1904 9212
rect 1132 8760 1904 8788
rect 2144 9212 2916 9240
rect 2144 8788 2832 9212
rect 2896 8788 2916 9212
rect 2144 8760 2916 8788
rect 3156 9212 3928 9240
rect 3156 8788 3844 9212
rect 3908 8788 3928 9212
rect 3156 8760 3928 8788
rect 4168 9212 4940 9240
rect 4168 8788 4856 9212
rect 4920 8788 4940 9212
rect 4168 8760 4940 8788
rect 5180 9212 5952 9240
rect 5180 8788 5868 9212
rect 5932 8788 5952 9212
rect 5180 8760 5952 8788
rect 6192 9212 6964 9240
rect 6192 8788 6880 9212
rect 6944 8788 6964 9212
rect 6192 8760 6964 8788
rect 7204 9212 7976 9240
rect 7204 8788 7892 9212
rect 7956 8788 7976 9212
rect 7204 8760 7976 8788
rect 8216 9212 8988 9240
rect 8216 8788 8904 9212
rect 8968 8788 8988 9212
rect 8216 8760 8988 8788
rect 9228 9212 10000 9240
rect 9228 8788 9916 9212
rect 9980 8788 10000 9212
rect 9228 8760 10000 8788
rect 10240 9212 11012 9240
rect 10240 8788 10928 9212
rect 10992 8788 11012 9212
rect 10240 8760 11012 8788
rect 11252 9212 12024 9240
rect 11252 8788 11940 9212
rect 12004 8788 12024 9212
rect 11252 8760 12024 8788
rect 12264 9212 13036 9240
rect 12264 8788 12952 9212
rect 13016 8788 13036 9212
rect 12264 8760 13036 8788
rect 13276 9212 14048 9240
rect 13276 8788 13964 9212
rect 14028 8788 14048 9212
rect 13276 8760 14048 8788
rect 14288 9212 15060 9240
rect 14288 8788 14976 9212
rect 15040 8788 15060 9212
rect 14288 8760 15060 8788
rect 15300 9212 16072 9240
rect 15300 8788 15988 9212
rect 16052 8788 16072 9212
rect 15300 8760 16072 8788
rect 16312 9212 17084 9240
rect 16312 8788 17000 9212
rect 17064 8788 17084 9212
rect 16312 8760 17084 8788
rect -17084 8492 -16312 8520
rect -17084 8068 -16396 8492
rect -16332 8068 -16312 8492
rect -17084 8040 -16312 8068
rect -16072 8492 -15300 8520
rect -16072 8068 -15384 8492
rect -15320 8068 -15300 8492
rect -16072 8040 -15300 8068
rect -15060 8492 -14288 8520
rect -15060 8068 -14372 8492
rect -14308 8068 -14288 8492
rect -15060 8040 -14288 8068
rect -14048 8492 -13276 8520
rect -14048 8068 -13360 8492
rect -13296 8068 -13276 8492
rect -14048 8040 -13276 8068
rect -13036 8492 -12264 8520
rect -13036 8068 -12348 8492
rect -12284 8068 -12264 8492
rect -13036 8040 -12264 8068
rect -12024 8492 -11252 8520
rect -12024 8068 -11336 8492
rect -11272 8068 -11252 8492
rect -12024 8040 -11252 8068
rect -11012 8492 -10240 8520
rect -11012 8068 -10324 8492
rect -10260 8068 -10240 8492
rect -11012 8040 -10240 8068
rect -10000 8492 -9228 8520
rect -10000 8068 -9312 8492
rect -9248 8068 -9228 8492
rect -10000 8040 -9228 8068
rect -8988 8492 -8216 8520
rect -8988 8068 -8300 8492
rect -8236 8068 -8216 8492
rect -8988 8040 -8216 8068
rect -7976 8492 -7204 8520
rect -7976 8068 -7288 8492
rect -7224 8068 -7204 8492
rect -7976 8040 -7204 8068
rect -6964 8492 -6192 8520
rect -6964 8068 -6276 8492
rect -6212 8068 -6192 8492
rect -6964 8040 -6192 8068
rect -5952 8492 -5180 8520
rect -5952 8068 -5264 8492
rect -5200 8068 -5180 8492
rect -5952 8040 -5180 8068
rect -4940 8492 -4168 8520
rect -4940 8068 -4252 8492
rect -4188 8068 -4168 8492
rect -4940 8040 -4168 8068
rect -3928 8492 -3156 8520
rect -3928 8068 -3240 8492
rect -3176 8068 -3156 8492
rect -3928 8040 -3156 8068
rect -2916 8492 -2144 8520
rect -2916 8068 -2228 8492
rect -2164 8068 -2144 8492
rect -2916 8040 -2144 8068
rect -1904 8492 -1132 8520
rect -1904 8068 -1216 8492
rect -1152 8068 -1132 8492
rect -1904 8040 -1132 8068
rect -892 8492 -120 8520
rect -892 8068 -204 8492
rect -140 8068 -120 8492
rect -892 8040 -120 8068
rect 120 8492 892 8520
rect 120 8068 808 8492
rect 872 8068 892 8492
rect 120 8040 892 8068
rect 1132 8492 1904 8520
rect 1132 8068 1820 8492
rect 1884 8068 1904 8492
rect 1132 8040 1904 8068
rect 2144 8492 2916 8520
rect 2144 8068 2832 8492
rect 2896 8068 2916 8492
rect 2144 8040 2916 8068
rect 3156 8492 3928 8520
rect 3156 8068 3844 8492
rect 3908 8068 3928 8492
rect 3156 8040 3928 8068
rect 4168 8492 4940 8520
rect 4168 8068 4856 8492
rect 4920 8068 4940 8492
rect 4168 8040 4940 8068
rect 5180 8492 5952 8520
rect 5180 8068 5868 8492
rect 5932 8068 5952 8492
rect 5180 8040 5952 8068
rect 6192 8492 6964 8520
rect 6192 8068 6880 8492
rect 6944 8068 6964 8492
rect 6192 8040 6964 8068
rect 7204 8492 7976 8520
rect 7204 8068 7892 8492
rect 7956 8068 7976 8492
rect 7204 8040 7976 8068
rect 8216 8492 8988 8520
rect 8216 8068 8904 8492
rect 8968 8068 8988 8492
rect 8216 8040 8988 8068
rect 9228 8492 10000 8520
rect 9228 8068 9916 8492
rect 9980 8068 10000 8492
rect 9228 8040 10000 8068
rect 10240 8492 11012 8520
rect 10240 8068 10928 8492
rect 10992 8068 11012 8492
rect 10240 8040 11012 8068
rect 11252 8492 12024 8520
rect 11252 8068 11940 8492
rect 12004 8068 12024 8492
rect 11252 8040 12024 8068
rect 12264 8492 13036 8520
rect 12264 8068 12952 8492
rect 13016 8068 13036 8492
rect 12264 8040 13036 8068
rect 13276 8492 14048 8520
rect 13276 8068 13964 8492
rect 14028 8068 14048 8492
rect 13276 8040 14048 8068
rect 14288 8492 15060 8520
rect 14288 8068 14976 8492
rect 15040 8068 15060 8492
rect 14288 8040 15060 8068
rect 15300 8492 16072 8520
rect 15300 8068 15988 8492
rect 16052 8068 16072 8492
rect 15300 8040 16072 8068
rect 16312 8492 17084 8520
rect 16312 8068 17000 8492
rect 17064 8068 17084 8492
rect 16312 8040 17084 8068
rect -17084 7772 -16312 7800
rect -17084 7348 -16396 7772
rect -16332 7348 -16312 7772
rect -17084 7320 -16312 7348
rect -16072 7772 -15300 7800
rect -16072 7348 -15384 7772
rect -15320 7348 -15300 7772
rect -16072 7320 -15300 7348
rect -15060 7772 -14288 7800
rect -15060 7348 -14372 7772
rect -14308 7348 -14288 7772
rect -15060 7320 -14288 7348
rect -14048 7772 -13276 7800
rect -14048 7348 -13360 7772
rect -13296 7348 -13276 7772
rect -14048 7320 -13276 7348
rect -13036 7772 -12264 7800
rect -13036 7348 -12348 7772
rect -12284 7348 -12264 7772
rect -13036 7320 -12264 7348
rect -12024 7772 -11252 7800
rect -12024 7348 -11336 7772
rect -11272 7348 -11252 7772
rect -12024 7320 -11252 7348
rect -11012 7772 -10240 7800
rect -11012 7348 -10324 7772
rect -10260 7348 -10240 7772
rect -11012 7320 -10240 7348
rect -10000 7772 -9228 7800
rect -10000 7348 -9312 7772
rect -9248 7348 -9228 7772
rect -10000 7320 -9228 7348
rect -8988 7772 -8216 7800
rect -8988 7348 -8300 7772
rect -8236 7348 -8216 7772
rect -8988 7320 -8216 7348
rect -7976 7772 -7204 7800
rect -7976 7348 -7288 7772
rect -7224 7348 -7204 7772
rect -7976 7320 -7204 7348
rect -6964 7772 -6192 7800
rect -6964 7348 -6276 7772
rect -6212 7348 -6192 7772
rect -6964 7320 -6192 7348
rect -5952 7772 -5180 7800
rect -5952 7348 -5264 7772
rect -5200 7348 -5180 7772
rect -5952 7320 -5180 7348
rect -4940 7772 -4168 7800
rect -4940 7348 -4252 7772
rect -4188 7348 -4168 7772
rect -4940 7320 -4168 7348
rect -3928 7772 -3156 7800
rect -3928 7348 -3240 7772
rect -3176 7348 -3156 7772
rect -3928 7320 -3156 7348
rect -2916 7772 -2144 7800
rect -2916 7348 -2228 7772
rect -2164 7348 -2144 7772
rect -2916 7320 -2144 7348
rect -1904 7772 -1132 7800
rect -1904 7348 -1216 7772
rect -1152 7348 -1132 7772
rect -1904 7320 -1132 7348
rect -892 7772 -120 7800
rect -892 7348 -204 7772
rect -140 7348 -120 7772
rect -892 7320 -120 7348
rect 120 7772 892 7800
rect 120 7348 808 7772
rect 872 7348 892 7772
rect 120 7320 892 7348
rect 1132 7772 1904 7800
rect 1132 7348 1820 7772
rect 1884 7348 1904 7772
rect 1132 7320 1904 7348
rect 2144 7772 2916 7800
rect 2144 7348 2832 7772
rect 2896 7348 2916 7772
rect 2144 7320 2916 7348
rect 3156 7772 3928 7800
rect 3156 7348 3844 7772
rect 3908 7348 3928 7772
rect 3156 7320 3928 7348
rect 4168 7772 4940 7800
rect 4168 7348 4856 7772
rect 4920 7348 4940 7772
rect 4168 7320 4940 7348
rect 5180 7772 5952 7800
rect 5180 7348 5868 7772
rect 5932 7348 5952 7772
rect 5180 7320 5952 7348
rect 6192 7772 6964 7800
rect 6192 7348 6880 7772
rect 6944 7348 6964 7772
rect 6192 7320 6964 7348
rect 7204 7772 7976 7800
rect 7204 7348 7892 7772
rect 7956 7348 7976 7772
rect 7204 7320 7976 7348
rect 8216 7772 8988 7800
rect 8216 7348 8904 7772
rect 8968 7348 8988 7772
rect 8216 7320 8988 7348
rect 9228 7772 10000 7800
rect 9228 7348 9916 7772
rect 9980 7348 10000 7772
rect 9228 7320 10000 7348
rect 10240 7772 11012 7800
rect 10240 7348 10928 7772
rect 10992 7348 11012 7772
rect 10240 7320 11012 7348
rect 11252 7772 12024 7800
rect 11252 7348 11940 7772
rect 12004 7348 12024 7772
rect 11252 7320 12024 7348
rect 12264 7772 13036 7800
rect 12264 7348 12952 7772
rect 13016 7348 13036 7772
rect 12264 7320 13036 7348
rect 13276 7772 14048 7800
rect 13276 7348 13964 7772
rect 14028 7348 14048 7772
rect 13276 7320 14048 7348
rect 14288 7772 15060 7800
rect 14288 7348 14976 7772
rect 15040 7348 15060 7772
rect 14288 7320 15060 7348
rect 15300 7772 16072 7800
rect 15300 7348 15988 7772
rect 16052 7348 16072 7772
rect 15300 7320 16072 7348
rect 16312 7772 17084 7800
rect 16312 7348 17000 7772
rect 17064 7348 17084 7772
rect 16312 7320 17084 7348
rect -17084 7052 -16312 7080
rect -17084 6628 -16396 7052
rect -16332 6628 -16312 7052
rect -17084 6600 -16312 6628
rect -16072 7052 -15300 7080
rect -16072 6628 -15384 7052
rect -15320 6628 -15300 7052
rect -16072 6600 -15300 6628
rect -15060 7052 -14288 7080
rect -15060 6628 -14372 7052
rect -14308 6628 -14288 7052
rect -15060 6600 -14288 6628
rect -14048 7052 -13276 7080
rect -14048 6628 -13360 7052
rect -13296 6628 -13276 7052
rect -14048 6600 -13276 6628
rect -13036 7052 -12264 7080
rect -13036 6628 -12348 7052
rect -12284 6628 -12264 7052
rect -13036 6600 -12264 6628
rect -12024 7052 -11252 7080
rect -12024 6628 -11336 7052
rect -11272 6628 -11252 7052
rect -12024 6600 -11252 6628
rect -11012 7052 -10240 7080
rect -11012 6628 -10324 7052
rect -10260 6628 -10240 7052
rect -11012 6600 -10240 6628
rect -10000 7052 -9228 7080
rect -10000 6628 -9312 7052
rect -9248 6628 -9228 7052
rect -10000 6600 -9228 6628
rect -8988 7052 -8216 7080
rect -8988 6628 -8300 7052
rect -8236 6628 -8216 7052
rect -8988 6600 -8216 6628
rect -7976 7052 -7204 7080
rect -7976 6628 -7288 7052
rect -7224 6628 -7204 7052
rect -7976 6600 -7204 6628
rect -6964 7052 -6192 7080
rect -6964 6628 -6276 7052
rect -6212 6628 -6192 7052
rect -6964 6600 -6192 6628
rect -5952 7052 -5180 7080
rect -5952 6628 -5264 7052
rect -5200 6628 -5180 7052
rect -5952 6600 -5180 6628
rect -4940 7052 -4168 7080
rect -4940 6628 -4252 7052
rect -4188 6628 -4168 7052
rect -4940 6600 -4168 6628
rect -3928 7052 -3156 7080
rect -3928 6628 -3240 7052
rect -3176 6628 -3156 7052
rect -3928 6600 -3156 6628
rect -2916 7052 -2144 7080
rect -2916 6628 -2228 7052
rect -2164 6628 -2144 7052
rect -2916 6600 -2144 6628
rect -1904 7052 -1132 7080
rect -1904 6628 -1216 7052
rect -1152 6628 -1132 7052
rect -1904 6600 -1132 6628
rect -892 7052 -120 7080
rect -892 6628 -204 7052
rect -140 6628 -120 7052
rect -892 6600 -120 6628
rect 120 7052 892 7080
rect 120 6628 808 7052
rect 872 6628 892 7052
rect 120 6600 892 6628
rect 1132 7052 1904 7080
rect 1132 6628 1820 7052
rect 1884 6628 1904 7052
rect 1132 6600 1904 6628
rect 2144 7052 2916 7080
rect 2144 6628 2832 7052
rect 2896 6628 2916 7052
rect 2144 6600 2916 6628
rect 3156 7052 3928 7080
rect 3156 6628 3844 7052
rect 3908 6628 3928 7052
rect 3156 6600 3928 6628
rect 4168 7052 4940 7080
rect 4168 6628 4856 7052
rect 4920 6628 4940 7052
rect 4168 6600 4940 6628
rect 5180 7052 5952 7080
rect 5180 6628 5868 7052
rect 5932 6628 5952 7052
rect 5180 6600 5952 6628
rect 6192 7052 6964 7080
rect 6192 6628 6880 7052
rect 6944 6628 6964 7052
rect 6192 6600 6964 6628
rect 7204 7052 7976 7080
rect 7204 6628 7892 7052
rect 7956 6628 7976 7052
rect 7204 6600 7976 6628
rect 8216 7052 8988 7080
rect 8216 6628 8904 7052
rect 8968 6628 8988 7052
rect 8216 6600 8988 6628
rect 9228 7052 10000 7080
rect 9228 6628 9916 7052
rect 9980 6628 10000 7052
rect 9228 6600 10000 6628
rect 10240 7052 11012 7080
rect 10240 6628 10928 7052
rect 10992 6628 11012 7052
rect 10240 6600 11012 6628
rect 11252 7052 12024 7080
rect 11252 6628 11940 7052
rect 12004 6628 12024 7052
rect 11252 6600 12024 6628
rect 12264 7052 13036 7080
rect 12264 6628 12952 7052
rect 13016 6628 13036 7052
rect 12264 6600 13036 6628
rect 13276 7052 14048 7080
rect 13276 6628 13964 7052
rect 14028 6628 14048 7052
rect 13276 6600 14048 6628
rect 14288 7052 15060 7080
rect 14288 6628 14976 7052
rect 15040 6628 15060 7052
rect 14288 6600 15060 6628
rect 15300 7052 16072 7080
rect 15300 6628 15988 7052
rect 16052 6628 16072 7052
rect 15300 6600 16072 6628
rect 16312 7052 17084 7080
rect 16312 6628 17000 7052
rect 17064 6628 17084 7052
rect 16312 6600 17084 6628
rect -17084 6332 -16312 6360
rect -17084 5908 -16396 6332
rect -16332 5908 -16312 6332
rect -17084 5880 -16312 5908
rect -16072 6332 -15300 6360
rect -16072 5908 -15384 6332
rect -15320 5908 -15300 6332
rect -16072 5880 -15300 5908
rect -15060 6332 -14288 6360
rect -15060 5908 -14372 6332
rect -14308 5908 -14288 6332
rect -15060 5880 -14288 5908
rect -14048 6332 -13276 6360
rect -14048 5908 -13360 6332
rect -13296 5908 -13276 6332
rect -14048 5880 -13276 5908
rect -13036 6332 -12264 6360
rect -13036 5908 -12348 6332
rect -12284 5908 -12264 6332
rect -13036 5880 -12264 5908
rect -12024 6332 -11252 6360
rect -12024 5908 -11336 6332
rect -11272 5908 -11252 6332
rect -12024 5880 -11252 5908
rect -11012 6332 -10240 6360
rect -11012 5908 -10324 6332
rect -10260 5908 -10240 6332
rect -11012 5880 -10240 5908
rect -10000 6332 -9228 6360
rect -10000 5908 -9312 6332
rect -9248 5908 -9228 6332
rect -10000 5880 -9228 5908
rect -8988 6332 -8216 6360
rect -8988 5908 -8300 6332
rect -8236 5908 -8216 6332
rect -8988 5880 -8216 5908
rect -7976 6332 -7204 6360
rect -7976 5908 -7288 6332
rect -7224 5908 -7204 6332
rect -7976 5880 -7204 5908
rect -6964 6332 -6192 6360
rect -6964 5908 -6276 6332
rect -6212 5908 -6192 6332
rect -6964 5880 -6192 5908
rect -5952 6332 -5180 6360
rect -5952 5908 -5264 6332
rect -5200 5908 -5180 6332
rect -5952 5880 -5180 5908
rect -4940 6332 -4168 6360
rect -4940 5908 -4252 6332
rect -4188 5908 -4168 6332
rect -4940 5880 -4168 5908
rect -3928 6332 -3156 6360
rect -3928 5908 -3240 6332
rect -3176 5908 -3156 6332
rect -3928 5880 -3156 5908
rect -2916 6332 -2144 6360
rect -2916 5908 -2228 6332
rect -2164 5908 -2144 6332
rect -2916 5880 -2144 5908
rect -1904 6332 -1132 6360
rect -1904 5908 -1216 6332
rect -1152 5908 -1132 6332
rect -1904 5880 -1132 5908
rect -892 6332 -120 6360
rect -892 5908 -204 6332
rect -140 5908 -120 6332
rect -892 5880 -120 5908
rect 120 6332 892 6360
rect 120 5908 808 6332
rect 872 5908 892 6332
rect 120 5880 892 5908
rect 1132 6332 1904 6360
rect 1132 5908 1820 6332
rect 1884 5908 1904 6332
rect 1132 5880 1904 5908
rect 2144 6332 2916 6360
rect 2144 5908 2832 6332
rect 2896 5908 2916 6332
rect 2144 5880 2916 5908
rect 3156 6332 3928 6360
rect 3156 5908 3844 6332
rect 3908 5908 3928 6332
rect 3156 5880 3928 5908
rect 4168 6332 4940 6360
rect 4168 5908 4856 6332
rect 4920 5908 4940 6332
rect 4168 5880 4940 5908
rect 5180 6332 5952 6360
rect 5180 5908 5868 6332
rect 5932 5908 5952 6332
rect 5180 5880 5952 5908
rect 6192 6332 6964 6360
rect 6192 5908 6880 6332
rect 6944 5908 6964 6332
rect 6192 5880 6964 5908
rect 7204 6332 7976 6360
rect 7204 5908 7892 6332
rect 7956 5908 7976 6332
rect 7204 5880 7976 5908
rect 8216 6332 8988 6360
rect 8216 5908 8904 6332
rect 8968 5908 8988 6332
rect 8216 5880 8988 5908
rect 9228 6332 10000 6360
rect 9228 5908 9916 6332
rect 9980 5908 10000 6332
rect 9228 5880 10000 5908
rect 10240 6332 11012 6360
rect 10240 5908 10928 6332
rect 10992 5908 11012 6332
rect 10240 5880 11012 5908
rect 11252 6332 12024 6360
rect 11252 5908 11940 6332
rect 12004 5908 12024 6332
rect 11252 5880 12024 5908
rect 12264 6332 13036 6360
rect 12264 5908 12952 6332
rect 13016 5908 13036 6332
rect 12264 5880 13036 5908
rect 13276 6332 14048 6360
rect 13276 5908 13964 6332
rect 14028 5908 14048 6332
rect 13276 5880 14048 5908
rect 14288 6332 15060 6360
rect 14288 5908 14976 6332
rect 15040 5908 15060 6332
rect 14288 5880 15060 5908
rect 15300 6332 16072 6360
rect 15300 5908 15988 6332
rect 16052 5908 16072 6332
rect 15300 5880 16072 5908
rect 16312 6332 17084 6360
rect 16312 5908 17000 6332
rect 17064 5908 17084 6332
rect 16312 5880 17084 5908
rect -17084 5612 -16312 5640
rect -17084 5188 -16396 5612
rect -16332 5188 -16312 5612
rect -17084 5160 -16312 5188
rect -16072 5612 -15300 5640
rect -16072 5188 -15384 5612
rect -15320 5188 -15300 5612
rect -16072 5160 -15300 5188
rect -15060 5612 -14288 5640
rect -15060 5188 -14372 5612
rect -14308 5188 -14288 5612
rect -15060 5160 -14288 5188
rect -14048 5612 -13276 5640
rect -14048 5188 -13360 5612
rect -13296 5188 -13276 5612
rect -14048 5160 -13276 5188
rect -13036 5612 -12264 5640
rect -13036 5188 -12348 5612
rect -12284 5188 -12264 5612
rect -13036 5160 -12264 5188
rect -12024 5612 -11252 5640
rect -12024 5188 -11336 5612
rect -11272 5188 -11252 5612
rect -12024 5160 -11252 5188
rect -11012 5612 -10240 5640
rect -11012 5188 -10324 5612
rect -10260 5188 -10240 5612
rect -11012 5160 -10240 5188
rect -10000 5612 -9228 5640
rect -10000 5188 -9312 5612
rect -9248 5188 -9228 5612
rect -10000 5160 -9228 5188
rect -8988 5612 -8216 5640
rect -8988 5188 -8300 5612
rect -8236 5188 -8216 5612
rect -8988 5160 -8216 5188
rect -7976 5612 -7204 5640
rect -7976 5188 -7288 5612
rect -7224 5188 -7204 5612
rect -7976 5160 -7204 5188
rect -6964 5612 -6192 5640
rect -6964 5188 -6276 5612
rect -6212 5188 -6192 5612
rect -6964 5160 -6192 5188
rect -5952 5612 -5180 5640
rect -5952 5188 -5264 5612
rect -5200 5188 -5180 5612
rect -5952 5160 -5180 5188
rect -4940 5612 -4168 5640
rect -4940 5188 -4252 5612
rect -4188 5188 -4168 5612
rect -4940 5160 -4168 5188
rect -3928 5612 -3156 5640
rect -3928 5188 -3240 5612
rect -3176 5188 -3156 5612
rect -3928 5160 -3156 5188
rect -2916 5612 -2144 5640
rect -2916 5188 -2228 5612
rect -2164 5188 -2144 5612
rect -2916 5160 -2144 5188
rect -1904 5612 -1132 5640
rect -1904 5188 -1216 5612
rect -1152 5188 -1132 5612
rect -1904 5160 -1132 5188
rect -892 5612 -120 5640
rect -892 5188 -204 5612
rect -140 5188 -120 5612
rect -892 5160 -120 5188
rect 120 5612 892 5640
rect 120 5188 808 5612
rect 872 5188 892 5612
rect 120 5160 892 5188
rect 1132 5612 1904 5640
rect 1132 5188 1820 5612
rect 1884 5188 1904 5612
rect 1132 5160 1904 5188
rect 2144 5612 2916 5640
rect 2144 5188 2832 5612
rect 2896 5188 2916 5612
rect 2144 5160 2916 5188
rect 3156 5612 3928 5640
rect 3156 5188 3844 5612
rect 3908 5188 3928 5612
rect 3156 5160 3928 5188
rect 4168 5612 4940 5640
rect 4168 5188 4856 5612
rect 4920 5188 4940 5612
rect 4168 5160 4940 5188
rect 5180 5612 5952 5640
rect 5180 5188 5868 5612
rect 5932 5188 5952 5612
rect 5180 5160 5952 5188
rect 6192 5612 6964 5640
rect 6192 5188 6880 5612
rect 6944 5188 6964 5612
rect 6192 5160 6964 5188
rect 7204 5612 7976 5640
rect 7204 5188 7892 5612
rect 7956 5188 7976 5612
rect 7204 5160 7976 5188
rect 8216 5612 8988 5640
rect 8216 5188 8904 5612
rect 8968 5188 8988 5612
rect 8216 5160 8988 5188
rect 9228 5612 10000 5640
rect 9228 5188 9916 5612
rect 9980 5188 10000 5612
rect 9228 5160 10000 5188
rect 10240 5612 11012 5640
rect 10240 5188 10928 5612
rect 10992 5188 11012 5612
rect 10240 5160 11012 5188
rect 11252 5612 12024 5640
rect 11252 5188 11940 5612
rect 12004 5188 12024 5612
rect 11252 5160 12024 5188
rect 12264 5612 13036 5640
rect 12264 5188 12952 5612
rect 13016 5188 13036 5612
rect 12264 5160 13036 5188
rect 13276 5612 14048 5640
rect 13276 5188 13964 5612
rect 14028 5188 14048 5612
rect 13276 5160 14048 5188
rect 14288 5612 15060 5640
rect 14288 5188 14976 5612
rect 15040 5188 15060 5612
rect 14288 5160 15060 5188
rect 15300 5612 16072 5640
rect 15300 5188 15988 5612
rect 16052 5188 16072 5612
rect 15300 5160 16072 5188
rect 16312 5612 17084 5640
rect 16312 5188 17000 5612
rect 17064 5188 17084 5612
rect 16312 5160 17084 5188
rect -17084 4892 -16312 4920
rect -17084 4468 -16396 4892
rect -16332 4468 -16312 4892
rect -17084 4440 -16312 4468
rect -16072 4892 -15300 4920
rect -16072 4468 -15384 4892
rect -15320 4468 -15300 4892
rect -16072 4440 -15300 4468
rect -15060 4892 -14288 4920
rect -15060 4468 -14372 4892
rect -14308 4468 -14288 4892
rect -15060 4440 -14288 4468
rect -14048 4892 -13276 4920
rect -14048 4468 -13360 4892
rect -13296 4468 -13276 4892
rect -14048 4440 -13276 4468
rect -13036 4892 -12264 4920
rect -13036 4468 -12348 4892
rect -12284 4468 -12264 4892
rect -13036 4440 -12264 4468
rect -12024 4892 -11252 4920
rect -12024 4468 -11336 4892
rect -11272 4468 -11252 4892
rect -12024 4440 -11252 4468
rect -11012 4892 -10240 4920
rect -11012 4468 -10324 4892
rect -10260 4468 -10240 4892
rect -11012 4440 -10240 4468
rect -10000 4892 -9228 4920
rect -10000 4468 -9312 4892
rect -9248 4468 -9228 4892
rect -10000 4440 -9228 4468
rect -8988 4892 -8216 4920
rect -8988 4468 -8300 4892
rect -8236 4468 -8216 4892
rect -8988 4440 -8216 4468
rect -7976 4892 -7204 4920
rect -7976 4468 -7288 4892
rect -7224 4468 -7204 4892
rect -7976 4440 -7204 4468
rect -6964 4892 -6192 4920
rect -6964 4468 -6276 4892
rect -6212 4468 -6192 4892
rect -6964 4440 -6192 4468
rect -5952 4892 -5180 4920
rect -5952 4468 -5264 4892
rect -5200 4468 -5180 4892
rect -5952 4440 -5180 4468
rect -4940 4892 -4168 4920
rect -4940 4468 -4252 4892
rect -4188 4468 -4168 4892
rect -4940 4440 -4168 4468
rect -3928 4892 -3156 4920
rect -3928 4468 -3240 4892
rect -3176 4468 -3156 4892
rect -3928 4440 -3156 4468
rect -2916 4892 -2144 4920
rect -2916 4468 -2228 4892
rect -2164 4468 -2144 4892
rect -2916 4440 -2144 4468
rect -1904 4892 -1132 4920
rect -1904 4468 -1216 4892
rect -1152 4468 -1132 4892
rect -1904 4440 -1132 4468
rect -892 4892 -120 4920
rect -892 4468 -204 4892
rect -140 4468 -120 4892
rect -892 4440 -120 4468
rect 120 4892 892 4920
rect 120 4468 808 4892
rect 872 4468 892 4892
rect 120 4440 892 4468
rect 1132 4892 1904 4920
rect 1132 4468 1820 4892
rect 1884 4468 1904 4892
rect 1132 4440 1904 4468
rect 2144 4892 2916 4920
rect 2144 4468 2832 4892
rect 2896 4468 2916 4892
rect 2144 4440 2916 4468
rect 3156 4892 3928 4920
rect 3156 4468 3844 4892
rect 3908 4468 3928 4892
rect 3156 4440 3928 4468
rect 4168 4892 4940 4920
rect 4168 4468 4856 4892
rect 4920 4468 4940 4892
rect 4168 4440 4940 4468
rect 5180 4892 5952 4920
rect 5180 4468 5868 4892
rect 5932 4468 5952 4892
rect 5180 4440 5952 4468
rect 6192 4892 6964 4920
rect 6192 4468 6880 4892
rect 6944 4468 6964 4892
rect 6192 4440 6964 4468
rect 7204 4892 7976 4920
rect 7204 4468 7892 4892
rect 7956 4468 7976 4892
rect 7204 4440 7976 4468
rect 8216 4892 8988 4920
rect 8216 4468 8904 4892
rect 8968 4468 8988 4892
rect 8216 4440 8988 4468
rect 9228 4892 10000 4920
rect 9228 4468 9916 4892
rect 9980 4468 10000 4892
rect 9228 4440 10000 4468
rect 10240 4892 11012 4920
rect 10240 4468 10928 4892
rect 10992 4468 11012 4892
rect 10240 4440 11012 4468
rect 11252 4892 12024 4920
rect 11252 4468 11940 4892
rect 12004 4468 12024 4892
rect 11252 4440 12024 4468
rect 12264 4892 13036 4920
rect 12264 4468 12952 4892
rect 13016 4468 13036 4892
rect 12264 4440 13036 4468
rect 13276 4892 14048 4920
rect 13276 4468 13964 4892
rect 14028 4468 14048 4892
rect 13276 4440 14048 4468
rect 14288 4892 15060 4920
rect 14288 4468 14976 4892
rect 15040 4468 15060 4892
rect 14288 4440 15060 4468
rect 15300 4892 16072 4920
rect 15300 4468 15988 4892
rect 16052 4468 16072 4892
rect 15300 4440 16072 4468
rect 16312 4892 17084 4920
rect 16312 4468 17000 4892
rect 17064 4468 17084 4892
rect 16312 4440 17084 4468
rect -17084 4172 -16312 4200
rect -17084 3748 -16396 4172
rect -16332 3748 -16312 4172
rect -17084 3720 -16312 3748
rect -16072 4172 -15300 4200
rect -16072 3748 -15384 4172
rect -15320 3748 -15300 4172
rect -16072 3720 -15300 3748
rect -15060 4172 -14288 4200
rect -15060 3748 -14372 4172
rect -14308 3748 -14288 4172
rect -15060 3720 -14288 3748
rect -14048 4172 -13276 4200
rect -14048 3748 -13360 4172
rect -13296 3748 -13276 4172
rect -14048 3720 -13276 3748
rect -13036 4172 -12264 4200
rect -13036 3748 -12348 4172
rect -12284 3748 -12264 4172
rect -13036 3720 -12264 3748
rect -12024 4172 -11252 4200
rect -12024 3748 -11336 4172
rect -11272 3748 -11252 4172
rect -12024 3720 -11252 3748
rect -11012 4172 -10240 4200
rect -11012 3748 -10324 4172
rect -10260 3748 -10240 4172
rect -11012 3720 -10240 3748
rect -10000 4172 -9228 4200
rect -10000 3748 -9312 4172
rect -9248 3748 -9228 4172
rect -10000 3720 -9228 3748
rect -8988 4172 -8216 4200
rect -8988 3748 -8300 4172
rect -8236 3748 -8216 4172
rect -8988 3720 -8216 3748
rect -7976 4172 -7204 4200
rect -7976 3748 -7288 4172
rect -7224 3748 -7204 4172
rect -7976 3720 -7204 3748
rect -6964 4172 -6192 4200
rect -6964 3748 -6276 4172
rect -6212 3748 -6192 4172
rect -6964 3720 -6192 3748
rect -5952 4172 -5180 4200
rect -5952 3748 -5264 4172
rect -5200 3748 -5180 4172
rect -5952 3720 -5180 3748
rect -4940 4172 -4168 4200
rect -4940 3748 -4252 4172
rect -4188 3748 -4168 4172
rect -4940 3720 -4168 3748
rect -3928 4172 -3156 4200
rect -3928 3748 -3240 4172
rect -3176 3748 -3156 4172
rect -3928 3720 -3156 3748
rect -2916 4172 -2144 4200
rect -2916 3748 -2228 4172
rect -2164 3748 -2144 4172
rect -2916 3720 -2144 3748
rect -1904 4172 -1132 4200
rect -1904 3748 -1216 4172
rect -1152 3748 -1132 4172
rect -1904 3720 -1132 3748
rect -892 4172 -120 4200
rect -892 3748 -204 4172
rect -140 3748 -120 4172
rect -892 3720 -120 3748
rect 120 4172 892 4200
rect 120 3748 808 4172
rect 872 3748 892 4172
rect 120 3720 892 3748
rect 1132 4172 1904 4200
rect 1132 3748 1820 4172
rect 1884 3748 1904 4172
rect 1132 3720 1904 3748
rect 2144 4172 2916 4200
rect 2144 3748 2832 4172
rect 2896 3748 2916 4172
rect 2144 3720 2916 3748
rect 3156 4172 3928 4200
rect 3156 3748 3844 4172
rect 3908 3748 3928 4172
rect 3156 3720 3928 3748
rect 4168 4172 4940 4200
rect 4168 3748 4856 4172
rect 4920 3748 4940 4172
rect 4168 3720 4940 3748
rect 5180 4172 5952 4200
rect 5180 3748 5868 4172
rect 5932 3748 5952 4172
rect 5180 3720 5952 3748
rect 6192 4172 6964 4200
rect 6192 3748 6880 4172
rect 6944 3748 6964 4172
rect 6192 3720 6964 3748
rect 7204 4172 7976 4200
rect 7204 3748 7892 4172
rect 7956 3748 7976 4172
rect 7204 3720 7976 3748
rect 8216 4172 8988 4200
rect 8216 3748 8904 4172
rect 8968 3748 8988 4172
rect 8216 3720 8988 3748
rect 9228 4172 10000 4200
rect 9228 3748 9916 4172
rect 9980 3748 10000 4172
rect 9228 3720 10000 3748
rect 10240 4172 11012 4200
rect 10240 3748 10928 4172
rect 10992 3748 11012 4172
rect 10240 3720 11012 3748
rect 11252 4172 12024 4200
rect 11252 3748 11940 4172
rect 12004 3748 12024 4172
rect 11252 3720 12024 3748
rect 12264 4172 13036 4200
rect 12264 3748 12952 4172
rect 13016 3748 13036 4172
rect 12264 3720 13036 3748
rect 13276 4172 14048 4200
rect 13276 3748 13964 4172
rect 14028 3748 14048 4172
rect 13276 3720 14048 3748
rect 14288 4172 15060 4200
rect 14288 3748 14976 4172
rect 15040 3748 15060 4172
rect 14288 3720 15060 3748
rect 15300 4172 16072 4200
rect 15300 3748 15988 4172
rect 16052 3748 16072 4172
rect 15300 3720 16072 3748
rect 16312 4172 17084 4200
rect 16312 3748 17000 4172
rect 17064 3748 17084 4172
rect 16312 3720 17084 3748
rect -17084 3452 -16312 3480
rect -17084 3028 -16396 3452
rect -16332 3028 -16312 3452
rect -17084 3000 -16312 3028
rect -16072 3452 -15300 3480
rect -16072 3028 -15384 3452
rect -15320 3028 -15300 3452
rect -16072 3000 -15300 3028
rect -15060 3452 -14288 3480
rect -15060 3028 -14372 3452
rect -14308 3028 -14288 3452
rect -15060 3000 -14288 3028
rect -14048 3452 -13276 3480
rect -14048 3028 -13360 3452
rect -13296 3028 -13276 3452
rect -14048 3000 -13276 3028
rect -13036 3452 -12264 3480
rect -13036 3028 -12348 3452
rect -12284 3028 -12264 3452
rect -13036 3000 -12264 3028
rect -12024 3452 -11252 3480
rect -12024 3028 -11336 3452
rect -11272 3028 -11252 3452
rect -12024 3000 -11252 3028
rect -11012 3452 -10240 3480
rect -11012 3028 -10324 3452
rect -10260 3028 -10240 3452
rect -11012 3000 -10240 3028
rect -10000 3452 -9228 3480
rect -10000 3028 -9312 3452
rect -9248 3028 -9228 3452
rect -10000 3000 -9228 3028
rect -8988 3452 -8216 3480
rect -8988 3028 -8300 3452
rect -8236 3028 -8216 3452
rect -8988 3000 -8216 3028
rect -7976 3452 -7204 3480
rect -7976 3028 -7288 3452
rect -7224 3028 -7204 3452
rect -7976 3000 -7204 3028
rect -6964 3452 -6192 3480
rect -6964 3028 -6276 3452
rect -6212 3028 -6192 3452
rect -6964 3000 -6192 3028
rect -5952 3452 -5180 3480
rect -5952 3028 -5264 3452
rect -5200 3028 -5180 3452
rect -5952 3000 -5180 3028
rect -4940 3452 -4168 3480
rect -4940 3028 -4252 3452
rect -4188 3028 -4168 3452
rect -4940 3000 -4168 3028
rect -3928 3452 -3156 3480
rect -3928 3028 -3240 3452
rect -3176 3028 -3156 3452
rect -3928 3000 -3156 3028
rect -2916 3452 -2144 3480
rect -2916 3028 -2228 3452
rect -2164 3028 -2144 3452
rect -2916 3000 -2144 3028
rect -1904 3452 -1132 3480
rect -1904 3028 -1216 3452
rect -1152 3028 -1132 3452
rect -1904 3000 -1132 3028
rect -892 3452 -120 3480
rect -892 3028 -204 3452
rect -140 3028 -120 3452
rect -892 3000 -120 3028
rect 120 3452 892 3480
rect 120 3028 808 3452
rect 872 3028 892 3452
rect 120 3000 892 3028
rect 1132 3452 1904 3480
rect 1132 3028 1820 3452
rect 1884 3028 1904 3452
rect 1132 3000 1904 3028
rect 2144 3452 2916 3480
rect 2144 3028 2832 3452
rect 2896 3028 2916 3452
rect 2144 3000 2916 3028
rect 3156 3452 3928 3480
rect 3156 3028 3844 3452
rect 3908 3028 3928 3452
rect 3156 3000 3928 3028
rect 4168 3452 4940 3480
rect 4168 3028 4856 3452
rect 4920 3028 4940 3452
rect 4168 3000 4940 3028
rect 5180 3452 5952 3480
rect 5180 3028 5868 3452
rect 5932 3028 5952 3452
rect 5180 3000 5952 3028
rect 6192 3452 6964 3480
rect 6192 3028 6880 3452
rect 6944 3028 6964 3452
rect 6192 3000 6964 3028
rect 7204 3452 7976 3480
rect 7204 3028 7892 3452
rect 7956 3028 7976 3452
rect 7204 3000 7976 3028
rect 8216 3452 8988 3480
rect 8216 3028 8904 3452
rect 8968 3028 8988 3452
rect 8216 3000 8988 3028
rect 9228 3452 10000 3480
rect 9228 3028 9916 3452
rect 9980 3028 10000 3452
rect 9228 3000 10000 3028
rect 10240 3452 11012 3480
rect 10240 3028 10928 3452
rect 10992 3028 11012 3452
rect 10240 3000 11012 3028
rect 11252 3452 12024 3480
rect 11252 3028 11940 3452
rect 12004 3028 12024 3452
rect 11252 3000 12024 3028
rect 12264 3452 13036 3480
rect 12264 3028 12952 3452
rect 13016 3028 13036 3452
rect 12264 3000 13036 3028
rect 13276 3452 14048 3480
rect 13276 3028 13964 3452
rect 14028 3028 14048 3452
rect 13276 3000 14048 3028
rect 14288 3452 15060 3480
rect 14288 3028 14976 3452
rect 15040 3028 15060 3452
rect 14288 3000 15060 3028
rect 15300 3452 16072 3480
rect 15300 3028 15988 3452
rect 16052 3028 16072 3452
rect 15300 3000 16072 3028
rect 16312 3452 17084 3480
rect 16312 3028 17000 3452
rect 17064 3028 17084 3452
rect 16312 3000 17084 3028
rect -17084 2732 -16312 2760
rect -17084 2308 -16396 2732
rect -16332 2308 -16312 2732
rect -17084 2280 -16312 2308
rect -16072 2732 -15300 2760
rect -16072 2308 -15384 2732
rect -15320 2308 -15300 2732
rect -16072 2280 -15300 2308
rect -15060 2732 -14288 2760
rect -15060 2308 -14372 2732
rect -14308 2308 -14288 2732
rect -15060 2280 -14288 2308
rect -14048 2732 -13276 2760
rect -14048 2308 -13360 2732
rect -13296 2308 -13276 2732
rect -14048 2280 -13276 2308
rect -13036 2732 -12264 2760
rect -13036 2308 -12348 2732
rect -12284 2308 -12264 2732
rect -13036 2280 -12264 2308
rect -12024 2732 -11252 2760
rect -12024 2308 -11336 2732
rect -11272 2308 -11252 2732
rect -12024 2280 -11252 2308
rect -11012 2732 -10240 2760
rect -11012 2308 -10324 2732
rect -10260 2308 -10240 2732
rect -11012 2280 -10240 2308
rect -10000 2732 -9228 2760
rect -10000 2308 -9312 2732
rect -9248 2308 -9228 2732
rect -10000 2280 -9228 2308
rect -8988 2732 -8216 2760
rect -8988 2308 -8300 2732
rect -8236 2308 -8216 2732
rect -8988 2280 -8216 2308
rect -7976 2732 -7204 2760
rect -7976 2308 -7288 2732
rect -7224 2308 -7204 2732
rect -7976 2280 -7204 2308
rect -6964 2732 -6192 2760
rect -6964 2308 -6276 2732
rect -6212 2308 -6192 2732
rect -6964 2280 -6192 2308
rect -5952 2732 -5180 2760
rect -5952 2308 -5264 2732
rect -5200 2308 -5180 2732
rect -5952 2280 -5180 2308
rect -4940 2732 -4168 2760
rect -4940 2308 -4252 2732
rect -4188 2308 -4168 2732
rect -4940 2280 -4168 2308
rect -3928 2732 -3156 2760
rect -3928 2308 -3240 2732
rect -3176 2308 -3156 2732
rect -3928 2280 -3156 2308
rect -2916 2732 -2144 2760
rect -2916 2308 -2228 2732
rect -2164 2308 -2144 2732
rect -2916 2280 -2144 2308
rect -1904 2732 -1132 2760
rect -1904 2308 -1216 2732
rect -1152 2308 -1132 2732
rect -1904 2280 -1132 2308
rect -892 2732 -120 2760
rect -892 2308 -204 2732
rect -140 2308 -120 2732
rect -892 2280 -120 2308
rect 120 2732 892 2760
rect 120 2308 808 2732
rect 872 2308 892 2732
rect 120 2280 892 2308
rect 1132 2732 1904 2760
rect 1132 2308 1820 2732
rect 1884 2308 1904 2732
rect 1132 2280 1904 2308
rect 2144 2732 2916 2760
rect 2144 2308 2832 2732
rect 2896 2308 2916 2732
rect 2144 2280 2916 2308
rect 3156 2732 3928 2760
rect 3156 2308 3844 2732
rect 3908 2308 3928 2732
rect 3156 2280 3928 2308
rect 4168 2732 4940 2760
rect 4168 2308 4856 2732
rect 4920 2308 4940 2732
rect 4168 2280 4940 2308
rect 5180 2732 5952 2760
rect 5180 2308 5868 2732
rect 5932 2308 5952 2732
rect 5180 2280 5952 2308
rect 6192 2732 6964 2760
rect 6192 2308 6880 2732
rect 6944 2308 6964 2732
rect 6192 2280 6964 2308
rect 7204 2732 7976 2760
rect 7204 2308 7892 2732
rect 7956 2308 7976 2732
rect 7204 2280 7976 2308
rect 8216 2732 8988 2760
rect 8216 2308 8904 2732
rect 8968 2308 8988 2732
rect 8216 2280 8988 2308
rect 9228 2732 10000 2760
rect 9228 2308 9916 2732
rect 9980 2308 10000 2732
rect 9228 2280 10000 2308
rect 10240 2732 11012 2760
rect 10240 2308 10928 2732
rect 10992 2308 11012 2732
rect 10240 2280 11012 2308
rect 11252 2732 12024 2760
rect 11252 2308 11940 2732
rect 12004 2308 12024 2732
rect 11252 2280 12024 2308
rect 12264 2732 13036 2760
rect 12264 2308 12952 2732
rect 13016 2308 13036 2732
rect 12264 2280 13036 2308
rect 13276 2732 14048 2760
rect 13276 2308 13964 2732
rect 14028 2308 14048 2732
rect 13276 2280 14048 2308
rect 14288 2732 15060 2760
rect 14288 2308 14976 2732
rect 15040 2308 15060 2732
rect 14288 2280 15060 2308
rect 15300 2732 16072 2760
rect 15300 2308 15988 2732
rect 16052 2308 16072 2732
rect 15300 2280 16072 2308
rect 16312 2732 17084 2760
rect 16312 2308 17000 2732
rect 17064 2308 17084 2732
rect 16312 2280 17084 2308
rect -17084 2012 -16312 2040
rect -17084 1588 -16396 2012
rect -16332 1588 -16312 2012
rect -17084 1560 -16312 1588
rect -16072 2012 -15300 2040
rect -16072 1588 -15384 2012
rect -15320 1588 -15300 2012
rect -16072 1560 -15300 1588
rect -15060 2012 -14288 2040
rect -15060 1588 -14372 2012
rect -14308 1588 -14288 2012
rect -15060 1560 -14288 1588
rect -14048 2012 -13276 2040
rect -14048 1588 -13360 2012
rect -13296 1588 -13276 2012
rect -14048 1560 -13276 1588
rect -13036 2012 -12264 2040
rect -13036 1588 -12348 2012
rect -12284 1588 -12264 2012
rect -13036 1560 -12264 1588
rect -12024 2012 -11252 2040
rect -12024 1588 -11336 2012
rect -11272 1588 -11252 2012
rect -12024 1560 -11252 1588
rect -11012 2012 -10240 2040
rect -11012 1588 -10324 2012
rect -10260 1588 -10240 2012
rect -11012 1560 -10240 1588
rect -10000 2012 -9228 2040
rect -10000 1588 -9312 2012
rect -9248 1588 -9228 2012
rect -10000 1560 -9228 1588
rect -8988 2012 -8216 2040
rect -8988 1588 -8300 2012
rect -8236 1588 -8216 2012
rect -8988 1560 -8216 1588
rect -7976 2012 -7204 2040
rect -7976 1588 -7288 2012
rect -7224 1588 -7204 2012
rect -7976 1560 -7204 1588
rect -6964 2012 -6192 2040
rect -6964 1588 -6276 2012
rect -6212 1588 -6192 2012
rect -6964 1560 -6192 1588
rect -5952 2012 -5180 2040
rect -5952 1588 -5264 2012
rect -5200 1588 -5180 2012
rect -5952 1560 -5180 1588
rect -4940 2012 -4168 2040
rect -4940 1588 -4252 2012
rect -4188 1588 -4168 2012
rect -4940 1560 -4168 1588
rect -3928 2012 -3156 2040
rect -3928 1588 -3240 2012
rect -3176 1588 -3156 2012
rect -3928 1560 -3156 1588
rect -2916 2012 -2144 2040
rect -2916 1588 -2228 2012
rect -2164 1588 -2144 2012
rect -2916 1560 -2144 1588
rect -1904 2012 -1132 2040
rect -1904 1588 -1216 2012
rect -1152 1588 -1132 2012
rect -1904 1560 -1132 1588
rect -892 2012 -120 2040
rect -892 1588 -204 2012
rect -140 1588 -120 2012
rect -892 1560 -120 1588
rect 120 2012 892 2040
rect 120 1588 808 2012
rect 872 1588 892 2012
rect 120 1560 892 1588
rect 1132 2012 1904 2040
rect 1132 1588 1820 2012
rect 1884 1588 1904 2012
rect 1132 1560 1904 1588
rect 2144 2012 2916 2040
rect 2144 1588 2832 2012
rect 2896 1588 2916 2012
rect 2144 1560 2916 1588
rect 3156 2012 3928 2040
rect 3156 1588 3844 2012
rect 3908 1588 3928 2012
rect 3156 1560 3928 1588
rect 4168 2012 4940 2040
rect 4168 1588 4856 2012
rect 4920 1588 4940 2012
rect 4168 1560 4940 1588
rect 5180 2012 5952 2040
rect 5180 1588 5868 2012
rect 5932 1588 5952 2012
rect 5180 1560 5952 1588
rect 6192 2012 6964 2040
rect 6192 1588 6880 2012
rect 6944 1588 6964 2012
rect 6192 1560 6964 1588
rect 7204 2012 7976 2040
rect 7204 1588 7892 2012
rect 7956 1588 7976 2012
rect 7204 1560 7976 1588
rect 8216 2012 8988 2040
rect 8216 1588 8904 2012
rect 8968 1588 8988 2012
rect 8216 1560 8988 1588
rect 9228 2012 10000 2040
rect 9228 1588 9916 2012
rect 9980 1588 10000 2012
rect 9228 1560 10000 1588
rect 10240 2012 11012 2040
rect 10240 1588 10928 2012
rect 10992 1588 11012 2012
rect 10240 1560 11012 1588
rect 11252 2012 12024 2040
rect 11252 1588 11940 2012
rect 12004 1588 12024 2012
rect 11252 1560 12024 1588
rect 12264 2012 13036 2040
rect 12264 1588 12952 2012
rect 13016 1588 13036 2012
rect 12264 1560 13036 1588
rect 13276 2012 14048 2040
rect 13276 1588 13964 2012
rect 14028 1588 14048 2012
rect 13276 1560 14048 1588
rect 14288 2012 15060 2040
rect 14288 1588 14976 2012
rect 15040 1588 15060 2012
rect 14288 1560 15060 1588
rect 15300 2012 16072 2040
rect 15300 1588 15988 2012
rect 16052 1588 16072 2012
rect 15300 1560 16072 1588
rect 16312 2012 17084 2040
rect 16312 1588 17000 2012
rect 17064 1588 17084 2012
rect 16312 1560 17084 1588
rect -17084 1292 -16312 1320
rect -17084 868 -16396 1292
rect -16332 868 -16312 1292
rect -17084 840 -16312 868
rect -16072 1292 -15300 1320
rect -16072 868 -15384 1292
rect -15320 868 -15300 1292
rect -16072 840 -15300 868
rect -15060 1292 -14288 1320
rect -15060 868 -14372 1292
rect -14308 868 -14288 1292
rect -15060 840 -14288 868
rect -14048 1292 -13276 1320
rect -14048 868 -13360 1292
rect -13296 868 -13276 1292
rect -14048 840 -13276 868
rect -13036 1292 -12264 1320
rect -13036 868 -12348 1292
rect -12284 868 -12264 1292
rect -13036 840 -12264 868
rect -12024 1292 -11252 1320
rect -12024 868 -11336 1292
rect -11272 868 -11252 1292
rect -12024 840 -11252 868
rect -11012 1292 -10240 1320
rect -11012 868 -10324 1292
rect -10260 868 -10240 1292
rect -11012 840 -10240 868
rect -10000 1292 -9228 1320
rect -10000 868 -9312 1292
rect -9248 868 -9228 1292
rect -10000 840 -9228 868
rect -8988 1292 -8216 1320
rect -8988 868 -8300 1292
rect -8236 868 -8216 1292
rect -8988 840 -8216 868
rect -7976 1292 -7204 1320
rect -7976 868 -7288 1292
rect -7224 868 -7204 1292
rect -7976 840 -7204 868
rect -6964 1292 -6192 1320
rect -6964 868 -6276 1292
rect -6212 868 -6192 1292
rect -6964 840 -6192 868
rect -5952 1292 -5180 1320
rect -5952 868 -5264 1292
rect -5200 868 -5180 1292
rect -5952 840 -5180 868
rect -4940 1292 -4168 1320
rect -4940 868 -4252 1292
rect -4188 868 -4168 1292
rect -4940 840 -4168 868
rect -3928 1292 -3156 1320
rect -3928 868 -3240 1292
rect -3176 868 -3156 1292
rect -3928 840 -3156 868
rect -2916 1292 -2144 1320
rect -2916 868 -2228 1292
rect -2164 868 -2144 1292
rect -2916 840 -2144 868
rect -1904 1292 -1132 1320
rect -1904 868 -1216 1292
rect -1152 868 -1132 1292
rect -1904 840 -1132 868
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect 1132 1292 1904 1320
rect 1132 868 1820 1292
rect 1884 868 1904 1292
rect 1132 840 1904 868
rect 2144 1292 2916 1320
rect 2144 868 2832 1292
rect 2896 868 2916 1292
rect 2144 840 2916 868
rect 3156 1292 3928 1320
rect 3156 868 3844 1292
rect 3908 868 3928 1292
rect 3156 840 3928 868
rect 4168 1292 4940 1320
rect 4168 868 4856 1292
rect 4920 868 4940 1292
rect 4168 840 4940 868
rect 5180 1292 5952 1320
rect 5180 868 5868 1292
rect 5932 868 5952 1292
rect 5180 840 5952 868
rect 6192 1292 6964 1320
rect 6192 868 6880 1292
rect 6944 868 6964 1292
rect 6192 840 6964 868
rect 7204 1292 7976 1320
rect 7204 868 7892 1292
rect 7956 868 7976 1292
rect 7204 840 7976 868
rect 8216 1292 8988 1320
rect 8216 868 8904 1292
rect 8968 868 8988 1292
rect 8216 840 8988 868
rect 9228 1292 10000 1320
rect 9228 868 9916 1292
rect 9980 868 10000 1292
rect 9228 840 10000 868
rect 10240 1292 11012 1320
rect 10240 868 10928 1292
rect 10992 868 11012 1292
rect 10240 840 11012 868
rect 11252 1292 12024 1320
rect 11252 868 11940 1292
rect 12004 868 12024 1292
rect 11252 840 12024 868
rect 12264 1292 13036 1320
rect 12264 868 12952 1292
rect 13016 868 13036 1292
rect 12264 840 13036 868
rect 13276 1292 14048 1320
rect 13276 868 13964 1292
rect 14028 868 14048 1292
rect 13276 840 14048 868
rect 14288 1292 15060 1320
rect 14288 868 14976 1292
rect 15040 868 15060 1292
rect 14288 840 15060 868
rect 15300 1292 16072 1320
rect 15300 868 15988 1292
rect 16052 868 16072 1292
rect 15300 840 16072 868
rect 16312 1292 17084 1320
rect 16312 868 17000 1292
rect 17064 868 17084 1292
rect 16312 840 17084 868
rect -17084 572 -16312 600
rect -17084 148 -16396 572
rect -16332 148 -16312 572
rect -17084 120 -16312 148
rect -16072 572 -15300 600
rect -16072 148 -15384 572
rect -15320 148 -15300 572
rect -16072 120 -15300 148
rect -15060 572 -14288 600
rect -15060 148 -14372 572
rect -14308 148 -14288 572
rect -15060 120 -14288 148
rect -14048 572 -13276 600
rect -14048 148 -13360 572
rect -13296 148 -13276 572
rect -14048 120 -13276 148
rect -13036 572 -12264 600
rect -13036 148 -12348 572
rect -12284 148 -12264 572
rect -13036 120 -12264 148
rect -12024 572 -11252 600
rect -12024 148 -11336 572
rect -11272 148 -11252 572
rect -12024 120 -11252 148
rect -11012 572 -10240 600
rect -11012 148 -10324 572
rect -10260 148 -10240 572
rect -11012 120 -10240 148
rect -10000 572 -9228 600
rect -10000 148 -9312 572
rect -9248 148 -9228 572
rect -10000 120 -9228 148
rect -8988 572 -8216 600
rect -8988 148 -8300 572
rect -8236 148 -8216 572
rect -8988 120 -8216 148
rect -7976 572 -7204 600
rect -7976 148 -7288 572
rect -7224 148 -7204 572
rect -7976 120 -7204 148
rect -6964 572 -6192 600
rect -6964 148 -6276 572
rect -6212 148 -6192 572
rect -6964 120 -6192 148
rect -5952 572 -5180 600
rect -5952 148 -5264 572
rect -5200 148 -5180 572
rect -5952 120 -5180 148
rect -4940 572 -4168 600
rect -4940 148 -4252 572
rect -4188 148 -4168 572
rect -4940 120 -4168 148
rect -3928 572 -3156 600
rect -3928 148 -3240 572
rect -3176 148 -3156 572
rect -3928 120 -3156 148
rect -2916 572 -2144 600
rect -2916 148 -2228 572
rect -2164 148 -2144 572
rect -2916 120 -2144 148
rect -1904 572 -1132 600
rect -1904 148 -1216 572
rect -1152 148 -1132 572
rect -1904 120 -1132 148
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect 1132 572 1904 600
rect 1132 148 1820 572
rect 1884 148 1904 572
rect 1132 120 1904 148
rect 2144 572 2916 600
rect 2144 148 2832 572
rect 2896 148 2916 572
rect 2144 120 2916 148
rect 3156 572 3928 600
rect 3156 148 3844 572
rect 3908 148 3928 572
rect 3156 120 3928 148
rect 4168 572 4940 600
rect 4168 148 4856 572
rect 4920 148 4940 572
rect 4168 120 4940 148
rect 5180 572 5952 600
rect 5180 148 5868 572
rect 5932 148 5952 572
rect 5180 120 5952 148
rect 6192 572 6964 600
rect 6192 148 6880 572
rect 6944 148 6964 572
rect 6192 120 6964 148
rect 7204 572 7976 600
rect 7204 148 7892 572
rect 7956 148 7976 572
rect 7204 120 7976 148
rect 8216 572 8988 600
rect 8216 148 8904 572
rect 8968 148 8988 572
rect 8216 120 8988 148
rect 9228 572 10000 600
rect 9228 148 9916 572
rect 9980 148 10000 572
rect 9228 120 10000 148
rect 10240 572 11012 600
rect 10240 148 10928 572
rect 10992 148 11012 572
rect 10240 120 11012 148
rect 11252 572 12024 600
rect 11252 148 11940 572
rect 12004 148 12024 572
rect 11252 120 12024 148
rect 12264 572 13036 600
rect 12264 148 12952 572
rect 13016 148 13036 572
rect 12264 120 13036 148
rect 13276 572 14048 600
rect 13276 148 13964 572
rect 14028 148 14048 572
rect 13276 120 14048 148
rect 14288 572 15060 600
rect 14288 148 14976 572
rect 15040 148 15060 572
rect 14288 120 15060 148
rect 15300 572 16072 600
rect 15300 148 15988 572
rect 16052 148 16072 572
rect 15300 120 16072 148
rect 16312 572 17084 600
rect 16312 148 17000 572
rect 17064 148 17084 572
rect 16312 120 17084 148
rect -17084 -148 -16312 -120
rect -17084 -572 -16396 -148
rect -16332 -572 -16312 -148
rect -17084 -600 -16312 -572
rect -16072 -148 -15300 -120
rect -16072 -572 -15384 -148
rect -15320 -572 -15300 -148
rect -16072 -600 -15300 -572
rect -15060 -148 -14288 -120
rect -15060 -572 -14372 -148
rect -14308 -572 -14288 -148
rect -15060 -600 -14288 -572
rect -14048 -148 -13276 -120
rect -14048 -572 -13360 -148
rect -13296 -572 -13276 -148
rect -14048 -600 -13276 -572
rect -13036 -148 -12264 -120
rect -13036 -572 -12348 -148
rect -12284 -572 -12264 -148
rect -13036 -600 -12264 -572
rect -12024 -148 -11252 -120
rect -12024 -572 -11336 -148
rect -11272 -572 -11252 -148
rect -12024 -600 -11252 -572
rect -11012 -148 -10240 -120
rect -11012 -572 -10324 -148
rect -10260 -572 -10240 -148
rect -11012 -600 -10240 -572
rect -10000 -148 -9228 -120
rect -10000 -572 -9312 -148
rect -9248 -572 -9228 -148
rect -10000 -600 -9228 -572
rect -8988 -148 -8216 -120
rect -8988 -572 -8300 -148
rect -8236 -572 -8216 -148
rect -8988 -600 -8216 -572
rect -7976 -148 -7204 -120
rect -7976 -572 -7288 -148
rect -7224 -572 -7204 -148
rect -7976 -600 -7204 -572
rect -6964 -148 -6192 -120
rect -6964 -572 -6276 -148
rect -6212 -572 -6192 -148
rect -6964 -600 -6192 -572
rect -5952 -148 -5180 -120
rect -5952 -572 -5264 -148
rect -5200 -572 -5180 -148
rect -5952 -600 -5180 -572
rect -4940 -148 -4168 -120
rect -4940 -572 -4252 -148
rect -4188 -572 -4168 -148
rect -4940 -600 -4168 -572
rect -3928 -148 -3156 -120
rect -3928 -572 -3240 -148
rect -3176 -572 -3156 -148
rect -3928 -600 -3156 -572
rect -2916 -148 -2144 -120
rect -2916 -572 -2228 -148
rect -2164 -572 -2144 -148
rect -2916 -600 -2144 -572
rect -1904 -148 -1132 -120
rect -1904 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -1904 -600 -1132 -572
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect 1132 -148 1904 -120
rect 1132 -572 1820 -148
rect 1884 -572 1904 -148
rect 1132 -600 1904 -572
rect 2144 -148 2916 -120
rect 2144 -572 2832 -148
rect 2896 -572 2916 -148
rect 2144 -600 2916 -572
rect 3156 -148 3928 -120
rect 3156 -572 3844 -148
rect 3908 -572 3928 -148
rect 3156 -600 3928 -572
rect 4168 -148 4940 -120
rect 4168 -572 4856 -148
rect 4920 -572 4940 -148
rect 4168 -600 4940 -572
rect 5180 -148 5952 -120
rect 5180 -572 5868 -148
rect 5932 -572 5952 -148
rect 5180 -600 5952 -572
rect 6192 -148 6964 -120
rect 6192 -572 6880 -148
rect 6944 -572 6964 -148
rect 6192 -600 6964 -572
rect 7204 -148 7976 -120
rect 7204 -572 7892 -148
rect 7956 -572 7976 -148
rect 7204 -600 7976 -572
rect 8216 -148 8988 -120
rect 8216 -572 8904 -148
rect 8968 -572 8988 -148
rect 8216 -600 8988 -572
rect 9228 -148 10000 -120
rect 9228 -572 9916 -148
rect 9980 -572 10000 -148
rect 9228 -600 10000 -572
rect 10240 -148 11012 -120
rect 10240 -572 10928 -148
rect 10992 -572 11012 -148
rect 10240 -600 11012 -572
rect 11252 -148 12024 -120
rect 11252 -572 11940 -148
rect 12004 -572 12024 -148
rect 11252 -600 12024 -572
rect 12264 -148 13036 -120
rect 12264 -572 12952 -148
rect 13016 -572 13036 -148
rect 12264 -600 13036 -572
rect 13276 -148 14048 -120
rect 13276 -572 13964 -148
rect 14028 -572 14048 -148
rect 13276 -600 14048 -572
rect 14288 -148 15060 -120
rect 14288 -572 14976 -148
rect 15040 -572 15060 -148
rect 14288 -600 15060 -572
rect 15300 -148 16072 -120
rect 15300 -572 15988 -148
rect 16052 -572 16072 -148
rect 15300 -600 16072 -572
rect 16312 -148 17084 -120
rect 16312 -572 17000 -148
rect 17064 -572 17084 -148
rect 16312 -600 17084 -572
rect -17084 -868 -16312 -840
rect -17084 -1292 -16396 -868
rect -16332 -1292 -16312 -868
rect -17084 -1320 -16312 -1292
rect -16072 -868 -15300 -840
rect -16072 -1292 -15384 -868
rect -15320 -1292 -15300 -868
rect -16072 -1320 -15300 -1292
rect -15060 -868 -14288 -840
rect -15060 -1292 -14372 -868
rect -14308 -1292 -14288 -868
rect -15060 -1320 -14288 -1292
rect -14048 -868 -13276 -840
rect -14048 -1292 -13360 -868
rect -13296 -1292 -13276 -868
rect -14048 -1320 -13276 -1292
rect -13036 -868 -12264 -840
rect -13036 -1292 -12348 -868
rect -12284 -1292 -12264 -868
rect -13036 -1320 -12264 -1292
rect -12024 -868 -11252 -840
rect -12024 -1292 -11336 -868
rect -11272 -1292 -11252 -868
rect -12024 -1320 -11252 -1292
rect -11012 -868 -10240 -840
rect -11012 -1292 -10324 -868
rect -10260 -1292 -10240 -868
rect -11012 -1320 -10240 -1292
rect -10000 -868 -9228 -840
rect -10000 -1292 -9312 -868
rect -9248 -1292 -9228 -868
rect -10000 -1320 -9228 -1292
rect -8988 -868 -8216 -840
rect -8988 -1292 -8300 -868
rect -8236 -1292 -8216 -868
rect -8988 -1320 -8216 -1292
rect -7976 -868 -7204 -840
rect -7976 -1292 -7288 -868
rect -7224 -1292 -7204 -868
rect -7976 -1320 -7204 -1292
rect -6964 -868 -6192 -840
rect -6964 -1292 -6276 -868
rect -6212 -1292 -6192 -868
rect -6964 -1320 -6192 -1292
rect -5952 -868 -5180 -840
rect -5952 -1292 -5264 -868
rect -5200 -1292 -5180 -868
rect -5952 -1320 -5180 -1292
rect -4940 -868 -4168 -840
rect -4940 -1292 -4252 -868
rect -4188 -1292 -4168 -868
rect -4940 -1320 -4168 -1292
rect -3928 -868 -3156 -840
rect -3928 -1292 -3240 -868
rect -3176 -1292 -3156 -868
rect -3928 -1320 -3156 -1292
rect -2916 -868 -2144 -840
rect -2916 -1292 -2228 -868
rect -2164 -1292 -2144 -868
rect -2916 -1320 -2144 -1292
rect -1904 -868 -1132 -840
rect -1904 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -1904 -1320 -1132 -1292
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect 1132 -868 1904 -840
rect 1132 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 1132 -1320 1904 -1292
rect 2144 -868 2916 -840
rect 2144 -1292 2832 -868
rect 2896 -1292 2916 -868
rect 2144 -1320 2916 -1292
rect 3156 -868 3928 -840
rect 3156 -1292 3844 -868
rect 3908 -1292 3928 -868
rect 3156 -1320 3928 -1292
rect 4168 -868 4940 -840
rect 4168 -1292 4856 -868
rect 4920 -1292 4940 -868
rect 4168 -1320 4940 -1292
rect 5180 -868 5952 -840
rect 5180 -1292 5868 -868
rect 5932 -1292 5952 -868
rect 5180 -1320 5952 -1292
rect 6192 -868 6964 -840
rect 6192 -1292 6880 -868
rect 6944 -1292 6964 -868
rect 6192 -1320 6964 -1292
rect 7204 -868 7976 -840
rect 7204 -1292 7892 -868
rect 7956 -1292 7976 -868
rect 7204 -1320 7976 -1292
rect 8216 -868 8988 -840
rect 8216 -1292 8904 -868
rect 8968 -1292 8988 -868
rect 8216 -1320 8988 -1292
rect 9228 -868 10000 -840
rect 9228 -1292 9916 -868
rect 9980 -1292 10000 -868
rect 9228 -1320 10000 -1292
rect 10240 -868 11012 -840
rect 10240 -1292 10928 -868
rect 10992 -1292 11012 -868
rect 10240 -1320 11012 -1292
rect 11252 -868 12024 -840
rect 11252 -1292 11940 -868
rect 12004 -1292 12024 -868
rect 11252 -1320 12024 -1292
rect 12264 -868 13036 -840
rect 12264 -1292 12952 -868
rect 13016 -1292 13036 -868
rect 12264 -1320 13036 -1292
rect 13276 -868 14048 -840
rect 13276 -1292 13964 -868
rect 14028 -1292 14048 -868
rect 13276 -1320 14048 -1292
rect 14288 -868 15060 -840
rect 14288 -1292 14976 -868
rect 15040 -1292 15060 -868
rect 14288 -1320 15060 -1292
rect 15300 -868 16072 -840
rect 15300 -1292 15988 -868
rect 16052 -1292 16072 -868
rect 15300 -1320 16072 -1292
rect 16312 -868 17084 -840
rect 16312 -1292 17000 -868
rect 17064 -1292 17084 -868
rect 16312 -1320 17084 -1292
rect -17084 -1588 -16312 -1560
rect -17084 -2012 -16396 -1588
rect -16332 -2012 -16312 -1588
rect -17084 -2040 -16312 -2012
rect -16072 -1588 -15300 -1560
rect -16072 -2012 -15384 -1588
rect -15320 -2012 -15300 -1588
rect -16072 -2040 -15300 -2012
rect -15060 -1588 -14288 -1560
rect -15060 -2012 -14372 -1588
rect -14308 -2012 -14288 -1588
rect -15060 -2040 -14288 -2012
rect -14048 -1588 -13276 -1560
rect -14048 -2012 -13360 -1588
rect -13296 -2012 -13276 -1588
rect -14048 -2040 -13276 -2012
rect -13036 -1588 -12264 -1560
rect -13036 -2012 -12348 -1588
rect -12284 -2012 -12264 -1588
rect -13036 -2040 -12264 -2012
rect -12024 -1588 -11252 -1560
rect -12024 -2012 -11336 -1588
rect -11272 -2012 -11252 -1588
rect -12024 -2040 -11252 -2012
rect -11012 -1588 -10240 -1560
rect -11012 -2012 -10324 -1588
rect -10260 -2012 -10240 -1588
rect -11012 -2040 -10240 -2012
rect -10000 -1588 -9228 -1560
rect -10000 -2012 -9312 -1588
rect -9248 -2012 -9228 -1588
rect -10000 -2040 -9228 -2012
rect -8988 -1588 -8216 -1560
rect -8988 -2012 -8300 -1588
rect -8236 -2012 -8216 -1588
rect -8988 -2040 -8216 -2012
rect -7976 -1588 -7204 -1560
rect -7976 -2012 -7288 -1588
rect -7224 -2012 -7204 -1588
rect -7976 -2040 -7204 -2012
rect -6964 -1588 -6192 -1560
rect -6964 -2012 -6276 -1588
rect -6212 -2012 -6192 -1588
rect -6964 -2040 -6192 -2012
rect -5952 -1588 -5180 -1560
rect -5952 -2012 -5264 -1588
rect -5200 -2012 -5180 -1588
rect -5952 -2040 -5180 -2012
rect -4940 -1588 -4168 -1560
rect -4940 -2012 -4252 -1588
rect -4188 -2012 -4168 -1588
rect -4940 -2040 -4168 -2012
rect -3928 -1588 -3156 -1560
rect -3928 -2012 -3240 -1588
rect -3176 -2012 -3156 -1588
rect -3928 -2040 -3156 -2012
rect -2916 -1588 -2144 -1560
rect -2916 -2012 -2228 -1588
rect -2164 -2012 -2144 -1588
rect -2916 -2040 -2144 -2012
rect -1904 -1588 -1132 -1560
rect -1904 -2012 -1216 -1588
rect -1152 -2012 -1132 -1588
rect -1904 -2040 -1132 -2012
rect -892 -1588 -120 -1560
rect -892 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect -892 -2040 -120 -2012
rect 120 -1588 892 -1560
rect 120 -2012 808 -1588
rect 872 -2012 892 -1588
rect 120 -2040 892 -2012
rect 1132 -1588 1904 -1560
rect 1132 -2012 1820 -1588
rect 1884 -2012 1904 -1588
rect 1132 -2040 1904 -2012
rect 2144 -1588 2916 -1560
rect 2144 -2012 2832 -1588
rect 2896 -2012 2916 -1588
rect 2144 -2040 2916 -2012
rect 3156 -1588 3928 -1560
rect 3156 -2012 3844 -1588
rect 3908 -2012 3928 -1588
rect 3156 -2040 3928 -2012
rect 4168 -1588 4940 -1560
rect 4168 -2012 4856 -1588
rect 4920 -2012 4940 -1588
rect 4168 -2040 4940 -2012
rect 5180 -1588 5952 -1560
rect 5180 -2012 5868 -1588
rect 5932 -2012 5952 -1588
rect 5180 -2040 5952 -2012
rect 6192 -1588 6964 -1560
rect 6192 -2012 6880 -1588
rect 6944 -2012 6964 -1588
rect 6192 -2040 6964 -2012
rect 7204 -1588 7976 -1560
rect 7204 -2012 7892 -1588
rect 7956 -2012 7976 -1588
rect 7204 -2040 7976 -2012
rect 8216 -1588 8988 -1560
rect 8216 -2012 8904 -1588
rect 8968 -2012 8988 -1588
rect 8216 -2040 8988 -2012
rect 9228 -1588 10000 -1560
rect 9228 -2012 9916 -1588
rect 9980 -2012 10000 -1588
rect 9228 -2040 10000 -2012
rect 10240 -1588 11012 -1560
rect 10240 -2012 10928 -1588
rect 10992 -2012 11012 -1588
rect 10240 -2040 11012 -2012
rect 11252 -1588 12024 -1560
rect 11252 -2012 11940 -1588
rect 12004 -2012 12024 -1588
rect 11252 -2040 12024 -2012
rect 12264 -1588 13036 -1560
rect 12264 -2012 12952 -1588
rect 13016 -2012 13036 -1588
rect 12264 -2040 13036 -2012
rect 13276 -1588 14048 -1560
rect 13276 -2012 13964 -1588
rect 14028 -2012 14048 -1588
rect 13276 -2040 14048 -2012
rect 14288 -1588 15060 -1560
rect 14288 -2012 14976 -1588
rect 15040 -2012 15060 -1588
rect 14288 -2040 15060 -2012
rect 15300 -1588 16072 -1560
rect 15300 -2012 15988 -1588
rect 16052 -2012 16072 -1588
rect 15300 -2040 16072 -2012
rect 16312 -1588 17084 -1560
rect 16312 -2012 17000 -1588
rect 17064 -2012 17084 -1588
rect 16312 -2040 17084 -2012
rect -17084 -2308 -16312 -2280
rect -17084 -2732 -16396 -2308
rect -16332 -2732 -16312 -2308
rect -17084 -2760 -16312 -2732
rect -16072 -2308 -15300 -2280
rect -16072 -2732 -15384 -2308
rect -15320 -2732 -15300 -2308
rect -16072 -2760 -15300 -2732
rect -15060 -2308 -14288 -2280
rect -15060 -2732 -14372 -2308
rect -14308 -2732 -14288 -2308
rect -15060 -2760 -14288 -2732
rect -14048 -2308 -13276 -2280
rect -14048 -2732 -13360 -2308
rect -13296 -2732 -13276 -2308
rect -14048 -2760 -13276 -2732
rect -13036 -2308 -12264 -2280
rect -13036 -2732 -12348 -2308
rect -12284 -2732 -12264 -2308
rect -13036 -2760 -12264 -2732
rect -12024 -2308 -11252 -2280
rect -12024 -2732 -11336 -2308
rect -11272 -2732 -11252 -2308
rect -12024 -2760 -11252 -2732
rect -11012 -2308 -10240 -2280
rect -11012 -2732 -10324 -2308
rect -10260 -2732 -10240 -2308
rect -11012 -2760 -10240 -2732
rect -10000 -2308 -9228 -2280
rect -10000 -2732 -9312 -2308
rect -9248 -2732 -9228 -2308
rect -10000 -2760 -9228 -2732
rect -8988 -2308 -8216 -2280
rect -8988 -2732 -8300 -2308
rect -8236 -2732 -8216 -2308
rect -8988 -2760 -8216 -2732
rect -7976 -2308 -7204 -2280
rect -7976 -2732 -7288 -2308
rect -7224 -2732 -7204 -2308
rect -7976 -2760 -7204 -2732
rect -6964 -2308 -6192 -2280
rect -6964 -2732 -6276 -2308
rect -6212 -2732 -6192 -2308
rect -6964 -2760 -6192 -2732
rect -5952 -2308 -5180 -2280
rect -5952 -2732 -5264 -2308
rect -5200 -2732 -5180 -2308
rect -5952 -2760 -5180 -2732
rect -4940 -2308 -4168 -2280
rect -4940 -2732 -4252 -2308
rect -4188 -2732 -4168 -2308
rect -4940 -2760 -4168 -2732
rect -3928 -2308 -3156 -2280
rect -3928 -2732 -3240 -2308
rect -3176 -2732 -3156 -2308
rect -3928 -2760 -3156 -2732
rect -2916 -2308 -2144 -2280
rect -2916 -2732 -2228 -2308
rect -2164 -2732 -2144 -2308
rect -2916 -2760 -2144 -2732
rect -1904 -2308 -1132 -2280
rect -1904 -2732 -1216 -2308
rect -1152 -2732 -1132 -2308
rect -1904 -2760 -1132 -2732
rect -892 -2308 -120 -2280
rect -892 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect -892 -2760 -120 -2732
rect 120 -2308 892 -2280
rect 120 -2732 808 -2308
rect 872 -2732 892 -2308
rect 120 -2760 892 -2732
rect 1132 -2308 1904 -2280
rect 1132 -2732 1820 -2308
rect 1884 -2732 1904 -2308
rect 1132 -2760 1904 -2732
rect 2144 -2308 2916 -2280
rect 2144 -2732 2832 -2308
rect 2896 -2732 2916 -2308
rect 2144 -2760 2916 -2732
rect 3156 -2308 3928 -2280
rect 3156 -2732 3844 -2308
rect 3908 -2732 3928 -2308
rect 3156 -2760 3928 -2732
rect 4168 -2308 4940 -2280
rect 4168 -2732 4856 -2308
rect 4920 -2732 4940 -2308
rect 4168 -2760 4940 -2732
rect 5180 -2308 5952 -2280
rect 5180 -2732 5868 -2308
rect 5932 -2732 5952 -2308
rect 5180 -2760 5952 -2732
rect 6192 -2308 6964 -2280
rect 6192 -2732 6880 -2308
rect 6944 -2732 6964 -2308
rect 6192 -2760 6964 -2732
rect 7204 -2308 7976 -2280
rect 7204 -2732 7892 -2308
rect 7956 -2732 7976 -2308
rect 7204 -2760 7976 -2732
rect 8216 -2308 8988 -2280
rect 8216 -2732 8904 -2308
rect 8968 -2732 8988 -2308
rect 8216 -2760 8988 -2732
rect 9228 -2308 10000 -2280
rect 9228 -2732 9916 -2308
rect 9980 -2732 10000 -2308
rect 9228 -2760 10000 -2732
rect 10240 -2308 11012 -2280
rect 10240 -2732 10928 -2308
rect 10992 -2732 11012 -2308
rect 10240 -2760 11012 -2732
rect 11252 -2308 12024 -2280
rect 11252 -2732 11940 -2308
rect 12004 -2732 12024 -2308
rect 11252 -2760 12024 -2732
rect 12264 -2308 13036 -2280
rect 12264 -2732 12952 -2308
rect 13016 -2732 13036 -2308
rect 12264 -2760 13036 -2732
rect 13276 -2308 14048 -2280
rect 13276 -2732 13964 -2308
rect 14028 -2732 14048 -2308
rect 13276 -2760 14048 -2732
rect 14288 -2308 15060 -2280
rect 14288 -2732 14976 -2308
rect 15040 -2732 15060 -2308
rect 14288 -2760 15060 -2732
rect 15300 -2308 16072 -2280
rect 15300 -2732 15988 -2308
rect 16052 -2732 16072 -2308
rect 15300 -2760 16072 -2732
rect 16312 -2308 17084 -2280
rect 16312 -2732 17000 -2308
rect 17064 -2732 17084 -2308
rect 16312 -2760 17084 -2732
rect -17084 -3028 -16312 -3000
rect -17084 -3452 -16396 -3028
rect -16332 -3452 -16312 -3028
rect -17084 -3480 -16312 -3452
rect -16072 -3028 -15300 -3000
rect -16072 -3452 -15384 -3028
rect -15320 -3452 -15300 -3028
rect -16072 -3480 -15300 -3452
rect -15060 -3028 -14288 -3000
rect -15060 -3452 -14372 -3028
rect -14308 -3452 -14288 -3028
rect -15060 -3480 -14288 -3452
rect -14048 -3028 -13276 -3000
rect -14048 -3452 -13360 -3028
rect -13296 -3452 -13276 -3028
rect -14048 -3480 -13276 -3452
rect -13036 -3028 -12264 -3000
rect -13036 -3452 -12348 -3028
rect -12284 -3452 -12264 -3028
rect -13036 -3480 -12264 -3452
rect -12024 -3028 -11252 -3000
rect -12024 -3452 -11336 -3028
rect -11272 -3452 -11252 -3028
rect -12024 -3480 -11252 -3452
rect -11012 -3028 -10240 -3000
rect -11012 -3452 -10324 -3028
rect -10260 -3452 -10240 -3028
rect -11012 -3480 -10240 -3452
rect -10000 -3028 -9228 -3000
rect -10000 -3452 -9312 -3028
rect -9248 -3452 -9228 -3028
rect -10000 -3480 -9228 -3452
rect -8988 -3028 -8216 -3000
rect -8988 -3452 -8300 -3028
rect -8236 -3452 -8216 -3028
rect -8988 -3480 -8216 -3452
rect -7976 -3028 -7204 -3000
rect -7976 -3452 -7288 -3028
rect -7224 -3452 -7204 -3028
rect -7976 -3480 -7204 -3452
rect -6964 -3028 -6192 -3000
rect -6964 -3452 -6276 -3028
rect -6212 -3452 -6192 -3028
rect -6964 -3480 -6192 -3452
rect -5952 -3028 -5180 -3000
rect -5952 -3452 -5264 -3028
rect -5200 -3452 -5180 -3028
rect -5952 -3480 -5180 -3452
rect -4940 -3028 -4168 -3000
rect -4940 -3452 -4252 -3028
rect -4188 -3452 -4168 -3028
rect -4940 -3480 -4168 -3452
rect -3928 -3028 -3156 -3000
rect -3928 -3452 -3240 -3028
rect -3176 -3452 -3156 -3028
rect -3928 -3480 -3156 -3452
rect -2916 -3028 -2144 -3000
rect -2916 -3452 -2228 -3028
rect -2164 -3452 -2144 -3028
rect -2916 -3480 -2144 -3452
rect -1904 -3028 -1132 -3000
rect -1904 -3452 -1216 -3028
rect -1152 -3452 -1132 -3028
rect -1904 -3480 -1132 -3452
rect -892 -3028 -120 -3000
rect -892 -3452 -204 -3028
rect -140 -3452 -120 -3028
rect -892 -3480 -120 -3452
rect 120 -3028 892 -3000
rect 120 -3452 808 -3028
rect 872 -3452 892 -3028
rect 120 -3480 892 -3452
rect 1132 -3028 1904 -3000
rect 1132 -3452 1820 -3028
rect 1884 -3452 1904 -3028
rect 1132 -3480 1904 -3452
rect 2144 -3028 2916 -3000
rect 2144 -3452 2832 -3028
rect 2896 -3452 2916 -3028
rect 2144 -3480 2916 -3452
rect 3156 -3028 3928 -3000
rect 3156 -3452 3844 -3028
rect 3908 -3452 3928 -3028
rect 3156 -3480 3928 -3452
rect 4168 -3028 4940 -3000
rect 4168 -3452 4856 -3028
rect 4920 -3452 4940 -3028
rect 4168 -3480 4940 -3452
rect 5180 -3028 5952 -3000
rect 5180 -3452 5868 -3028
rect 5932 -3452 5952 -3028
rect 5180 -3480 5952 -3452
rect 6192 -3028 6964 -3000
rect 6192 -3452 6880 -3028
rect 6944 -3452 6964 -3028
rect 6192 -3480 6964 -3452
rect 7204 -3028 7976 -3000
rect 7204 -3452 7892 -3028
rect 7956 -3452 7976 -3028
rect 7204 -3480 7976 -3452
rect 8216 -3028 8988 -3000
rect 8216 -3452 8904 -3028
rect 8968 -3452 8988 -3028
rect 8216 -3480 8988 -3452
rect 9228 -3028 10000 -3000
rect 9228 -3452 9916 -3028
rect 9980 -3452 10000 -3028
rect 9228 -3480 10000 -3452
rect 10240 -3028 11012 -3000
rect 10240 -3452 10928 -3028
rect 10992 -3452 11012 -3028
rect 10240 -3480 11012 -3452
rect 11252 -3028 12024 -3000
rect 11252 -3452 11940 -3028
rect 12004 -3452 12024 -3028
rect 11252 -3480 12024 -3452
rect 12264 -3028 13036 -3000
rect 12264 -3452 12952 -3028
rect 13016 -3452 13036 -3028
rect 12264 -3480 13036 -3452
rect 13276 -3028 14048 -3000
rect 13276 -3452 13964 -3028
rect 14028 -3452 14048 -3028
rect 13276 -3480 14048 -3452
rect 14288 -3028 15060 -3000
rect 14288 -3452 14976 -3028
rect 15040 -3452 15060 -3028
rect 14288 -3480 15060 -3452
rect 15300 -3028 16072 -3000
rect 15300 -3452 15988 -3028
rect 16052 -3452 16072 -3028
rect 15300 -3480 16072 -3452
rect 16312 -3028 17084 -3000
rect 16312 -3452 17000 -3028
rect 17064 -3452 17084 -3028
rect 16312 -3480 17084 -3452
rect -17084 -3748 -16312 -3720
rect -17084 -4172 -16396 -3748
rect -16332 -4172 -16312 -3748
rect -17084 -4200 -16312 -4172
rect -16072 -3748 -15300 -3720
rect -16072 -4172 -15384 -3748
rect -15320 -4172 -15300 -3748
rect -16072 -4200 -15300 -4172
rect -15060 -3748 -14288 -3720
rect -15060 -4172 -14372 -3748
rect -14308 -4172 -14288 -3748
rect -15060 -4200 -14288 -4172
rect -14048 -3748 -13276 -3720
rect -14048 -4172 -13360 -3748
rect -13296 -4172 -13276 -3748
rect -14048 -4200 -13276 -4172
rect -13036 -3748 -12264 -3720
rect -13036 -4172 -12348 -3748
rect -12284 -4172 -12264 -3748
rect -13036 -4200 -12264 -4172
rect -12024 -3748 -11252 -3720
rect -12024 -4172 -11336 -3748
rect -11272 -4172 -11252 -3748
rect -12024 -4200 -11252 -4172
rect -11012 -3748 -10240 -3720
rect -11012 -4172 -10324 -3748
rect -10260 -4172 -10240 -3748
rect -11012 -4200 -10240 -4172
rect -10000 -3748 -9228 -3720
rect -10000 -4172 -9312 -3748
rect -9248 -4172 -9228 -3748
rect -10000 -4200 -9228 -4172
rect -8988 -3748 -8216 -3720
rect -8988 -4172 -8300 -3748
rect -8236 -4172 -8216 -3748
rect -8988 -4200 -8216 -4172
rect -7976 -3748 -7204 -3720
rect -7976 -4172 -7288 -3748
rect -7224 -4172 -7204 -3748
rect -7976 -4200 -7204 -4172
rect -6964 -3748 -6192 -3720
rect -6964 -4172 -6276 -3748
rect -6212 -4172 -6192 -3748
rect -6964 -4200 -6192 -4172
rect -5952 -3748 -5180 -3720
rect -5952 -4172 -5264 -3748
rect -5200 -4172 -5180 -3748
rect -5952 -4200 -5180 -4172
rect -4940 -3748 -4168 -3720
rect -4940 -4172 -4252 -3748
rect -4188 -4172 -4168 -3748
rect -4940 -4200 -4168 -4172
rect -3928 -3748 -3156 -3720
rect -3928 -4172 -3240 -3748
rect -3176 -4172 -3156 -3748
rect -3928 -4200 -3156 -4172
rect -2916 -3748 -2144 -3720
rect -2916 -4172 -2228 -3748
rect -2164 -4172 -2144 -3748
rect -2916 -4200 -2144 -4172
rect -1904 -3748 -1132 -3720
rect -1904 -4172 -1216 -3748
rect -1152 -4172 -1132 -3748
rect -1904 -4200 -1132 -4172
rect -892 -3748 -120 -3720
rect -892 -4172 -204 -3748
rect -140 -4172 -120 -3748
rect -892 -4200 -120 -4172
rect 120 -3748 892 -3720
rect 120 -4172 808 -3748
rect 872 -4172 892 -3748
rect 120 -4200 892 -4172
rect 1132 -3748 1904 -3720
rect 1132 -4172 1820 -3748
rect 1884 -4172 1904 -3748
rect 1132 -4200 1904 -4172
rect 2144 -3748 2916 -3720
rect 2144 -4172 2832 -3748
rect 2896 -4172 2916 -3748
rect 2144 -4200 2916 -4172
rect 3156 -3748 3928 -3720
rect 3156 -4172 3844 -3748
rect 3908 -4172 3928 -3748
rect 3156 -4200 3928 -4172
rect 4168 -3748 4940 -3720
rect 4168 -4172 4856 -3748
rect 4920 -4172 4940 -3748
rect 4168 -4200 4940 -4172
rect 5180 -3748 5952 -3720
rect 5180 -4172 5868 -3748
rect 5932 -4172 5952 -3748
rect 5180 -4200 5952 -4172
rect 6192 -3748 6964 -3720
rect 6192 -4172 6880 -3748
rect 6944 -4172 6964 -3748
rect 6192 -4200 6964 -4172
rect 7204 -3748 7976 -3720
rect 7204 -4172 7892 -3748
rect 7956 -4172 7976 -3748
rect 7204 -4200 7976 -4172
rect 8216 -3748 8988 -3720
rect 8216 -4172 8904 -3748
rect 8968 -4172 8988 -3748
rect 8216 -4200 8988 -4172
rect 9228 -3748 10000 -3720
rect 9228 -4172 9916 -3748
rect 9980 -4172 10000 -3748
rect 9228 -4200 10000 -4172
rect 10240 -3748 11012 -3720
rect 10240 -4172 10928 -3748
rect 10992 -4172 11012 -3748
rect 10240 -4200 11012 -4172
rect 11252 -3748 12024 -3720
rect 11252 -4172 11940 -3748
rect 12004 -4172 12024 -3748
rect 11252 -4200 12024 -4172
rect 12264 -3748 13036 -3720
rect 12264 -4172 12952 -3748
rect 13016 -4172 13036 -3748
rect 12264 -4200 13036 -4172
rect 13276 -3748 14048 -3720
rect 13276 -4172 13964 -3748
rect 14028 -4172 14048 -3748
rect 13276 -4200 14048 -4172
rect 14288 -3748 15060 -3720
rect 14288 -4172 14976 -3748
rect 15040 -4172 15060 -3748
rect 14288 -4200 15060 -4172
rect 15300 -3748 16072 -3720
rect 15300 -4172 15988 -3748
rect 16052 -4172 16072 -3748
rect 15300 -4200 16072 -4172
rect 16312 -3748 17084 -3720
rect 16312 -4172 17000 -3748
rect 17064 -4172 17084 -3748
rect 16312 -4200 17084 -4172
rect -17084 -4468 -16312 -4440
rect -17084 -4892 -16396 -4468
rect -16332 -4892 -16312 -4468
rect -17084 -4920 -16312 -4892
rect -16072 -4468 -15300 -4440
rect -16072 -4892 -15384 -4468
rect -15320 -4892 -15300 -4468
rect -16072 -4920 -15300 -4892
rect -15060 -4468 -14288 -4440
rect -15060 -4892 -14372 -4468
rect -14308 -4892 -14288 -4468
rect -15060 -4920 -14288 -4892
rect -14048 -4468 -13276 -4440
rect -14048 -4892 -13360 -4468
rect -13296 -4892 -13276 -4468
rect -14048 -4920 -13276 -4892
rect -13036 -4468 -12264 -4440
rect -13036 -4892 -12348 -4468
rect -12284 -4892 -12264 -4468
rect -13036 -4920 -12264 -4892
rect -12024 -4468 -11252 -4440
rect -12024 -4892 -11336 -4468
rect -11272 -4892 -11252 -4468
rect -12024 -4920 -11252 -4892
rect -11012 -4468 -10240 -4440
rect -11012 -4892 -10324 -4468
rect -10260 -4892 -10240 -4468
rect -11012 -4920 -10240 -4892
rect -10000 -4468 -9228 -4440
rect -10000 -4892 -9312 -4468
rect -9248 -4892 -9228 -4468
rect -10000 -4920 -9228 -4892
rect -8988 -4468 -8216 -4440
rect -8988 -4892 -8300 -4468
rect -8236 -4892 -8216 -4468
rect -8988 -4920 -8216 -4892
rect -7976 -4468 -7204 -4440
rect -7976 -4892 -7288 -4468
rect -7224 -4892 -7204 -4468
rect -7976 -4920 -7204 -4892
rect -6964 -4468 -6192 -4440
rect -6964 -4892 -6276 -4468
rect -6212 -4892 -6192 -4468
rect -6964 -4920 -6192 -4892
rect -5952 -4468 -5180 -4440
rect -5952 -4892 -5264 -4468
rect -5200 -4892 -5180 -4468
rect -5952 -4920 -5180 -4892
rect -4940 -4468 -4168 -4440
rect -4940 -4892 -4252 -4468
rect -4188 -4892 -4168 -4468
rect -4940 -4920 -4168 -4892
rect -3928 -4468 -3156 -4440
rect -3928 -4892 -3240 -4468
rect -3176 -4892 -3156 -4468
rect -3928 -4920 -3156 -4892
rect -2916 -4468 -2144 -4440
rect -2916 -4892 -2228 -4468
rect -2164 -4892 -2144 -4468
rect -2916 -4920 -2144 -4892
rect -1904 -4468 -1132 -4440
rect -1904 -4892 -1216 -4468
rect -1152 -4892 -1132 -4468
rect -1904 -4920 -1132 -4892
rect -892 -4468 -120 -4440
rect -892 -4892 -204 -4468
rect -140 -4892 -120 -4468
rect -892 -4920 -120 -4892
rect 120 -4468 892 -4440
rect 120 -4892 808 -4468
rect 872 -4892 892 -4468
rect 120 -4920 892 -4892
rect 1132 -4468 1904 -4440
rect 1132 -4892 1820 -4468
rect 1884 -4892 1904 -4468
rect 1132 -4920 1904 -4892
rect 2144 -4468 2916 -4440
rect 2144 -4892 2832 -4468
rect 2896 -4892 2916 -4468
rect 2144 -4920 2916 -4892
rect 3156 -4468 3928 -4440
rect 3156 -4892 3844 -4468
rect 3908 -4892 3928 -4468
rect 3156 -4920 3928 -4892
rect 4168 -4468 4940 -4440
rect 4168 -4892 4856 -4468
rect 4920 -4892 4940 -4468
rect 4168 -4920 4940 -4892
rect 5180 -4468 5952 -4440
rect 5180 -4892 5868 -4468
rect 5932 -4892 5952 -4468
rect 5180 -4920 5952 -4892
rect 6192 -4468 6964 -4440
rect 6192 -4892 6880 -4468
rect 6944 -4892 6964 -4468
rect 6192 -4920 6964 -4892
rect 7204 -4468 7976 -4440
rect 7204 -4892 7892 -4468
rect 7956 -4892 7976 -4468
rect 7204 -4920 7976 -4892
rect 8216 -4468 8988 -4440
rect 8216 -4892 8904 -4468
rect 8968 -4892 8988 -4468
rect 8216 -4920 8988 -4892
rect 9228 -4468 10000 -4440
rect 9228 -4892 9916 -4468
rect 9980 -4892 10000 -4468
rect 9228 -4920 10000 -4892
rect 10240 -4468 11012 -4440
rect 10240 -4892 10928 -4468
rect 10992 -4892 11012 -4468
rect 10240 -4920 11012 -4892
rect 11252 -4468 12024 -4440
rect 11252 -4892 11940 -4468
rect 12004 -4892 12024 -4468
rect 11252 -4920 12024 -4892
rect 12264 -4468 13036 -4440
rect 12264 -4892 12952 -4468
rect 13016 -4892 13036 -4468
rect 12264 -4920 13036 -4892
rect 13276 -4468 14048 -4440
rect 13276 -4892 13964 -4468
rect 14028 -4892 14048 -4468
rect 13276 -4920 14048 -4892
rect 14288 -4468 15060 -4440
rect 14288 -4892 14976 -4468
rect 15040 -4892 15060 -4468
rect 14288 -4920 15060 -4892
rect 15300 -4468 16072 -4440
rect 15300 -4892 15988 -4468
rect 16052 -4892 16072 -4468
rect 15300 -4920 16072 -4892
rect 16312 -4468 17084 -4440
rect 16312 -4892 17000 -4468
rect 17064 -4892 17084 -4468
rect 16312 -4920 17084 -4892
rect -17084 -5188 -16312 -5160
rect -17084 -5612 -16396 -5188
rect -16332 -5612 -16312 -5188
rect -17084 -5640 -16312 -5612
rect -16072 -5188 -15300 -5160
rect -16072 -5612 -15384 -5188
rect -15320 -5612 -15300 -5188
rect -16072 -5640 -15300 -5612
rect -15060 -5188 -14288 -5160
rect -15060 -5612 -14372 -5188
rect -14308 -5612 -14288 -5188
rect -15060 -5640 -14288 -5612
rect -14048 -5188 -13276 -5160
rect -14048 -5612 -13360 -5188
rect -13296 -5612 -13276 -5188
rect -14048 -5640 -13276 -5612
rect -13036 -5188 -12264 -5160
rect -13036 -5612 -12348 -5188
rect -12284 -5612 -12264 -5188
rect -13036 -5640 -12264 -5612
rect -12024 -5188 -11252 -5160
rect -12024 -5612 -11336 -5188
rect -11272 -5612 -11252 -5188
rect -12024 -5640 -11252 -5612
rect -11012 -5188 -10240 -5160
rect -11012 -5612 -10324 -5188
rect -10260 -5612 -10240 -5188
rect -11012 -5640 -10240 -5612
rect -10000 -5188 -9228 -5160
rect -10000 -5612 -9312 -5188
rect -9248 -5612 -9228 -5188
rect -10000 -5640 -9228 -5612
rect -8988 -5188 -8216 -5160
rect -8988 -5612 -8300 -5188
rect -8236 -5612 -8216 -5188
rect -8988 -5640 -8216 -5612
rect -7976 -5188 -7204 -5160
rect -7976 -5612 -7288 -5188
rect -7224 -5612 -7204 -5188
rect -7976 -5640 -7204 -5612
rect -6964 -5188 -6192 -5160
rect -6964 -5612 -6276 -5188
rect -6212 -5612 -6192 -5188
rect -6964 -5640 -6192 -5612
rect -5952 -5188 -5180 -5160
rect -5952 -5612 -5264 -5188
rect -5200 -5612 -5180 -5188
rect -5952 -5640 -5180 -5612
rect -4940 -5188 -4168 -5160
rect -4940 -5612 -4252 -5188
rect -4188 -5612 -4168 -5188
rect -4940 -5640 -4168 -5612
rect -3928 -5188 -3156 -5160
rect -3928 -5612 -3240 -5188
rect -3176 -5612 -3156 -5188
rect -3928 -5640 -3156 -5612
rect -2916 -5188 -2144 -5160
rect -2916 -5612 -2228 -5188
rect -2164 -5612 -2144 -5188
rect -2916 -5640 -2144 -5612
rect -1904 -5188 -1132 -5160
rect -1904 -5612 -1216 -5188
rect -1152 -5612 -1132 -5188
rect -1904 -5640 -1132 -5612
rect -892 -5188 -120 -5160
rect -892 -5612 -204 -5188
rect -140 -5612 -120 -5188
rect -892 -5640 -120 -5612
rect 120 -5188 892 -5160
rect 120 -5612 808 -5188
rect 872 -5612 892 -5188
rect 120 -5640 892 -5612
rect 1132 -5188 1904 -5160
rect 1132 -5612 1820 -5188
rect 1884 -5612 1904 -5188
rect 1132 -5640 1904 -5612
rect 2144 -5188 2916 -5160
rect 2144 -5612 2832 -5188
rect 2896 -5612 2916 -5188
rect 2144 -5640 2916 -5612
rect 3156 -5188 3928 -5160
rect 3156 -5612 3844 -5188
rect 3908 -5612 3928 -5188
rect 3156 -5640 3928 -5612
rect 4168 -5188 4940 -5160
rect 4168 -5612 4856 -5188
rect 4920 -5612 4940 -5188
rect 4168 -5640 4940 -5612
rect 5180 -5188 5952 -5160
rect 5180 -5612 5868 -5188
rect 5932 -5612 5952 -5188
rect 5180 -5640 5952 -5612
rect 6192 -5188 6964 -5160
rect 6192 -5612 6880 -5188
rect 6944 -5612 6964 -5188
rect 6192 -5640 6964 -5612
rect 7204 -5188 7976 -5160
rect 7204 -5612 7892 -5188
rect 7956 -5612 7976 -5188
rect 7204 -5640 7976 -5612
rect 8216 -5188 8988 -5160
rect 8216 -5612 8904 -5188
rect 8968 -5612 8988 -5188
rect 8216 -5640 8988 -5612
rect 9228 -5188 10000 -5160
rect 9228 -5612 9916 -5188
rect 9980 -5612 10000 -5188
rect 9228 -5640 10000 -5612
rect 10240 -5188 11012 -5160
rect 10240 -5612 10928 -5188
rect 10992 -5612 11012 -5188
rect 10240 -5640 11012 -5612
rect 11252 -5188 12024 -5160
rect 11252 -5612 11940 -5188
rect 12004 -5612 12024 -5188
rect 11252 -5640 12024 -5612
rect 12264 -5188 13036 -5160
rect 12264 -5612 12952 -5188
rect 13016 -5612 13036 -5188
rect 12264 -5640 13036 -5612
rect 13276 -5188 14048 -5160
rect 13276 -5612 13964 -5188
rect 14028 -5612 14048 -5188
rect 13276 -5640 14048 -5612
rect 14288 -5188 15060 -5160
rect 14288 -5612 14976 -5188
rect 15040 -5612 15060 -5188
rect 14288 -5640 15060 -5612
rect 15300 -5188 16072 -5160
rect 15300 -5612 15988 -5188
rect 16052 -5612 16072 -5188
rect 15300 -5640 16072 -5612
rect 16312 -5188 17084 -5160
rect 16312 -5612 17000 -5188
rect 17064 -5612 17084 -5188
rect 16312 -5640 17084 -5612
rect -17084 -5908 -16312 -5880
rect -17084 -6332 -16396 -5908
rect -16332 -6332 -16312 -5908
rect -17084 -6360 -16312 -6332
rect -16072 -5908 -15300 -5880
rect -16072 -6332 -15384 -5908
rect -15320 -6332 -15300 -5908
rect -16072 -6360 -15300 -6332
rect -15060 -5908 -14288 -5880
rect -15060 -6332 -14372 -5908
rect -14308 -6332 -14288 -5908
rect -15060 -6360 -14288 -6332
rect -14048 -5908 -13276 -5880
rect -14048 -6332 -13360 -5908
rect -13296 -6332 -13276 -5908
rect -14048 -6360 -13276 -6332
rect -13036 -5908 -12264 -5880
rect -13036 -6332 -12348 -5908
rect -12284 -6332 -12264 -5908
rect -13036 -6360 -12264 -6332
rect -12024 -5908 -11252 -5880
rect -12024 -6332 -11336 -5908
rect -11272 -6332 -11252 -5908
rect -12024 -6360 -11252 -6332
rect -11012 -5908 -10240 -5880
rect -11012 -6332 -10324 -5908
rect -10260 -6332 -10240 -5908
rect -11012 -6360 -10240 -6332
rect -10000 -5908 -9228 -5880
rect -10000 -6332 -9312 -5908
rect -9248 -6332 -9228 -5908
rect -10000 -6360 -9228 -6332
rect -8988 -5908 -8216 -5880
rect -8988 -6332 -8300 -5908
rect -8236 -6332 -8216 -5908
rect -8988 -6360 -8216 -6332
rect -7976 -5908 -7204 -5880
rect -7976 -6332 -7288 -5908
rect -7224 -6332 -7204 -5908
rect -7976 -6360 -7204 -6332
rect -6964 -5908 -6192 -5880
rect -6964 -6332 -6276 -5908
rect -6212 -6332 -6192 -5908
rect -6964 -6360 -6192 -6332
rect -5952 -5908 -5180 -5880
rect -5952 -6332 -5264 -5908
rect -5200 -6332 -5180 -5908
rect -5952 -6360 -5180 -6332
rect -4940 -5908 -4168 -5880
rect -4940 -6332 -4252 -5908
rect -4188 -6332 -4168 -5908
rect -4940 -6360 -4168 -6332
rect -3928 -5908 -3156 -5880
rect -3928 -6332 -3240 -5908
rect -3176 -6332 -3156 -5908
rect -3928 -6360 -3156 -6332
rect -2916 -5908 -2144 -5880
rect -2916 -6332 -2228 -5908
rect -2164 -6332 -2144 -5908
rect -2916 -6360 -2144 -6332
rect -1904 -5908 -1132 -5880
rect -1904 -6332 -1216 -5908
rect -1152 -6332 -1132 -5908
rect -1904 -6360 -1132 -6332
rect -892 -5908 -120 -5880
rect -892 -6332 -204 -5908
rect -140 -6332 -120 -5908
rect -892 -6360 -120 -6332
rect 120 -5908 892 -5880
rect 120 -6332 808 -5908
rect 872 -6332 892 -5908
rect 120 -6360 892 -6332
rect 1132 -5908 1904 -5880
rect 1132 -6332 1820 -5908
rect 1884 -6332 1904 -5908
rect 1132 -6360 1904 -6332
rect 2144 -5908 2916 -5880
rect 2144 -6332 2832 -5908
rect 2896 -6332 2916 -5908
rect 2144 -6360 2916 -6332
rect 3156 -5908 3928 -5880
rect 3156 -6332 3844 -5908
rect 3908 -6332 3928 -5908
rect 3156 -6360 3928 -6332
rect 4168 -5908 4940 -5880
rect 4168 -6332 4856 -5908
rect 4920 -6332 4940 -5908
rect 4168 -6360 4940 -6332
rect 5180 -5908 5952 -5880
rect 5180 -6332 5868 -5908
rect 5932 -6332 5952 -5908
rect 5180 -6360 5952 -6332
rect 6192 -5908 6964 -5880
rect 6192 -6332 6880 -5908
rect 6944 -6332 6964 -5908
rect 6192 -6360 6964 -6332
rect 7204 -5908 7976 -5880
rect 7204 -6332 7892 -5908
rect 7956 -6332 7976 -5908
rect 7204 -6360 7976 -6332
rect 8216 -5908 8988 -5880
rect 8216 -6332 8904 -5908
rect 8968 -6332 8988 -5908
rect 8216 -6360 8988 -6332
rect 9228 -5908 10000 -5880
rect 9228 -6332 9916 -5908
rect 9980 -6332 10000 -5908
rect 9228 -6360 10000 -6332
rect 10240 -5908 11012 -5880
rect 10240 -6332 10928 -5908
rect 10992 -6332 11012 -5908
rect 10240 -6360 11012 -6332
rect 11252 -5908 12024 -5880
rect 11252 -6332 11940 -5908
rect 12004 -6332 12024 -5908
rect 11252 -6360 12024 -6332
rect 12264 -5908 13036 -5880
rect 12264 -6332 12952 -5908
rect 13016 -6332 13036 -5908
rect 12264 -6360 13036 -6332
rect 13276 -5908 14048 -5880
rect 13276 -6332 13964 -5908
rect 14028 -6332 14048 -5908
rect 13276 -6360 14048 -6332
rect 14288 -5908 15060 -5880
rect 14288 -6332 14976 -5908
rect 15040 -6332 15060 -5908
rect 14288 -6360 15060 -6332
rect 15300 -5908 16072 -5880
rect 15300 -6332 15988 -5908
rect 16052 -6332 16072 -5908
rect 15300 -6360 16072 -6332
rect 16312 -5908 17084 -5880
rect 16312 -6332 17000 -5908
rect 17064 -6332 17084 -5908
rect 16312 -6360 17084 -6332
rect -17084 -6628 -16312 -6600
rect -17084 -7052 -16396 -6628
rect -16332 -7052 -16312 -6628
rect -17084 -7080 -16312 -7052
rect -16072 -6628 -15300 -6600
rect -16072 -7052 -15384 -6628
rect -15320 -7052 -15300 -6628
rect -16072 -7080 -15300 -7052
rect -15060 -6628 -14288 -6600
rect -15060 -7052 -14372 -6628
rect -14308 -7052 -14288 -6628
rect -15060 -7080 -14288 -7052
rect -14048 -6628 -13276 -6600
rect -14048 -7052 -13360 -6628
rect -13296 -7052 -13276 -6628
rect -14048 -7080 -13276 -7052
rect -13036 -6628 -12264 -6600
rect -13036 -7052 -12348 -6628
rect -12284 -7052 -12264 -6628
rect -13036 -7080 -12264 -7052
rect -12024 -6628 -11252 -6600
rect -12024 -7052 -11336 -6628
rect -11272 -7052 -11252 -6628
rect -12024 -7080 -11252 -7052
rect -11012 -6628 -10240 -6600
rect -11012 -7052 -10324 -6628
rect -10260 -7052 -10240 -6628
rect -11012 -7080 -10240 -7052
rect -10000 -6628 -9228 -6600
rect -10000 -7052 -9312 -6628
rect -9248 -7052 -9228 -6628
rect -10000 -7080 -9228 -7052
rect -8988 -6628 -8216 -6600
rect -8988 -7052 -8300 -6628
rect -8236 -7052 -8216 -6628
rect -8988 -7080 -8216 -7052
rect -7976 -6628 -7204 -6600
rect -7976 -7052 -7288 -6628
rect -7224 -7052 -7204 -6628
rect -7976 -7080 -7204 -7052
rect -6964 -6628 -6192 -6600
rect -6964 -7052 -6276 -6628
rect -6212 -7052 -6192 -6628
rect -6964 -7080 -6192 -7052
rect -5952 -6628 -5180 -6600
rect -5952 -7052 -5264 -6628
rect -5200 -7052 -5180 -6628
rect -5952 -7080 -5180 -7052
rect -4940 -6628 -4168 -6600
rect -4940 -7052 -4252 -6628
rect -4188 -7052 -4168 -6628
rect -4940 -7080 -4168 -7052
rect -3928 -6628 -3156 -6600
rect -3928 -7052 -3240 -6628
rect -3176 -7052 -3156 -6628
rect -3928 -7080 -3156 -7052
rect -2916 -6628 -2144 -6600
rect -2916 -7052 -2228 -6628
rect -2164 -7052 -2144 -6628
rect -2916 -7080 -2144 -7052
rect -1904 -6628 -1132 -6600
rect -1904 -7052 -1216 -6628
rect -1152 -7052 -1132 -6628
rect -1904 -7080 -1132 -7052
rect -892 -6628 -120 -6600
rect -892 -7052 -204 -6628
rect -140 -7052 -120 -6628
rect -892 -7080 -120 -7052
rect 120 -6628 892 -6600
rect 120 -7052 808 -6628
rect 872 -7052 892 -6628
rect 120 -7080 892 -7052
rect 1132 -6628 1904 -6600
rect 1132 -7052 1820 -6628
rect 1884 -7052 1904 -6628
rect 1132 -7080 1904 -7052
rect 2144 -6628 2916 -6600
rect 2144 -7052 2832 -6628
rect 2896 -7052 2916 -6628
rect 2144 -7080 2916 -7052
rect 3156 -6628 3928 -6600
rect 3156 -7052 3844 -6628
rect 3908 -7052 3928 -6628
rect 3156 -7080 3928 -7052
rect 4168 -6628 4940 -6600
rect 4168 -7052 4856 -6628
rect 4920 -7052 4940 -6628
rect 4168 -7080 4940 -7052
rect 5180 -6628 5952 -6600
rect 5180 -7052 5868 -6628
rect 5932 -7052 5952 -6628
rect 5180 -7080 5952 -7052
rect 6192 -6628 6964 -6600
rect 6192 -7052 6880 -6628
rect 6944 -7052 6964 -6628
rect 6192 -7080 6964 -7052
rect 7204 -6628 7976 -6600
rect 7204 -7052 7892 -6628
rect 7956 -7052 7976 -6628
rect 7204 -7080 7976 -7052
rect 8216 -6628 8988 -6600
rect 8216 -7052 8904 -6628
rect 8968 -7052 8988 -6628
rect 8216 -7080 8988 -7052
rect 9228 -6628 10000 -6600
rect 9228 -7052 9916 -6628
rect 9980 -7052 10000 -6628
rect 9228 -7080 10000 -7052
rect 10240 -6628 11012 -6600
rect 10240 -7052 10928 -6628
rect 10992 -7052 11012 -6628
rect 10240 -7080 11012 -7052
rect 11252 -6628 12024 -6600
rect 11252 -7052 11940 -6628
rect 12004 -7052 12024 -6628
rect 11252 -7080 12024 -7052
rect 12264 -6628 13036 -6600
rect 12264 -7052 12952 -6628
rect 13016 -7052 13036 -6628
rect 12264 -7080 13036 -7052
rect 13276 -6628 14048 -6600
rect 13276 -7052 13964 -6628
rect 14028 -7052 14048 -6628
rect 13276 -7080 14048 -7052
rect 14288 -6628 15060 -6600
rect 14288 -7052 14976 -6628
rect 15040 -7052 15060 -6628
rect 14288 -7080 15060 -7052
rect 15300 -6628 16072 -6600
rect 15300 -7052 15988 -6628
rect 16052 -7052 16072 -6628
rect 15300 -7080 16072 -7052
rect 16312 -6628 17084 -6600
rect 16312 -7052 17000 -6628
rect 17064 -7052 17084 -6628
rect 16312 -7080 17084 -7052
rect -17084 -7348 -16312 -7320
rect -17084 -7772 -16396 -7348
rect -16332 -7772 -16312 -7348
rect -17084 -7800 -16312 -7772
rect -16072 -7348 -15300 -7320
rect -16072 -7772 -15384 -7348
rect -15320 -7772 -15300 -7348
rect -16072 -7800 -15300 -7772
rect -15060 -7348 -14288 -7320
rect -15060 -7772 -14372 -7348
rect -14308 -7772 -14288 -7348
rect -15060 -7800 -14288 -7772
rect -14048 -7348 -13276 -7320
rect -14048 -7772 -13360 -7348
rect -13296 -7772 -13276 -7348
rect -14048 -7800 -13276 -7772
rect -13036 -7348 -12264 -7320
rect -13036 -7772 -12348 -7348
rect -12284 -7772 -12264 -7348
rect -13036 -7800 -12264 -7772
rect -12024 -7348 -11252 -7320
rect -12024 -7772 -11336 -7348
rect -11272 -7772 -11252 -7348
rect -12024 -7800 -11252 -7772
rect -11012 -7348 -10240 -7320
rect -11012 -7772 -10324 -7348
rect -10260 -7772 -10240 -7348
rect -11012 -7800 -10240 -7772
rect -10000 -7348 -9228 -7320
rect -10000 -7772 -9312 -7348
rect -9248 -7772 -9228 -7348
rect -10000 -7800 -9228 -7772
rect -8988 -7348 -8216 -7320
rect -8988 -7772 -8300 -7348
rect -8236 -7772 -8216 -7348
rect -8988 -7800 -8216 -7772
rect -7976 -7348 -7204 -7320
rect -7976 -7772 -7288 -7348
rect -7224 -7772 -7204 -7348
rect -7976 -7800 -7204 -7772
rect -6964 -7348 -6192 -7320
rect -6964 -7772 -6276 -7348
rect -6212 -7772 -6192 -7348
rect -6964 -7800 -6192 -7772
rect -5952 -7348 -5180 -7320
rect -5952 -7772 -5264 -7348
rect -5200 -7772 -5180 -7348
rect -5952 -7800 -5180 -7772
rect -4940 -7348 -4168 -7320
rect -4940 -7772 -4252 -7348
rect -4188 -7772 -4168 -7348
rect -4940 -7800 -4168 -7772
rect -3928 -7348 -3156 -7320
rect -3928 -7772 -3240 -7348
rect -3176 -7772 -3156 -7348
rect -3928 -7800 -3156 -7772
rect -2916 -7348 -2144 -7320
rect -2916 -7772 -2228 -7348
rect -2164 -7772 -2144 -7348
rect -2916 -7800 -2144 -7772
rect -1904 -7348 -1132 -7320
rect -1904 -7772 -1216 -7348
rect -1152 -7772 -1132 -7348
rect -1904 -7800 -1132 -7772
rect -892 -7348 -120 -7320
rect -892 -7772 -204 -7348
rect -140 -7772 -120 -7348
rect -892 -7800 -120 -7772
rect 120 -7348 892 -7320
rect 120 -7772 808 -7348
rect 872 -7772 892 -7348
rect 120 -7800 892 -7772
rect 1132 -7348 1904 -7320
rect 1132 -7772 1820 -7348
rect 1884 -7772 1904 -7348
rect 1132 -7800 1904 -7772
rect 2144 -7348 2916 -7320
rect 2144 -7772 2832 -7348
rect 2896 -7772 2916 -7348
rect 2144 -7800 2916 -7772
rect 3156 -7348 3928 -7320
rect 3156 -7772 3844 -7348
rect 3908 -7772 3928 -7348
rect 3156 -7800 3928 -7772
rect 4168 -7348 4940 -7320
rect 4168 -7772 4856 -7348
rect 4920 -7772 4940 -7348
rect 4168 -7800 4940 -7772
rect 5180 -7348 5952 -7320
rect 5180 -7772 5868 -7348
rect 5932 -7772 5952 -7348
rect 5180 -7800 5952 -7772
rect 6192 -7348 6964 -7320
rect 6192 -7772 6880 -7348
rect 6944 -7772 6964 -7348
rect 6192 -7800 6964 -7772
rect 7204 -7348 7976 -7320
rect 7204 -7772 7892 -7348
rect 7956 -7772 7976 -7348
rect 7204 -7800 7976 -7772
rect 8216 -7348 8988 -7320
rect 8216 -7772 8904 -7348
rect 8968 -7772 8988 -7348
rect 8216 -7800 8988 -7772
rect 9228 -7348 10000 -7320
rect 9228 -7772 9916 -7348
rect 9980 -7772 10000 -7348
rect 9228 -7800 10000 -7772
rect 10240 -7348 11012 -7320
rect 10240 -7772 10928 -7348
rect 10992 -7772 11012 -7348
rect 10240 -7800 11012 -7772
rect 11252 -7348 12024 -7320
rect 11252 -7772 11940 -7348
rect 12004 -7772 12024 -7348
rect 11252 -7800 12024 -7772
rect 12264 -7348 13036 -7320
rect 12264 -7772 12952 -7348
rect 13016 -7772 13036 -7348
rect 12264 -7800 13036 -7772
rect 13276 -7348 14048 -7320
rect 13276 -7772 13964 -7348
rect 14028 -7772 14048 -7348
rect 13276 -7800 14048 -7772
rect 14288 -7348 15060 -7320
rect 14288 -7772 14976 -7348
rect 15040 -7772 15060 -7348
rect 14288 -7800 15060 -7772
rect 15300 -7348 16072 -7320
rect 15300 -7772 15988 -7348
rect 16052 -7772 16072 -7348
rect 15300 -7800 16072 -7772
rect 16312 -7348 17084 -7320
rect 16312 -7772 17000 -7348
rect 17064 -7772 17084 -7348
rect 16312 -7800 17084 -7772
rect -17084 -8068 -16312 -8040
rect -17084 -8492 -16396 -8068
rect -16332 -8492 -16312 -8068
rect -17084 -8520 -16312 -8492
rect -16072 -8068 -15300 -8040
rect -16072 -8492 -15384 -8068
rect -15320 -8492 -15300 -8068
rect -16072 -8520 -15300 -8492
rect -15060 -8068 -14288 -8040
rect -15060 -8492 -14372 -8068
rect -14308 -8492 -14288 -8068
rect -15060 -8520 -14288 -8492
rect -14048 -8068 -13276 -8040
rect -14048 -8492 -13360 -8068
rect -13296 -8492 -13276 -8068
rect -14048 -8520 -13276 -8492
rect -13036 -8068 -12264 -8040
rect -13036 -8492 -12348 -8068
rect -12284 -8492 -12264 -8068
rect -13036 -8520 -12264 -8492
rect -12024 -8068 -11252 -8040
rect -12024 -8492 -11336 -8068
rect -11272 -8492 -11252 -8068
rect -12024 -8520 -11252 -8492
rect -11012 -8068 -10240 -8040
rect -11012 -8492 -10324 -8068
rect -10260 -8492 -10240 -8068
rect -11012 -8520 -10240 -8492
rect -10000 -8068 -9228 -8040
rect -10000 -8492 -9312 -8068
rect -9248 -8492 -9228 -8068
rect -10000 -8520 -9228 -8492
rect -8988 -8068 -8216 -8040
rect -8988 -8492 -8300 -8068
rect -8236 -8492 -8216 -8068
rect -8988 -8520 -8216 -8492
rect -7976 -8068 -7204 -8040
rect -7976 -8492 -7288 -8068
rect -7224 -8492 -7204 -8068
rect -7976 -8520 -7204 -8492
rect -6964 -8068 -6192 -8040
rect -6964 -8492 -6276 -8068
rect -6212 -8492 -6192 -8068
rect -6964 -8520 -6192 -8492
rect -5952 -8068 -5180 -8040
rect -5952 -8492 -5264 -8068
rect -5200 -8492 -5180 -8068
rect -5952 -8520 -5180 -8492
rect -4940 -8068 -4168 -8040
rect -4940 -8492 -4252 -8068
rect -4188 -8492 -4168 -8068
rect -4940 -8520 -4168 -8492
rect -3928 -8068 -3156 -8040
rect -3928 -8492 -3240 -8068
rect -3176 -8492 -3156 -8068
rect -3928 -8520 -3156 -8492
rect -2916 -8068 -2144 -8040
rect -2916 -8492 -2228 -8068
rect -2164 -8492 -2144 -8068
rect -2916 -8520 -2144 -8492
rect -1904 -8068 -1132 -8040
rect -1904 -8492 -1216 -8068
rect -1152 -8492 -1132 -8068
rect -1904 -8520 -1132 -8492
rect -892 -8068 -120 -8040
rect -892 -8492 -204 -8068
rect -140 -8492 -120 -8068
rect -892 -8520 -120 -8492
rect 120 -8068 892 -8040
rect 120 -8492 808 -8068
rect 872 -8492 892 -8068
rect 120 -8520 892 -8492
rect 1132 -8068 1904 -8040
rect 1132 -8492 1820 -8068
rect 1884 -8492 1904 -8068
rect 1132 -8520 1904 -8492
rect 2144 -8068 2916 -8040
rect 2144 -8492 2832 -8068
rect 2896 -8492 2916 -8068
rect 2144 -8520 2916 -8492
rect 3156 -8068 3928 -8040
rect 3156 -8492 3844 -8068
rect 3908 -8492 3928 -8068
rect 3156 -8520 3928 -8492
rect 4168 -8068 4940 -8040
rect 4168 -8492 4856 -8068
rect 4920 -8492 4940 -8068
rect 4168 -8520 4940 -8492
rect 5180 -8068 5952 -8040
rect 5180 -8492 5868 -8068
rect 5932 -8492 5952 -8068
rect 5180 -8520 5952 -8492
rect 6192 -8068 6964 -8040
rect 6192 -8492 6880 -8068
rect 6944 -8492 6964 -8068
rect 6192 -8520 6964 -8492
rect 7204 -8068 7976 -8040
rect 7204 -8492 7892 -8068
rect 7956 -8492 7976 -8068
rect 7204 -8520 7976 -8492
rect 8216 -8068 8988 -8040
rect 8216 -8492 8904 -8068
rect 8968 -8492 8988 -8068
rect 8216 -8520 8988 -8492
rect 9228 -8068 10000 -8040
rect 9228 -8492 9916 -8068
rect 9980 -8492 10000 -8068
rect 9228 -8520 10000 -8492
rect 10240 -8068 11012 -8040
rect 10240 -8492 10928 -8068
rect 10992 -8492 11012 -8068
rect 10240 -8520 11012 -8492
rect 11252 -8068 12024 -8040
rect 11252 -8492 11940 -8068
rect 12004 -8492 12024 -8068
rect 11252 -8520 12024 -8492
rect 12264 -8068 13036 -8040
rect 12264 -8492 12952 -8068
rect 13016 -8492 13036 -8068
rect 12264 -8520 13036 -8492
rect 13276 -8068 14048 -8040
rect 13276 -8492 13964 -8068
rect 14028 -8492 14048 -8068
rect 13276 -8520 14048 -8492
rect 14288 -8068 15060 -8040
rect 14288 -8492 14976 -8068
rect 15040 -8492 15060 -8068
rect 14288 -8520 15060 -8492
rect 15300 -8068 16072 -8040
rect 15300 -8492 15988 -8068
rect 16052 -8492 16072 -8068
rect 15300 -8520 16072 -8492
rect 16312 -8068 17084 -8040
rect 16312 -8492 17000 -8068
rect 17064 -8492 17084 -8068
rect 16312 -8520 17084 -8492
rect -17084 -8788 -16312 -8760
rect -17084 -9212 -16396 -8788
rect -16332 -9212 -16312 -8788
rect -17084 -9240 -16312 -9212
rect -16072 -8788 -15300 -8760
rect -16072 -9212 -15384 -8788
rect -15320 -9212 -15300 -8788
rect -16072 -9240 -15300 -9212
rect -15060 -8788 -14288 -8760
rect -15060 -9212 -14372 -8788
rect -14308 -9212 -14288 -8788
rect -15060 -9240 -14288 -9212
rect -14048 -8788 -13276 -8760
rect -14048 -9212 -13360 -8788
rect -13296 -9212 -13276 -8788
rect -14048 -9240 -13276 -9212
rect -13036 -8788 -12264 -8760
rect -13036 -9212 -12348 -8788
rect -12284 -9212 -12264 -8788
rect -13036 -9240 -12264 -9212
rect -12024 -8788 -11252 -8760
rect -12024 -9212 -11336 -8788
rect -11272 -9212 -11252 -8788
rect -12024 -9240 -11252 -9212
rect -11012 -8788 -10240 -8760
rect -11012 -9212 -10324 -8788
rect -10260 -9212 -10240 -8788
rect -11012 -9240 -10240 -9212
rect -10000 -8788 -9228 -8760
rect -10000 -9212 -9312 -8788
rect -9248 -9212 -9228 -8788
rect -10000 -9240 -9228 -9212
rect -8988 -8788 -8216 -8760
rect -8988 -9212 -8300 -8788
rect -8236 -9212 -8216 -8788
rect -8988 -9240 -8216 -9212
rect -7976 -8788 -7204 -8760
rect -7976 -9212 -7288 -8788
rect -7224 -9212 -7204 -8788
rect -7976 -9240 -7204 -9212
rect -6964 -8788 -6192 -8760
rect -6964 -9212 -6276 -8788
rect -6212 -9212 -6192 -8788
rect -6964 -9240 -6192 -9212
rect -5952 -8788 -5180 -8760
rect -5952 -9212 -5264 -8788
rect -5200 -9212 -5180 -8788
rect -5952 -9240 -5180 -9212
rect -4940 -8788 -4168 -8760
rect -4940 -9212 -4252 -8788
rect -4188 -9212 -4168 -8788
rect -4940 -9240 -4168 -9212
rect -3928 -8788 -3156 -8760
rect -3928 -9212 -3240 -8788
rect -3176 -9212 -3156 -8788
rect -3928 -9240 -3156 -9212
rect -2916 -8788 -2144 -8760
rect -2916 -9212 -2228 -8788
rect -2164 -9212 -2144 -8788
rect -2916 -9240 -2144 -9212
rect -1904 -8788 -1132 -8760
rect -1904 -9212 -1216 -8788
rect -1152 -9212 -1132 -8788
rect -1904 -9240 -1132 -9212
rect -892 -8788 -120 -8760
rect -892 -9212 -204 -8788
rect -140 -9212 -120 -8788
rect -892 -9240 -120 -9212
rect 120 -8788 892 -8760
rect 120 -9212 808 -8788
rect 872 -9212 892 -8788
rect 120 -9240 892 -9212
rect 1132 -8788 1904 -8760
rect 1132 -9212 1820 -8788
rect 1884 -9212 1904 -8788
rect 1132 -9240 1904 -9212
rect 2144 -8788 2916 -8760
rect 2144 -9212 2832 -8788
rect 2896 -9212 2916 -8788
rect 2144 -9240 2916 -9212
rect 3156 -8788 3928 -8760
rect 3156 -9212 3844 -8788
rect 3908 -9212 3928 -8788
rect 3156 -9240 3928 -9212
rect 4168 -8788 4940 -8760
rect 4168 -9212 4856 -8788
rect 4920 -9212 4940 -8788
rect 4168 -9240 4940 -9212
rect 5180 -8788 5952 -8760
rect 5180 -9212 5868 -8788
rect 5932 -9212 5952 -8788
rect 5180 -9240 5952 -9212
rect 6192 -8788 6964 -8760
rect 6192 -9212 6880 -8788
rect 6944 -9212 6964 -8788
rect 6192 -9240 6964 -9212
rect 7204 -8788 7976 -8760
rect 7204 -9212 7892 -8788
rect 7956 -9212 7976 -8788
rect 7204 -9240 7976 -9212
rect 8216 -8788 8988 -8760
rect 8216 -9212 8904 -8788
rect 8968 -9212 8988 -8788
rect 8216 -9240 8988 -9212
rect 9228 -8788 10000 -8760
rect 9228 -9212 9916 -8788
rect 9980 -9212 10000 -8788
rect 9228 -9240 10000 -9212
rect 10240 -8788 11012 -8760
rect 10240 -9212 10928 -8788
rect 10992 -9212 11012 -8788
rect 10240 -9240 11012 -9212
rect 11252 -8788 12024 -8760
rect 11252 -9212 11940 -8788
rect 12004 -9212 12024 -8788
rect 11252 -9240 12024 -9212
rect 12264 -8788 13036 -8760
rect 12264 -9212 12952 -8788
rect 13016 -9212 13036 -8788
rect 12264 -9240 13036 -9212
rect 13276 -8788 14048 -8760
rect 13276 -9212 13964 -8788
rect 14028 -9212 14048 -8788
rect 13276 -9240 14048 -9212
rect 14288 -8788 15060 -8760
rect 14288 -9212 14976 -8788
rect 15040 -9212 15060 -8788
rect 14288 -9240 15060 -9212
rect 15300 -8788 16072 -8760
rect 15300 -9212 15988 -8788
rect 16052 -9212 16072 -8788
rect 15300 -9240 16072 -9212
rect 16312 -8788 17084 -8760
rect 16312 -9212 17000 -8788
rect 17064 -9212 17084 -8788
rect 16312 -9240 17084 -9212
rect -17084 -9508 -16312 -9480
rect -17084 -9932 -16396 -9508
rect -16332 -9932 -16312 -9508
rect -17084 -9960 -16312 -9932
rect -16072 -9508 -15300 -9480
rect -16072 -9932 -15384 -9508
rect -15320 -9932 -15300 -9508
rect -16072 -9960 -15300 -9932
rect -15060 -9508 -14288 -9480
rect -15060 -9932 -14372 -9508
rect -14308 -9932 -14288 -9508
rect -15060 -9960 -14288 -9932
rect -14048 -9508 -13276 -9480
rect -14048 -9932 -13360 -9508
rect -13296 -9932 -13276 -9508
rect -14048 -9960 -13276 -9932
rect -13036 -9508 -12264 -9480
rect -13036 -9932 -12348 -9508
rect -12284 -9932 -12264 -9508
rect -13036 -9960 -12264 -9932
rect -12024 -9508 -11252 -9480
rect -12024 -9932 -11336 -9508
rect -11272 -9932 -11252 -9508
rect -12024 -9960 -11252 -9932
rect -11012 -9508 -10240 -9480
rect -11012 -9932 -10324 -9508
rect -10260 -9932 -10240 -9508
rect -11012 -9960 -10240 -9932
rect -10000 -9508 -9228 -9480
rect -10000 -9932 -9312 -9508
rect -9248 -9932 -9228 -9508
rect -10000 -9960 -9228 -9932
rect -8988 -9508 -8216 -9480
rect -8988 -9932 -8300 -9508
rect -8236 -9932 -8216 -9508
rect -8988 -9960 -8216 -9932
rect -7976 -9508 -7204 -9480
rect -7976 -9932 -7288 -9508
rect -7224 -9932 -7204 -9508
rect -7976 -9960 -7204 -9932
rect -6964 -9508 -6192 -9480
rect -6964 -9932 -6276 -9508
rect -6212 -9932 -6192 -9508
rect -6964 -9960 -6192 -9932
rect -5952 -9508 -5180 -9480
rect -5952 -9932 -5264 -9508
rect -5200 -9932 -5180 -9508
rect -5952 -9960 -5180 -9932
rect -4940 -9508 -4168 -9480
rect -4940 -9932 -4252 -9508
rect -4188 -9932 -4168 -9508
rect -4940 -9960 -4168 -9932
rect -3928 -9508 -3156 -9480
rect -3928 -9932 -3240 -9508
rect -3176 -9932 -3156 -9508
rect -3928 -9960 -3156 -9932
rect -2916 -9508 -2144 -9480
rect -2916 -9932 -2228 -9508
rect -2164 -9932 -2144 -9508
rect -2916 -9960 -2144 -9932
rect -1904 -9508 -1132 -9480
rect -1904 -9932 -1216 -9508
rect -1152 -9932 -1132 -9508
rect -1904 -9960 -1132 -9932
rect -892 -9508 -120 -9480
rect -892 -9932 -204 -9508
rect -140 -9932 -120 -9508
rect -892 -9960 -120 -9932
rect 120 -9508 892 -9480
rect 120 -9932 808 -9508
rect 872 -9932 892 -9508
rect 120 -9960 892 -9932
rect 1132 -9508 1904 -9480
rect 1132 -9932 1820 -9508
rect 1884 -9932 1904 -9508
rect 1132 -9960 1904 -9932
rect 2144 -9508 2916 -9480
rect 2144 -9932 2832 -9508
rect 2896 -9932 2916 -9508
rect 2144 -9960 2916 -9932
rect 3156 -9508 3928 -9480
rect 3156 -9932 3844 -9508
rect 3908 -9932 3928 -9508
rect 3156 -9960 3928 -9932
rect 4168 -9508 4940 -9480
rect 4168 -9932 4856 -9508
rect 4920 -9932 4940 -9508
rect 4168 -9960 4940 -9932
rect 5180 -9508 5952 -9480
rect 5180 -9932 5868 -9508
rect 5932 -9932 5952 -9508
rect 5180 -9960 5952 -9932
rect 6192 -9508 6964 -9480
rect 6192 -9932 6880 -9508
rect 6944 -9932 6964 -9508
rect 6192 -9960 6964 -9932
rect 7204 -9508 7976 -9480
rect 7204 -9932 7892 -9508
rect 7956 -9932 7976 -9508
rect 7204 -9960 7976 -9932
rect 8216 -9508 8988 -9480
rect 8216 -9932 8904 -9508
rect 8968 -9932 8988 -9508
rect 8216 -9960 8988 -9932
rect 9228 -9508 10000 -9480
rect 9228 -9932 9916 -9508
rect 9980 -9932 10000 -9508
rect 9228 -9960 10000 -9932
rect 10240 -9508 11012 -9480
rect 10240 -9932 10928 -9508
rect 10992 -9932 11012 -9508
rect 10240 -9960 11012 -9932
rect 11252 -9508 12024 -9480
rect 11252 -9932 11940 -9508
rect 12004 -9932 12024 -9508
rect 11252 -9960 12024 -9932
rect 12264 -9508 13036 -9480
rect 12264 -9932 12952 -9508
rect 13016 -9932 13036 -9508
rect 12264 -9960 13036 -9932
rect 13276 -9508 14048 -9480
rect 13276 -9932 13964 -9508
rect 14028 -9932 14048 -9508
rect 13276 -9960 14048 -9932
rect 14288 -9508 15060 -9480
rect 14288 -9932 14976 -9508
rect 15040 -9932 15060 -9508
rect 14288 -9960 15060 -9932
rect 15300 -9508 16072 -9480
rect 15300 -9932 15988 -9508
rect 16052 -9932 16072 -9508
rect 15300 -9960 16072 -9932
rect 16312 -9508 17084 -9480
rect 16312 -9932 17000 -9508
rect 17064 -9932 17084 -9508
rect 16312 -9960 17084 -9932
rect -17084 -10228 -16312 -10200
rect -17084 -10652 -16396 -10228
rect -16332 -10652 -16312 -10228
rect -17084 -10680 -16312 -10652
rect -16072 -10228 -15300 -10200
rect -16072 -10652 -15384 -10228
rect -15320 -10652 -15300 -10228
rect -16072 -10680 -15300 -10652
rect -15060 -10228 -14288 -10200
rect -15060 -10652 -14372 -10228
rect -14308 -10652 -14288 -10228
rect -15060 -10680 -14288 -10652
rect -14048 -10228 -13276 -10200
rect -14048 -10652 -13360 -10228
rect -13296 -10652 -13276 -10228
rect -14048 -10680 -13276 -10652
rect -13036 -10228 -12264 -10200
rect -13036 -10652 -12348 -10228
rect -12284 -10652 -12264 -10228
rect -13036 -10680 -12264 -10652
rect -12024 -10228 -11252 -10200
rect -12024 -10652 -11336 -10228
rect -11272 -10652 -11252 -10228
rect -12024 -10680 -11252 -10652
rect -11012 -10228 -10240 -10200
rect -11012 -10652 -10324 -10228
rect -10260 -10652 -10240 -10228
rect -11012 -10680 -10240 -10652
rect -10000 -10228 -9228 -10200
rect -10000 -10652 -9312 -10228
rect -9248 -10652 -9228 -10228
rect -10000 -10680 -9228 -10652
rect -8988 -10228 -8216 -10200
rect -8988 -10652 -8300 -10228
rect -8236 -10652 -8216 -10228
rect -8988 -10680 -8216 -10652
rect -7976 -10228 -7204 -10200
rect -7976 -10652 -7288 -10228
rect -7224 -10652 -7204 -10228
rect -7976 -10680 -7204 -10652
rect -6964 -10228 -6192 -10200
rect -6964 -10652 -6276 -10228
rect -6212 -10652 -6192 -10228
rect -6964 -10680 -6192 -10652
rect -5952 -10228 -5180 -10200
rect -5952 -10652 -5264 -10228
rect -5200 -10652 -5180 -10228
rect -5952 -10680 -5180 -10652
rect -4940 -10228 -4168 -10200
rect -4940 -10652 -4252 -10228
rect -4188 -10652 -4168 -10228
rect -4940 -10680 -4168 -10652
rect -3928 -10228 -3156 -10200
rect -3928 -10652 -3240 -10228
rect -3176 -10652 -3156 -10228
rect -3928 -10680 -3156 -10652
rect -2916 -10228 -2144 -10200
rect -2916 -10652 -2228 -10228
rect -2164 -10652 -2144 -10228
rect -2916 -10680 -2144 -10652
rect -1904 -10228 -1132 -10200
rect -1904 -10652 -1216 -10228
rect -1152 -10652 -1132 -10228
rect -1904 -10680 -1132 -10652
rect -892 -10228 -120 -10200
rect -892 -10652 -204 -10228
rect -140 -10652 -120 -10228
rect -892 -10680 -120 -10652
rect 120 -10228 892 -10200
rect 120 -10652 808 -10228
rect 872 -10652 892 -10228
rect 120 -10680 892 -10652
rect 1132 -10228 1904 -10200
rect 1132 -10652 1820 -10228
rect 1884 -10652 1904 -10228
rect 1132 -10680 1904 -10652
rect 2144 -10228 2916 -10200
rect 2144 -10652 2832 -10228
rect 2896 -10652 2916 -10228
rect 2144 -10680 2916 -10652
rect 3156 -10228 3928 -10200
rect 3156 -10652 3844 -10228
rect 3908 -10652 3928 -10228
rect 3156 -10680 3928 -10652
rect 4168 -10228 4940 -10200
rect 4168 -10652 4856 -10228
rect 4920 -10652 4940 -10228
rect 4168 -10680 4940 -10652
rect 5180 -10228 5952 -10200
rect 5180 -10652 5868 -10228
rect 5932 -10652 5952 -10228
rect 5180 -10680 5952 -10652
rect 6192 -10228 6964 -10200
rect 6192 -10652 6880 -10228
rect 6944 -10652 6964 -10228
rect 6192 -10680 6964 -10652
rect 7204 -10228 7976 -10200
rect 7204 -10652 7892 -10228
rect 7956 -10652 7976 -10228
rect 7204 -10680 7976 -10652
rect 8216 -10228 8988 -10200
rect 8216 -10652 8904 -10228
rect 8968 -10652 8988 -10228
rect 8216 -10680 8988 -10652
rect 9228 -10228 10000 -10200
rect 9228 -10652 9916 -10228
rect 9980 -10652 10000 -10228
rect 9228 -10680 10000 -10652
rect 10240 -10228 11012 -10200
rect 10240 -10652 10928 -10228
rect 10992 -10652 11012 -10228
rect 10240 -10680 11012 -10652
rect 11252 -10228 12024 -10200
rect 11252 -10652 11940 -10228
rect 12004 -10652 12024 -10228
rect 11252 -10680 12024 -10652
rect 12264 -10228 13036 -10200
rect 12264 -10652 12952 -10228
rect 13016 -10652 13036 -10228
rect 12264 -10680 13036 -10652
rect 13276 -10228 14048 -10200
rect 13276 -10652 13964 -10228
rect 14028 -10652 14048 -10228
rect 13276 -10680 14048 -10652
rect 14288 -10228 15060 -10200
rect 14288 -10652 14976 -10228
rect 15040 -10652 15060 -10228
rect 14288 -10680 15060 -10652
rect 15300 -10228 16072 -10200
rect 15300 -10652 15988 -10228
rect 16052 -10652 16072 -10228
rect 15300 -10680 16072 -10652
rect 16312 -10228 17084 -10200
rect 16312 -10652 17000 -10228
rect 17064 -10652 17084 -10228
rect 16312 -10680 17084 -10652
rect -17084 -10948 -16312 -10920
rect -17084 -11372 -16396 -10948
rect -16332 -11372 -16312 -10948
rect -17084 -11400 -16312 -11372
rect -16072 -10948 -15300 -10920
rect -16072 -11372 -15384 -10948
rect -15320 -11372 -15300 -10948
rect -16072 -11400 -15300 -11372
rect -15060 -10948 -14288 -10920
rect -15060 -11372 -14372 -10948
rect -14308 -11372 -14288 -10948
rect -15060 -11400 -14288 -11372
rect -14048 -10948 -13276 -10920
rect -14048 -11372 -13360 -10948
rect -13296 -11372 -13276 -10948
rect -14048 -11400 -13276 -11372
rect -13036 -10948 -12264 -10920
rect -13036 -11372 -12348 -10948
rect -12284 -11372 -12264 -10948
rect -13036 -11400 -12264 -11372
rect -12024 -10948 -11252 -10920
rect -12024 -11372 -11336 -10948
rect -11272 -11372 -11252 -10948
rect -12024 -11400 -11252 -11372
rect -11012 -10948 -10240 -10920
rect -11012 -11372 -10324 -10948
rect -10260 -11372 -10240 -10948
rect -11012 -11400 -10240 -11372
rect -10000 -10948 -9228 -10920
rect -10000 -11372 -9312 -10948
rect -9248 -11372 -9228 -10948
rect -10000 -11400 -9228 -11372
rect -8988 -10948 -8216 -10920
rect -8988 -11372 -8300 -10948
rect -8236 -11372 -8216 -10948
rect -8988 -11400 -8216 -11372
rect -7976 -10948 -7204 -10920
rect -7976 -11372 -7288 -10948
rect -7224 -11372 -7204 -10948
rect -7976 -11400 -7204 -11372
rect -6964 -10948 -6192 -10920
rect -6964 -11372 -6276 -10948
rect -6212 -11372 -6192 -10948
rect -6964 -11400 -6192 -11372
rect -5952 -10948 -5180 -10920
rect -5952 -11372 -5264 -10948
rect -5200 -11372 -5180 -10948
rect -5952 -11400 -5180 -11372
rect -4940 -10948 -4168 -10920
rect -4940 -11372 -4252 -10948
rect -4188 -11372 -4168 -10948
rect -4940 -11400 -4168 -11372
rect -3928 -10948 -3156 -10920
rect -3928 -11372 -3240 -10948
rect -3176 -11372 -3156 -10948
rect -3928 -11400 -3156 -11372
rect -2916 -10948 -2144 -10920
rect -2916 -11372 -2228 -10948
rect -2164 -11372 -2144 -10948
rect -2916 -11400 -2144 -11372
rect -1904 -10948 -1132 -10920
rect -1904 -11372 -1216 -10948
rect -1152 -11372 -1132 -10948
rect -1904 -11400 -1132 -11372
rect -892 -10948 -120 -10920
rect -892 -11372 -204 -10948
rect -140 -11372 -120 -10948
rect -892 -11400 -120 -11372
rect 120 -10948 892 -10920
rect 120 -11372 808 -10948
rect 872 -11372 892 -10948
rect 120 -11400 892 -11372
rect 1132 -10948 1904 -10920
rect 1132 -11372 1820 -10948
rect 1884 -11372 1904 -10948
rect 1132 -11400 1904 -11372
rect 2144 -10948 2916 -10920
rect 2144 -11372 2832 -10948
rect 2896 -11372 2916 -10948
rect 2144 -11400 2916 -11372
rect 3156 -10948 3928 -10920
rect 3156 -11372 3844 -10948
rect 3908 -11372 3928 -10948
rect 3156 -11400 3928 -11372
rect 4168 -10948 4940 -10920
rect 4168 -11372 4856 -10948
rect 4920 -11372 4940 -10948
rect 4168 -11400 4940 -11372
rect 5180 -10948 5952 -10920
rect 5180 -11372 5868 -10948
rect 5932 -11372 5952 -10948
rect 5180 -11400 5952 -11372
rect 6192 -10948 6964 -10920
rect 6192 -11372 6880 -10948
rect 6944 -11372 6964 -10948
rect 6192 -11400 6964 -11372
rect 7204 -10948 7976 -10920
rect 7204 -11372 7892 -10948
rect 7956 -11372 7976 -10948
rect 7204 -11400 7976 -11372
rect 8216 -10948 8988 -10920
rect 8216 -11372 8904 -10948
rect 8968 -11372 8988 -10948
rect 8216 -11400 8988 -11372
rect 9228 -10948 10000 -10920
rect 9228 -11372 9916 -10948
rect 9980 -11372 10000 -10948
rect 9228 -11400 10000 -11372
rect 10240 -10948 11012 -10920
rect 10240 -11372 10928 -10948
rect 10992 -11372 11012 -10948
rect 10240 -11400 11012 -11372
rect 11252 -10948 12024 -10920
rect 11252 -11372 11940 -10948
rect 12004 -11372 12024 -10948
rect 11252 -11400 12024 -11372
rect 12264 -10948 13036 -10920
rect 12264 -11372 12952 -10948
rect 13016 -11372 13036 -10948
rect 12264 -11400 13036 -11372
rect 13276 -10948 14048 -10920
rect 13276 -11372 13964 -10948
rect 14028 -11372 14048 -10948
rect 13276 -11400 14048 -11372
rect 14288 -10948 15060 -10920
rect 14288 -11372 14976 -10948
rect 15040 -11372 15060 -10948
rect 14288 -11400 15060 -11372
rect 15300 -10948 16072 -10920
rect 15300 -11372 15988 -10948
rect 16052 -11372 16072 -10948
rect 15300 -11400 16072 -11372
rect 16312 -10948 17084 -10920
rect 16312 -11372 17000 -10948
rect 17064 -11372 17084 -10948
rect 16312 -11400 17084 -11372
<< via3 >>
rect -16396 10948 -16332 11372
rect -15384 10948 -15320 11372
rect -14372 10948 -14308 11372
rect -13360 10948 -13296 11372
rect -12348 10948 -12284 11372
rect -11336 10948 -11272 11372
rect -10324 10948 -10260 11372
rect -9312 10948 -9248 11372
rect -8300 10948 -8236 11372
rect -7288 10948 -7224 11372
rect -6276 10948 -6212 11372
rect -5264 10948 -5200 11372
rect -4252 10948 -4188 11372
rect -3240 10948 -3176 11372
rect -2228 10948 -2164 11372
rect -1216 10948 -1152 11372
rect -204 10948 -140 11372
rect 808 10948 872 11372
rect 1820 10948 1884 11372
rect 2832 10948 2896 11372
rect 3844 10948 3908 11372
rect 4856 10948 4920 11372
rect 5868 10948 5932 11372
rect 6880 10948 6944 11372
rect 7892 10948 7956 11372
rect 8904 10948 8968 11372
rect 9916 10948 9980 11372
rect 10928 10948 10992 11372
rect 11940 10948 12004 11372
rect 12952 10948 13016 11372
rect 13964 10948 14028 11372
rect 14976 10948 15040 11372
rect 15988 10948 16052 11372
rect 17000 10948 17064 11372
rect -16396 10228 -16332 10652
rect -15384 10228 -15320 10652
rect -14372 10228 -14308 10652
rect -13360 10228 -13296 10652
rect -12348 10228 -12284 10652
rect -11336 10228 -11272 10652
rect -10324 10228 -10260 10652
rect -9312 10228 -9248 10652
rect -8300 10228 -8236 10652
rect -7288 10228 -7224 10652
rect -6276 10228 -6212 10652
rect -5264 10228 -5200 10652
rect -4252 10228 -4188 10652
rect -3240 10228 -3176 10652
rect -2228 10228 -2164 10652
rect -1216 10228 -1152 10652
rect -204 10228 -140 10652
rect 808 10228 872 10652
rect 1820 10228 1884 10652
rect 2832 10228 2896 10652
rect 3844 10228 3908 10652
rect 4856 10228 4920 10652
rect 5868 10228 5932 10652
rect 6880 10228 6944 10652
rect 7892 10228 7956 10652
rect 8904 10228 8968 10652
rect 9916 10228 9980 10652
rect 10928 10228 10992 10652
rect 11940 10228 12004 10652
rect 12952 10228 13016 10652
rect 13964 10228 14028 10652
rect 14976 10228 15040 10652
rect 15988 10228 16052 10652
rect 17000 10228 17064 10652
rect -16396 9508 -16332 9932
rect -15384 9508 -15320 9932
rect -14372 9508 -14308 9932
rect -13360 9508 -13296 9932
rect -12348 9508 -12284 9932
rect -11336 9508 -11272 9932
rect -10324 9508 -10260 9932
rect -9312 9508 -9248 9932
rect -8300 9508 -8236 9932
rect -7288 9508 -7224 9932
rect -6276 9508 -6212 9932
rect -5264 9508 -5200 9932
rect -4252 9508 -4188 9932
rect -3240 9508 -3176 9932
rect -2228 9508 -2164 9932
rect -1216 9508 -1152 9932
rect -204 9508 -140 9932
rect 808 9508 872 9932
rect 1820 9508 1884 9932
rect 2832 9508 2896 9932
rect 3844 9508 3908 9932
rect 4856 9508 4920 9932
rect 5868 9508 5932 9932
rect 6880 9508 6944 9932
rect 7892 9508 7956 9932
rect 8904 9508 8968 9932
rect 9916 9508 9980 9932
rect 10928 9508 10992 9932
rect 11940 9508 12004 9932
rect 12952 9508 13016 9932
rect 13964 9508 14028 9932
rect 14976 9508 15040 9932
rect 15988 9508 16052 9932
rect 17000 9508 17064 9932
rect -16396 8788 -16332 9212
rect -15384 8788 -15320 9212
rect -14372 8788 -14308 9212
rect -13360 8788 -13296 9212
rect -12348 8788 -12284 9212
rect -11336 8788 -11272 9212
rect -10324 8788 -10260 9212
rect -9312 8788 -9248 9212
rect -8300 8788 -8236 9212
rect -7288 8788 -7224 9212
rect -6276 8788 -6212 9212
rect -5264 8788 -5200 9212
rect -4252 8788 -4188 9212
rect -3240 8788 -3176 9212
rect -2228 8788 -2164 9212
rect -1216 8788 -1152 9212
rect -204 8788 -140 9212
rect 808 8788 872 9212
rect 1820 8788 1884 9212
rect 2832 8788 2896 9212
rect 3844 8788 3908 9212
rect 4856 8788 4920 9212
rect 5868 8788 5932 9212
rect 6880 8788 6944 9212
rect 7892 8788 7956 9212
rect 8904 8788 8968 9212
rect 9916 8788 9980 9212
rect 10928 8788 10992 9212
rect 11940 8788 12004 9212
rect 12952 8788 13016 9212
rect 13964 8788 14028 9212
rect 14976 8788 15040 9212
rect 15988 8788 16052 9212
rect 17000 8788 17064 9212
rect -16396 8068 -16332 8492
rect -15384 8068 -15320 8492
rect -14372 8068 -14308 8492
rect -13360 8068 -13296 8492
rect -12348 8068 -12284 8492
rect -11336 8068 -11272 8492
rect -10324 8068 -10260 8492
rect -9312 8068 -9248 8492
rect -8300 8068 -8236 8492
rect -7288 8068 -7224 8492
rect -6276 8068 -6212 8492
rect -5264 8068 -5200 8492
rect -4252 8068 -4188 8492
rect -3240 8068 -3176 8492
rect -2228 8068 -2164 8492
rect -1216 8068 -1152 8492
rect -204 8068 -140 8492
rect 808 8068 872 8492
rect 1820 8068 1884 8492
rect 2832 8068 2896 8492
rect 3844 8068 3908 8492
rect 4856 8068 4920 8492
rect 5868 8068 5932 8492
rect 6880 8068 6944 8492
rect 7892 8068 7956 8492
rect 8904 8068 8968 8492
rect 9916 8068 9980 8492
rect 10928 8068 10992 8492
rect 11940 8068 12004 8492
rect 12952 8068 13016 8492
rect 13964 8068 14028 8492
rect 14976 8068 15040 8492
rect 15988 8068 16052 8492
rect 17000 8068 17064 8492
rect -16396 7348 -16332 7772
rect -15384 7348 -15320 7772
rect -14372 7348 -14308 7772
rect -13360 7348 -13296 7772
rect -12348 7348 -12284 7772
rect -11336 7348 -11272 7772
rect -10324 7348 -10260 7772
rect -9312 7348 -9248 7772
rect -8300 7348 -8236 7772
rect -7288 7348 -7224 7772
rect -6276 7348 -6212 7772
rect -5264 7348 -5200 7772
rect -4252 7348 -4188 7772
rect -3240 7348 -3176 7772
rect -2228 7348 -2164 7772
rect -1216 7348 -1152 7772
rect -204 7348 -140 7772
rect 808 7348 872 7772
rect 1820 7348 1884 7772
rect 2832 7348 2896 7772
rect 3844 7348 3908 7772
rect 4856 7348 4920 7772
rect 5868 7348 5932 7772
rect 6880 7348 6944 7772
rect 7892 7348 7956 7772
rect 8904 7348 8968 7772
rect 9916 7348 9980 7772
rect 10928 7348 10992 7772
rect 11940 7348 12004 7772
rect 12952 7348 13016 7772
rect 13964 7348 14028 7772
rect 14976 7348 15040 7772
rect 15988 7348 16052 7772
rect 17000 7348 17064 7772
rect -16396 6628 -16332 7052
rect -15384 6628 -15320 7052
rect -14372 6628 -14308 7052
rect -13360 6628 -13296 7052
rect -12348 6628 -12284 7052
rect -11336 6628 -11272 7052
rect -10324 6628 -10260 7052
rect -9312 6628 -9248 7052
rect -8300 6628 -8236 7052
rect -7288 6628 -7224 7052
rect -6276 6628 -6212 7052
rect -5264 6628 -5200 7052
rect -4252 6628 -4188 7052
rect -3240 6628 -3176 7052
rect -2228 6628 -2164 7052
rect -1216 6628 -1152 7052
rect -204 6628 -140 7052
rect 808 6628 872 7052
rect 1820 6628 1884 7052
rect 2832 6628 2896 7052
rect 3844 6628 3908 7052
rect 4856 6628 4920 7052
rect 5868 6628 5932 7052
rect 6880 6628 6944 7052
rect 7892 6628 7956 7052
rect 8904 6628 8968 7052
rect 9916 6628 9980 7052
rect 10928 6628 10992 7052
rect 11940 6628 12004 7052
rect 12952 6628 13016 7052
rect 13964 6628 14028 7052
rect 14976 6628 15040 7052
rect 15988 6628 16052 7052
rect 17000 6628 17064 7052
rect -16396 5908 -16332 6332
rect -15384 5908 -15320 6332
rect -14372 5908 -14308 6332
rect -13360 5908 -13296 6332
rect -12348 5908 -12284 6332
rect -11336 5908 -11272 6332
rect -10324 5908 -10260 6332
rect -9312 5908 -9248 6332
rect -8300 5908 -8236 6332
rect -7288 5908 -7224 6332
rect -6276 5908 -6212 6332
rect -5264 5908 -5200 6332
rect -4252 5908 -4188 6332
rect -3240 5908 -3176 6332
rect -2228 5908 -2164 6332
rect -1216 5908 -1152 6332
rect -204 5908 -140 6332
rect 808 5908 872 6332
rect 1820 5908 1884 6332
rect 2832 5908 2896 6332
rect 3844 5908 3908 6332
rect 4856 5908 4920 6332
rect 5868 5908 5932 6332
rect 6880 5908 6944 6332
rect 7892 5908 7956 6332
rect 8904 5908 8968 6332
rect 9916 5908 9980 6332
rect 10928 5908 10992 6332
rect 11940 5908 12004 6332
rect 12952 5908 13016 6332
rect 13964 5908 14028 6332
rect 14976 5908 15040 6332
rect 15988 5908 16052 6332
rect 17000 5908 17064 6332
rect -16396 5188 -16332 5612
rect -15384 5188 -15320 5612
rect -14372 5188 -14308 5612
rect -13360 5188 -13296 5612
rect -12348 5188 -12284 5612
rect -11336 5188 -11272 5612
rect -10324 5188 -10260 5612
rect -9312 5188 -9248 5612
rect -8300 5188 -8236 5612
rect -7288 5188 -7224 5612
rect -6276 5188 -6212 5612
rect -5264 5188 -5200 5612
rect -4252 5188 -4188 5612
rect -3240 5188 -3176 5612
rect -2228 5188 -2164 5612
rect -1216 5188 -1152 5612
rect -204 5188 -140 5612
rect 808 5188 872 5612
rect 1820 5188 1884 5612
rect 2832 5188 2896 5612
rect 3844 5188 3908 5612
rect 4856 5188 4920 5612
rect 5868 5188 5932 5612
rect 6880 5188 6944 5612
rect 7892 5188 7956 5612
rect 8904 5188 8968 5612
rect 9916 5188 9980 5612
rect 10928 5188 10992 5612
rect 11940 5188 12004 5612
rect 12952 5188 13016 5612
rect 13964 5188 14028 5612
rect 14976 5188 15040 5612
rect 15988 5188 16052 5612
rect 17000 5188 17064 5612
rect -16396 4468 -16332 4892
rect -15384 4468 -15320 4892
rect -14372 4468 -14308 4892
rect -13360 4468 -13296 4892
rect -12348 4468 -12284 4892
rect -11336 4468 -11272 4892
rect -10324 4468 -10260 4892
rect -9312 4468 -9248 4892
rect -8300 4468 -8236 4892
rect -7288 4468 -7224 4892
rect -6276 4468 -6212 4892
rect -5264 4468 -5200 4892
rect -4252 4468 -4188 4892
rect -3240 4468 -3176 4892
rect -2228 4468 -2164 4892
rect -1216 4468 -1152 4892
rect -204 4468 -140 4892
rect 808 4468 872 4892
rect 1820 4468 1884 4892
rect 2832 4468 2896 4892
rect 3844 4468 3908 4892
rect 4856 4468 4920 4892
rect 5868 4468 5932 4892
rect 6880 4468 6944 4892
rect 7892 4468 7956 4892
rect 8904 4468 8968 4892
rect 9916 4468 9980 4892
rect 10928 4468 10992 4892
rect 11940 4468 12004 4892
rect 12952 4468 13016 4892
rect 13964 4468 14028 4892
rect 14976 4468 15040 4892
rect 15988 4468 16052 4892
rect 17000 4468 17064 4892
rect -16396 3748 -16332 4172
rect -15384 3748 -15320 4172
rect -14372 3748 -14308 4172
rect -13360 3748 -13296 4172
rect -12348 3748 -12284 4172
rect -11336 3748 -11272 4172
rect -10324 3748 -10260 4172
rect -9312 3748 -9248 4172
rect -8300 3748 -8236 4172
rect -7288 3748 -7224 4172
rect -6276 3748 -6212 4172
rect -5264 3748 -5200 4172
rect -4252 3748 -4188 4172
rect -3240 3748 -3176 4172
rect -2228 3748 -2164 4172
rect -1216 3748 -1152 4172
rect -204 3748 -140 4172
rect 808 3748 872 4172
rect 1820 3748 1884 4172
rect 2832 3748 2896 4172
rect 3844 3748 3908 4172
rect 4856 3748 4920 4172
rect 5868 3748 5932 4172
rect 6880 3748 6944 4172
rect 7892 3748 7956 4172
rect 8904 3748 8968 4172
rect 9916 3748 9980 4172
rect 10928 3748 10992 4172
rect 11940 3748 12004 4172
rect 12952 3748 13016 4172
rect 13964 3748 14028 4172
rect 14976 3748 15040 4172
rect 15988 3748 16052 4172
rect 17000 3748 17064 4172
rect -16396 3028 -16332 3452
rect -15384 3028 -15320 3452
rect -14372 3028 -14308 3452
rect -13360 3028 -13296 3452
rect -12348 3028 -12284 3452
rect -11336 3028 -11272 3452
rect -10324 3028 -10260 3452
rect -9312 3028 -9248 3452
rect -8300 3028 -8236 3452
rect -7288 3028 -7224 3452
rect -6276 3028 -6212 3452
rect -5264 3028 -5200 3452
rect -4252 3028 -4188 3452
rect -3240 3028 -3176 3452
rect -2228 3028 -2164 3452
rect -1216 3028 -1152 3452
rect -204 3028 -140 3452
rect 808 3028 872 3452
rect 1820 3028 1884 3452
rect 2832 3028 2896 3452
rect 3844 3028 3908 3452
rect 4856 3028 4920 3452
rect 5868 3028 5932 3452
rect 6880 3028 6944 3452
rect 7892 3028 7956 3452
rect 8904 3028 8968 3452
rect 9916 3028 9980 3452
rect 10928 3028 10992 3452
rect 11940 3028 12004 3452
rect 12952 3028 13016 3452
rect 13964 3028 14028 3452
rect 14976 3028 15040 3452
rect 15988 3028 16052 3452
rect 17000 3028 17064 3452
rect -16396 2308 -16332 2732
rect -15384 2308 -15320 2732
rect -14372 2308 -14308 2732
rect -13360 2308 -13296 2732
rect -12348 2308 -12284 2732
rect -11336 2308 -11272 2732
rect -10324 2308 -10260 2732
rect -9312 2308 -9248 2732
rect -8300 2308 -8236 2732
rect -7288 2308 -7224 2732
rect -6276 2308 -6212 2732
rect -5264 2308 -5200 2732
rect -4252 2308 -4188 2732
rect -3240 2308 -3176 2732
rect -2228 2308 -2164 2732
rect -1216 2308 -1152 2732
rect -204 2308 -140 2732
rect 808 2308 872 2732
rect 1820 2308 1884 2732
rect 2832 2308 2896 2732
rect 3844 2308 3908 2732
rect 4856 2308 4920 2732
rect 5868 2308 5932 2732
rect 6880 2308 6944 2732
rect 7892 2308 7956 2732
rect 8904 2308 8968 2732
rect 9916 2308 9980 2732
rect 10928 2308 10992 2732
rect 11940 2308 12004 2732
rect 12952 2308 13016 2732
rect 13964 2308 14028 2732
rect 14976 2308 15040 2732
rect 15988 2308 16052 2732
rect 17000 2308 17064 2732
rect -16396 1588 -16332 2012
rect -15384 1588 -15320 2012
rect -14372 1588 -14308 2012
rect -13360 1588 -13296 2012
rect -12348 1588 -12284 2012
rect -11336 1588 -11272 2012
rect -10324 1588 -10260 2012
rect -9312 1588 -9248 2012
rect -8300 1588 -8236 2012
rect -7288 1588 -7224 2012
rect -6276 1588 -6212 2012
rect -5264 1588 -5200 2012
rect -4252 1588 -4188 2012
rect -3240 1588 -3176 2012
rect -2228 1588 -2164 2012
rect -1216 1588 -1152 2012
rect -204 1588 -140 2012
rect 808 1588 872 2012
rect 1820 1588 1884 2012
rect 2832 1588 2896 2012
rect 3844 1588 3908 2012
rect 4856 1588 4920 2012
rect 5868 1588 5932 2012
rect 6880 1588 6944 2012
rect 7892 1588 7956 2012
rect 8904 1588 8968 2012
rect 9916 1588 9980 2012
rect 10928 1588 10992 2012
rect 11940 1588 12004 2012
rect 12952 1588 13016 2012
rect 13964 1588 14028 2012
rect 14976 1588 15040 2012
rect 15988 1588 16052 2012
rect 17000 1588 17064 2012
rect -16396 868 -16332 1292
rect -15384 868 -15320 1292
rect -14372 868 -14308 1292
rect -13360 868 -13296 1292
rect -12348 868 -12284 1292
rect -11336 868 -11272 1292
rect -10324 868 -10260 1292
rect -9312 868 -9248 1292
rect -8300 868 -8236 1292
rect -7288 868 -7224 1292
rect -6276 868 -6212 1292
rect -5264 868 -5200 1292
rect -4252 868 -4188 1292
rect -3240 868 -3176 1292
rect -2228 868 -2164 1292
rect -1216 868 -1152 1292
rect -204 868 -140 1292
rect 808 868 872 1292
rect 1820 868 1884 1292
rect 2832 868 2896 1292
rect 3844 868 3908 1292
rect 4856 868 4920 1292
rect 5868 868 5932 1292
rect 6880 868 6944 1292
rect 7892 868 7956 1292
rect 8904 868 8968 1292
rect 9916 868 9980 1292
rect 10928 868 10992 1292
rect 11940 868 12004 1292
rect 12952 868 13016 1292
rect 13964 868 14028 1292
rect 14976 868 15040 1292
rect 15988 868 16052 1292
rect 17000 868 17064 1292
rect -16396 148 -16332 572
rect -15384 148 -15320 572
rect -14372 148 -14308 572
rect -13360 148 -13296 572
rect -12348 148 -12284 572
rect -11336 148 -11272 572
rect -10324 148 -10260 572
rect -9312 148 -9248 572
rect -8300 148 -8236 572
rect -7288 148 -7224 572
rect -6276 148 -6212 572
rect -5264 148 -5200 572
rect -4252 148 -4188 572
rect -3240 148 -3176 572
rect -2228 148 -2164 572
rect -1216 148 -1152 572
rect -204 148 -140 572
rect 808 148 872 572
rect 1820 148 1884 572
rect 2832 148 2896 572
rect 3844 148 3908 572
rect 4856 148 4920 572
rect 5868 148 5932 572
rect 6880 148 6944 572
rect 7892 148 7956 572
rect 8904 148 8968 572
rect 9916 148 9980 572
rect 10928 148 10992 572
rect 11940 148 12004 572
rect 12952 148 13016 572
rect 13964 148 14028 572
rect 14976 148 15040 572
rect 15988 148 16052 572
rect 17000 148 17064 572
rect -16396 -572 -16332 -148
rect -15384 -572 -15320 -148
rect -14372 -572 -14308 -148
rect -13360 -572 -13296 -148
rect -12348 -572 -12284 -148
rect -11336 -572 -11272 -148
rect -10324 -572 -10260 -148
rect -9312 -572 -9248 -148
rect -8300 -572 -8236 -148
rect -7288 -572 -7224 -148
rect -6276 -572 -6212 -148
rect -5264 -572 -5200 -148
rect -4252 -572 -4188 -148
rect -3240 -572 -3176 -148
rect -2228 -572 -2164 -148
rect -1216 -572 -1152 -148
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect 1820 -572 1884 -148
rect 2832 -572 2896 -148
rect 3844 -572 3908 -148
rect 4856 -572 4920 -148
rect 5868 -572 5932 -148
rect 6880 -572 6944 -148
rect 7892 -572 7956 -148
rect 8904 -572 8968 -148
rect 9916 -572 9980 -148
rect 10928 -572 10992 -148
rect 11940 -572 12004 -148
rect 12952 -572 13016 -148
rect 13964 -572 14028 -148
rect 14976 -572 15040 -148
rect 15988 -572 16052 -148
rect 17000 -572 17064 -148
rect -16396 -1292 -16332 -868
rect -15384 -1292 -15320 -868
rect -14372 -1292 -14308 -868
rect -13360 -1292 -13296 -868
rect -12348 -1292 -12284 -868
rect -11336 -1292 -11272 -868
rect -10324 -1292 -10260 -868
rect -9312 -1292 -9248 -868
rect -8300 -1292 -8236 -868
rect -7288 -1292 -7224 -868
rect -6276 -1292 -6212 -868
rect -5264 -1292 -5200 -868
rect -4252 -1292 -4188 -868
rect -3240 -1292 -3176 -868
rect -2228 -1292 -2164 -868
rect -1216 -1292 -1152 -868
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect 1820 -1292 1884 -868
rect 2832 -1292 2896 -868
rect 3844 -1292 3908 -868
rect 4856 -1292 4920 -868
rect 5868 -1292 5932 -868
rect 6880 -1292 6944 -868
rect 7892 -1292 7956 -868
rect 8904 -1292 8968 -868
rect 9916 -1292 9980 -868
rect 10928 -1292 10992 -868
rect 11940 -1292 12004 -868
rect 12952 -1292 13016 -868
rect 13964 -1292 14028 -868
rect 14976 -1292 15040 -868
rect 15988 -1292 16052 -868
rect 17000 -1292 17064 -868
rect -16396 -2012 -16332 -1588
rect -15384 -2012 -15320 -1588
rect -14372 -2012 -14308 -1588
rect -13360 -2012 -13296 -1588
rect -12348 -2012 -12284 -1588
rect -11336 -2012 -11272 -1588
rect -10324 -2012 -10260 -1588
rect -9312 -2012 -9248 -1588
rect -8300 -2012 -8236 -1588
rect -7288 -2012 -7224 -1588
rect -6276 -2012 -6212 -1588
rect -5264 -2012 -5200 -1588
rect -4252 -2012 -4188 -1588
rect -3240 -2012 -3176 -1588
rect -2228 -2012 -2164 -1588
rect -1216 -2012 -1152 -1588
rect -204 -2012 -140 -1588
rect 808 -2012 872 -1588
rect 1820 -2012 1884 -1588
rect 2832 -2012 2896 -1588
rect 3844 -2012 3908 -1588
rect 4856 -2012 4920 -1588
rect 5868 -2012 5932 -1588
rect 6880 -2012 6944 -1588
rect 7892 -2012 7956 -1588
rect 8904 -2012 8968 -1588
rect 9916 -2012 9980 -1588
rect 10928 -2012 10992 -1588
rect 11940 -2012 12004 -1588
rect 12952 -2012 13016 -1588
rect 13964 -2012 14028 -1588
rect 14976 -2012 15040 -1588
rect 15988 -2012 16052 -1588
rect 17000 -2012 17064 -1588
rect -16396 -2732 -16332 -2308
rect -15384 -2732 -15320 -2308
rect -14372 -2732 -14308 -2308
rect -13360 -2732 -13296 -2308
rect -12348 -2732 -12284 -2308
rect -11336 -2732 -11272 -2308
rect -10324 -2732 -10260 -2308
rect -9312 -2732 -9248 -2308
rect -8300 -2732 -8236 -2308
rect -7288 -2732 -7224 -2308
rect -6276 -2732 -6212 -2308
rect -5264 -2732 -5200 -2308
rect -4252 -2732 -4188 -2308
rect -3240 -2732 -3176 -2308
rect -2228 -2732 -2164 -2308
rect -1216 -2732 -1152 -2308
rect -204 -2732 -140 -2308
rect 808 -2732 872 -2308
rect 1820 -2732 1884 -2308
rect 2832 -2732 2896 -2308
rect 3844 -2732 3908 -2308
rect 4856 -2732 4920 -2308
rect 5868 -2732 5932 -2308
rect 6880 -2732 6944 -2308
rect 7892 -2732 7956 -2308
rect 8904 -2732 8968 -2308
rect 9916 -2732 9980 -2308
rect 10928 -2732 10992 -2308
rect 11940 -2732 12004 -2308
rect 12952 -2732 13016 -2308
rect 13964 -2732 14028 -2308
rect 14976 -2732 15040 -2308
rect 15988 -2732 16052 -2308
rect 17000 -2732 17064 -2308
rect -16396 -3452 -16332 -3028
rect -15384 -3452 -15320 -3028
rect -14372 -3452 -14308 -3028
rect -13360 -3452 -13296 -3028
rect -12348 -3452 -12284 -3028
rect -11336 -3452 -11272 -3028
rect -10324 -3452 -10260 -3028
rect -9312 -3452 -9248 -3028
rect -8300 -3452 -8236 -3028
rect -7288 -3452 -7224 -3028
rect -6276 -3452 -6212 -3028
rect -5264 -3452 -5200 -3028
rect -4252 -3452 -4188 -3028
rect -3240 -3452 -3176 -3028
rect -2228 -3452 -2164 -3028
rect -1216 -3452 -1152 -3028
rect -204 -3452 -140 -3028
rect 808 -3452 872 -3028
rect 1820 -3452 1884 -3028
rect 2832 -3452 2896 -3028
rect 3844 -3452 3908 -3028
rect 4856 -3452 4920 -3028
rect 5868 -3452 5932 -3028
rect 6880 -3452 6944 -3028
rect 7892 -3452 7956 -3028
rect 8904 -3452 8968 -3028
rect 9916 -3452 9980 -3028
rect 10928 -3452 10992 -3028
rect 11940 -3452 12004 -3028
rect 12952 -3452 13016 -3028
rect 13964 -3452 14028 -3028
rect 14976 -3452 15040 -3028
rect 15988 -3452 16052 -3028
rect 17000 -3452 17064 -3028
rect -16396 -4172 -16332 -3748
rect -15384 -4172 -15320 -3748
rect -14372 -4172 -14308 -3748
rect -13360 -4172 -13296 -3748
rect -12348 -4172 -12284 -3748
rect -11336 -4172 -11272 -3748
rect -10324 -4172 -10260 -3748
rect -9312 -4172 -9248 -3748
rect -8300 -4172 -8236 -3748
rect -7288 -4172 -7224 -3748
rect -6276 -4172 -6212 -3748
rect -5264 -4172 -5200 -3748
rect -4252 -4172 -4188 -3748
rect -3240 -4172 -3176 -3748
rect -2228 -4172 -2164 -3748
rect -1216 -4172 -1152 -3748
rect -204 -4172 -140 -3748
rect 808 -4172 872 -3748
rect 1820 -4172 1884 -3748
rect 2832 -4172 2896 -3748
rect 3844 -4172 3908 -3748
rect 4856 -4172 4920 -3748
rect 5868 -4172 5932 -3748
rect 6880 -4172 6944 -3748
rect 7892 -4172 7956 -3748
rect 8904 -4172 8968 -3748
rect 9916 -4172 9980 -3748
rect 10928 -4172 10992 -3748
rect 11940 -4172 12004 -3748
rect 12952 -4172 13016 -3748
rect 13964 -4172 14028 -3748
rect 14976 -4172 15040 -3748
rect 15988 -4172 16052 -3748
rect 17000 -4172 17064 -3748
rect -16396 -4892 -16332 -4468
rect -15384 -4892 -15320 -4468
rect -14372 -4892 -14308 -4468
rect -13360 -4892 -13296 -4468
rect -12348 -4892 -12284 -4468
rect -11336 -4892 -11272 -4468
rect -10324 -4892 -10260 -4468
rect -9312 -4892 -9248 -4468
rect -8300 -4892 -8236 -4468
rect -7288 -4892 -7224 -4468
rect -6276 -4892 -6212 -4468
rect -5264 -4892 -5200 -4468
rect -4252 -4892 -4188 -4468
rect -3240 -4892 -3176 -4468
rect -2228 -4892 -2164 -4468
rect -1216 -4892 -1152 -4468
rect -204 -4892 -140 -4468
rect 808 -4892 872 -4468
rect 1820 -4892 1884 -4468
rect 2832 -4892 2896 -4468
rect 3844 -4892 3908 -4468
rect 4856 -4892 4920 -4468
rect 5868 -4892 5932 -4468
rect 6880 -4892 6944 -4468
rect 7892 -4892 7956 -4468
rect 8904 -4892 8968 -4468
rect 9916 -4892 9980 -4468
rect 10928 -4892 10992 -4468
rect 11940 -4892 12004 -4468
rect 12952 -4892 13016 -4468
rect 13964 -4892 14028 -4468
rect 14976 -4892 15040 -4468
rect 15988 -4892 16052 -4468
rect 17000 -4892 17064 -4468
rect -16396 -5612 -16332 -5188
rect -15384 -5612 -15320 -5188
rect -14372 -5612 -14308 -5188
rect -13360 -5612 -13296 -5188
rect -12348 -5612 -12284 -5188
rect -11336 -5612 -11272 -5188
rect -10324 -5612 -10260 -5188
rect -9312 -5612 -9248 -5188
rect -8300 -5612 -8236 -5188
rect -7288 -5612 -7224 -5188
rect -6276 -5612 -6212 -5188
rect -5264 -5612 -5200 -5188
rect -4252 -5612 -4188 -5188
rect -3240 -5612 -3176 -5188
rect -2228 -5612 -2164 -5188
rect -1216 -5612 -1152 -5188
rect -204 -5612 -140 -5188
rect 808 -5612 872 -5188
rect 1820 -5612 1884 -5188
rect 2832 -5612 2896 -5188
rect 3844 -5612 3908 -5188
rect 4856 -5612 4920 -5188
rect 5868 -5612 5932 -5188
rect 6880 -5612 6944 -5188
rect 7892 -5612 7956 -5188
rect 8904 -5612 8968 -5188
rect 9916 -5612 9980 -5188
rect 10928 -5612 10992 -5188
rect 11940 -5612 12004 -5188
rect 12952 -5612 13016 -5188
rect 13964 -5612 14028 -5188
rect 14976 -5612 15040 -5188
rect 15988 -5612 16052 -5188
rect 17000 -5612 17064 -5188
rect -16396 -6332 -16332 -5908
rect -15384 -6332 -15320 -5908
rect -14372 -6332 -14308 -5908
rect -13360 -6332 -13296 -5908
rect -12348 -6332 -12284 -5908
rect -11336 -6332 -11272 -5908
rect -10324 -6332 -10260 -5908
rect -9312 -6332 -9248 -5908
rect -8300 -6332 -8236 -5908
rect -7288 -6332 -7224 -5908
rect -6276 -6332 -6212 -5908
rect -5264 -6332 -5200 -5908
rect -4252 -6332 -4188 -5908
rect -3240 -6332 -3176 -5908
rect -2228 -6332 -2164 -5908
rect -1216 -6332 -1152 -5908
rect -204 -6332 -140 -5908
rect 808 -6332 872 -5908
rect 1820 -6332 1884 -5908
rect 2832 -6332 2896 -5908
rect 3844 -6332 3908 -5908
rect 4856 -6332 4920 -5908
rect 5868 -6332 5932 -5908
rect 6880 -6332 6944 -5908
rect 7892 -6332 7956 -5908
rect 8904 -6332 8968 -5908
rect 9916 -6332 9980 -5908
rect 10928 -6332 10992 -5908
rect 11940 -6332 12004 -5908
rect 12952 -6332 13016 -5908
rect 13964 -6332 14028 -5908
rect 14976 -6332 15040 -5908
rect 15988 -6332 16052 -5908
rect 17000 -6332 17064 -5908
rect -16396 -7052 -16332 -6628
rect -15384 -7052 -15320 -6628
rect -14372 -7052 -14308 -6628
rect -13360 -7052 -13296 -6628
rect -12348 -7052 -12284 -6628
rect -11336 -7052 -11272 -6628
rect -10324 -7052 -10260 -6628
rect -9312 -7052 -9248 -6628
rect -8300 -7052 -8236 -6628
rect -7288 -7052 -7224 -6628
rect -6276 -7052 -6212 -6628
rect -5264 -7052 -5200 -6628
rect -4252 -7052 -4188 -6628
rect -3240 -7052 -3176 -6628
rect -2228 -7052 -2164 -6628
rect -1216 -7052 -1152 -6628
rect -204 -7052 -140 -6628
rect 808 -7052 872 -6628
rect 1820 -7052 1884 -6628
rect 2832 -7052 2896 -6628
rect 3844 -7052 3908 -6628
rect 4856 -7052 4920 -6628
rect 5868 -7052 5932 -6628
rect 6880 -7052 6944 -6628
rect 7892 -7052 7956 -6628
rect 8904 -7052 8968 -6628
rect 9916 -7052 9980 -6628
rect 10928 -7052 10992 -6628
rect 11940 -7052 12004 -6628
rect 12952 -7052 13016 -6628
rect 13964 -7052 14028 -6628
rect 14976 -7052 15040 -6628
rect 15988 -7052 16052 -6628
rect 17000 -7052 17064 -6628
rect -16396 -7772 -16332 -7348
rect -15384 -7772 -15320 -7348
rect -14372 -7772 -14308 -7348
rect -13360 -7772 -13296 -7348
rect -12348 -7772 -12284 -7348
rect -11336 -7772 -11272 -7348
rect -10324 -7772 -10260 -7348
rect -9312 -7772 -9248 -7348
rect -8300 -7772 -8236 -7348
rect -7288 -7772 -7224 -7348
rect -6276 -7772 -6212 -7348
rect -5264 -7772 -5200 -7348
rect -4252 -7772 -4188 -7348
rect -3240 -7772 -3176 -7348
rect -2228 -7772 -2164 -7348
rect -1216 -7772 -1152 -7348
rect -204 -7772 -140 -7348
rect 808 -7772 872 -7348
rect 1820 -7772 1884 -7348
rect 2832 -7772 2896 -7348
rect 3844 -7772 3908 -7348
rect 4856 -7772 4920 -7348
rect 5868 -7772 5932 -7348
rect 6880 -7772 6944 -7348
rect 7892 -7772 7956 -7348
rect 8904 -7772 8968 -7348
rect 9916 -7772 9980 -7348
rect 10928 -7772 10992 -7348
rect 11940 -7772 12004 -7348
rect 12952 -7772 13016 -7348
rect 13964 -7772 14028 -7348
rect 14976 -7772 15040 -7348
rect 15988 -7772 16052 -7348
rect 17000 -7772 17064 -7348
rect -16396 -8492 -16332 -8068
rect -15384 -8492 -15320 -8068
rect -14372 -8492 -14308 -8068
rect -13360 -8492 -13296 -8068
rect -12348 -8492 -12284 -8068
rect -11336 -8492 -11272 -8068
rect -10324 -8492 -10260 -8068
rect -9312 -8492 -9248 -8068
rect -8300 -8492 -8236 -8068
rect -7288 -8492 -7224 -8068
rect -6276 -8492 -6212 -8068
rect -5264 -8492 -5200 -8068
rect -4252 -8492 -4188 -8068
rect -3240 -8492 -3176 -8068
rect -2228 -8492 -2164 -8068
rect -1216 -8492 -1152 -8068
rect -204 -8492 -140 -8068
rect 808 -8492 872 -8068
rect 1820 -8492 1884 -8068
rect 2832 -8492 2896 -8068
rect 3844 -8492 3908 -8068
rect 4856 -8492 4920 -8068
rect 5868 -8492 5932 -8068
rect 6880 -8492 6944 -8068
rect 7892 -8492 7956 -8068
rect 8904 -8492 8968 -8068
rect 9916 -8492 9980 -8068
rect 10928 -8492 10992 -8068
rect 11940 -8492 12004 -8068
rect 12952 -8492 13016 -8068
rect 13964 -8492 14028 -8068
rect 14976 -8492 15040 -8068
rect 15988 -8492 16052 -8068
rect 17000 -8492 17064 -8068
rect -16396 -9212 -16332 -8788
rect -15384 -9212 -15320 -8788
rect -14372 -9212 -14308 -8788
rect -13360 -9212 -13296 -8788
rect -12348 -9212 -12284 -8788
rect -11336 -9212 -11272 -8788
rect -10324 -9212 -10260 -8788
rect -9312 -9212 -9248 -8788
rect -8300 -9212 -8236 -8788
rect -7288 -9212 -7224 -8788
rect -6276 -9212 -6212 -8788
rect -5264 -9212 -5200 -8788
rect -4252 -9212 -4188 -8788
rect -3240 -9212 -3176 -8788
rect -2228 -9212 -2164 -8788
rect -1216 -9212 -1152 -8788
rect -204 -9212 -140 -8788
rect 808 -9212 872 -8788
rect 1820 -9212 1884 -8788
rect 2832 -9212 2896 -8788
rect 3844 -9212 3908 -8788
rect 4856 -9212 4920 -8788
rect 5868 -9212 5932 -8788
rect 6880 -9212 6944 -8788
rect 7892 -9212 7956 -8788
rect 8904 -9212 8968 -8788
rect 9916 -9212 9980 -8788
rect 10928 -9212 10992 -8788
rect 11940 -9212 12004 -8788
rect 12952 -9212 13016 -8788
rect 13964 -9212 14028 -8788
rect 14976 -9212 15040 -8788
rect 15988 -9212 16052 -8788
rect 17000 -9212 17064 -8788
rect -16396 -9932 -16332 -9508
rect -15384 -9932 -15320 -9508
rect -14372 -9932 -14308 -9508
rect -13360 -9932 -13296 -9508
rect -12348 -9932 -12284 -9508
rect -11336 -9932 -11272 -9508
rect -10324 -9932 -10260 -9508
rect -9312 -9932 -9248 -9508
rect -8300 -9932 -8236 -9508
rect -7288 -9932 -7224 -9508
rect -6276 -9932 -6212 -9508
rect -5264 -9932 -5200 -9508
rect -4252 -9932 -4188 -9508
rect -3240 -9932 -3176 -9508
rect -2228 -9932 -2164 -9508
rect -1216 -9932 -1152 -9508
rect -204 -9932 -140 -9508
rect 808 -9932 872 -9508
rect 1820 -9932 1884 -9508
rect 2832 -9932 2896 -9508
rect 3844 -9932 3908 -9508
rect 4856 -9932 4920 -9508
rect 5868 -9932 5932 -9508
rect 6880 -9932 6944 -9508
rect 7892 -9932 7956 -9508
rect 8904 -9932 8968 -9508
rect 9916 -9932 9980 -9508
rect 10928 -9932 10992 -9508
rect 11940 -9932 12004 -9508
rect 12952 -9932 13016 -9508
rect 13964 -9932 14028 -9508
rect 14976 -9932 15040 -9508
rect 15988 -9932 16052 -9508
rect 17000 -9932 17064 -9508
rect -16396 -10652 -16332 -10228
rect -15384 -10652 -15320 -10228
rect -14372 -10652 -14308 -10228
rect -13360 -10652 -13296 -10228
rect -12348 -10652 -12284 -10228
rect -11336 -10652 -11272 -10228
rect -10324 -10652 -10260 -10228
rect -9312 -10652 -9248 -10228
rect -8300 -10652 -8236 -10228
rect -7288 -10652 -7224 -10228
rect -6276 -10652 -6212 -10228
rect -5264 -10652 -5200 -10228
rect -4252 -10652 -4188 -10228
rect -3240 -10652 -3176 -10228
rect -2228 -10652 -2164 -10228
rect -1216 -10652 -1152 -10228
rect -204 -10652 -140 -10228
rect 808 -10652 872 -10228
rect 1820 -10652 1884 -10228
rect 2832 -10652 2896 -10228
rect 3844 -10652 3908 -10228
rect 4856 -10652 4920 -10228
rect 5868 -10652 5932 -10228
rect 6880 -10652 6944 -10228
rect 7892 -10652 7956 -10228
rect 8904 -10652 8968 -10228
rect 9916 -10652 9980 -10228
rect 10928 -10652 10992 -10228
rect 11940 -10652 12004 -10228
rect 12952 -10652 13016 -10228
rect 13964 -10652 14028 -10228
rect 14976 -10652 15040 -10228
rect 15988 -10652 16052 -10228
rect 17000 -10652 17064 -10228
rect -16396 -11372 -16332 -10948
rect -15384 -11372 -15320 -10948
rect -14372 -11372 -14308 -10948
rect -13360 -11372 -13296 -10948
rect -12348 -11372 -12284 -10948
rect -11336 -11372 -11272 -10948
rect -10324 -11372 -10260 -10948
rect -9312 -11372 -9248 -10948
rect -8300 -11372 -8236 -10948
rect -7288 -11372 -7224 -10948
rect -6276 -11372 -6212 -10948
rect -5264 -11372 -5200 -10948
rect -4252 -11372 -4188 -10948
rect -3240 -11372 -3176 -10948
rect -2228 -11372 -2164 -10948
rect -1216 -11372 -1152 -10948
rect -204 -11372 -140 -10948
rect 808 -11372 872 -10948
rect 1820 -11372 1884 -10948
rect 2832 -11372 2896 -10948
rect 3844 -11372 3908 -10948
rect 4856 -11372 4920 -10948
rect 5868 -11372 5932 -10948
rect 6880 -11372 6944 -10948
rect 7892 -11372 7956 -10948
rect 8904 -11372 8968 -10948
rect 9916 -11372 9980 -10948
rect 10928 -11372 10992 -10948
rect 11940 -11372 12004 -10948
rect 12952 -11372 13016 -10948
rect 13964 -11372 14028 -10948
rect 14976 -11372 15040 -10948
rect 15988 -11372 16052 -10948
rect 17000 -11372 17064 -10948
<< mimcap >>
rect -17044 11320 -16644 11360
rect -17044 11000 -17004 11320
rect -16684 11000 -16644 11320
rect -17044 10960 -16644 11000
rect -16032 11320 -15632 11360
rect -16032 11000 -15992 11320
rect -15672 11000 -15632 11320
rect -16032 10960 -15632 11000
rect -15020 11320 -14620 11360
rect -15020 11000 -14980 11320
rect -14660 11000 -14620 11320
rect -15020 10960 -14620 11000
rect -14008 11320 -13608 11360
rect -14008 11000 -13968 11320
rect -13648 11000 -13608 11320
rect -14008 10960 -13608 11000
rect -12996 11320 -12596 11360
rect -12996 11000 -12956 11320
rect -12636 11000 -12596 11320
rect -12996 10960 -12596 11000
rect -11984 11320 -11584 11360
rect -11984 11000 -11944 11320
rect -11624 11000 -11584 11320
rect -11984 10960 -11584 11000
rect -10972 11320 -10572 11360
rect -10972 11000 -10932 11320
rect -10612 11000 -10572 11320
rect -10972 10960 -10572 11000
rect -9960 11320 -9560 11360
rect -9960 11000 -9920 11320
rect -9600 11000 -9560 11320
rect -9960 10960 -9560 11000
rect -8948 11320 -8548 11360
rect -8948 11000 -8908 11320
rect -8588 11000 -8548 11320
rect -8948 10960 -8548 11000
rect -7936 11320 -7536 11360
rect -7936 11000 -7896 11320
rect -7576 11000 -7536 11320
rect -7936 10960 -7536 11000
rect -6924 11320 -6524 11360
rect -6924 11000 -6884 11320
rect -6564 11000 -6524 11320
rect -6924 10960 -6524 11000
rect -5912 11320 -5512 11360
rect -5912 11000 -5872 11320
rect -5552 11000 -5512 11320
rect -5912 10960 -5512 11000
rect -4900 11320 -4500 11360
rect -4900 11000 -4860 11320
rect -4540 11000 -4500 11320
rect -4900 10960 -4500 11000
rect -3888 11320 -3488 11360
rect -3888 11000 -3848 11320
rect -3528 11000 -3488 11320
rect -3888 10960 -3488 11000
rect -2876 11320 -2476 11360
rect -2876 11000 -2836 11320
rect -2516 11000 -2476 11320
rect -2876 10960 -2476 11000
rect -1864 11320 -1464 11360
rect -1864 11000 -1824 11320
rect -1504 11000 -1464 11320
rect -1864 10960 -1464 11000
rect -852 11320 -452 11360
rect -852 11000 -812 11320
rect -492 11000 -452 11320
rect -852 10960 -452 11000
rect 160 11320 560 11360
rect 160 11000 200 11320
rect 520 11000 560 11320
rect 160 10960 560 11000
rect 1172 11320 1572 11360
rect 1172 11000 1212 11320
rect 1532 11000 1572 11320
rect 1172 10960 1572 11000
rect 2184 11320 2584 11360
rect 2184 11000 2224 11320
rect 2544 11000 2584 11320
rect 2184 10960 2584 11000
rect 3196 11320 3596 11360
rect 3196 11000 3236 11320
rect 3556 11000 3596 11320
rect 3196 10960 3596 11000
rect 4208 11320 4608 11360
rect 4208 11000 4248 11320
rect 4568 11000 4608 11320
rect 4208 10960 4608 11000
rect 5220 11320 5620 11360
rect 5220 11000 5260 11320
rect 5580 11000 5620 11320
rect 5220 10960 5620 11000
rect 6232 11320 6632 11360
rect 6232 11000 6272 11320
rect 6592 11000 6632 11320
rect 6232 10960 6632 11000
rect 7244 11320 7644 11360
rect 7244 11000 7284 11320
rect 7604 11000 7644 11320
rect 7244 10960 7644 11000
rect 8256 11320 8656 11360
rect 8256 11000 8296 11320
rect 8616 11000 8656 11320
rect 8256 10960 8656 11000
rect 9268 11320 9668 11360
rect 9268 11000 9308 11320
rect 9628 11000 9668 11320
rect 9268 10960 9668 11000
rect 10280 11320 10680 11360
rect 10280 11000 10320 11320
rect 10640 11000 10680 11320
rect 10280 10960 10680 11000
rect 11292 11320 11692 11360
rect 11292 11000 11332 11320
rect 11652 11000 11692 11320
rect 11292 10960 11692 11000
rect 12304 11320 12704 11360
rect 12304 11000 12344 11320
rect 12664 11000 12704 11320
rect 12304 10960 12704 11000
rect 13316 11320 13716 11360
rect 13316 11000 13356 11320
rect 13676 11000 13716 11320
rect 13316 10960 13716 11000
rect 14328 11320 14728 11360
rect 14328 11000 14368 11320
rect 14688 11000 14728 11320
rect 14328 10960 14728 11000
rect 15340 11320 15740 11360
rect 15340 11000 15380 11320
rect 15700 11000 15740 11320
rect 15340 10960 15740 11000
rect 16352 11320 16752 11360
rect 16352 11000 16392 11320
rect 16712 11000 16752 11320
rect 16352 10960 16752 11000
rect -17044 10600 -16644 10640
rect -17044 10280 -17004 10600
rect -16684 10280 -16644 10600
rect -17044 10240 -16644 10280
rect -16032 10600 -15632 10640
rect -16032 10280 -15992 10600
rect -15672 10280 -15632 10600
rect -16032 10240 -15632 10280
rect -15020 10600 -14620 10640
rect -15020 10280 -14980 10600
rect -14660 10280 -14620 10600
rect -15020 10240 -14620 10280
rect -14008 10600 -13608 10640
rect -14008 10280 -13968 10600
rect -13648 10280 -13608 10600
rect -14008 10240 -13608 10280
rect -12996 10600 -12596 10640
rect -12996 10280 -12956 10600
rect -12636 10280 -12596 10600
rect -12996 10240 -12596 10280
rect -11984 10600 -11584 10640
rect -11984 10280 -11944 10600
rect -11624 10280 -11584 10600
rect -11984 10240 -11584 10280
rect -10972 10600 -10572 10640
rect -10972 10280 -10932 10600
rect -10612 10280 -10572 10600
rect -10972 10240 -10572 10280
rect -9960 10600 -9560 10640
rect -9960 10280 -9920 10600
rect -9600 10280 -9560 10600
rect -9960 10240 -9560 10280
rect -8948 10600 -8548 10640
rect -8948 10280 -8908 10600
rect -8588 10280 -8548 10600
rect -8948 10240 -8548 10280
rect -7936 10600 -7536 10640
rect -7936 10280 -7896 10600
rect -7576 10280 -7536 10600
rect -7936 10240 -7536 10280
rect -6924 10600 -6524 10640
rect -6924 10280 -6884 10600
rect -6564 10280 -6524 10600
rect -6924 10240 -6524 10280
rect -5912 10600 -5512 10640
rect -5912 10280 -5872 10600
rect -5552 10280 -5512 10600
rect -5912 10240 -5512 10280
rect -4900 10600 -4500 10640
rect -4900 10280 -4860 10600
rect -4540 10280 -4500 10600
rect -4900 10240 -4500 10280
rect -3888 10600 -3488 10640
rect -3888 10280 -3848 10600
rect -3528 10280 -3488 10600
rect -3888 10240 -3488 10280
rect -2876 10600 -2476 10640
rect -2876 10280 -2836 10600
rect -2516 10280 -2476 10600
rect -2876 10240 -2476 10280
rect -1864 10600 -1464 10640
rect -1864 10280 -1824 10600
rect -1504 10280 -1464 10600
rect -1864 10240 -1464 10280
rect -852 10600 -452 10640
rect -852 10280 -812 10600
rect -492 10280 -452 10600
rect -852 10240 -452 10280
rect 160 10600 560 10640
rect 160 10280 200 10600
rect 520 10280 560 10600
rect 160 10240 560 10280
rect 1172 10600 1572 10640
rect 1172 10280 1212 10600
rect 1532 10280 1572 10600
rect 1172 10240 1572 10280
rect 2184 10600 2584 10640
rect 2184 10280 2224 10600
rect 2544 10280 2584 10600
rect 2184 10240 2584 10280
rect 3196 10600 3596 10640
rect 3196 10280 3236 10600
rect 3556 10280 3596 10600
rect 3196 10240 3596 10280
rect 4208 10600 4608 10640
rect 4208 10280 4248 10600
rect 4568 10280 4608 10600
rect 4208 10240 4608 10280
rect 5220 10600 5620 10640
rect 5220 10280 5260 10600
rect 5580 10280 5620 10600
rect 5220 10240 5620 10280
rect 6232 10600 6632 10640
rect 6232 10280 6272 10600
rect 6592 10280 6632 10600
rect 6232 10240 6632 10280
rect 7244 10600 7644 10640
rect 7244 10280 7284 10600
rect 7604 10280 7644 10600
rect 7244 10240 7644 10280
rect 8256 10600 8656 10640
rect 8256 10280 8296 10600
rect 8616 10280 8656 10600
rect 8256 10240 8656 10280
rect 9268 10600 9668 10640
rect 9268 10280 9308 10600
rect 9628 10280 9668 10600
rect 9268 10240 9668 10280
rect 10280 10600 10680 10640
rect 10280 10280 10320 10600
rect 10640 10280 10680 10600
rect 10280 10240 10680 10280
rect 11292 10600 11692 10640
rect 11292 10280 11332 10600
rect 11652 10280 11692 10600
rect 11292 10240 11692 10280
rect 12304 10600 12704 10640
rect 12304 10280 12344 10600
rect 12664 10280 12704 10600
rect 12304 10240 12704 10280
rect 13316 10600 13716 10640
rect 13316 10280 13356 10600
rect 13676 10280 13716 10600
rect 13316 10240 13716 10280
rect 14328 10600 14728 10640
rect 14328 10280 14368 10600
rect 14688 10280 14728 10600
rect 14328 10240 14728 10280
rect 15340 10600 15740 10640
rect 15340 10280 15380 10600
rect 15700 10280 15740 10600
rect 15340 10240 15740 10280
rect 16352 10600 16752 10640
rect 16352 10280 16392 10600
rect 16712 10280 16752 10600
rect 16352 10240 16752 10280
rect -17044 9880 -16644 9920
rect -17044 9560 -17004 9880
rect -16684 9560 -16644 9880
rect -17044 9520 -16644 9560
rect -16032 9880 -15632 9920
rect -16032 9560 -15992 9880
rect -15672 9560 -15632 9880
rect -16032 9520 -15632 9560
rect -15020 9880 -14620 9920
rect -15020 9560 -14980 9880
rect -14660 9560 -14620 9880
rect -15020 9520 -14620 9560
rect -14008 9880 -13608 9920
rect -14008 9560 -13968 9880
rect -13648 9560 -13608 9880
rect -14008 9520 -13608 9560
rect -12996 9880 -12596 9920
rect -12996 9560 -12956 9880
rect -12636 9560 -12596 9880
rect -12996 9520 -12596 9560
rect -11984 9880 -11584 9920
rect -11984 9560 -11944 9880
rect -11624 9560 -11584 9880
rect -11984 9520 -11584 9560
rect -10972 9880 -10572 9920
rect -10972 9560 -10932 9880
rect -10612 9560 -10572 9880
rect -10972 9520 -10572 9560
rect -9960 9880 -9560 9920
rect -9960 9560 -9920 9880
rect -9600 9560 -9560 9880
rect -9960 9520 -9560 9560
rect -8948 9880 -8548 9920
rect -8948 9560 -8908 9880
rect -8588 9560 -8548 9880
rect -8948 9520 -8548 9560
rect -7936 9880 -7536 9920
rect -7936 9560 -7896 9880
rect -7576 9560 -7536 9880
rect -7936 9520 -7536 9560
rect -6924 9880 -6524 9920
rect -6924 9560 -6884 9880
rect -6564 9560 -6524 9880
rect -6924 9520 -6524 9560
rect -5912 9880 -5512 9920
rect -5912 9560 -5872 9880
rect -5552 9560 -5512 9880
rect -5912 9520 -5512 9560
rect -4900 9880 -4500 9920
rect -4900 9560 -4860 9880
rect -4540 9560 -4500 9880
rect -4900 9520 -4500 9560
rect -3888 9880 -3488 9920
rect -3888 9560 -3848 9880
rect -3528 9560 -3488 9880
rect -3888 9520 -3488 9560
rect -2876 9880 -2476 9920
rect -2876 9560 -2836 9880
rect -2516 9560 -2476 9880
rect -2876 9520 -2476 9560
rect -1864 9880 -1464 9920
rect -1864 9560 -1824 9880
rect -1504 9560 -1464 9880
rect -1864 9520 -1464 9560
rect -852 9880 -452 9920
rect -852 9560 -812 9880
rect -492 9560 -452 9880
rect -852 9520 -452 9560
rect 160 9880 560 9920
rect 160 9560 200 9880
rect 520 9560 560 9880
rect 160 9520 560 9560
rect 1172 9880 1572 9920
rect 1172 9560 1212 9880
rect 1532 9560 1572 9880
rect 1172 9520 1572 9560
rect 2184 9880 2584 9920
rect 2184 9560 2224 9880
rect 2544 9560 2584 9880
rect 2184 9520 2584 9560
rect 3196 9880 3596 9920
rect 3196 9560 3236 9880
rect 3556 9560 3596 9880
rect 3196 9520 3596 9560
rect 4208 9880 4608 9920
rect 4208 9560 4248 9880
rect 4568 9560 4608 9880
rect 4208 9520 4608 9560
rect 5220 9880 5620 9920
rect 5220 9560 5260 9880
rect 5580 9560 5620 9880
rect 5220 9520 5620 9560
rect 6232 9880 6632 9920
rect 6232 9560 6272 9880
rect 6592 9560 6632 9880
rect 6232 9520 6632 9560
rect 7244 9880 7644 9920
rect 7244 9560 7284 9880
rect 7604 9560 7644 9880
rect 7244 9520 7644 9560
rect 8256 9880 8656 9920
rect 8256 9560 8296 9880
rect 8616 9560 8656 9880
rect 8256 9520 8656 9560
rect 9268 9880 9668 9920
rect 9268 9560 9308 9880
rect 9628 9560 9668 9880
rect 9268 9520 9668 9560
rect 10280 9880 10680 9920
rect 10280 9560 10320 9880
rect 10640 9560 10680 9880
rect 10280 9520 10680 9560
rect 11292 9880 11692 9920
rect 11292 9560 11332 9880
rect 11652 9560 11692 9880
rect 11292 9520 11692 9560
rect 12304 9880 12704 9920
rect 12304 9560 12344 9880
rect 12664 9560 12704 9880
rect 12304 9520 12704 9560
rect 13316 9880 13716 9920
rect 13316 9560 13356 9880
rect 13676 9560 13716 9880
rect 13316 9520 13716 9560
rect 14328 9880 14728 9920
rect 14328 9560 14368 9880
rect 14688 9560 14728 9880
rect 14328 9520 14728 9560
rect 15340 9880 15740 9920
rect 15340 9560 15380 9880
rect 15700 9560 15740 9880
rect 15340 9520 15740 9560
rect 16352 9880 16752 9920
rect 16352 9560 16392 9880
rect 16712 9560 16752 9880
rect 16352 9520 16752 9560
rect -17044 9160 -16644 9200
rect -17044 8840 -17004 9160
rect -16684 8840 -16644 9160
rect -17044 8800 -16644 8840
rect -16032 9160 -15632 9200
rect -16032 8840 -15992 9160
rect -15672 8840 -15632 9160
rect -16032 8800 -15632 8840
rect -15020 9160 -14620 9200
rect -15020 8840 -14980 9160
rect -14660 8840 -14620 9160
rect -15020 8800 -14620 8840
rect -14008 9160 -13608 9200
rect -14008 8840 -13968 9160
rect -13648 8840 -13608 9160
rect -14008 8800 -13608 8840
rect -12996 9160 -12596 9200
rect -12996 8840 -12956 9160
rect -12636 8840 -12596 9160
rect -12996 8800 -12596 8840
rect -11984 9160 -11584 9200
rect -11984 8840 -11944 9160
rect -11624 8840 -11584 9160
rect -11984 8800 -11584 8840
rect -10972 9160 -10572 9200
rect -10972 8840 -10932 9160
rect -10612 8840 -10572 9160
rect -10972 8800 -10572 8840
rect -9960 9160 -9560 9200
rect -9960 8840 -9920 9160
rect -9600 8840 -9560 9160
rect -9960 8800 -9560 8840
rect -8948 9160 -8548 9200
rect -8948 8840 -8908 9160
rect -8588 8840 -8548 9160
rect -8948 8800 -8548 8840
rect -7936 9160 -7536 9200
rect -7936 8840 -7896 9160
rect -7576 8840 -7536 9160
rect -7936 8800 -7536 8840
rect -6924 9160 -6524 9200
rect -6924 8840 -6884 9160
rect -6564 8840 -6524 9160
rect -6924 8800 -6524 8840
rect -5912 9160 -5512 9200
rect -5912 8840 -5872 9160
rect -5552 8840 -5512 9160
rect -5912 8800 -5512 8840
rect -4900 9160 -4500 9200
rect -4900 8840 -4860 9160
rect -4540 8840 -4500 9160
rect -4900 8800 -4500 8840
rect -3888 9160 -3488 9200
rect -3888 8840 -3848 9160
rect -3528 8840 -3488 9160
rect -3888 8800 -3488 8840
rect -2876 9160 -2476 9200
rect -2876 8840 -2836 9160
rect -2516 8840 -2476 9160
rect -2876 8800 -2476 8840
rect -1864 9160 -1464 9200
rect -1864 8840 -1824 9160
rect -1504 8840 -1464 9160
rect -1864 8800 -1464 8840
rect -852 9160 -452 9200
rect -852 8840 -812 9160
rect -492 8840 -452 9160
rect -852 8800 -452 8840
rect 160 9160 560 9200
rect 160 8840 200 9160
rect 520 8840 560 9160
rect 160 8800 560 8840
rect 1172 9160 1572 9200
rect 1172 8840 1212 9160
rect 1532 8840 1572 9160
rect 1172 8800 1572 8840
rect 2184 9160 2584 9200
rect 2184 8840 2224 9160
rect 2544 8840 2584 9160
rect 2184 8800 2584 8840
rect 3196 9160 3596 9200
rect 3196 8840 3236 9160
rect 3556 8840 3596 9160
rect 3196 8800 3596 8840
rect 4208 9160 4608 9200
rect 4208 8840 4248 9160
rect 4568 8840 4608 9160
rect 4208 8800 4608 8840
rect 5220 9160 5620 9200
rect 5220 8840 5260 9160
rect 5580 8840 5620 9160
rect 5220 8800 5620 8840
rect 6232 9160 6632 9200
rect 6232 8840 6272 9160
rect 6592 8840 6632 9160
rect 6232 8800 6632 8840
rect 7244 9160 7644 9200
rect 7244 8840 7284 9160
rect 7604 8840 7644 9160
rect 7244 8800 7644 8840
rect 8256 9160 8656 9200
rect 8256 8840 8296 9160
rect 8616 8840 8656 9160
rect 8256 8800 8656 8840
rect 9268 9160 9668 9200
rect 9268 8840 9308 9160
rect 9628 8840 9668 9160
rect 9268 8800 9668 8840
rect 10280 9160 10680 9200
rect 10280 8840 10320 9160
rect 10640 8840 10680 9160
rect 10280 8800 10680 8840
rect 11292 9160 11692 9200
rect 11292 8840 11332 9160
rect 11652 8840 11692 9160
rect 11292 8800 11692 8840
rect 12304 9160 12704 9200
rect 12304 8840 12344 9160
rect 12664 8840 12704 9160
rect 12304 8800 12704 8840
rect 13316 9160 13716 9200
rect 13316 8840 13356 9160
rect 13676 8840 13716 9160
rect 13316 8800 13716 8840
rect 14328 9160 14728 9200
rect 14328 8840 14368 9160
rect 14688 8840 14728 9160
rect 14328 8800 14728 8840
rect 15340 9160 15740 9200
rect 15340 8840 15380 9160
rect 15700 8840 15740 9160
rect 15340 8800 15740 8840
rect 16352 9160 16752 9200
rect 16352 8840 16392 9160
rect 16712 8840 16752 9160
rect 16352 8800 16752 8840
rect -17044 8440 -16644 8480
rect -17044 8120 -17004 8440
rect -16684 8120 -16644 8440
rect -17044 8080 -16644 8120
rect -16032 8440 -15632 8480
rect -16032 8120 -15992 8440
rect -15672 8120 -15632 8440
rect -16032 8080 -15632 8120
rect -15020 8440 -14620 8480
rect -15020 8120 -14980 8440
rect -14660 8120 -14620 8440
rect -15020 8080 -14620 8120
rect -14008 8440 -13608 8480
rect -14008 8120 -13968 8440
rect -13648 8120 -13608 8440
rect -14008 8080 -13608 8120
rect -12996 8440 -12596 8480
rect -12996 8120 -12956 8440
rect -12636 8120 -12596 8440
rect -12996 8080 -12596 8120
rect -11984 8440 -11584 8480
rect -11984 8120 -11944 8440
rect -11624 8120 -11584 8440
rect -11984 8080 -11584 8120
rect -10972 8440 -10572 8480
rect -10972 8120 -10932 8440
rect -10612 8120 -10572 8440
rect -10972 8080 -10572 8120
rect -9960 8440 -9560 8480
rect -9960 8120 -9920 8440
rect -9600 8120 -9560 8440
rect -9960 8080 -9560 8120
rect -8948 8440 -8548 8480
rect -8948 8120 -8908 8440
rect -8588 8120 -8548 8440
rect -8948 8080 -8548 8120
rect -7936 8440 -7536 8480
rect -7936 8120 -7896 8440
rect -7576 8120 -7536 8440
rect -7936 8080 -7536 8120
rect -6924 8440 -6524 8480
rect -6924 8120 -6884 8440
rect -6564 8120 -6524 8440
rect -6924 8080 -6524 8120
rect -5912 8440 -5512 8480
rect -5912 8120 -5872 8440
rect -5552 8120 -5512 8440
rect -5912 8080 -5512 8120
rect -4900 8440 -4500 8480
rect -4900 8120 -4860 8440
rect -4540 8120 -4500 8440
rect -4900 8080 -4500 8120
rect -3888 8440 -3488 8480
rect -3888 8120 -3848 8440
rect -3528 8120 -3488 8440
rect -3888 8080 -3488 8120
rect -2876 8440 -2476 8480
rect -2876 8120 -2836 8440
rect -2516 8120 -2476 8440
rect -2876 8080 -2476 8120
rect -1864 8440 -1464 8480
rect -1864 8120 -1824 8440
rect -1504 8120 -1464 8440
rect -1864 8080 -1464 8120
rect -852 8440 -452 8480
rect -852 8120 -812 8440
rect -492 8120 -452 8440
rect -852 8080 -452 8120
rect 160 8440 560 8480
rect 160 8120 200 8440
rect 520 8120 560 8440
rect 160 8080 560 8120
rect 1172 8440 1572 8480
rect 1172 8120 1212 8440
rect 1532 8120 1572 8440
rect 1172 8080 1572 8120
rect 2184 8440 2584 8480
rect 2184 8120 2224 8440
rect 2544 8120 2584 8440
rect 2184 8080 2584 8120
rect 3196 8440 3596 8480
rect 3196 8120 3236 8440
rect 3556 8120 3596 8440
rect 3196 8080 3596 8120
rect 4208 8440 4608 8480
rect 4208 8120 4248 8440
rect 4568 8120 4608 8440
rect 4208 8080 4608 8120
rect 5220 8440 5620 8480
rect 5220 8120 5260 8440
rect 5580 8120 5620 8440
rect 5220 8080 5620 8120
rect 6232 8440 6632 8480
rect 6232 8120 6272 8440
rect 6592 8120 6632 8440
rect 6232 8080 6632 8120
rect 7244 8440 7644 8480
rect 7244 8120 7284 8440
rect 7604 8120 7644 8440
rect 7244 8080 7644 8120
rect 8256 8440 8656 8480
rect 8256 8120 8296 8440
rect 8616 8120 8656 8440
rect 8256 8080 8656 8120
rect 9268 8440 9668 8480
rect 9268 8120 9308 8440
rect 9628 8120 9668 8440
rect 9268 8080 9668 8120
rect 10280 8440 10680 8480
rect 10280 8120 10320 8440
rect 10640 8120 10680 8440
rect 10280 8080 10680 8120
rect 11292 8440 11692 8480
rect 11292 8120 11332 8440
rect 11652 8120 11692 8440
rect 11292 8080 11692 8120
rect 12304 8440 12704 8480
rect 12304 8120 12344 8440
rect 12664 8120 12704 8440
rect 12304 8080 12704 8120
rect 13316 8440 13716 8480
rect 13316 8120 13356 8440
rect 13676 8120 13716 8440
rect 13316 8080 13716 8120
rect 14328 8440 14728 8480
rect 14328 8120 14368 8440
rect 14688 8120 14728 8440
rect 14328 8080 14728 8120
rect 15340 8440 15740 8480
rect 15340 8120 15380 8440
rect 15700 8120 15740 8440
rect 15340 8080 15740 8120
rect 16352 8440 16752 8480
rect 16352 8120 16392 8440
rect 16712 8120 16752 8440
rect 16352 8080 16752 8120
rect -17044 7720 -16644 7760
rect -17044 7400 -17004 7720
rect -16684 7400 -16644 7720
rect -17044 7360 -16644 7400
rect -16032 7720 -15632 7760
rect -16032 7400 -15992 7720
rect -15672 7400 -15632 7720
rect -16032 7360 -15632 7400
rect -15020 7720 -14620 7760
rect -15020 7400 -14980 7720
rect -14660 7400 -14620 7720
rect -15020 7360 -14620 7400
rect -14008 7720 -13608 7760
rect -14008 7400 -13968 7720
rect -13648 7400 -13608 7720
rect -14008 7360 -13608 7400
rect -12996 7720 -12596 7760
rect -12996 7400 -12956 7720
rect -12636 7400 -12596 7720
rect -12996 7360 -12596 7400
rect -11984 7720 -11584 7760
rect -11984 7400 -11944 7720
rect -11624 7400 -11584 7720
rect -11984 7360 -11584 7400
rect -10972 7720 -10572 7760
rect -10972 7400 -10932 7720
rect -10612 7400 -10572 7720
rect -10972 7360 -10572 7400
rect -9960 7720 -9560 7760
rect -9960 7400 -9920 7720
rect -9600 7400 -9560 7720
rect -9960 7360 -9560 7400
rect -8948 7720 -8548 7760
rect -8948 7400 -8908 7720
rect -8588 7400 -8548 7720
rect -8948 7360 -8548 7400
rect -7936 7720 -7536 7760
rect -7936 7400 -7896 7720
rect -7576 7400 -7536 7720
rect -7936 7360 -7536 7400
rect -6924 7720 -6524 7760
rect -6924 7400 -6884 7720
rect -6564 7400 -6524 7720
rect -6924 7360 -6524 7400
rect -5912 7720 -5512 7760
rect -5912 7400 -5872 7720
rect -5552 7400 -5512 7720
rect -5912 7360 -5512 7400
rect -4900 7720 -4500 7760
rect -4900 7400 -4860 7720
rect -4540 7400 -4500 7720
rect -4900 7360 -4500 7400
rect -3888 7720 -3488 7760
rect -3888 7400 -3848 7720
rect -3528 7400 -3488 7720
rect -3888 7360 -3488 7400
rect -2876 7720 -2476 7760
rect -2876 7400 -2836 7720
rect -2516 7400 -2476 7720
rect -2876 7360 -2476 7400
rect -1864 7720 -1464 7760
rect -1864 7400 -1824 7720
rect -1504 7400 -1464 7720
rect -1864 7360 -1464 7400
rect -852 7720 -452 7760
rect -852 7400 -812 7720
rect -492 7400 -452 7720
rect -852 7360 -452 7400
rect 160 7720 560 7760
rect 160 7400 200 7720
rect 520 7400 560 7720
rect 160 7360 560 7400
rect 1172 7720 1572 7760
rect 1172 7400 1212 7720
rect 1532 7400 1572 7720
rect 1172 7360 1572 7400
rect 2184 7720 2584 7760
rect 2184 7400 2224 7720
rect 2544 7400 2584 7720
rect 2184 7360 2584 7400
rect 3196 7720 3596 7760
rect 3196 7400 3236 7720
rect 3556 7400 3596 7720
rect 3196 7360 3596 7400
rect 4208 7720 4608 7760
rect 4208 7400 4248 7720
rect 4568 7400 4608 7720
rect 4208 7360 4608 7400
rect 5220 7720 5620 7760
rect 5220 7400 5260 7720
rect 5580 7400 5620 7720
rect 5220 7360 5620 7400
rect 6232 7720 6632 7760
rect 6232 7400 6272 7720
rect 6592 7400 6632 7720
rect 6232 7360 6632 7400
rect 7244 7720 7644 7760
rect 7244 7400 7284 7720
rect 7604 7400 7644 7720
rect 7244 7360 7644 7400
rect 8256 7720 8656 7760
rect 8256 7400 8296 7720
rect 8616 7400 8656 7720
rect 8256 7360 8656 7400
rect 9268 7720 9668 7760
rect 9268 7400 9308 7720
rect 9628 7400 9668 7720
rect 9268 7360 9668 7400
rect 10280 7720 10680 7760
rect 10280 7400 10320 7720
rect 10640 7400 10680 7720
rect 10280 7360 10680 7400
rect 11292 7720 11692 7760
rect 11292 7400 11332 7720
rect 11652 7400 11692 7720
rect 11292 7360 11692 7400
rect 12304 7720 12704 7760
rect 12304 7400 12344 7720
rect 12664 7400 12704 7720
rect 12304 7360 12704 7400
rect 13316 7720 13716 7760
rect 13316 7400 13356 7720
rect 13676 7400 13716 7720
rect 13316 7360 13716 7400
rect 14328 7720 14728 7760
rect 14328 7400 14368 7720
rect 14688 7400 14728 7720
rect 14328 7360 14728 7400
rect 15340 7720 15740 7760
rect 15340 7400 15380 7720
rect 15700 7400 15740 7720
rect 15340 7360 15740 7400
rect 16352 7720 16752 7760
rect 16352 7400 16392 7720
rect 16712 7400 16752 7720
rect 16352 7360 16752 7400
rect -17044 7000 -16644 7040
rect -17044 6680 -17004 7000
rect -16684 6680 -16644 7000
rect -17044 6640 -16644 6680
rect -16032 7000 -15632 7040
rect -16032 6680 -15992 7000
rect -15672 6680 -15632 7000
rect -16032 6640 -15632 6680
rect -15020 7000 -14620 7040
rect -15020 6680 -14980 7000
rect -14660 6680 -14620 7000
rect -15020 6640 -14620 6680
rect -14008 7000 -13608 7040
rect -14008 6680 -13968 7000
rect -13648 6680 -13608 7000
rect -14008 6640 -13608 6680
rect -12996 7000 -12596 7040
rect -12996 6680 -12956 7000
rect -12636 6680 -12596 7000
rect -12996 6640 -12596 6680
rect -11984 7000 -11584 7040
rect -11984 6680 -11944 7000
rect -11624 6680 -11584 7000
rect -11984 6640 -11584 6680
rect -10972 7000 -10572 7040
rect -10972 6680 -10932 7000
rect -10612 6680 -10572 7000
rect -10972 6640 -10572 6680
rect -9960 7000 -9560 7040
rect -9960 6680 -9920 7000
rect -9600 6680 -9560 7000
rect -9960 6640 -9560 6680
rect -8948 7000 -8548 7040
rect -8948 6680 -8908 7000
rect -8588 6680 -8548 7000
rect -8948 6640 -8548 6680
rect -7936 7000 -7536 7040
rect -7936 6680 -7896 7000
rect -7576 6680 -7536 7000
rect -7936 6640 -7536 6680
rect -6924 7000 -6524 7040
rect -6924 6680 -6884 7000
rect -6564 6680 -6524 7000
rect -6924 6640 -6524 6680
rect -5912 7000 -5512 7040
rect -5912 6680 -5872 7000
rect -5552 6680 -5512 7000
rect -5912 6640 -5512 6680
rect -4900 7000 -4500 7040
rect -4900 6680 -4860 7000
rect -4540 6680 -4500 7000
rect -4900 6640 -4500 6680
rect -3888 7000 -3488 7040
rect -3888 6680 -3848 7000
rect -3528 6680 -3488 7000
rect -3888 6640 -3488 6680
rect -2876 7000 -2476 7040
rect -2876 6680 -2836 7000
rect -2516 6680 -2476 7000
rect -2876 6640 -2476 6680
rect -1864 7000 -1464 7040
rect -1864 6680 -1824 7000
rect -1504 6680 -1464 7000
rect -1864 6640 -1464 6680
rect -852 7000 -452 7040
rect -852 6680 -812 7000
rect -492 6680 -452 7000
rect -852 6640 -452 6680
rect 160 7000 560 7040
rect 160 6680 200 7000
rect 520 6680 560 7000
rect 160 6640 560 6680
rect 1172 7000 1572 7040
rect 1172 6680 1212 7000
rect 1532 6680 1572 7000
rect 1172 6640 1572 6680
rect 2184 7000 2584 7040
rect 2184 6680 2224 7000
rect 2544 6680 2584 7000
rect 2184 6640 2584 6680
rect 3196 7000 3596 7040
rect 3196 6680 3236 7000
rect 3556 6680 3596 7000
rect 3196 6640 3596 6680
rect 4208 7000 4608 7040
rect 4208 6680 4248 7000
rect 4568 6680 4608 7000
rect 4208 6640 4608 6680
rect 5220 7000 5620 7040
rect 5220 6680 5260 7000
rect 5580 6680 5620 7000
rect 5220 6640 5620 6680
rect 6232 7000 6632 7040
rect 6232 6680 6272 7000
rect 6592 6680 6632 7000
rect 6232 6640 6632 6680
rect 7244 7000 7644 7040
rect 7244 6680 7284 7000
rect 7604 6680 7644 7000
rect 7244 6640 7644 6680
rect 8256 7000 8656 7040
rect 8256 6680 8296 7000
rect 8616 6680 8656 7000
rect 8256 6640 8656 6680
rect 9268 7000 9668 7040
rect 9268 6680 9308 7000
rect 9628 6680 9668 7000
rect 9268 6640 9668 6680
rect 10280 7000 10680 7040
rect 10280 6680 10320 7000
rect 10640 6680 10680 7000
rect 10280 6640 10680 6680
rect 11292 7000 11692 7040
rect 11292 6680 11332 7000
rect 11652 6680 11692 7000
rect 11292 6640 11692 6680
rect 12304 7000 12704 7040
rect 12304 6680 12344 7000
rect 12664 6680 12704 7000
rect 12304 6640 12704 6680
rect 13316 7000 13716 7040
rect 13316 6680 13356 7000
rect 13676 6680 13716 7000
rect 13316 6640 13716 6680
rect 14328 7000 14728 7040
rect 14328 6680 14368 7000
rect 14688 6680 14728 7000
rect 14328 6640 14728 6680
rect 15340 7000 15740 7040
rect 15340 6680 15380 7000
rect 15700 6680 15740 7000
rect 15340 6640 15740 6680
rect 16352 7000 16752 7040
rect 16352 6680 16392 7000
rect 16712 6680 16752 7000
rect 16352 6640 16752 6680
rect -17044 6280 -16644 6320
rect -17044 5960 -17004 6280
rect -16684 5960 -16644 6280
rect -17044 5920 -16644 5960
rect -16032 6280 -15632 6320
rect -16032 5960 -15992 6280
rect -15672 5960 -15632 6280
rect -16032 5920 -15632 5960
rect -15020 6280 -14620 6320
rect -15020 5960 -14980 6280
rect -14660 5960 -14620 6280
rect -15020 5920 -14620 5960
rect -14008 6280 -13608 6320
rect -14008 5960 -13968 6280
rect -13648 5960 -13608 6280
rect -14008 5920 -13608 5960
rect -12996 6280 -12596 6320
rect -12996 5960 -12956 6280
rect -12636 5960 -12596 6280
rect -12996 5920 -12596 5960
rect -11984 6280 -11584 6320
rect -11984 5960 -11944 6280
rect -11624 5960 -11584 6280
rect -11984 5920 -11584 5960
rect -10972 6280 -10572 6320
rect -10972 5960 -10932 6280
rect -10612 5960 -10572 6280
rect -10972 5920 -10572 5960
rect -9960 6280 -9560 6320
rect -9960 5960 -9920 6280
rect -9600 5960 -9560 6280
rect -9960 5920 -9560 5960
rect -8948 6280 -8548 6320
rect -8948 5960 -8908 6280
rect -8588 5960 -8548 6280
rect -8948 5920 -8548 5960
rect -7936 6280 -7536 6320
rect -7936 5960 -7896 6280
rect -7576 5960 -7536 6280
rect -7936 5920 -7536 5960
rect -6924 6280 -6524 6320
rect -6924 5960 -6884 6280
rect -6564 5960 -6524 6280
rect -6924 5920 -6524 5960
rect -5912 6280 -5512 6320
rect -5912 5960 -5872 6280
rect -5552 5960 -5512 6280
rect -5912 5920 -5512 5960
rect -4900 6280 -4500 6320
rect -4900 5960 -4860 6280
rect -4540 5960 -4500 6280
rect -4900 5920 -4500 5960
rect -3888 6280 -3488 6320
rect -3888 5960 -3848 6280
rect -3528 5960 -3488 6280
rect -3888 5920 -3488 5960
rect -2876 6280 -2476 6320
rect -2876 5960 -2836 6280
rect -2516 5960 -2476 6280
rect -2876 5920 -2476 5960
rect -1864 6280 -1464 6320
rect -1864 5960 -1824 6280
rect -1504 5960 -1464 6280
rect -1864 5920 -1464 5960
rect -852 6280 -452 6320
rect -852 5960 -812 6280
rect -492 5960 -452 6280
rect -852 5920 -452 5960
rect 160 6280 560 6320
rect 160 5960 200 6280
rect 520 5960 560 6280
rect 160 5920 560 5960
rect 1172 6280 1572 6320
rect 1172 5960 1212 6280
rect 1532 5960 1572 6280
rect 1172 5920 1572 5960
rect 2184 6280 2584 6320
rect 2184 5960 2224 6280
rect 2544 5960 2584 6280
rect 2184 5920 2584 5960
rect 3196 6280 3596 6320
rect 3196 5960 3236 6280
rect 3556 5960 3596 6280
rect 3196 5920 3596 5960
rect 4208 6280 4608 6320
rect 4208 5960 4248 6280
rect 4568 5960 4608 6280
rect 4208 5920 4608 5960
rect 5220 6280 5620 6320
rect 5220 5960 5260 6280
rect 5580 5960 5620 6280
rect 5220 5920 5620 5960
rect 6232 6280 6632 6320
rect 6232 5960 6272 6280
rect 6592 5960 6632 6280
rect 6232 5920 6632 5960
rect 7244 6280 7644 6320
rect 7244 5960 7284 6280
rect 7604 5960 7644 6280
rect 7244 5920 7644 5960
rect 8256 6280 8656 6320
rect 8256 5960 8296 6280
rect 8616 5960 8656 6280
rect 8256 5920 8656 5960
rect 9268 6280 9668 6320
rect 9268 5960 9308 6280
rect 9628 5960 9668 6280
rect 9268 5920 9668 5960
rect 10280 6280 10680 6320
rect 10280 5960 10320 6280
rect 10640 5960 10680 6280
rect 10280 5920 10680 5960
rect 11292 6280 11692 6320
rect 11292 5960 11332 6280
rect 11652 5960 11692 6280
rect 11292 5920 11692 5960
rect 12304 6280 12704 6320
rect 12304 5960 12344 6280
rect 12664 5960 12704 6280
rect 12304 5920 12704 5960
rect 13316 6280 13716 6320
rect 13316 5960 13356 6280
rect 13676 5960 13716 6280
rect 13316 5920 13716 5960
rect 14328 6280 14728 6320
rect 14328 5960 14368 6280
rect 14688 5960 14728 6280
rect 14328 5920 14728 5960
rect 15340 6280 15740 6320
rect 15340 5960 15380 6280
rect 15700 5960 15740 6280
rect 15340 5920 15740 5960
rect 16352 6280 16752 6320
rect 16352 5960 16392 6280
rect 16712 5960 16752 6280
rect 16352 5920 16752 5960
rect -17044 5560 -16644 5600
rect -17044 5240 -17004 5560
rect -16684 5240 -16644 5560
rect -17044 5200 -16644 5240
rect -16032 5560 -15632 5600
rect -16032 5240 -15992 5560
rect -15672 5240 -15632 5560
rect -16032 5200 -15632 5240
rect -15020 5560 -14620 5600
rect -15020 5240 -14980 5560
rect -14660 5240 -14620 5560
rect -15020 5200 -14620 5240
rect -14008 5560 -13608 5600
rect -14008 5240 -13968 5560
rect -13648 5240 -13608 5560
rect -14008 5200 -13608 5240
rect -12996 5560 -12596 5600
rect -12996 5240 -12956 5560
rect -12636 5240 -12596 5560
rect -12996 5200 -12596 5240
rect -11984 5560 -11584 5600
rect -11984 5240 -11944 5560
rect -11624 5240 -11584 5560
rect -11984 5200 -11584 5240
rect -10972 5560 -10572 5600
rect -10972 5240 -10932 5560
rect -10612 5240 -10572 5560
rect -10972 5200 -10572 5240
rect -9960 5560 -9560 5600
rect -9960 5240 -9920 5560
rect -9600 5240 -9560 5560
rect -9960 5200 -9560 5240
rect -8948 5560 -8548 5600
rect -8948 5240 -8908 5560
rect -8588 5240 -8548 5560
rect -8948 5200 -8548 5240
rect -7936 5560 -7536 5600
rect -7936 5240 -7896 5560
rect -7576 5240 -7536 5560
rect -7936 5200 -7536 5240
rect -6924 5560 -6524 5600
rect -6924 5240 -6884 5560
rect -6564 5240 -6524 5560
rect -6924 5200 -6524 5240
rect -5912 5560 -5512 5600
rect -5912 5240 -5872 5560
rect -5552 5240 -5512 5560
rect -5912 5200 -5512 5240
rect -4900 5560 -4500 5600
rect -4900 5240 -4860 5560
rect -4540 5240 -4500 5560
rect -4900 5200 -4500 5240
rect -3888 5560 -3488 5600
rect -3888 5240 -3848 5560
rect -3528 5240 -3488 5560
rect -3888 5200 -3488 5240
rect -2876 5560 -2476 5600
rect -2876 5240 -2836 5560
rect -2516 5240 -2476 5560
rect -2876 5200 -2476 5240
rect -1864 5560 -1464 5600
rect -1864 5240 -1824 5560
rect -1504 5240 -1464 5560
rect -1864 5200 -1464 5240
rect -852 5560 -452 5600
rect -852 5240 -812 5560
rect -492 5240 -452 5560
rect -852 5200 -452 5240
rect 160 5560 560 5600
rect 160 5240 200 5560
rect 520 5240 560 5560
rect 160 5200 560 5240
rect 1172 5560 1572 5600
rect 1172 5240 1212 5560
rect 1532 5240 1572 5560
rect 1172 5200 1572 5240
rect 2184 5560 2584 5600
rect 2184 5240 2224 5560
rect 2544 5240 2584 5560
rect 2184 5200 2584 5240
rect 3196 5560 3596 5600
rect 3196 5240 3236 5560
rect 3556 5240 3596 5560
rect 3196 5200 3596 5240
rect 4208 5560 4608 5600
rect 4208 5240 4248 5560
rect 4568 5240 4608 5560
rect 4208 5200 4608 5240
rect 5220 5560 5620 5600
rect 5220 5240 5260 5560
rect 5580 5240 5620 5560
rect 5220 5200 5620 5240
rect 6232 5560 6632 5600
rect 6232 5240 6272 5560
rect 6592 5240 6632 5560
rect 6232 5200 6632 5240
rect 7244 5560 7644 5600
rect 7244 5240 7284 5560
rect 7604 5240 7644 5560
rect 7244 5200 7644 5240
rect 8256 5560 8656 5600
rect 8256 5240 8296 5560
rect 8616 5240 8656 5560
rect 8256 5200 8656 5240
rect 9268 5560 9668 5600
rect 9268 5240 9308 5560
rect 9628 5240 9668 5560
rect 9268 5200 9668 5240
rect 10280 5560 10680 5600
rect 10280 5240 10320 5560
rect 10640 5240 10680 5560
rect 10280 5200 10680 5240
rect 11292 5560 11692 5600
rect 11292 5240 11332 5560
rect 11652 5240 11692 5560
rect 11292 5200 11692 5240
rect 12304 5560 12704 5600
rect 12304 5240 12344 5560
rect 12664 5240 12704 5560
rect 12304 5200 12704 5240
rect 13316 5560 13716 5600
rect 13316 5240 13356 5560
rect 13676 5240 13716 5560
rect 13316 5200 13716 5240
rect 14328 5560 14728 5600
rect 14328 5240 14368 5560
rect 14688 5240 14728 5560
rect 14328 5200 14728 5240
rect 15340 5560 15740 5600
rect 15340 5240 15380 5560
rect 15700 5240 15740 5560
rect 15340 5200 15740 5240
rect 16352 5560 16752 5600
rect 16352 5240 16392 5560
rect 16712 5240 16752 5560
rect 16352 5200 16752 5240
rect -17044 4840 -16644 4880
rect -17044 4520 -17004 4840
rect -16684 4520 -16644 4840
rect -17044 4480 -16644 4520
rect -16032 4840 -15632 4880
rect -16032 4520 -15992 4840
rect -15672 4520 -15632 4840
rect -16032 4480 -15632 4520
rect -15020 4840 -14620 4880
rect -15020 4520 -14980 4840
rect -14660 4520 -14620 4840
rect -15020 4480 -14620 4520
rect -14008 4840 -13608 4880
rect -14008 4520 -13968 4840
rect -13648 4520 -13608 4840
rect -14008 4480 -13608 4520
rect -12996 4840 -12596 4880
rect -12996 4520 -12956 4840
rect -12636 4520 -12596 4840
rect -12996 4480 -12596 4520
rect -11984 4840 -11584 4880
rect -11984 4520 -11944 4840
rect -11624 4520 -11584 4840
rect -11984 4480 -11584 4520
rect -10972 4840 -10572 4880
rect -10972 4520 -10932 4840
rect -10612 4520 -10572 4840
rect -10972 4480 -10572 4520
rect -9960 4840 -9560 4880
rect -9960 4520 -9920 4840
rect -9600 4520 -9560 4840
rect -9960 4480 -9560 4520
rect -8948 4840 -8548 4880
rect -8948 4520 -8908 4840
rect -8588 4520 -8548 4840
rect -8948 4480 -8548 4520
rect -7936 4840 -7536 4880
rect -7936 4520 -7896 4840
rect -7576 4520 -7536 4840
rect -7936 4480 -7536 4520
rect -6924 4840 -6524 4880
rect -6924 4520 -6884 4840
rect -6564 4520 -6524 4840
rect -6924 4480 -6524 4520
rect -5912 4840 -5512 4880
rect -5912 4520 -5872 4840
rect -5552 4520 -5512 4840
rect -5912 4480 -5512 4520
rect -4900 4840 -4500 4880
rect -4900 4520 -4860 4840
rect -4540 4520 -4500 4840
rect -4900 4480 -4500 4520
rect -3888 4840 -3488 4880
rect -3888 4520 -3848 4840
rect -3528 4520 -3488 4840
rect -3888 4480 -3488 4520
rect -2876 4840 -2476 4880
rect -2876 4520 -2836 4840
rect -2516 4520 -2476 4840
rect -2876 4480 -2476 4520
rect -1864 4840 -1464 4880
rect -1864 4520 -1824 4840
rect -1504 4520 -1464 4840
rect -1864 4480 -1464 4520
rect -852 4840 -452 4880
rect -852 4520 -812 4840
rect -492 4520 -452 4840
rect -852 4480 -452 4520
rect 160 4840 560 4880
rect 160 4520 200 4840
rect 520 4520 560 4840
rect 160 4480 560 4520
rect 1172 4840 1572 4880
rect 1172 4520 1212 4840
rect 1532 4520 1572 4840
rect 1172 4480 1572 4520
rect 2184 4840 2584 4880
rect 2184 4520 2224 4840
rect 2544 4520 2584 4840
rect 2184 4480 2584 4520
rect 3196 4840 3596 4880
rect 3196 4520 3236 4840
rect 3556 4520 3596 4840
rect 3196 4480 3596 4520
rect 4208 4840 4608 4880
rect 4208 4520 4248 4840
rect 4568 4520 4608 4840
rect 4208 4480 4608 4520
rect 5220 4840 5620 4880
rect 5220 4520 5260 4840
rect 5580 4520 5620 4840
rect 5220 4480 5620 4520
rect 6232 4840 6632 4880
rect 6232 4520 6272 4840
rect 6592 4520 6632 4840
rect 6232 4480 6632 4520
rect 7244 4840 7644 4880
rect 7244 4520 7284 4840
rect 7604 4520 7644 4840
rect 7244 4480 7644 4520
rect 8256 4840 8656 4880
rect 8256 4520 8296 4840
rect 8616 4520 8656 4840
rect 8256 4480 8656 4520
rect 9268 4840 9668 4880
rect 9268 4520 9308 4840
rect 9628 4520 9668 4840
rect 9268 4480 9668 4520
rect 10280 4840 10680 4880
rect 10280 4520 10320 4840
rect 10640 4520 10680 4840
rect 10280 4480 10680 4520
rect 11292 4840 11692 4880
rect 11292 4520 11332 4840
rect 11652 4520 11692 4840
rect 11292 4480 11692 4520
rect 12304 4840 12704 4880
rect 12304 4520 12344 4840
rect 12664 4520 12704 4840
rect 12304 4480 12704 4520
rect 13316 4840 13716 4880
rect 13316 4520 13356 4840
rect 13676 4520 13716 4840
rect 13316 4480 13716 4520
rect 14328 4840 14728 4880
rect 14328 4520 14368 4840
rect 14688 4520 14728 4840
rect 14328 4480 14728 4520
rect 15340 4840 15740 4880
rect 15340 4520 15380 4840
rect 15700 4520 15740 4840
rect 15340 4480 15740 4520
rect 16352 4840 16752 4880
rect 16352 4520 16392 4840
rect 16712 4520 16752 4840
rect 16352 4480 16752 4520
rect -17044 4120 -16644 4160
rect -17044 3800 -17004 4120
rect -16684 3800 -16644 4120
rect -17044 3760 -16644 3800
rect -16032 4120 -15632 4160
rect -16032 3800 -15992 4120
rect -15672 3800 -15632 4120
rect -16032 3760 -15632 3800
rect -15020 4120 -14620 4160
rect -15020 3800 -14980 4120
rect -14660 3800 -14620 4120
rect -15020 3760 -14620 3800
rect -14008 4120 -13608 4160
rect -14008 3800 -13968 4120
rect -13648 3800 -13608 4120
rect -14008 3760 -13608 3800
rect -12996 4120 -12596 4160
rect -12996 3800 -12956 4120
rect -12636 3800 -12596 4120
rect -12996 3760 -12596 3800
rect -11984 4120 -11584 4160
rect -11984 3800 -11944 4120
rect -11624 3800 -11584 4120
rect -11984 3760 -11584 3800
rect -10972 4120 -10572 4160
rect -10972 3800 -10932 4120
rect -10612 3800 -10572 4120
rect -10972 3760 -10572 3800
rect -9960 4120 -9560 4160
rect -9960 3800 -9920 4120
rect -9600 3800 -9560 4120
rect -9960 3760 -9560 3800
rect -8948 4120 -8548 4160
rect -8948 3800 -8908 4120
rect -8588 3800 -8548 4120
rect -8948 3760 -8548 3800
rect -7936 4120 -7536 4160
rect -7936 3800 -7896 4120
rect -7576 3800 -7536 4120
rect -7936 3760 -7536 3800
rect -6924 4120 -6524 4160
rect -6924 3800 -6884 4120
rect -6564 3800 -6524 4120
rect -6924 3760 -6524 3800
rect -5912 4120 -5512 4160
rect -5912 3800 -5872 4120
rect -5552 3800 -5512 4120
rect -5912 3760 -5512 3800
rect -4900 4120 -4500 4160
rect -4900 3800 -4860 4120
rect -4540 3800 -4500 4120
rect -4900 3760 -4500 3800
rect -3888 4120 -3488 4160
rect -3888 3800 -3848 4120
rect -3528 3800 -3488 4120
rect -3888 3760 -3488 3800
rect -2876 4120 -2476 4160
rect -2876 3800 -2836 4120
rect -2516 3800 -2476 4120
rect -2876 3760 -2476 3800
rect -1864 4120 -1464 4160
rect -1864 3800 -1824 4120
rect -1504 3800 -1464 4120
rect -1864 3760 -1464 3800
rect -852 4120 -452 4160
rect -852 3800 -812 4120
rect -492 3800 -452 4120
rect -852 3760 -452 3800
rect 160 4120 560 4160
rect 160 3800 200 4120
rect 520 3800 560 4120
rect 160 3760 560 3800
rect 1172 4120 1572 4160
rect 1172 3800 1212 4120
rect 1532 3800 1572 4120
rect 1172 3760 1572 3800
rect 2184 4120 2584 4160
rect 2184 3800 2224 4120
rect 2544 3800 2584 4120
rect 2184 3760 2584 3800
rect 3196 4120 3596 4160
rect 3196 3800 3236 4120
rect 3556 3800 3596 4120
rect 3196 3760 3596 3800
rect 4208 4120 4608 4160
rect 4208 3800 4248 4120
rect 4568 3800 4608 4120
rect 4208 3760 4608 3800
rect 5220 4120 5620 4160
rect 5220 3800 5260 4120
rect 5580 3800 5620 4120
rect 5220 3760 5620 3800
rect 6232 4120 6632 4160
rect 6232 3800 6272 4120
rect 6592 3800 6632 4120
rect 6232 3760 6632 3800
rect 7244 4120 7644 4160
rect 7244 3800 7284 4120
rect 7604 3800 7644 4120
rect 7244 3760 7644 3800
rect 8256 4120 8656 4160
rect 8256 3800 8296 4120
rect 8616 3800 8656 4120
rect 8256 3760 8656 3800
rect 9268 4120 9668 4160
rect 9268 3800 9308 4120
rect 9628 3800 9668 4120
rect 9268 3760 9668 3800
rect 10280 4120 10680 4160
rect 10280 3800 10320 4120
rect 10640 3800 10680 4120
rect 10280 3760 10680 3800
rect 11292 4120 11692 4160
rect 11292 3800 11332 4120
rect 11652 3800 11692 4120
rect 11292 3760 11692 3800
rect 12304 4120 12704 4160
rect 12304 3800 12344 4120
rect 12664 3800 12704 4120
rect 12304 3760 12704 3800
rect 13316 4120 13716 4160
rect 13316 3800 13356 4120
rect 13676 3800 13716 4120
rect 13316 3760 13716 3800
rect 14328 4120 14728 4160
rect 14328 3800 14368 4120
rect 14688 3800 14728 4120
rect 14328 3760 14728 3800
rect 15340 4120 15740 4160
rect 15340 3800 15380 4120
rect 15700 3800 15740 4120
rect 15340 3760 15740 3800
rect 16352 4120 16752 4160
rect 16352 3800 16392 4120
rect 16712 3800 16752 4120
rect 16352 3760 16752 3800
rect -17044 3400 -16644 3440
rect -17044 3080 -17004 3400
rect -16684 3080 -16644 3400
rect -17044 3040 -16644 3080
rect -16032 3400 -15632 3440
rect -16032 3080 -15992 3400
rect -15672 3080 -15632 3400
rect -16032 3040 -15632 3080
rect -15020 3400 -14620 3440
rect -15020 3080 -14980 3400
rect -14660 3080 -14620 3400
rect -15020 3040 -14620 3080
rect -14008 3400 -13608 3440
rect -14008 3080 -13968 3400
rect -13648 3080 -13608 3400
rect -14008 3040 -13608 3080
rect -12996 3400 -12596 3440
rect -12996 3080 -12956 3400
rect -12636 3080 -12596 3400
rect -12996 3040 -12596 3080
rect -11984 3400 -11584 3440
rect -11984 3080 -11944 3400
rect -11624 3080 -11584 3400
rect -11984 3040 -11584 3080
rect -10972 3400 -10572 3440
rect -10972 3080 -10932 3400
rect -10612 3080 -10572 3400
rect -10972 3040 -10572 3080
rect -9960 3400 -9560 3440
rect -9960 3080 -9920 3400
rect -9600 3080 -9560 3400
rect -9960 3040 -9560 3080
rect -8948 3400 -8548 3440
rect -8948 3080 -8908 3400
rect -8588 3080 -8548 3400
rect -8948 3040 -8548 3080
rect -7936 3400 -7536 3440
rect -7936 3080 -7896 3400
rect -7576 3080 -7536 3400
rect -7936 3040 -7536 3080
rect -6924 3400 -6524 3440
rect -6924 3080 -6884 3400
rect -6564 3080 -6524 3400
rect -6924 3040 -6524 3080
rect -5912 3400 -5512 3440
rect -5912 3080 -5872 3400
rect -5552 3080 -5512 3400
rect -5912 3040 -5512 3080
rect -4900 3400 -4500 3440
rect -4900 3080 -4860 3400
rect -4540 3080 -4500 3400
rect -4900 3040 -4500 3080
rect -3888 3400 -3488 3440
rect -3888 3080 -3848 3400
rect -3528 3080 -3488 3400
rect -3888 3040 -3488 3080
rect -2876 3400 -2476 3440
rect -2876 3080 -2836 3400
rect -2516 3080 -2476 3400
rect -2876 3040 -2476 3080
rect -1864 3400 -1464 3440
rect -1864 3080 -1824 3400
rect -1504 3080 -1464 3400
rect -1864 3040 -1464 3080
rect -852 3400 -452 3440
rect -852 3080 -812 3400
rect -492 3080 -452 3400
rect -852 3040 -452 3080
rect 160 3400 560 3440
rect 160 3080 200 3400
rect 520 3080 560 3400
rect 160 3040 560 3080
rect 1172 3400 1572 3440
rect 1172 3080 1212 3400
rect 1532 3080 1572 3400
rect 1172 3040 1572 3080
rect 2184 3400 2584 3440
rect 2184 3080 2224 3400
rect 2544 3080 2584 3400
rect 2184 3040 2584 3080
rect 3196 3400 3596 3440
rect 3196 3080 3236 3400
rect 3556 3080 3596 3400
rect 3196 3040 3596 3080
rect 4208 3400 4608 3440
rect 4208 3080 4248 3400
rect 4568 3080 4608 3400
rect 4208 3040 4608 3080
rect 5220 3400 5620 3440
rect 5220 3080 5260 3400
rect 5580 3080 5620 3400
rect 5220 3040 5620 3080
rect 6232 3400 6632 3440
rect 6232 3080 6272 3400
rect 6592 3080 6632 3400
rect 6232 3040 6632 3080
rect 7244 3400 7644 3440
rect 7244 3080 7284 3400
rect 7604 3080 7644 3400
rect 7244 3040 7644 3080
rect 8256 3400 8656 3440
rect 8256 3080 8296 3400
rect 8616 3080 8656 3400
rect 8256 3040 8656 3080
rect 9268 3400 9668 3440
rect 9268 3080 9308 3400
rect 9628 3080 9668 3400
rect 9268 3040 9668 3080
rect 10280 3400 10680 3440
rect 10280 3080 10320 3400
rect 10640 3080 10680 3400
rect 10280 3040 10680 3080
rect 11292 3400 11692 3440
rect 11292 3080 11332 3400
rect 11652 3080 11692 3400
rect 11292 3040 11692 3080
rect 12304 3400 12704 3440
rect 12304 3080 12344 3400
rect 12664 3080 12704 3400
rect 12304 3040 12704 3080
rect 13316 3400 13716 3440
rect 13316 3080 13356 3400
rect 13676 3080 13716 3400
rect 13316 3040 13716 3080
rect 14328 3400 14728 3440
rect 14328 3080 14368 3400
rect 14688 3080 14728 3400
rect 14328 3040 14728 3080
rect 15340 3400 15740 3440
rect 15340 3080 15380 3400
rect 15700 3080 15740 3400
rect 15340 3040 15740 3080
rect 16352 3400 16752 3440
rect 16352 3080 16392 3400
rect 16712 3080 16752 3400
rect 16352 3040 16752 3080
rect -17044 2680 -16644 2720
rect -17044 2360 -17004 2680
rect -16684 2360 -16644 2680
rect -17044 2320 -16644 2360
rect -16032 2680 -15632 2720
rect -16032 2360 -15992 2680
rect -15672 2360 -15632 2680
rect -16032 2320 -15632 2360
rect -15020 2680 -14620 2720
rect -15020 2360 -14980 2680
rect -14660 2360 -14620 2680
rect -15020 2320 -14620 2360
rect -14008 2680 -13608 2720
rect -14008 2360 -13968 2680
rect -13648 2360 -13608 2680
rect -14008 2320 -13608 2360
rect -12996 2680 -12596 2720
rect -12996 2360 -12956 2680
rect -12636 2360 -12596 2680
rect -12996 2320 -12596 2360
rect -11984 2680 -11584 2720
rect -11984 2360 -11944 2680
rect -11624 2360 -11584 2680
rect -11984 2320 -11584 2360
rect -10972 2680 -10572 2720
rect -10972 2360 -10932 2680
rect -10612 2360 -10572 2680
rect -10972 2320 -10572 2360
rect -9960 2680 -9560 2720
rect -9960 2360 -9920 2680
rect -9600 2360 -9560 2680
rect -9960 2320 -9560 2360
rect -8948 2680 -8548 2720
rect -8948 2360 -8908 2680
rect -8588 2360 -8548 2680
rect -8948 2320 -8548 2360
rect -7936 2680 -7536 2720
rect -7936 2360 -7896 2680
rect -7576 2360 -7536 2680
rect -7936 2320 -7536 2360
rect -6924 2680 -6524 2720
rect -6924 2360 -6884 2680
rect -6564 2360 -6524 2680
rect -6924 2320 -6524 2360
rect -5912 2680 -5512 2720
rect -5912 2360 -5872 2680
rect -5552 2360 -5512 2680
rect -5912 2320 -5512 2360
rect -4900 2680 -4500 2720
rect -4900 2360 -4860 2680
rect -4540 2360 -4500 2680
rect -4900 2320 -4500 2360
rect -3888 2680 -3488 2720
rect -3888 2360 -3848 2680
rect -3528 2360 -3488 2680
rect -3888 2320 -3488 2360
rect -2876 2680 -2476 2720
rect -2876 2360 -2836 2680
rect -2516 2360 -2476 2680
rect -2876 2320 -2476 2360
rect -1864 2680 -1464 2720
rect -1864 2360 -1824 2680
rect -1504 2360 -1464 2680
rect -1864 2320 -1464 2360
rect -852 2680 -452 2720
rect -852 2360 -812 2680
rect -492 2360 -452 2680
rect -852 2320 -452 2360
rect 160 2680 560 2720
rect 160 2360 200 2680
rect 520 2360 560 2680
rect 160 2320 560 2360
rect 1172 2680 1572 2720
rect 1172 2360 1212 2680
rect 1532 2360 1572 2680
rect 1172 2320 1572 2360
rect 2184 2680 2584 2720
rect 2184 2360 2224 2680
rect 2544 2360 2584 2680
rect 2184 2320 2584 2360
rect 3196 2680 3596 2720
rect 3196 2360 3236 2680
rect 3556 2360 3596 2680
rect 3196 2320 3596 2360
rect 4208 2680 4608 2720
rect 4208 2360 4248 2680
rect 4568 2360 4608 2680
rect 4208 2320 4608 2360
rect 5220 2680 5620 2720
rect 5220 2360 5260 2680
rect 5580 2360 5620 2680
rect 5220 2320 5620 2360
rect 6232 2680 6632 2720
rect 6232 2360 6272 2680
rect 6592 2360 6632 2680
rect 6232 2320 6632 2360
rect 7244 2680 7644 2720
rect 7244 2360 7284 2680
rect 7604 2360 7644 2680
rect 7244 2320 7644 2360
rect 8256 2680 8656 2720
rect 8256 2360 8296 2680
rect 8616 2360 8656 2680
rect 8256 2320 8656 2360
rect 9268 2680 9668 2720
rect 9268 2360 9308 2680
rect 9628 2360 9668 2680
rect 9268 2320 9668 2360
rect 10280 2680 10680 2720
rect 10280 2360 10320 2680
rect 10640 2360 10680 2680
rect 10280 2320 10680 2360
rect 11292 2680 11692 2720
rect 11292 2360 11332 2680
rect 11652 2360 11692 2680
rect 11292 2320 11692 2360
rect 12304 2680 12704 2720
rect 12304 2360 12344 2680
rect 12664 2360 12704 2680
rect 12304 2320 12704 2360
rect 13316 2680 13716 2720
rect 13316 2360 13356 2680
rect 13676 2360 13716 2680
rect 13316 2320 13716 2360
rect 14328 2680 14728 2720
rect 14328 2360 14368 2680
rect 14688 2360 14728 2680
rect 14328 2320 14728 2360
rect 15340 2680 15740 2720
rect 15340 2360 15380 2680
rect 15700 2360 15740 2680
rect 15340 2320 15740 2360
rect 16352 2680 16752 2720
rect 16352 2360 16392 2680
rect 16712 2360 16752 2680
rect 16352 2320 16752 2360
rect -17044 1960 -16644 2000
rect -17044 1640 -17004 1960
rect -16684 1640 -16644 1960
rect -17044 1600 -16644 1640
rect -16032 1960 -15632 2000
rect -16032 1640 -15992 1960
rect -15672 1640 -15632 1960
rect -16032 1600 -15632 1640
rect -15020 1960 -14620 2000
rect -15020 1640 -14980 1960
rect -14660 1640 -14620 1960
rect -15020 1600 -14620 1640
rect -14008 1960 -13608 2000
rect -14008 1640 -13968 1960
rect -13648 1640 -13608 1960
rect -14008 1600 -13608 1640
rect -12996 1960 -12596 2000
rect -12996 1640 -12956 1960
rect -12636 1640 -12596 1960
rect -12996 1600 -12596 1640
rect -11984 1960 -11584 2000
rect -11984 1640 -11944 1960
rect -11624 1640 -11584 1960
rect -11984 1600 -11584 1640
rect -10972 1960 -10572 2000
rect -10972 1640 -10932 1960
rect -10612 1640 -10572 1960
rect -10972 1600 -10572 1640
rect -9960 1960 -9560 2000
rect -9960 1640 -9920 1960
rect -9600 1640 -9560 1960
rect -9960 1600 -9560 1640
rect -8948 1960 -8548 2000
rect -8948 1640 -8908 1960
rect -8588 1640 -8548 1960
rect -8948 1600 -8548 1640
rect -7936 1960 -7536 2000
rect -7936 1640 -7896 1960
rect -7576 1640 -7536 1960
rect -7936 1600 -7536 1640
rect -6924 1960 -6524 2000
rect -6924 1640 -6884 1960
rect -6564 1640 -6524 1960
rect -6924 1600 -6524 1640
rect -5912 1960 -5512 2000
rect -5912 1640 -5872 1960
rect -5552 1640 -5512 1960
rect -5912 1600 -5512 1640
rect -4900 1960 -4500 2000
rect -4900 1640 -4860 1960
rect -4540 1640 -4500 1960
rect -4900 1600 -4500 1640
rect -3888 1960 -3488 2000
rect -3888 1640 -3848 1960
rect -3528 1640 -3488 1960
rect -3888 1600 -3488 1640
rect -2876 1960 -2476 2000
rect -2876 1640 -2836 1960
rect -2516 1640 -2476 1960
rect -2876 1600 -2476 1640
rect -1864 1960 -1464 2000
rect -1864 1640 -1824 1960
rect -1504 1640 -1464 1960
rect -1864 1600 -1464 1640
rect -852 1960 -452 2000
rect -852 1640 -812 1960
rect -492 1640 -452 1960
rect -852 1600 -452 1640
rect 160 1960 560 2000
rect 160 1640 200 1960
rect 520 1640 560 1960
rect 160 1600 560 1640
rect 1172 1960 1572 2000
rect 1172 1640 1212 1960
rect 1532 1640 1572 1960
rect 1172 1600 1572 1640
rect 2184 1960 2584 2000
rect 2184 1640 2224 1960
rect 2544 1640 2584 1960
rect 2184 1600 2584 1640
rect 3196 1960 3596 2000
rect 3196 1640 3236 1960
rect 3556 1640 3596 1960
rect 3196 1600 3596 1640
rect 4208 1960 4608 2000
rect 4208 1640 4248 1960
rect 4568 1640 4608 1960
rect 4208 1600 4608 1640
rect 5220 1960 5620 2000
rect 5220 1640 5260 1960
rect 5580 1640 5620 1960
rect 5220 1600 5620 1640
rect 6232 1960 6632 2000
rect 6232 1640 6272 1960
rect 6592 1640 6632 1960
rect 6232 1600 6632 1640
rect 7244 1960 7644 2000
rect 7244 1640 7284 1960
rect 7604 1640 7644 1960
rect 7244 1600 7644 1640
rect 8256 1960 8656 2000
rect 8256 1640 8296 1960
rect 8616 1640 8656 1960
rect 8256 1600 8656 1640
rect 9268 1960 9668 2000
rect 9268 1640 9308 1960
rect 9628 1640 9668 1960
rect 9268 1600 9668 1640
rect 10280 1960 10680 2000
rect 10280 1640 10320 1960
rect 10640 1640 10680 1960
rect 10280 1600 10680 1640
rect 11292 1960 11692 2000
rect 11292 1640 11332 1960
rect 11652 1640 11692 1960
rect 11292 1600 11692 1640
rect 12304 1960 12704 2000
rect 12304 1640 12344 1960
rect 12664 1640 12704 1960
rect 12304 1600 12704 1640
rect 13316 1960 13716 2000
rect 13316 1640 13356 1960
rect 13676 1640 13716 1960
rect 13316 1600 13716 1640
rect 14328 1960 14728 2000
rect 14328 1640 14368 1960
rect 14688 1640 14728 1960
rect 14328 1600 14728 1640
rect 15340 1960 15740 2000
rect 15340 1640 15380 1960
rect 15700 1640 15740 1960
rect 15340 1600 15740 1640
rect 16352 1960 16752 2000
rect 16352 1640 16392 1960
rect 16712 1640 16752 1960
rect 16352 1600 16752 1640
rect -17044 1240 -16644 1280
rect -17044 920 -17004 1240
rect -16684 920 -16644 1240
rect -17044 880 -16644 920
rect -16032 1240 -15632 1280
rect -16032 920 -15992 1240
rect -15672 920 -15632 1240
rect -16032 880 -15632 920
rect -15020 1240 -14620 1280
rect -15020 920 -14980 1240
rect -14660 920 -14620 1240
rect -15020 880 -14620 920
rect -14008 1240 -13608 1280
rect -14008 920 -13968 1240
rect -13648 920 -13608 1240
rect -14008 880 -13608 920
rect -12996 1240 -12596 1280
rect -12996 920 -12956 1240
rect -12636 920 -12596 1240
rect -12996 880 -12596 920
rect -11984 1240 -11584 1280
rect -11984 920 -11944 1240
rect -11624 920 -11584 1240
rect -11984 880 -11584 920
rect -10972 1240 -10572 1280
rect -10972 920 -10932 1240
rect -10612 920 -10572 1240
rect -10972 880 -10572 920
rect -9960 1240 -9560 1280
rect -9960 920 -9920 1240
rect -9600 920 -9560 1240
rect -9960 880 -9560 920
rect -8948 1240 -8548 1280
rect -8948 920 -8908 1240
rect -8588 920 -8548 1240
rect -8948 880 -8548 920
rect -7936 1240 -7536 1280
rect -7936 920 -7896 1240
rect -7576 920 -7536 1240
rect -7936 880 -7536 920
rect -6924 1240 -6524 1280
rect -6924 920 -6884 1240
rect -6564 920 -6524 1240
rect -6924 880 -6524 920
rect -5912 1240 -5512 1280
rect -5912 920 -5872 1240
rect -5552 920 -5512 1240
rect -5912 880 -5512 920
rect -4900 1240 -4500 1280
rect -4900 920 -4860 1240
rect -4540 920 -4500 1240
rect -4900 880 -4500 920
rect -3888 1240 -3488 1280
rect -3888 920 -3848 1240
rect -3528 920 -3488 1240
rect -3888 880 -3488 920
rect -2876 1240 -2476 1280
rect -2876 920 -2836 1240
rect -2516 920 -2476 1240
rect -2876 880 -2476 920
rect -1864 1240 -1464 1280
rect -1864 920 -1824 1240
rect -1504 920 -1464 1240
rect -1864 880 -1464 920
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect 1172 1240 1572 1280
rect 1172 920 1212 1240
rect 1532 920 1572 1240
rect 1172 880 1572 920
rect 2184 1240 2584 1280
rect 2184 920 2224 1240
rect 2544 920 2584 1240
rect 2184 880 2584 920
rect 3196 1240 3596 1280
rect 3196 920 3236 1240
rect 3556 920 3596 1240
rect 3196 880 3596 920
rect 4208 1240 4608 1280
rect 4208 920 4248 1240
rect 4568 920 4608 1240
rect 4208 880 4608 920
rect 5220 1240 5620 1280
rect 5220 920 5260 1240
rect 5580 920 5620 1240
rect 5220 880 5620 920
rect 6232 1240 6632 1280
rect 6232 920 6272 1240
rect 6592 920 6632 1240
rect 6232 880 6632 920
rect 7244 1240 7644 1280
rect 7244 920 7284 1240
rect 7604 920 7644 1240
rect 7244 880 7644 920
rect 8256 1240 8656 1280
rect 8256 920 8296 1240
rect 8616 920 8656 1240
rect 8256 880 8656 920
rect 9268 1240 9668 1280
rect 9268 920 9308 1240
rect 9628 920 9668 1240
rect 9268 880 9668 920
rect 10280 1240 10680 1280
rect 10280 920 10320 1240
rect 10640 920 10680 1240
rect 10280 880 10680 920
rect 11292 1240 11692 1280
rect 11292 920 11332 1240
rect 11652 920 11692 1240
rect 11292 880 11692 920
rect 12304 1240 12704 1280
rect 12304 920 12344 1240
rect 12664 920 12704 1240
rect 12304 880 12704 920
rect 13316 1240 13716 1280
rect 13316 920 13356 1240
rect 13676 920 13716 1240
rect 13316 880 13716 920
rect 14328 1240 14728 1280
rect 14328 920 14368 1240
rect 14688 920 14728 1240
rect 14328 880 14728 920
rect 15340 1240 15740 1280
rect 15340 920 15380 1240
rect 15700 920 15740 1240
rect 15340 880 15740 920
rect 16352 1240 16752 1280
rect 16352 920 16392 1240
rect 16712 920 16752 1240
rect 16352 880 16752 920
rect -17044 520 -16644 560
rect -17044 200 -17004 520
rect -16684 200 -16644 520
rect -17044 160 -16644 200
rect -16032 520 -15632 560
rect -16032 200 -15992 520
rect -15672 200 -15632 520
rect -16032 160 -15632 200
rect -15020 520 -14620 560
rect -15020 200 -14980 520
rect -14660 200 -14620 520
rect -15020 160 -14620 200
rect -14008 520 -13608 560
rect -14008 200 -13968 520
rect -13648 200 -13608 520
rect -14008 160 -13608 200
rect -12996 520 -12596 560
rect -12996 200 -12956 520
rect -12636 200 -12596 520
rect -12996 160 -12596 200
rect -11984 520 -11584 560
rect -11984 200 -11944 520
rect -11624 200 -11584 520
rect -11984 160 -11584 200
rect -10972 520 -10572 560
rect -10972 200 -10932 520
rect -10612 200 -10572 520
rect -10972 160 -10572 200
rect -9960 520 -9560 560
rect -9960 200 -9920 520
rect -9600 200 -9560 520
rect -9960 160 -9560 200
rect -8948 520 -8548 560
rect -8948 200 -8908 520
rect -8588 200 -8548 520
rect -8948 160 -8548 200
rect -7936 520 -7536 560
rect -7936 200 -7896 520
rect -7576 200 -7536 520
rect -7936 160 -7536 200
rect -6924 520 -6524 560
rect -6924 200 -6884 520
rect -6564 200 -6524 520
rect -6924 160 -6524 200
rect -5912 520 -5512 560
rect -5912 200 -5872 520
rect -5552 200 -5512 520
rect -5912 160 -5512 200
rect -4900 520 -4500 560
rect -4900 200 -4860 520
rect -4540 200 -4500 520
rect -4900 160 -4500 200
rect -3888 520 -3488 560
rect -3888 200 -3848 520
rect -3528 200 -3488 520
rect -3888 160 -3488 200
rect -2876 520 -2476 560
rect -2876 200 -2836 520
rect -2516 200 -2476 520
rect -2876 160 -2476 200
rect -1864 520 -1464 560
rect -1864 200 -1824 520
rect -1504 200 -1464 520
rect -1864 160 -1464 200
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect 1172 520 1572 560
rect 1172 200 1212 520
rect 1532 200 1572 520
rect 1172 160 1572 200
rect 2184 520 2584 560
rect 2184 200 2224 520
rect 2544 200 2584 520
rect 2184 160 2584 200
rect 3196 520 3596 560
rect 3196 200 3236 520
rect 3556 200 3596 520
rect 3196 160 3596 200
rect 4208 520 4608 560
rect 4208 200 4248 520
rect 4568 200 4608 520
rect 4208 160 4608 200
rect 5220 520 5620 560
rect 5220 200 5260 520
rect 5580 200 5620 520
rect 5220 160 5620 200
rect 6232 520 6632 560
rect 6232 200 6272 520
rect 6592 200 6632 520
rect 6232 160 6632 200
rect 7244 520 7644 560
rect 7244 200 7284 520
rect 7604 200 7644 520
rect 7244 160 7644 200
rect 8256 520 8656 560
rect 8256 200 8296 520
rect 8616 200 8656 520
rect 8256 160 8656 200
rect 9268 520 9668 560
rect 9268 200 9308 520
rect 9628 200 9668 520
rect 9268 160 9668 200
rect 10280 520 10680 560
rect 10280 200 10320 520
rect 10640 200 10680 520
rect 10280 160 10680 200
rect 11292 520 11692 560
rect 11292 200 11332 520
rect 11652 200 11692 520
rect 11292 160 11692 200
rect 12304 520 12704 560
rect 12304 200 12344 520
rect 12664 200 12704 520
rect 12304 160 12704 200
rect 13316 520 13716 560
rect 13316 200 13356 520
rect 13676 200 13716 520
rect 13316 160 13716 200
rect 14328 520 14728 560
rect 14328 200 14368 520
rect 14688 200 14728 520
rect 14328 160 14728 200
rect 15340 520 15740 560
rect 15340 200 15380 520
rect 15700 200 15740 520
rect 15340 160 15740 200
rect 16352 520 16752 560
rect 16352 200 16392 520
rect 16712 200 16752 520
rect 16352 160 16752 200
rect -17044 -200 -16644 -160
rect -17044 -520 -17004 -200
rect -16684 -520 -16644 -200
rect -17044 -560 -16644 -520
rect -16032 -200 -15632 -160
rect -16032 -520 -15992 -200
rect -15672 -520 -15632 -200
rect -16032 -560 -15632 -520
rect -15020 -200 -14620 -160
rect -15020 -520 -14980 -200
rect -14660 -520 -14620 -200
rect -15020 -560 -14620 -520
rect -14008 -200 -13608 -160
rect -14008 -520 -13968 -200
rect -13648 -520 -13608 -200
rect -14008 -560 -13608 -520
rect -12996 -200 -12596 -160
rect -12996 -520 -12956 -200
rect -12636 -520 -12596 -200
rect -12996 -560 -12596 -520
rect -11984 -200 -11584 -160
rect -11984 -520 -11944 -200
rect -11624 -520 -11584 -200
rect -11984 -560 -11584 -520
rect -10972 -200 -10572 -160
rect -10972 -520 -10932 -200
rect -10612 -520 -10572 -200
rect -10972 -560 -10572 -520
rect -9960 -200 -9560 -160
rect -9960 -520 -9920 -200
rect -9600 -520 -9560 -200
rect -9960 -560 -9560 -520
rect -8948 -200 -8548 -160
rect -8948 -520 -8908 -200
rect -8588 -520 -8548 -200
rect -8948 -560 -8548 -520
rect -7936 -200 -7536 -160
rect -7936 -520 -7896 -200
rect -7576 -520 -7536 -200
rect -7936 -560 -7536 -520
rect -6924 -200 -6524 -160
rect -6924 -520 -6884 -200
rect -6564 -520 -6524 -200
rect -6924 -560 -6524 -520
rect -5912 -200 -5512 -160
rect -5912 -520 -5872 -200
rect -5552 -520 -5512 -200
rect -5912 -560 -5512 -520
rect -4900 -200 -4500 -160
rect -4900 -520 -4860 -200
rect -4540 -520 -4500 -200
rect -4900 -560 -4500 -520
rect -3888 -200 -3488 -160
rect -3888 -520 -3848 -200
rect -3528 -520 -3488 -200
rect -3888 -560 -3488 -520
rect -2876 -200 -2476 -160
rect -2876 -520 -2836 -200
rect -2516 -520 -2476 -200
rect -2876 -560 -2476 -520
rect -1864 -200 -1464 -160
rect -1864 -520 -1824 -200
rect -1504 -520 -1464 -200
rect -1864 -560 -1464 -520
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect 1172 -200 1572 -160
rect 1172 -520 1212 -200
rect 1532 -520 1572 -200
rect 1172 -560 1572 -520
rect 2184 -200 2584 -160
rect 2184 -520 2224 -200
rect 2544 -520 2584 -200
rect 2184 -560 2584 -520
rect 3196 -200 3596 -160
rect 3196 -520 3236 -200
rect 3556 -520 3596 -200
rect 3196 -560 3596 -520
rect 4208 -200 4608 -160
rect 4208 -520 4248 -200
rect 4568 -520 4608 -200
rect 4208 -560 4608 -520
rect 5220 -200 5620 -160
rect 5220 -520 5260 -200
rect 5580 -520 5620 -200
rect 5220 -560 5620 -520
rect 6232 -200 6632 -160
rect 6232 -520 6272 -200
rect 6592 -520 6632 -200
rect 6232 -560 6632 -520
rect 7244 -200 7644 -160
rect 7244 -520 7284 -200
rect 7604 -520 7644 -200
rect 7244 -560 7644 -520
rect 8256 -200 8656 -160
rect 8256 -520 8296 -200
rect 8616 -520 8656 -200
rect 8256 -560 8656 -520
rect 9268 -200 9668 -160
rect 9268 -520 9308 -200
rect 9628 -520 9668 -200
rect 9268 -560 9668 -520
rect 10280 -200 10680 -160
rect 10280 -520 10320 -200
rect 10640 -520 10680 -200
rect 10280 -560 10680 -520
rect 11292 -200 11692 -160
rect 11292 -520 11332 -200
rect 11652 -520 11692 -200
rect 11292 -560 11692 -520
rect 12304 -200 12704 -160
rect 12304 -520 12344 -200
rect 12664 -520 12704 -200
rect 12304 -560 12704 -520
rect 13316 -200 13716 -160
rect 13316 -520 13356 -200
rect 13676 -520 13716 -200
rect 13316 -560 13716 -520
rect 14328 -200 14728 -160
rect 14328 -520 14368 -200
rect 14688 -520 14728 -200
rect 14328 -560 14728 -520
rect 15340 -200 15740 -160
rect 15340 -520 15380 -200
rect 15700 -520 15740 -200
rect 15340 -560 15740 -520
rect 16352 -200 16752 -160
rect 16352 -520 16392 -200
rect 16712 -520 16752 -200
rect 16352 -560 16752 -520
rect -17044 -920 -16644 -880
rect -17044 -1240 -17004 -920
rect -16684 -1240 -16644 -920
rect -17044 -1280 -16644 -1240
rect -16032 -920 -15632 -880
rect -16032 -1240 -15992 -920
rect -15672 -1240 -15632 -920
rect -16032 -1280 -15632 -1240
rect -15020 -920 -14620 -880
rect -15020 -1240 -14980 -920
rect -14660 -1240 -14620 -920
rect -15020 -1280 -14620 -1240
rect -14008 -920 -13608 -880
rect -14008 -1240 -13968 -920
rect -13648 -1240 -13608 -920
rect -14008 -1280 -13608 -1240
rect -12996 -920 -12596 -880
rect -12996 -1240 -12956 -920
rect -12636 -1240 -12596 -920
rect -12996 -1280 -12596 -1240
rect -11984 -920 -11584 -880
rect -11984 -1240 -11944 -920
rect -11624 -1240 -11584 -920
rect -11984 -1280 -11584 -1240
rect -10972 -920 -10572 -880
rect -10972 -1240 -10932 -920
rect -10612 -1240 -10572 -920
rect -10972 -1280 -10572 -1240
rect -9960 -920 -9560 -880
rect -9960 -1240 -9920 -920
rect -9600 -1240 -9560 -920
rect -9960 -1280 -9560 -1240
rect -8948 -920 -8548 -880
rect -8948 -1240 -8908 -920
rect -8588 -1240 -8548 -920
rect -8948 -1280 -8548 -1240
rect -7936 -920 -7536 -880
rect -7936 -1240 -7896 -920
rect -7576 -1240 -7536 -920
rect -7936 -1280 -7536 -1240
rect -6924 -920 -6524 -880
rect -6924 -1240 -6884 -920
rect -6564 -1240 -6524 -920
rect -6924 -1280 -6524 -1240
rect -5912 -920 -5512 -880
rect -5912 -1240 -5872 -920
rect -5552 -1240 -5512 -920
rect -5912 -1280 -5512 -1240
rect -4900 -920 -4500 -880
rect -4900 -1240 -4860 -920
rect -4540 -1240 -4500 -920
rect -4900 -1280 -4500 -1240
rect -3888 -920 -3488 -880
rect -3888 -1240 -3848 -920
rect -3528 -1240 -3488 -920
rect -3888 -1280 -3488 -1240
rect -2876 -920 -2476 -880
rect -2876 -1240 -2836 -920
rect -2516 -1240 -2476 -920
rect -2876 -1280 -2476 -1240
rect -1864 -920 -1464 -880
rect -1864 -1240 -1824 -920
rect -1504 -1240 -1464 -920
rect -1864 -1280 -1464 -1240
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect 1172 -920 1572 -880
rect 1172 -1240 1212 -920
rect 1532 -1240 1572 -920
rect 1172 -1280 1572 -1240
rect 2184 -920 2584 -880
rect 2184 -1240 2224 -920
rect 2544 -1240 2584 -920
rect 2184 -1280 2584 -1240
rect 3196 -920 3596 -880
rect 3196 -1240 3236 -920
rect 3556 -1240 3596 -920
rect 3196 -1280 3596 -1240
rect 4208 -920 4608 -880
rect 4208 -1240 4248 -920
rect 4568 -1240 4608 -920
rect 4208 -1280 4608 -1240
rect 5220 -920 5620 -880
rect 5220 -1240 5260 -920
rect 5580 -1240 5620 -920
rect 5220 -1280 5620 -1240
rect 6232 -920 6632 -880
rect 6232 -1240 6272 -920
rect 6592 -1240 6632 -920
rect 6232 -1280 6632 -1240
rect 7244 -920 7644 -880
rect 7244 -1240 7284 -920
rect 7604 -1240 7644 -920
rect 7244 -1280 7644 -1240
rect 8256 -920 8656 -880
rect 8256 -1240 8296 -920
rect 8616 -1240 8656 -920
rect 8256 -1280 8656 -1240
rect 9268 -920 9668 -880
rect 9268 -1240 9308 -920
rect 9628 -1240 9668 -920
rect 9268 -1280 9668 -1240
rect 10280 -920 10680 -880
rect 10280 -1240 10320 -920
rect 10640 -1240 10680 -920
rect 10280 -1280 10680 -1240
rect 11292 -920 11692 -880
rect 11292 -1240 11332 -920
rect 11652 -1240 11692 -920
rect 11292 -1280 11692 -1240
rect 12304 -920 12704 -880
rect 12304 -1240 12344 -920
rect 12664 -1240 12704 -920
rect 12304 -1280 12704 -1240
rect 13316 -920 13716 -880
rect 13316 -1240 13356 -920
rect 13676 -1240 13716 -920
rect 13316 -1280 13716 -1240
rect 14328 -920 14728 -880
rect 14328 -1240 14368 -920
rect 14688 -1240 14728 -920
rect 14328 -1280 14728 -1240
rect 15340 -920 15740 -880
rect 15340 -1240 15380 -920
rect 15700 -1240 15740 -920
rect 15340 -1280 15740 -1240
rect 16352 -920 16752 -880
rect 16352 -1240 16392 -920
rect 16712 -1240 16752 -920
rect 16352 -1280 16752 -1240
rect -17044 -1640 -16644 -1600
rect -17044 -1960 -17004 -1640
rect -16684 -1960 -16644 -1640
rect -17044 -2000 -16644 -1960
rect -16032 -1640 -15632 -1600
rect -16032 -1960 -15992 -1640
rect -15672 -1960 -15632 -1640
rect -16032 -2000 -15632 -1960
rect -15020 -1640 -14620 -1600
rect -15020 -1960 -14980 -1640
rect -14660 -1960 -14620 -1640
rect -15020 -2000 -14620 -1960
rect -14008 -1640 -13608 -1600
rect -14008 -1960 -13968 -1640
rect -13648 -1960 -13608 -1640
rect -14008 -2000 -13608 -1960
rect -12996 -1640 -12596 -1600
rect -12996 -1960 -12956 -1640
rect -12636 -1960 -12596 -1640
rect -12996 -2000 -12596 -1960
rect -11984 -1640 -11584 -1600
rect -11984 -1960 -11944 -1640
rect -11624 -1960 -11584 -1640
rect -11984 -2000 -11584 -1960
rect -10972 -1640 -10572 -1600
rect -10972 -1960 -10932 -1640
rect -10612 -1960 -10572 -1640
rect -10972 -2000 -10572 -1960
rect -9960 -1640 -9560 -1600
rect -9960 -1960 -9920 -1640
rect -9600 -1960 -9560 -1640
rect -9960 -2000 -9560 -1960
rect -8948 -1640 -8548 -1600
rect -8948 -1960 -8908 -1640
rect -8588 -1960 -8548 -1640
rect -8948 -2000 -8548 -1960
rect -7936 -1640 -7536 -1600
rect -7936 -1960 -7896 -1640
rect -7576 -1960 -7536 -1640
rect -7936 -2000 -7536 -1960
rect -6924 -1640 -6524 -1600
rect -6924 -1960 -6884 -1640
rect -6564 -1960 -6524 -1640
rect -6924 -2000 -6524 -1960
rect -5912 -1640 -5512 -1600
rect -5912 -1960 -5872 -1640
rect -5552 -1960 -5512 -1640
rect -5912 -2000 -5512 -1960
rect -4900 -1640 -4500 -1600
rect -4900 -1960 -4860 -1640
rect -4540 -1960 -4500 -1640
rect -4900 -2000 -4500 -1960
rect -3888 -1640 -3488 -1600
rect -3888 -1960 -3848 -1640
rect -3528 -1960 -3488 -1640
rect -3888 -2000 -3488 -1960
rect -2876 -1640 -2476 -1600
rect -2876 -1960 -2836 -1640
rect -2516 -1960 -2476 -1640
rect -2876 -2000 -2476 -1960
rect -1864 -1640 -1464 -1600
rect -1864 -1960 -1824 -1640
rect -1504 -1960 -1464 -1640
rect -1864 -2000 -1464 -1960
rect -852 -1640 -452 -1600
rect -852 -1960 -812 -1640
rect -492 -1960 -452 -1640
rect -852 -2000 -452 -1960
rect 160 -1640 560 -1600
rect 160 -1960 200 -1640
rect 520 -1960 560 -1640
rect 160 -2000 560 -1960
rect 1172 -1640 1572 -1600
rect 1172 -1960 1212 -1640
rect 1532 -1960 1572 -1640
rect 1172 -2000 1572 -1960
rect 2184 -1640 2584 -1600
rect 2184 -1960 2224 -1640
rect 2544 -1960 2584 -1640
rect 2184 -2000 2584 -1960
rect 3196 -1640 3596 -1600
rect 3196 -1960 3236 -1640
rect 3556 -1960 3596 -1640
rect 3196 -2000 3596 -1960
rect 4208 -1640 4608 -1600
rect 4208 -1960 4248 -1640
rect 4568 -1960 4608 -1640
rect 4208 -2000 4608 -1960
rect 5220 -1640 5620 -1600
rect 5220 -1960 5260 -1640
rect 5580 -1960 5620 -1640
rect 5220 -2000 5620 -1960
rect 6232 -1640 6632 -1600
rect 6232 -1960 6272 -1640
rect 6592 -1960 6632 -1640
rect 6232 -2000 6632 -1960
rect 7244 -1640 7644 -1600
rect 7244 -1960 7284 -1640
rect 7604 -1960 7644 -1640
rect 7244 -2000 7644 -1960
rect 8256 -1640 8656 -1600
rect 8256 -1960 8296 -1640
rect 8616 -1960 8656 -1640
rect 8256 -2000 8656 -1960
rect 9268 -1640 9668 -1600
rect 9268 -1960 9308 -1640
rect 9628 -1960 9668 -1640
rect 9268 -2000 9668 -1960
rect 10280 -1640 10680 -1600
rect 10280 -1960 10320 -1640
rect 10640 -1960 10680 -1640
rect 10280 -2000 10680 -1960
rect 11292 -1640 11692 -1600
rect 11292 -1960 11332 -1640
rect 11652 -1960 11692 -1640
rect 11292 -2000 11692 -1960
rect 12304 -1640 12704 -1600
rect 12304 -1960 12344 -1640
rect 12664 -1960 12704 -1640
rect 12304 -2000 12704 -1960
rect 13316 -1640 13716 -1600
rect 13316 -1960 13356 -1640
rect 13676 -1960 13716 -1640
rect 13316 -2000 13716 -1960
rect 14328 -1640 14728 -1600
rect 14328 -1960 14368 -1640
rect 14688 -1960 14728 -1640
rect 14328 -2000 14728 -1960
rect 15340 -1640 15740 -1600
rect 15340 -1960 15380 -1640
rect 15700 -1960 15740 -1640
rect 15340 -2000 15740 -1960
rect 16352 -1640 16752 -1600
rect 16352 -1960 16392 -1640
rect 16712 -1960 16752 -1640
rect 16352 -2000 16752 -1960
rect -17044 -2360 -16644 -2320
rect -17044 -2680 -17004 -2360
rect -16684 -2680 -16644 -2360
rect -17044 -2720 -16644 -2680
rect -16032 -2360 -15632 -2320
rect -16032 -2680 -15992 -2360
rect -15672 -2680 -15632 -2360
rect -16032 -2720 -15632 -2680
rect -15020 -2360 -14620 -2320
rect -15020 -2680 -14980 -2360
rect -14660 -2680 -14620 -2360
rect -15020 -2720 -14620 -2680
rect -14008 -2360 -13608 -2320
rect -14008 -2680 -13968 -2360
rect -13648 -2680 -13608 -2360
rect -14008 -2720 -13608 -2680
rect -12996 -2360 -12596 -2320
rect -12996 -2680 -12956 -2360
rect -12636 -2680 -12596 -2360
rect -12996 -2720 -12596 -2680
rect -11984 -2360 -11584 -2320
rect -11984 -2680 -11944 -2360
rect -11624 -2680 -11584 -2360
rect -11984 -2720 -11584 -2680
rect -10972 -2360 -10572 -2320
rect -10972 -2680 -10932 -2360
rect -10612 -2680 -10572 -2360
rect -10972 -2720 -10572 -2680
rect -9960 -2360 -9560 -2320
rect -9960 -2680 -9920 -2360
rect -9600 -2680 -9560 -2360
rect -9960 -2720 -9560 -2680
rect -8948 -2360 -8548 -2320
rect -8948 -2680 -8908 -2360
rect -8588 -2680 -8548 -2360
rect -8948 -2720 -8548 -2680
rect -7936 -2360 -7536 -2320
rect -7936 -2680 -7896 -2360
rect -7576 -2680 -7536 -2360
rect -7936 -2720 -7536 -2680
rect -6924 -2360 -6524 -2320
rect -6924 -2680 -6884 -2360
rect -6564 -2680 -6524 -2360
rect -6924 -2720 -6524 -2680
rect -5912 -2360 -5512 -2320
rect -5912 -2680 -5872 -2360
rect -5552 -2680 -5512 -2360
rect -5912 -2720 -5512 -2680
rect -4900 -2360 -4500 -2320
rect -4900 -2680 -4860 -2360
rect -4540 -2680 -4500 -2360
rect -4900 -2720 -4500 -2680
rect -3888 -2360 -3488 -2320
rect -3888 -2680 -3848 -2360
rect -3528 -2680 -3488 -2360
rect -3888 -2720 -3488 -2680
rect -2876 -2360 -2476 -2320
rect -2876 -2680 -2836 -2360
rect -2516 -2680 -2476 -2360
rect -2876 -2720 -2476 -2680
rect -1864 -2360 -1464 -2320
rect -1864 -2680 -1824 -2360
rect -1504 -2680 -1464 -2360
rect -1864 -2720 -1464 -2680
rect -852 -2360 -452 -2320
rect -852 -2680 -812 -2360
rect -492 -2680 -452 -2360
rect -852 -2720 -452 -2680
rect 160 -2360 560 -2320
rect 160 -2680 200 -2360
rect 520 -2680 560 -2360
rect 160 -2720 560 -2680
rect 1172 -2360 1572 -2320
rect 1172 -2680 1212 -2360
rect 1532 -2680 1572 -2360
rect 1172 -2720 1572 -2680
rect 2184 -2360 2584 -2320
rect 2184 -2680 2224 -2360
rect 2544 -2680 2584 -2360
rect 2184 -2720 2584 -2680
rect 3196 -2360 3596 -2320
rect 3196 -2680 3236 -2360
rect 3556 -2680 3596 -2360
rect 3196 -2720 3596 -2680
rect 4208 -2360 4608 -2320
rect 4208 -2680 4248 -2360
rect 4568 -2680 4608 -2360
rect 4208 -2720 4608 -2680
rect 5220 -2360 5620 -2320
rect 5220 -2680 5260 -2360
rect 5580 -2680 5620 -2360
rect 5220 -2720 5620 -2680
rect 6232 -2360 6632 -2320
rect 6232 -2680 6272 -2360
rect 6592 -2680 6632 -2360
rect 6232 -2720 6632 -2680
rect 7244 -2360 7644 -2320
rect 7244 -2680 7284 -2360
rect 7604 -2680 7644 -2360
rect 7244 -2720 7644 -2680
rect 8256 -2360 8656 -2320
rect 8256 -2680 8296 -2360
rect 8616 -2680 8656 -2360
rect 8256 -2720 8656 -2680
rect 9268 -2360 9668 -2320
rect 9268 -2680 9308 -2360
rect 9628 -2680 9668 -2360
rect 9268 -2720 9668 -2680
rect 10280 -2360 10680 -2320
rect 10280 -2680 10320 -2360
rect 10640 -2680 10680 -2360
rect 10280 -2720 10680 -2680
rect 11292 -2360 11692 -2320
rect 11292 -2680 11332 -2360
rect 11652 -2680 11692 -2360
rect 11292 -2720 11692 -2680
rect 12304 -2360 12704 -2320
rect 12304 -2680 12344 -2360
rect 12664 -2680 12704 -2360
rect 12304 -2720 12704 -2680
rect 13316 -2360 13716 -2320
rect 13316 -2680 13356 -2360
rect 13676 -2680 13716 -2360
rect 13316 -2720 13716 -2680
rect 14328 -2360 14728 -2320
rect 14328 -2680 14368 -2360
rect 14688 -2680 14728 -2360
rect 14328 -2720 14728 -2680
rect 15340 -2360 15740 -2320
rect 15340 -2680 15380 -2360
rect 15700 -2680 15740 -2360
rect 15340 -2720 15740 -2680
rect 16352 -2360 16752 -2320
rect 16352 -2680 16392 -2360
rect 16712 -2680 16752 -2360
rect 16352 -2720 16752 -2680
rect -17044 -3080 -16644 -3040
rect -17044 -3400 -17004 -3080
rect -16684 -3400 -16644 -3080
rect -17044 -3440 -16644 -3400
rect -16032 -3080 -15632 -3040
rect -16032 -3400 -15992 -3080
rect -15672 -3400 -15632 -3080
rect -16032 -3440 -15632 -3400
rect -15020 -3080 -14620 -3040
rect -15020 -3400 -14980 -3080
rect -14660 -3400 -14620 -3080
rect -15020 -3440 -14620 -3400
rect -14008 -3080 -13608 -3040
rect -14008 -3400 -13968 -3080
rect -13648 -3400 -13608 -3080
rect -14008 -3440 -13608 -3400
rect -12996 -3080 -12596 -3040
rect -12996 -3400 -12956 -3080
rect -12636 -3400 -12596 -3080
rect -12996 -3440 -12596 -3400
rect -11984 -3080 -11584 -3040
rect -11984 -3400 -11944 -3080
rect -11624 -3400 -11584 -3080
rect -11984 -3440 -11584 -3400
rect -10972 -3080 -10572 -3040
rect -10972 -3400 -10932 -3080
rect -10612 -3400 -10572 -3080
rect -10972 -3440 -10572 -3400
rect -9960 -3080 -9560 -3040
rect -9960 -3400 -9920 -3080
rect -9600 -3400 -9560 -3080
rect -9960 -3440 -9560 -3400
rect -8948 -3080 -8548 -3040
rect -8948 -3400 -8908 -3080
rect -8588 -3400 -8548 -3080
rect -8948 -3440 -8548 -3400
rect -7936 -3080 -7536 -3040
rect -7936 -3400 -7896 -3080
rect -7576 -3400 -7536 -3080
rect -7936 -3440 -7536 -3400
rect -6924 -3080 -6524 -3040
rect -6924 -3400 -6884 -3080
rect -6564 -3400 -6524 -3080
rect -6924 -3440 -6524 -3400
rect -5912 -3080 -5512 -3040
rect -5912 -3400 -5872 -3080
rect -5552 -3400 -5512 -3080
rect -5912 -3440 -5512 -3400
rect -4900 -3080 -4500 -3040
rect -4900 -3400 -4860 -3080
rect -4540 -3400 -4500 -3080
rect -4900 -3440 -4500 -3400
rect -3888 -3080 -3488 -3040
rect -3888 -3400 -3848 -3080
rect -3528 -3400 -3488 -3080
rect -3888 -3440 -3488 -3400
rect -2876 -3080 -2476 -3040
rect -2876 -3400 -2836 -3080
rect -2516 -3400 -2476 -3080
rect -2876 -3440 -2476 -3400
rect -1864 -3080 -1464 -3040
rect -1864 -3400 -1824 -3080
rect -1504 -3400 -1464 -3080
rect -1864 -3440 -1464 -3400
rect -852 -3080 -452 -3040
rect -852 -3400 -812 -3080
rect -492 -3400 -452 -3080
rect -852 -3440 -452 -3400
rect 160 -3080 560 -3040
rect 160 -3400 200 -3080
rect 520 -3400 560 -3080
rect 160 -3440 560 -3400
rect 1172 -3080 1572 -3040
rect 1172 -3400 1212 -3080
rect 1532 -3400 1572 -3080
rect 1172 -3440 1572 -3400
rect 2184 -3080 2584 -3040
rect 2184 -3400 2224 -3080
rect 2544 -3400 2584 -3080
rect 2184 -3440 2584 -3400
rect 3196 -3080 3596 -3040
rect 3196 -3400 3236 -3080
rect 3556 -3400 3596 -3080
rect 3196 -3440 3596 -3400
rect 4208 -3080 4608 -3040
rect 4208 -3400 4248 -3080
rect 4568 -3400 4608 -3080
rect 4208 -3440 4608 -3400
rect 5220 -3080 5620 -3040
rect 5220 -3400 5260 -3080
rect 5580 -3400 5620 -3080
rect 5220 -3440 5620 -3400
rect 6232 -3080 6632 -3040
rect 6232 -3400 6272 -3080
rect 6592 -3400 6632 -3080
rect 6232 -3440 6632 -3400
rect 7244 -3080 7644 -3040
rect 7244 -3400 7284 -3080
rect 7604 -3400 7644 -3080
rect 7244 -3440 7644 -3400
rect 8256 -3080 8656 -3040
rect 8256 -3400 8296 -3080
rect 8616 -3400 8656 -3080
rect 8256 -3440 8656 -3400
rect 9268 -3080 9668 -3040
rect 9268 -3400 9308 -3080
rect 9628 -3400 9668 -3080
rect 9268 -3440 9668 -3400
rect 10280 -3080 10680 -3040
rect 10280 -3400 10320 -3080
rect 10640 -3400 10680 -3080
rect 10280 -3440 10680 -3400
rect 11292 -3080 11692 -3040
rect 11292 -3400 11332 -3080
rect 11652 -3400 11692 -3080
rect 11292 -3440 11692 -3400
rect 12304 -3080 12704 -3040
rect 12304 -3400 12344 -3080
rect 12664 -3400 12704 -3080
rect 12304 -3440 12704 -3400
rect 13316 -3080 13716 -3040
rect 13316 -3400 13356 -3080
rect 13676 -3400 13716 -3080
rect 13316 -3440 13716 -3400
rect 14328 -3080 14728 -3040
rect 14328 -3400 14368 -3080
rect 14688 -3400 14728 -3080
rect 14328 -3440 14728 -3400
rect 15340 -3080 15740 -3040
rect 15340 -3400 15380 -3080
rect 15700 -3400 15740 -3080
rect 15340 -3440 15740 -3400
rect 16352 -3080 16752 -3040
rect 16352 -3400 16392 -3080
rect 16712 -3400 16752 -3080
rect 16352 -3440 16752 -3400
rect -17044 -3800 -16644 -3760
rect -17044 -4120 -17004 -3800
rect -16684 -4120 -16644 -3800
rect -17044 -4160 -16644 -4120
rect -16032 -3800 -15632 -3760
rect -16032 -4120 -15992 -3800
rect -15672 -4120 -15632 -3800
rect -16032 -4160 -15632 -4120
rect -15020 -3800 -14620 -3760
rect -15020 -4120 -14980 -3800
rect -14660 -4120 -14620 -3800
rect -15020 -4160 -14620 -4120
rect -14008 -3800 -13608 -3760
rect -14008 -4120 -13968 -3800
rect -13648 -4120 -13608 -3800
rect -14008 -4160 -13608 -4120
rect -12996 -3800 -12596 -3760
rect -12996 -4120 -12956 -3800
rect -12636 -4120 -12596 -3800
rect -12996 -4160 -12596 -4120
rect -11984 -3800 -11584 -3760
rect -11984 -4120 -11944 -3800
rect -11624 -4120 -11584 -3800
rect -11984 -4160 -11584 -4120
rect -10972 -3800 -10572 -3760
rect -10972 -4120 -10932 -3800
rect -10612 -4120 -10572 -3800
rect -10972 -4160 -10572 -4120
rect -9960 -3800 -9560 -3760
rect -9960 -4120 -9920 -3800
rect -9600 -4120 -9560 -3800
rect -9960 -4160 -9560 -4120
rect -8948 -3800 -8548 -3760
rect -8948 -4120 -8908 -3800
rect -8588 -4120 -8548 -3800
rect -8948 -4160 -8548 -4120
rect -7936 -3800 -7536 -3760
rect -7936 -4120 -7896 -3800
rect -7576 -4120 -7536 -3800
rect -7936 -4160 -7536 -4120
rect -6924 -3800 -6524 -3760
rect -6924 -4120 -6884 -3800
rect -6564 -4120 -6524 -3800
rect -6924 -4160 -6524 -4120
rect -5912 -3800 -5512 -3760
rect -5912 -4120 -5872 -3800
rect -5552 -4120 -5512 -3800
rect -5912 -4160 -5512 -4120
rect -4900 -3800 -4500 -3760
rect -4900 -4120 -4860 -3800
rect -4540 -4120 -4500 -3800
rect -4900 -4160 -4500 -4120
rect -3888 -3800 -3488 -3760
rect -3888 -4120 -3848 -3800
rect -3528 -4120 -3488 -3800
rect -3888 -4160 -3488 -4120
rect -2876 -3800 -2476 -3760
rect -2876 -4120 -2836 -3800
rect -2516 -4120 -2476 -3800
rect -2876 -4160 -2476 -4120
rect -1864 -3800 -1464 -3760
rect -1864 -4120 -1824 -3800
rect -1504 -4120 -1464 -3800
rect -1864 -4160 -1464 -4120
rect -852 -3800 -452 -3760
rect -852 -4120 -812 -3800
rect -492 -4120 -452 -3800
rect -852 -4160 -452 -4120
rect 160 -3800 560 -3760
rect 160 -4120 200 -3800
rect 520 -4120 560 -3800
rect 160 -4160 560 -4120
rect 1172 -3800 1572 -3760
rect 1172 -4120 1212 -3800
rect 1532 -4120 1572 -3800
rect 1172 -4160 1572 -4120
rect 2184 -3800 2584 -3760
rect 2184 -4120 2224 -3800
rect 2544 -4120 2584 -3800
rect 2184 -4160 2584 -4120
rect 3196 -3800 3596 -3760
rect 3196 -4120 3236 -3800
rect 3556 -4120 3596 -3800
rect 3196 -4160 3596 -4120
rect 4208 -3800 4608 -3760
rect 4208 -4120 4248 -3800
rect 4568 -4120 4608 -3800
rect 4208 -4160 4608 -4120
rect 5220 -3800 5620 -3760
rect 5220 -4120 5260 -3800
rect 5580 -4120 5620 -3800
rect 5220 -4160 5620 -4120
rect 6232 -3800 6632 -3760
rect 6232 -4120 6272 -3800
rect 6592 -4120 6632 -3800
rect 6232 -4160 6632 -4120
rect 7244 -3800 7644 -3760
rect 7244 -4120 7284 -3800
rect 7604 -4120 7644 -3800
rect 7244 -4160 7644 -4120
rect 8256 -3800 8656 -3760
rect 8256 -4120 8296 -3800
rect 8616 -4120 8656 -3800
rect 8256 -4160 8656 -4120
rect 9268 -3800 9668 -3760
rect 9268 -4120 9308 -3800
rect 9628 -4120 9668 -3800
rect 9268 -4160 9668 -4120
rect 10280 -3800 10680 -3760
rect 10280 -4120 10320 -3800
rect 10640 -4120 10680 -3800
rect 10280 -4160 10680 -4120
rect 11292 -3800 11692 -3760
rect 11292 -4120 11332 -3800
rect 11652 -4120 11692 -3800
rect 11292 -4160 11692 -4120
rect 12304 -3800 12704 -3760
rect 12304 -4120 12344 -3800
rect 12664 -4120 12704 -3800
rect 12304 -4160 12704 -4120
rect 13316 -3800 13716 -3760
rect 13316 -4120 13356 -3800
rect 13676 -4120 13716 -3800
rect 13316 -4160 13716 -4120
rect 14328 -3800 14728 -3760
rect 14328 -4120 14368 -3800
rect 14688 -4120 14728 -3800
rect 14328 -4160 14728 -4120
rect 15340 -3800 15740 -3760
rect 15340 -4120 15380 -3800
rect 15700 -4120 15740 -3800
rect 15340 -4160 15740 -4120
rect 16352 -3800 16752 -3760
rect 16352 -4120 16392 -3800
rect 16712 -4120 16752 -3800
rect 16352 -4160 16752 -4120
rect -17044 -4520 -16644 -4480
rect -17044 -4840 -17004 -4520
rect -16684 -4840 -16644 -4520
rect -17044 -4880 -16644 -4840
rect -16032 -4520 -15632 -4480
rect -16032 -4840 -15992 -4520
rect -15672 -4840 -15632 -4520
rect -16032 -4880 -15632 -4840
rect -15020 -4520 -14620 -4480
rect -15020 -4840 -14980 -4520
rect -14660 -4840 -14620 -4520
rect -15020 -4880 -14620 -4840
rect -14008 -4520 -13608 -4480
rect -14008 -4840 -13968 -4520
rect -13648 -4840 -13608 -4520
rect -14008 -4880 -13608 -4840
rect -12996 -4520 -12596 -4480
rect -12996 -4840 -12956 -4520
rect -12636 -4840 -12596 -4520
rect -12996 -4880 -12596 -4840
rect -11984 -4520 -11584 -4480
rect -11984 -4840 -11944 -4520
rect -11624 -4840 -11584 -4520
rect -11984 -4880 -11584 -4840
rect -10972 -4520 -10572 -4480
rect -10972 -4840 -10932 -4520
rect -10612 -4840 -10572 -4520
rect -10972 -4880 -10572 -4840
rect -9960 -4520 -9560 -4480
rect -9960 -4840 -9920 -4520
rect -9600 -4840 -9560 -4520
rect -9960 -4880 -9560 -4840
rect -8948 -4520 -8548 -4480
rect -8948 -4840 -8908 -4520
rect -8588 -4840 -8548 -4520
rect -8948 -4880 -8548 -4840
rect -7936 -4520 -7536 -4480
rect -7936 -4840 -7896 -4520
rect -7576 -4840 -7536 -4520
rect -7936 -4880 -7536 -4840
rect -6924 -4520 -6524 -4480
rect -6924 -4840 -6884 -4520
rect -6564 -4840 -6524 -4520
rect -6924 -4880 -6524 -4840
rect -5912 -4520 -5512 -4480
rect -5912 -4840 -5872 -4520
rect -5552 -4840 -5512 -4520
rect -5912 -4880 -5512 -4840
rect -4900 -4520 -4500 -4480
rect -4900 -4840 -4860 -4520
rect -4540 -4840 -4500 -4520
rect -4900 -4880 -4500 -4840
rect -3888 -4520 -3488 -4480
rect -3888 -4840 -3848 -4520
rect -3528 -4840 -3488 -4520
rect -3888 -4880 -3488 -4840
rect -2876 -4520 -2476 -4480
rect -2876 -4840 -2836 -4520
rect -2516 -4840 -2476 -4520
rect -2876 -4880 -2476 -4840
rect -1864 -4520 -1464 -4480
rect -1864 -4840 -1824 -4520
rect -1504 -4840 -1464 -4520
rect -1864 -4880 -1464 -4840
rect -852 -4520 -452 -4480
rect -852 -4840 -812 -4520
rect -492 -4840 -452 -4520
rect -852 -4880 -452 -4840
rect 160 -4520 560 -4480
rect 160 -4840 200 -4520
rect 520 -4840 560 -4520
rect 160 -4880 560 -4840
rect 1172 -4520 1572 -4480
rect 1172 -4840 1212 -4520
rect 1532 -4840 1572 -4520
rect 1172 -4880 1572 -4840
rect 2184 -4520 2584 -4480
rect 2184 -4840 2224 -4520
rect 2544 -4840 2584 -4520
rect 2184 -4880 2584 -4840
rect 3196 -4520 3596 -4480
rect 3196 -4840 3236 -4520
rect 3556 -4840 3596 -4520
rect 3196 -4880 3596 -4840
rect 4208 -4520 4608 -4480
rect 4208 -4840 4248 -4520
rect 4568 -4840 4608 -4520
rect 4208 -4880 4608 -4840
rect 5220 -4520 5620 -4480
rect 5220 -4840 5260 -4520
rect 5580 -4840 5620 -4520
rect 5220 -4880 5620 -4840
rect 6232 -4520 6632 -4480
rect 6232 -4840 6272 -4520
rect 6592 -4840 6632 -4520
rect 6232 -4880 6632 -4840
rect 7244 -4520 7644 -4480
rect 7244 -4840 7284 -4520
rect 7604 -4840 7644 -4520
rect 7244 -4880 7644 -4840
rect 8256 -4520 8656 -4480
rect 8256 -4840 8296 -4520
rect 8616 -4840 8656 -4520
rect 8256 -4880 8656 -4840
rect 9268 -4520 9668 -4480
rect 9268 -4840 9308 -4520
rect 9628 -4840 9668 -4520
rect 9268 -4880 9668 -4840
rect 10280 -4520 10680 -4480
rect 10280 -4840 10320 -4520
rect 10640 -4840 10680 -4520
rect 10280 -4880 10680 -4840
rect 11292 -4520 11692 -4480
rect 11292 -4840 11332 -4520
rect 11652 -4840 11692 -4520
rect 11292 -4880 11692 -4840
rect 12304 -4520 12704 -4480
rect 12304 -4840 12344 -4520
rect 12664 -4840 12704 -4520
rect 12304 -4880 12704 -4840
rect 13316 -4520 13716 -4480
rect 13316 -4840 13356 -4520
rect 13676 -4840 13716 -4520
rect 13316 -4880 13716 -4840
rect 14328 -4520 14728 -4480
rect 14328 -4840 14368 -4520
rect 14688 -4840 14728 -4520
rect 14328 -4880 14728 -4840
rect 15340 -4520 15740 -4480
rect 15340 -4840 15380 -4520
rect 15700 -4840 15740 -4520
rect 15340 -4880 15740 -4840
rect 16352 -4520 16752 -4480
rect 16352 -4840 16392 -4520
rect 16712 -4840 16752 -4520
rect 16352 -4880 16752 -4840
rect -17044 -5240 -16644 -5200
rect -17044 -5560 -17004 -5240
rect -16684 -5560 -16644 -5240
rect -17044 -5600 -16644 -5560
rect -16032 -5240 -15632 -5200
rect -16032 -5560 -15992 -5240
rect -15672 -5560 -15632 -5240
rect -16032 -5600 -15632 -5560
rect -15020 -5240 -14620 -5200
rect -15020 -5560 -14980 -5240
rect -14660 -5560 -14620 -5240
rect -15020 -5600 -14620 -5560
rect -14008 -5240 -13608 -5200
rect -14008 -5560 -13968 -5240
rect -13648 -5560 -13608 -5240
rect -14008 -5600 -13608 -5560
rect -12996 -5240 -12596 -5200
rect -12996 -5560 -12956 -5240
rect -12636 -5560 -12596 -5240
rect -12996 -5600 -12596 -5560
rect -11984 -5240 -11584 -5200
rect -11984 -5560 -11944 -5240
rect -11624 -5560 -11584 -5240
rect -11984 -5600 -11584 -5560
rect -10972 -5240 -10572 -5200
rect -10972 -5560 -10932 -5240
rect -10612 -5560 -10572 -5240
rect -10972 -5600 -10572 -5560
rect -9960 -5240 -9560 -5200
rect -9960 -5560 -9920 -5240
rect -9600 -5560 -9560 -5240
rect -9960 -5600 -9560 -5560
rect -8948 -5240 -8548 -5200
rect -8948 -5560 -8908 -5240
rect -8588 -5560 -8548 -5240
rect -8948 -5600 -8548 -5560
rect -7936 -5240 -7536 -5200
rect -7936 -5560 -7896 -5240
rect -7576 -5560 -7536 -5240
rect -7936 -5600 -7536 -5560
rect -6924 -5240 -6524 -5200
rect -6924 -5560 -6884 -5240
rect -6564 -5560 -6524 -5240
rect -6924 -5600 -6524 -5560
rect -5912 -5240 -5512 -5200
rect -5912 -5560 -5872 -5240
rect -5552 -5560 -5512 -5240
rect -5912 -5600 -5512 -5560
rect -4900 -5240 -4500 -5200
rect -4900 -5560 -4860 -5240
rect -4540 -5560 -4500 -5240
rect -4900 -5600 -4500 -5560
rect -3888 -5240 -3488 -5200
rect -3888 -5560 -3848 -5240
rect -3528 -5560 -3488 -5240
rect -3888 -5600 -3488 -5560
rect -2876 -5240 -2476 -5200
rect -2876 -5560 -2836 -5240
rect -2516 -5560 -2476 -5240
rect -2876 -5600 -2476 -5560
rect -1864 -5240 -1464 -5200
rect -1864 -5560 -1824 -5240
rect -1504 -5560 -1464 -5240
rect -1864 -5600 -1464 -5560
rect -852 -5240 -452 -5200
rect -852 -5560 -812 -5240
rect -492 -5560 -452 -5240
rect -852 -5600 -452 -5560
rect 160 -5240 560 -5200
rect 160 -5560 200 -5240
rect 520 -5560 560 -5240
rect 160 -5600 560 -5560
rect 1172 -5240 1572 -5200
rect 1172 -5560 1212 -5240
rect 1532 -5560 1572 -5240
rect 1172 -5600 1572 -5560
rect 2184 -5240 2584 -5200
rect 2184 -5560 2224 -5240
rect 2544 -5560 2584 -5240
rect 2184 -5600 2584 -5560
rect 3196 -5240 3596 -5200
rect 3196 -5560 3236 -5240
rect 3556 -5560 3596 -5240
rect 3196 -5600 3596 -5560
rect 4208 -5240 4608 -5200
rect 4208 -5560 4248 -5240
rect 4568 -5560 4608 -5240
rect 4208 -5600 4608 -5560
rect 5220 -5240 5620 -5200
rect 5220 -5560 5260 -5240
rect 5580 -5560 5620 -5240
rect 5220 -5600 5620 -5560
rect 6232 -5240 6632 -5200
rect 6232 -5560 6272 -5240
rect 6592 -5560 6632 -5240
rect 6232 -5600 6632 -5560
rect 7244 -5240 7644 -5200
rect 7244 -5560 7284 -5240
rect 7604 -5560 7644 -5240
rect 7244 -5600 7644 -5560
rect 8256 -5240 8656 -5200
rect 8256 -5560 8296 -5240
rect 8616 -5560 8656 -5240
rect 8256 -5600 8656 -5560
rect 9268 -5240 9668 -5200
rect 9268 -5560 9308 -5240
rect 9628 -5560 9668 -5240
rect 9268 -5600 9668 -5560
rect 10280 -5240 10680 -5200
rect 10280 -5560 10320 -5240
rect 10640 -5560 10680 -5240
rect 10280 -5600 10680 -5560
rect 11292 -5240 11692 -5200
rect 11292 -5560 11332 -5240
rect 11652 -5560 11692 -5240
rect 11292 -5600 11692 -5560
rect 12304 -5240 12704 -5200
rect 12304 -5560 12344 -5240
rect 12664 -5560 12704 -5240
rect 12304 -5600 12704 -5560
rect 13316 -5240 13716 -5200
rect 13316 -5560 13356 -5240
rect 13676 -5560 13716 -5240
rect 13316 -5600 13716 -5560
rect 14328 -5240 14728 -5200
rect 14328 -5560 14368 -5240
rect 14688 -5560 14728 -5240
rect 14328 -5600 14728 -5560
rect 15340 -5240 15740 -5200
rect 15340 -5560 15380 -5240
rect 15700 -5560 15740 -5240
rect 15340 -5600 15740 -5560
rect 16352 -5240 16752 -5200
rect 16352 -5560 16392 -5240
rect 16712 -5560 16752 -5240
rect 16352 -5600 16752 -5560
rect -17044 -5960 -16644 -5920
rect -17044 -6280 -17004 -5960
rect -16684 -6280 -16644 -5960
rect -17044 -6320 -16644 -6280
rect -16032 -5960 -15632 -5920
rect -16032 -6280 -15992 -5960
rect -15672 -6280 -15632 -5960
rect -16032 -6320 -15632 -6280
rect -15020 -5960 -14620 -5920
rect -15020 -6280 -14980 -5960
rect -14660 -6280 -14620 -5960
rect -15020 -6320 -14620 -6280
rect -14008 -5960 -13608 -5920
rect -14008 -6280 -13968 -5960
rect -13648 -6280 -13608 -5960
rect -14008 -6320 -13608 -6280
rect -12996 -5960 -12596 -5920
rect -12996 -6280 -12956 -5960
rect -12636 -6280 -12596 -5960
rect -12996 -6320 -12596 -6280
rect -11984 -5960 -11584 -5920
rect -11984 -6280 -11944 -5960
rect -11624 -6280 -11584 -5960
rect -11984 -6320 -11584 -6280
rect -10972 -5960 -10572 -5920
rect -10972 -6280 -10932 -5960
rect -10612 -6280 -10572 -5960
rect -10972 -6320 -10572 -6280
rect -9960 -5960 -9560 -5920
rect -9960 -6280 -9920 -5960
rect -9600 -6280 -9560 -5960
rect -9960 -6320 -9560 -6280
rect -8948 -5960 -8548 -5920
rect -8948 -6280 -8908 -5960
rect -8588 -6280 -8548 -5960
rect -8948 -6320 -8548 -6280
rect -7936 -5960 -7536 -5920
rect -7936 -6280 -7896 -5960
rect -7576 -6280 -7536 -5960
rect -7936 -6320 -7536 -6280
rect -6924 -5960 -6524 -5920
rect -6924 -6280 -6884 -5960
rect -6564 -6280 -6524 -5960
rect -6924 -6320 -6524 -6280
rect -5912 -5960 -5512 -5920
rect -5912 -6280 -5872 -5960
rect -5552 -6280 -5512 -5960
rect -5912 -6320 -5512 -6280
rect -4900 -5960 -4500 -5920
rect -4900 -6280 -4860 -5960
rect -4540 -6280 -4500 -5960
rect -4900 -6320 -4500 -6280
rect -3888 -5960 -3488 -5920
rect -3888 -6280 -3848 -5960
rect -3528 -6280 -3488 -5960
rect -3888 -6320 -3488 -6280
rect -2876 -5960 -2476 -5920
rect -2876 -6280 -2836 -5960
rect -2516 -6280 -2476 -5960
rect -2876 -6320 -2476 -6280
rect -1864 -5960 -1464 -5920
rect -1864 -6280 -1824 -5960
rect -1504 -6280 -1464 -5960
rect -1864 -6320 -1464 -6280
rect -852 -5960 -452 -5920
rect -852 -6280 -812 -5960
rect -492 -6280 -452 -5960
rect -852 -6320 -452 -6280
rect 160 -5960 560 -5920
rect 160 -6280 200 -5960
rect 520 -6280 560 -5960
rect 160 -6320 560 -6280
rect 1172 -5960 1572 -5920
rect 1172 -6280 1212 -5960
rect 1532 -6280 1572 -5960
rect 1172 -6320 1572 -6280
rect 2184 -5960 2584 -5920
rect 2184 -6280 2224 -5960
rect 2544 -6280 2584 -5960
rect 2184 -6320 2584 -6280
rect 3196 -5960 3596 -5920
rect 3196 -6280 3236 -5960
rect 3556 -6280 3596 -5960
rect 3196 -6320 3596 -6280
rect 4208 -5960 4608 -5920
rect 4208 -6280 4248 -5960
rect 4568 -6280 4608 -5960
rect 4208 -6320 4608 -6280
rect 5220 -5960 5620 -5920
rect 5220 -6280 5260 -5960
rect 5580 -6280 5620 -5960
rect 5220 -6320 5620 -6280
rect 6232 -5960 6632 -5920
rect 6232 -6280 6272 -5960
rect 6592 -6280 6632 -5960
rect 6232 -6320 6632 -6280
rect 7244 -5960 7644 -5920
rect 7244 -6280 7284 -5960
rect 7604 -6280 7644 -5960
rect 7244 -6320 7644 -6280
rect 8256 -5960 8656 -5920
rect 8256 -6280 8296 -5960
rect 8616 -6280 8656 -5960
rect 8256 -6320 8656 -6280
rect 9268 -5960 9668 -5920
rect 9268 -6280 9308 -5960
rect 9628 -6280 9668 -5960
rect 9268 -6320 9668 -6280
rect 10280 -5960 10680 -5920
rect 10280 -6280 10320 -5960
rect 10640 -6280 10680 -5960
rect 10280 -6320 10680 -6280
rect 11292 -5960 11692 -5920
rect 11292 -6280 11332 -5960
rect 11652 -6280 11692 -5960
rect 11292 -6320 11692 -6280
rect 12304 -5960 12704 -5920
rect 12304 -6280 12344 -5960
rect 12664 -6280 12704 -5960
rect 12304 -6320 12704 -6280
rect 13316 -5960 13716 -5920
rect 13316 -6280 13356 -5960
rect 13676 -6280 13716 -5960
rect 13316 -6320 13716 -6280
rect 14328 -5960 14728 -5920
rect 14328 -6280 14368 -5960
rect 14688 -6280 14728 -5960
rect 14328 -6320 14728 -6280
rect 15340 -5960 15740 -5920
rect 15340 -6280 15380 -5960
rect 15700 -6280 15740 -5960
rect 15340 -6320 15740 -6280
rect 16352 -5960 16752 -5920
rect 16352 -6280 16392 -5960
rect 16712 -6280 16752 -5960
rect 16352 -6320 16752 -6280
rect -17044 -6680 -16644 -6640
rect -17044 -7000 -17004 -6680
rect -16684 -7000 -16644 -6680
rect -17044 -7040 -16644 -7000
rect -16032 -6680 -15632 -6640
rect -16032 -7000 -15992 -6680
rect -15672 -7000 -15632 -6680
rect -16032 -7040 -15632 -7000
rect -15020 -6680 -14620 -6640
rect -15020 -7000 -14980 -6680
rect -14660 -7000 -14620 -6680
rect -15020 -7040 -14620 -7000
rect -14008 -6680 -13608 -6640
rect -14008 -7000 -13968 -6680
rect -13648 -7000 -13608 -6680
rect -14008 -7040 -13608 -7000
rect -12996 -6680 -12596 -6640
rect -12996 -7000 -12956 -6680
rect -12636 -7000 -12596 -6680
rect -12996 -7040 -12596 -7000
rect -11984 -6680 -11584 -6640
rect -11984 -7000 -11944 -6680
rect -11624 -7000 -11584 -6680
rect -11984 -7040 -11584 -7000
rect -10972 -6680 -10572 -6640
rect -10972 -7000 -10932 -6680
rect -10612 -7000 -10572 -6680
rect -10972 -7040 -10572 -7000
rect -9960 -6680 -9560 -6640
rect -9960 -7000 -9920 -6680
rect -9600 -7000 -9560 -6680
rect -9960 -7040 -9560 -7000
rect -8948 -6680 -8548 -6640
rect -8948 -7000 -8908 -6680
rect -8588 -7000 -8548 -6680
rect -8948 -7040 -8548 -7000
rect -7936 -6680 -7536 -6640
rect -7936 -7000 -7896 -6680
rect -7576 -7000 -7536 -6680
rect -7936 -7040 -7536 -7000
rect -6924 -6680 -6524 -6640
rect -6924 -7000 -6884 -6680
rect -6564 -7000 -6524 -6680
rect -6924 -7040 -6524 -7000
rect -5912 -6680 -5512 -6640
rect -5912 -7000 -5872 -6680
rect -5552 -7000 -5512 -6680
rect -5912 -7040 -5512 -7000
rect -4900 -6680 -4500 -6640
rect -4900 -7000 -4860 -6680
rect -4540 -7000 -4500 -6680
rect -4900 -7040 -4500 -7000
rect -3888 -6680 -3488 -6640
rect -3888 -7000 -3848 -6680
rect -3528 -7000 -3488 -6680
rect -3888 -7040 -3488 -7000
rect -2876 -6680 -2476 -6640
rect -2876 -7000 -2836 -6680
rect -2516 -7000 -2476 -6680
rect -2876 -7040 -2476 -7000
rect -1864 -6680 -1464 -6640
rect -1864 -7000 -1824 -6680
rect -1504 -7000 -1464 -6680
rect -1864 -7040 -1464 -7000
rect -852 -6680 -452 -6640
rect -852 -7000 -812 -6680
rect -492 -7000 -452 -6680
rect -852 -7040 -452 -7000
rect 160 -6680 560 -6640
rect 160 -7000 200 -6680
rect 520 -7000 560 -6680
rect 160 -7040 560 -7000
rect 1172 -6680 1572 -6640
rect 1172 -7000 1212 -6680
rect 1532 -7000 1572 -6680
rect 1172 -7040 1572 -7000
rect 2184 -6680 2584 -6640
rect 2184 -7000 2224 -6680
rect 2544 -7000 2584 -6680
rect 2184 -7040 2584 -7000
rect 3196 -6680 3596 -6640
rect 3196 -7000 3236 -6680
rect 3556 -7000 3596 -6680
rect 3196 -7040 3596 -7000
rect 4208 -6680 4608 -6640
rect 4208 -7000 4248 -6680
rect 4568 -7000 4608 -6680
rect 4208 -7040 4608 -7000
rect 5220 -6680 5620 -6640
rect 5220 -7000 5260 -6680
rect 5580 -7000 5620 -6680
rect 5220 -7040 5620 -7000
rect 6232 -6680 6632 -6640
rect 6232 -7000 6272 -6680
rect 6592 -7000 6632 -6680
rect 6232 -7040 6632 -7000
rect 7244 -6680 7644 -6640
rect 7244 -7000 7284 -6680
rect 7604 -7000 7644 -6680
rect 7244 -7040 7644 -7000
rect 8256 -6680 8656 -6640
rect 8256 -7000 8296 -6680
rect 8616 -7000 8656 -6680
rect 8256 -7040 8656 -7000
rect 9268 -6680 9668 -6640
rect 9268 -7000 9308 -6680
rect 9628 -7000 9668 -6680
rect 9268 -7040 9668 -7000
rect 10280 -6680 10680 -6640
rect 10280 -7000 10320 -6680
rect 10640 -7000 10680 -6680
rect 10280 -7040 10680 -7000
rect 11292 -6680 11692 -6640
rect 11292 -7000 11332 -6680
rect 11652 -7000 11692 -6680
rect 11292 -7040 11692 -7000
rect 12304 -6680 12704 -6640
rect 12304 -7000 12344 -6680
rect 12664 -7000 12704 -6680
rect 12304 -7040 12704 -7000
rect 13316 -6680 13716 -6640
rect 13316 -7000 13356 -6680
rect 13676 -7000 13716 -6680
rect 13316 -7040 13716 -7000
rect 14328 -6680 14728 -6640
rect 14328 -7000 14368 -6680
rect 14688 -7000 14728 -6680
rect 14328 -7040 14728 -7000
rect 15340 -6680 15740 -6640
rect 15340 -7000 15380 -6680
rect 15700 -7000 15740 -6680
rect 15340 -7040 15740 -7000
rect 16352 -6680 16752 -6640
rect 16352 -7000 16392 -6680
rect 16712 -7000 16752 -6680
rect 16352 -7040 16752 -7000
rect -17044 -7400 -16644 -7360
rect -17044 -7720 -17004 -7400
rect -16684 -7720 -16644 -7400
rect -17044 -7760 -16644 -7720
rect -16032 -7400 -15632 -7360
rect -16032 -7720 -15992 -7400
rect -15672 -7720 -15632 -7400
rect -16032 -7760 -15632 -7720
rect -15020 -7400 -14620 -7360
rect -15020 -7720 -14980 -7400
rect -14660 -7720 -14620 -7400
rect -15020 -7760 -14620 -7720
rect -14008 -7400 -13608 -7360
rect -14008 -7720 -13968 -7400
rect -13648 -7720 -13608 -7400
rect -14008 -7760 -13608 -7720
rect -12996 -7400 -12596 -7360
rect -12996 -7720 -12956 -7400
rect -12636 -7720 -12596 -7400
rect -12996 -7760 -12596 -7720
rect -11984 -7400 -11584 -7360
rect -11984 -7720 -11944 -7400
rect -11624 -7720 -11584 -7400
rect -11984 -7760 -11584 -7720
rect -10972 -7400 -10572 -7360
rect -10972 -7720 -10932 -7400
rect -10612 -7720 -10572 -7400
rect -10972 -7760 -10572 -7720
rect -9960 -7400 -9560 -7360
rect -9960 -7720 -9920 -7400
rect -9600 -7720 -9560 -7400
rect -9960 -7760 -9560 -7720
rect -8948 -7400 -8548 -7360
rect -8948 -7720 -8908 -7400
rect -8588 -7720 -8548 -7400
rect -8948 -7760 -8548 -7720
rect -7936 -7400 -7536 -7360
rect -7936 -7720 -7896 -7400
rect -7576 -7720 -7536 -7400
rect -7936 -7760 -7536 -7720
rect -6924 -7400 -6524 -7360
rect -6924 -7720 -6884 -7400
rect -6564 -7720 -6524 -7400
rect -6924 -7760 -6524 -7720
rect -5912 -7400 -5512 -7360
rect -5912 -7720 -5872 -7400
rect -5552 -7720 -5512 -7400
rect -5912 -7760 -5512 -7720
rect -4900 -7400 -4500 -7360
rect -4900 -7720 -4860 -7400
rect -4540 -7720 -4500 -7400
rect -4900 -7760 -4500 -7720
rect -3888 -7400 -3488 -7360
rect -3888 -7720 -3848 -7400
rect -3528 -7720 -3488 -7400
rect -3888 -7760 -3488 -7720
rect -2876 -7400 -2476 -7360
rect -2876 -7720 -2836 -7400
rect -2516 -7720 -2476 -7400
rect -2876 -7760 -2476 -7720
rect -1864 -7400 -1464 -7360
rect -1864 -7720 -1824 -7400
rect -1504 -7720 -1464 -7400
rect -1864 -7760 -1464 -7720
rect -852 -7400 -452 -7360
rect -852 -7720 -812 -7400
rect -492 -7720 -452 -7400
rect -852 -7760 -452 -7720
rect 160 -7400 560 -7360
rect 160 -7720 200 -7400
rect 520 -7720 560 -7400
rect 160 -7760 560 -7720
rect 1172 -7400 1572 -7360
rect 1172 -7720 1212 -7400
rect 1532 -7720 1572 -7400
rect 1172 -7760 1572 -7720
rect 2184 -7400 2584 -7360
rect 2184 -7720 2224 -7400
rect 2544 -7720 2584 -7400
rect 2184 -7760 2584 -7720
rect 3196 -7400 3596 -7360
rect 3196 -7720 3236 -7400
rect 3556 -7720 3596 -7400
rect 3196 -7760 3596 -7720
rect 4208 -7400 4608 -7360
rect 4208 -7720 4248 -7400
rect 4568 -7720 4608 -7400
rect 4208 -7760 4608 -7720
rect 5220 -7400 5620 -7360
rect 5220 -7720 5260 -7400
rect 5580 -7720 5620 -7400
rect 5220 -7760 5620 -7720
rect 6232 -7400 6632 -7360
rect 6232 -7720 6272 -7400
rect 6592 -7720 6632 -7400
rect 6232 -7760 6632 -7720
rect 7244 -7400 7644 -7360
rect 7244 -7720 7284 -7400
rect 7604 -7720 7644 -7400
rect 7244 -7760 7644 -7720
rect 8256 -7400 8656 -7360
rect 8256 -7720 8296 -7400
rect 8616 -7720 8656 -7400
rect 8256 -7760 8656 -7720
rect 9268 -7400 9668 -7360
rect 9268 -7720 9308 -7400
rect 9628 -7720 9668 -7400
rect 9268 -7760 9668 -7720
rect 10280 -7400 10680 -7360
rect 10280 -7720 10320 -7400
rect 10640 -7720 10680 -7400
rect 10280 -7760 10680 -7720
rect 11292 -7400 11692 -7360
rect 11292 -7720 11332 -7400
rect 11652 -7720 11692 -7400
rect 11292 -7760 11692 -7720
rect 12304 -7400 12704 -7360
rect 12304 -7720 12344 -7400
rect 12664 -7720 12704 -7400
rect 12304 -7760 12704 -7720
rect 13316 -7400 13716 -7360
rect 13316 -7720 13356 -7400
rect 13676 -7720 13716 -7400
rect 13316 -7760 13716 -7720
rect 14328 -7400 14728 -7360
rect 14328 -7720 14368 -7400
rect 14688 -7720 14728 -7400
rect 14328 -7760 14728 -7720
rect 15340 -7400 15740 -7360
rect 15340 -7720 15380 -7400
rect 15700 -7720 15740 -7400
rect 15340 -7760 15740 -7720
rect 16352 -7400 16752 -7360
rect 16352 -7720 16392 -7400
rect 16712 -7720 16752 -7400
rect 16352 -7760 16752 -7720
rect -17044 -8120 -16644 -8080
rect -17044 -8440 -17004 -8120
rect -16684 -8440 -16644 -8120
rect -17044 -8480 -16644 -8440
rect -16032 -8120 -15632 -8080
rect -16032 -8440 -15992 -8120
rect -15672 -8440 -15632 -8120
rect -16032 -8480 -15632 -8440
rect -15020 -8120 -14620 -8080
rect -15020 -8440 -14980 -8120
rect -14660 -8440 -14620 -8120
rect -15020 -8480 -14620 -8440
rect -14008 -8120 -13608 -8080
rect -14008 -8440 -13968 -8120
rect -13648 -8440 -13608 -8120
rect -14008 -8480 -13608 -8440
rect -12996 -8120 -12596 -8080
rect -12996 -8440 -12956 -8120
rect -12636 -8440 -12596 -8120
rect -12996 -8480 -12596 -8440
rect -11984 -8120 -11584 -8080
rect -11984 -8440 -11944 -8120
rect -11624 -8440 -11584 -8120
rect -11984 -8480 -11584 -8440
rect -10972 -8120 -10572 -8080
rect -10972 -8440 -10932 -8120
rect -10612 -8440 -10572 -8120
rect -10972 -8480 -10572 -8440
rect -9960 -8120 -9560 -8080
rect -9960 -8440 -9920 -8120
rect -9600 -8440 -9560 -8120
rect -9960 -8480 -9560 -8440
rect -8948 -8120 -8548 -8080
rect -8948 -8440 -8908 -8120
rect -8588 -8440 -8548 -8120
rect -8948 -8480 -8548 -8440
rect -7936 -8120 -7536 -8080
rect -7936 -8440 -7896 -8120
rect -7576 -8440 -7536 -8120
rect -7936 -8480 -7536 -8440
rect -6924 -8120 -6524 -8080
rect -6924 -8440 -6884 -8120
rect -6564 -8440 -6524 -8120
rect -6924 -8480 -6524 -8440
rect -5912 -8120 -5512 -8080
rect -5912 -8440 -5872 -8120
rect -5552 -8440 -5512 -8120
rect -5912 -8480 -5512 -8440
rect -4900 -8120 -4500 -8080
rect -4900 -8440 -4860 -8120
rect -4540 -8440 -4500 -8120
rect -4900 -8480 -4500 -8440
rect -3888 -8120 -3488 -8080
rect -3888 -8440 -3848 -8120
rect -3528 -8440 -3488 -8120
rect -3888 -8480 -3488 -8440
rect -2876 -8120 -2476 -8080
rect -2876 -8440 -2836 -8120
rect -2516 -8440 -2476 -8120
rect -2876 -8480 -2476 -8440
rect -1864 -8120 -1464 -8080
rect -1864 -8440 -1824 -8120
rect -1504 -8440 -1464 -8120
rect -1864 -8480 -1464 -8440
rect -852 -8120 -452 -8080
rect -852 -8440 -812 -8120
rect -492 -8440 -452 -8120
rect -852 -8480 -452 -8440
rect 160 -8120 560 -8080
rect 160 -8440 200 -8120
rect 520 -8440 560 -8120
rect 160 -8480 560 -8440
rect 1172 -8120 1572 -8080
rect 1172 -8440 1212 -8120
rect 1532 -8440 1572 -8120
rect 1172 -8480 1572 -8440
rect 2184 -8120 2584 -8080
rect 2184 -8440 2224 -8120
rect 2544 -8440 2584 -8120
rect 2184 -8480 2584 -8440
rect 3196 -8120 3596 -8080
rect 3196 -8440 3236 -8120
rect 3556 -8440 3596 -8120
rect 3196 -8480 3596 -8440
rect 4208 -8120 4608 -8080
rect 4208 -8440 4248 -8120
rect 4568 -8440 4608 -8120
rect 4208 -8480 4608 -8440
rect 5220 -8120 5620 -8080
rect 5220 -8440 5260 -8120
rect 5580 -8440 5620 -8120
rect 5220 -8480 5620 -8440
rect 6232 -8120 6632 -8080
rect 6232 -8440 6272 -8120
rect 6592 -8440 6632 -8120
rect 6232 -8480 6632 -8440
rect 7244 -8120 7644 -8080
rect 7244 -8440 7284 -8120
rect 7604 -8440 7644 -8120
rect 7244 -8480 7644 -8440
rect 8256 -8120 8656 -8080
rect 8256 -8440 8296 -8120
rect 8616 -8440 8656 -8120
rect 8256 -8480 8656 -8440
rect 9268 -8120 9668 -8080
rect 9268 -8440 9308 -8120
rect 9628 -8440 9668 -8120
rect 9268 -8480 9668 -8440
rect 10280 -8120 10680 -8080
rect 10280 -8440 10320 -8120
rect 10640 -8440 10680 -8120
rect 10280 -8480 10680 -8440
rect 11292 -8120 11692 -8080
rect 11292 -8440 11332 -8120
rect 11652 -8440 11692 -8120
rect 11292 -8480 11692 -8440
rect 12304 -8120 12704 -8080
rect 12304 -8440 12344 -8120
rect 12664 -8440 12704 -8120
rect 12304 -8480 12704 -8440
rect 13316 -8120 13716 -8080
rect 13316 -8440 13356 -8120
rect 13676 -8440 13716 -8120
rect 13316 -8480 13716 -8440
rect 14328 -8120 14728 -8080
rect 14328 -8440 14368 -8120
rect 14688 -8440 14728 -8120
rect 14328 -8480 14728 -8440
rect 15340 -8120 15740 -8080
rect 15340 -8440 15380 -8120
rect 15700 -8440 15740 -8120
rect 15340 -8480 15740 -8440
rect 16352 -8120 16752 -8080
rect 16352 -8440 16392 -8120
rect 16712 -8440 16752 -8120
rect 16352 -8480 16752 -8440
rect -17044 -8840 -16644 -8800
rect -17044 -9160 -17004 -8840
rect -16684 -9160 -16644 -8840
rect -17044 -9200 -16644 -9160
rect -16032 -8840 -15632 -8800
rect -16032 -9160 -15992 -8840
rect -15672 -9160 -15632 -8840
rect -16032 -9200 -15632 -9160
rect -15020 -8840 -14620 -8800
rect -15020 -9160 -14980 -8840
rect -14660 -9160 -14620 -8840
rect -15020 -9200 -14620 -9160
rect -14008 -8840 -13608 -8800
rect -14008 -9160 -13968 -8840
rect -13648 -9160 -13608 -8840
rect -14008 -9200 -13608 -9160
rect -12996 -8840 -12596 -8800
rect -12996 -9160 -12956 -8840
rect -12636 -9160 -12596 -8840
rect -12996 -9200 -12596 -9160
rect -11984 -8840 -11584 -8800
rect -11984 -9160 -11944 -8840
rect -11624 -9160 -11584 -8840
rect -11984 -9200 -11584 -9160
rect -10972 -8840 -10572 -8800
rect -10972 -9160 -10932 -8840
rect -10612 -9160 -10572 -8840
rect -10972 -9200 -10572 -9160
rect -9960 -8840 -9560 -8800
rect -9960 -9160 -9920 -8840
rect -9600 -9160 -9560 -8840
rect -9960 -9200 -9560 -9160
rect -8948 -8840 -8548 -8800
rect -8948 -9160 -8908 -8840
rect -8588 -9160 -8548 -8840
rect -8948 -9200 -8548 -9160
rect -7936 -8840 -7536 -8800
rect -7936 -9160 -7896 -8840
rect -7576 -9160 -7536 -8840
rect -7936 -9200 -7536 -9160
rect -6924 -8840 -6524 -8800
rect -6924 -9160 -6884 -8840
rect -6564 -9160 -6524 -8840
rect -6924 -9200 -6524 -9160
rect -5912 -8840 -5512 -8800
rect -5912 -9160 -5872 -8840
rect -5552 -9160 -5512 -8840
rect -5912 -9200 -5512 -9160
rect -4900 -8840 -4500 -8800
rect -4900 -9160 -4860 -8840
rect -4540 -9160 -4500 -8840
rect -4900 -9200 -4500 -9160
rect -3888 -8840 -3488 -8800
rect -3888 -9160 -3848 -8840
rect -3528 -9160 -3488 -8840
rect -3888 -9200 -3488 -9160
rect -2876 -8840 -2476 -8800
rect -2876 -9160 -2836 -8840
rect -2516 -9160 -2476 -8840
rect -2876 -9200 -2476 -9160
rect -1864 -8840 -1464 -8800
rect -1864 -9160 -1824 -8840
rect -1504 -9160 -1464 -8840
rect -1864 -9200 -1464 -9160
rect -852 -8840 -452 -8800
rect -852 -9160 -812 -8840
rect -492 -9160 -452 -8840
rect -852 -9200 -452 -9160
rect 160 -8840 560 -8800
rect 160 -9160 200 -8840
rect 520 -9160 560 -8840
rect 160 -9200 560 -9160
rect 1172 -8840 1572 -8800
rect 1172 -9160 1212 -8840
rect 1532 -9160 1572 -8840
rect 1172 -9200 1572 -9160
rect 2184 -8840 2584 -8800
rect 2184 -9160 2224 -8840
rect 2544 -9160 2584 -8840
rect 2184 -9200 2584 -9160
rect 3196 -8840 3596 -8800
rect 3196 -9160 3236 -8840
rect 3556 -9160 3596 -8840
rect 3196 -9200 3596 -9160
rect 4208 -8840 4608 -8800
rect 4208 -9160 4248 -8840
rect 4568 -9160 4608 -8840
rect 4208 -9200 4608 -9160
rect 5220 -8840 5620 -8800
rect 5220 -9160 5260 -8840
rect 5580 -9160 5620 -8840
rect 5220 -9200 5620 -9160
rect 6232 -8840 6632 -8800
rect 6232 -9160 6272 -8840
rect 6592 -9160 6632 -8840
rect 6232 -9200 6632 -9160
rect 7244 -8840 7644 -8800
rect 7244 -9160 7284 -8840
rect 7604 -9160 7644 -8840
rect 7244 -9200 7644 -9160
rect 8256 -8840 8656 -8800
rect 8256 -9160 8296 -8840
rect 8616 -9160 8656 -8840
rect 8256 -9200 8656 -9160
rect 9268 -8840 9668 -8800
rect 9268 -9160 9308 -8840
rect 9628 -9160 9668 -8840
rect 9268 -9200 9668 -9160
rect 10280 -8840 10680 -8800
rect 10280 -9160 10320 -8840
rect 10640 -9160 10680 -8840
rect 10280 -9200 10680 -9160
rect 11292 -8840 11692 -8800
rect 11292 -9160 11332 -8840
rect 11652 -9160 11692 -8840
rect 11292 -9200 11692 -9160
rect 12304 -8840 12704 -8800
rect 12304 -9160 12344 -8840
rect 12664 -9160 12704 -8840
rect 12304 -9200 12704 -9160
rect 13316 -8840 13716 -8800
rect 13316 -9160 13356 -8840
rect 13676 -9160 13716 -8840
rect 13316 -9200 13716 -9160
rect 14328 -8840 14728 -8800
rect 14328 -9160 14368 -8840
rect 14688 -9160 14728 -8840
rect 14328 -9200 14728 -9160
rect 15340 -8840 15740 -8800
rect 15340 -9160 15380 -8840
rect 15700 -9160 15740 -8840
rect 15340 -9200 15740 -9160
rect 16352 -8840 16752 -8800
rect 16352 -9160 16392 -8840
rect 16712 -9160 16752 -8840
rect 16352 -9200 16752 -9160
rect -17044 -9560 -16644 -9520
rect -17044 -9880 -17004 -9560
rect -16684 -9880 -16644 -9560
rect -17044 -9920 -16644 -9880
rect -16032 -9560 -15632 -9520
rect -16032 -9880 -15992 -9560
rect -15672 -9880 -15632 -9560
rect -16032 -9920 -15632 -9880
rect -15020 -9560 -14620 -9520
rect -15020 -9880 -14980 -9560
rect -14660 -9880 -14620 -9560
rect -15020 -9920 -14620 -9880
rect -14008 -9560 -13608 -9520
rect -14008 -9880 -13968 -9560
rect -13648 -9880 -13608 -9560
rect -14008 -9920 -13608 -9880
rect -12996 -9560 -12596 -9520
rect -12996 -9880 -12956 -9560
rect -12636 -9880 -12596 -9560
rect -12996 -9920 -12596 -9880
rect -11984 -9560 -11584 -9520
rect -11984 -9880 -11944 -9560
rect -11624 -9880 -11584 -9560
rect -11984 -9920 -11584 -9880
rect -10972 -9560 -10572 -9520
rect -10972 -9880 -10932 -9560
rect -10612 -9880 -10572 -9560
rect -10972 -9920 -10572 -9880
rect -9960 -9560 -9560 -9520
rect -9960 -9880 -9920 -9560
rect -9600 -9880 -9560 -9560
rect -9960 -9920 -9560 -9880
rect -8948 -9560 -8548 -9520
rect -8948 -9880 -8908 -9560
rect -8588 -9880 -8548 -9560
rect -8948 -9920 -8548 -9880
rect -7936 -9560 -7536 -9520
rect -7936 -9880 -7896 -9560
rect -7576 -9880 -7536 -9560
rect -7936 -9920 -7536 -9880
rect -6924 -9560 -6524 -9520
rect -6924 -9880 -6884 -9560
rect -6564 -9880 -6524 -9560
rect -6924 -9920 -6524 -9880
rect -5912 -9560 -5512 -9520
rect -5912 -9880 -5872 -9560
rect -5552 -9880 -5512 -9560
rect -5912 -9920 -5512 -9880
rect -4900 -9560 -4500 -9520
rect -4900 -9880 -4860 -9560
rect -4540 -9880 -4500 -9560
rect -4900 -9920 -4500 -9880
rect -3888 -9560 -3488 -9520
rect -3888 -9880 -3848 -9560
rect -3528 -9880 -3488 -9560
rect -3888 -9920 -3488 -9880
rect -2876 -9560 -2476 -9520
rect -2876 -9880 -2836 -9560
rect -2516 -9880 -2476 -9560
rect -2876 -9920 -2476 -9880
rect -1864 -9560 -1464 -9520
rect -1864 -9880 -1824 -9560
rect -1504 -9880 -1464 -9560
rect -1864 -9920 -1464 -9880
rect -852 -9560 -452 -9520
rect -852 -9880 -812 -9560
rect -492 -9880 -452 -9560
rect -852 -9920 -452 -9880
rect 160 -9560 560 -9520
rect 160 -9880 200 -9560
rect 520 -9880 560 -9560
rect 160 -9920 560 -9880
rect 1172 -9560 1572 -9520
rect 1172 -9880 1212 -9560
rect 1532 -9880 1572 -9560
rect 1172 -9920 1572 -9880
rect 2184 -9560 2584 -9520
rect 2184 -9880 2224 -9560
rect 2544 -9880 2584 -9560
rect 2184 -9920 2584 -9880
rect 3196 -9560 3596 -9520
rect 3196 -9880 3236 -9560
rect 3556 -9880 3596 -9560
rect 3196 -9920 3596 -9880
rect 4208 -9560 4608 -9520
rect 4208 -9880 4248 -9560
rect 4568 -9880 4608 -9560
rect 4208 -9920 4608 -9880
rect 5220 -9560 5620 -9520
rect 5220 -9880 5260 -9560
rect 5580 -9880 5620 -9560
rect 5220 -9920 5620 -9880
rect 6232 -9560 6632 -9520
rect 6232 -9880 6272 -9560
rect 6592 -9880 6632 -9560
rect 6232 -9920 6632 -9880
rect 7244 -9560 7644 -9520
rect 7244 -9880 7284 -9560
rect 7604 -9880 7644 -9560
rect 7244 -9920 7644 -9880
rect 8256 -9560 8656 -9520
rect 8256 -9880 8296 -9560
rect 8616 -9880 8656 -9560
rect 8256 -9920 8656 -9880
rect 9268 -9560 9668 -9520
rect 9268 -9880 9308 -9560
rect 9628 -9880 9668 -9560
rect 9268 -9920 9668 -9880
rect 10280 -9560 10680 -9520
rect 10280 -9880 10320 -9560
rect 10640 -9880 10680 -9560
rect 10280 -9920 10680 -9880
rect 11292 -9560 11692 -9520
rect 11292 -9880 11332 -9560
rect 11652 -9880 11692 -9560
rect 11292 -9920 11692 -9880
rect 12304 -9560 12704 -9520
rect 12304 -9880 12344 -9560
rect 12664 -9880 12704 -9560
rect 12304 -9920 12704 -9880
rect 13316 -9560 13716 -9520
rect 13316 -9880 13356 -9560
rect 13676 -9880 13716 -9560
rect 13316 -9920 13716 -9880
rect 14328 -9560 14728 -9520
rect 14328 -9880 14368 -9560
rect 14688 -9880 14728 -9560
rect 14328 -9920 14728 -9880
rect 15340 -9560 15740 -9520
rect 15340 -9880 15380 -9560
rect 15700 -9880 15740 -9560
rect 15340 -9920 15740 -9880
rect 16352 -9560 16752 -9520
rect 16352 -9880 16392 -9560
rect 16712 -9880 16752 -9560
rect 16352 -9920 16752 -9880
rect -17044 -10280 -16644 -10240
rect -17044 -10600 -17004 -10280
rect -16684 -10600 -16644 -10280
rect -17044 -10640 -16644 -10600
rect -16032 -10280 -15632 -10240
rect -16032 -10600 -15992 -10280
rect -15672 -10600 -15632 -10280
rect -16032 -10640 -15632 -10600
rect -15020 -10280 -14620 -10240
rect -15020 -10600 -14980 -10280
rect -14660 -10600 -14620 -10280
rect -15020 -10640 -14620 -10600
rect -14008 -10280 -13608 -10240
rect -14008 -10600 -13968 -10280
rect -13648 -10600 -13608 -10280
rect -14008 -10640 -13608 -10600
rect -12996 -10280 -12596 -10240
rect -12996 -10600 -12956 -10280
rect -12636 -10600 -12596 -10280
rect -12996 -10640 -12596 -10600
rect -11984 -10280 -11584 -10240
rect -11984 -10600 -11944 -10280
rect -11624 -10600 -11584 -10280
rect -11984 -10640 -11584 -10600
rect -10972 -10280 -10572 -10240
rect -10972 -10600 -10932 -10280
rect -10612 -10600 -10572 -10280
rect -10972 -10640 -10572 -10600
rect -9960 -10280 -9560 -10240
rect -9960 -10600 -9920 -10280
rect -9600 -10600 -9560 -10280
rect -9960 -10640 -9560 -10600
rect -8948 -10280 -8548 -10240
rect -8948 -10600 -8908 -10280
rect -8588 -10600 -8548 -10280
rect -8948 -10640 -8548 -10600
rect -7936 -10280 -7536 -10240
rect -7936 -10600 -7896 -10280
rect -7576 -10600 -7536 -10280
rect -7936 -10640 -7536 -10600
rect -6924 -10280 -6524 -10240
rect -6924 -10600 -6884 -10280
rect -6564 -10600 -6524 -10280
rect -6924 -10640 -6524 -10600
rect -5912 -10280 -5512 -10240
rect -5912 -10600 -5872 -10280
rect -5552 -10600 -5512 -10280
rect -5912 -10640 -5512 -10600
rect -4900 -10280 -4500 -10240
rect -4900 -10600 -4860 -10280
rect -4540 -10600 -4500 -10280
rect -4900 -10640 -4500 -10600
rect -3888 -10280 -3488 -10240
rect -3888 -10600 -3848 -10280
rect -3528 -10600 -3488 -10280
rect -3888 -10640 -3488 -10600
rect -2876 -10280 -2476 -10240
rect -2876 -10600 -2836 -10280
rect -2516 -10600 -2476 -10280
rect -2876 -10640 -2476 -10600
rect -1864 -10280 -1464 -10240
rect -1864 -10600 -1824 -10280
rect -1504 -10600 -1464 -10280
rect -1864 -10640 -1464 -10600
rect -852 -10280 -452 -10240
rect -852 -10600 -812 -10280
rect -492 -10600 -452 -10280
rect -852 -10640 -452 -10600
rect 160 -10280 560 -10240
rect 160 -10600 200 -10280
rect 520 -10600 560 -10280
rect 160 -10640 560 -10600
rect 1172 -10280 1572 -10240
rect 1172 -10600 1212 -10280
rect 1532 -10600 1572 -10280
rect 1172 -10640 1572 -10600
rect 2184 -10280 2584 -10240
rect 2184 -10600 2224 -10280
rect 2544 -10600 2584 -10280
rect 2184 -10640 2584 -10600
rect 3196 -10280 3596 -10240
rect 3196 -10600 3236 -10280
rect 3556 -10600 3596 -10280
rect 3196 -10640 3596 -10600
rect 4208 -10280 4608 -10240
rect 4208 -10600 4248 -10280
rect 4568 -10600 4608 -10280
rect 4208 -10640 4608 -10600
rect 5220 -10280 5620 -10240
rect 5220 -10600 5260 -10280
rect 5580 -10600 5620 -10280
rect 5220 -10640 5620 -10600
rect 6232 -10280 6632 -10240
rect 6232 -10600 6272 -10280
rect 6592 -10600 6632 -10280
rect 6232 -10640 6632 -10600
rect 7244 -10280 7644 -10240
rect 7244 -10600 7284 -10280
rect 7604 -10600 7644 -10280
rect 7244 -10640 7644 -10600
rect 8256 -10280 8656 -10240
rect 8256 -10600 8296 -10280
rect 8616 -10600 8656 -10280
rect 8256 -10640 8656 -10600
rect 9268 -10280 9668 -10240
rect 9268 -10600 9308 -10280
rect 9628 -10600 9668 -10280
rect 9268 -10640 9668 -10600
rect 10280 -10280 10680 -10240
rect 10280 -10600 10320 -10280
rect 10640 -10600 10680 -10280
rect 10280 -10640 10680 -10600
rect 11292 -10280 11692 -10240
rect 11292 -10600 11332 -10280
rect 11652 -10600 11692 -10280
rect 11292 -10640 11692 -10600
rect 12304 -10280 12704 -10240
rect 12304 -10600 12344 -10280
rect 12664 -10600 12704 -10280
rect 12304 -10640 12704 -10600
rect 13316 -10280 13716 -10240
rect 13316 -10600 13356 -10280
rect 13676 -10600 13716 -10280
rect 13316 -10640 13716 -10600
rect 14328 -10280 14728 -10240
rect 14328 -10600 14368 -10280
rect 14688 -10600 14728 -10280
rect 14328 -10640 14728 -10600
rect 15340 -10280 15740 -10240
rect 15340 -10600 15380 -10280
rect 15700 -10600 15740 -10280
rect 15340 -10640 15740 -10600
rect 16352 -10280 16752 -10240
rect 16352 -10600 16392 -10280
rect 16712 -10600 16752 -10280
rect 16352 -10640 16752 -10600
rect -17044 -11000 -16644 -10960
rect -17044 -11320 -17004 -11000
rect -16684 -11320 -16644 -11000
rect -17044 -11360 -16644 -11320
rect -16032 -11000 -15632 -10960
rect -16032 -11320 -15992 -11000
rect -15672 -11320 -15632 -11000
rect -16032 -11360 -15632 -11320
rect -15020 -11000 -14620 -10960
rect -15020 -11320 -14980 -11000
rect -14660 -11320 -14620 -11000
rect -15020 -11360 -14620 -11320
rect -14008 -11000 -13608 -10960
rect -14008 -11320 -13968 -11000
rect -13648 -11320 -13608 -11000
rect -14008 -11360 -13608 -11320
rect -12996 -11000 -12596 -10960
rect -12996 -11320 -12956 -11000
rect -12636 -11320 -12596 -11000
rect -12996 -11360 -12596 -11320
rect -11984 -11000 -11584 -10960
rect -11984 -11320 -11944 -11000
rect -11624 -11320 -11584 -11000
rect -11984 -11360 -11584 -11320
rect -10972 -11000 -10572 -10960
rect -10972 -11320 -10932 -11000
rect -10612 -11320 -10572 -11000
rect -10972 -11360 -10572 -11320
rect -9960 -11000 -9560 -10960
rect -9960 -11320 -9920 -11000
rect -9600 -11320 -9560 -11000
rect -9960 -11360 -9560 -11320
rect -8948 -11000 -8548 -10960
rect -8948 -11320 -8908 -11000
rect -8588 -11320 -8548 -11000
rect -8948 -11360 -8548 -11320
rect -7936 -11000 -7536 -10960
rect -7936 -11320 -7896 -11000
rect -7576 -11320 -7536 -11000
rect -7936 -11360 -7536 -11320
rect -6924 -11000 -6524 -10960
rect -6924 -11320 -6884 -11000
rect -6564 -11320 -6524 -11000
rect -6924 -11360 -6524 -11320
rect -5912 -11000 -5512 -10960
rect -5912 -11320 -5872 -11000
rect -5552 -11320 -5512 -11000
rect -5912 -11360 -5512 -11320
rect -4900 -11000 -4500 -10960
rect -4900 -11320 -4860 -11000
rect -4540 -11320 -4500 -11000
rect -4900 -11360 -4500 -11320
rect -3888 -11000 -3488 -10960
rect -3888 -11320 -3848 -11000
rect -3528 -11320 -3488 -11000
rect -3888 -11360 -3488 -11320
rect -2876 -11000 -2476 -10960
rect -2876 -11320 -2836 -11000
rect -2516 -11320 -2476 -11000
rect -2876 -11360 -2476 -11320
rect -1864 -11000 -1464 -10960
rect -1864 -11320 -1824 -11000
rect -1504 -11320 -1464 -11000
rect -1864 -11360 -1464 -11320
rect -852 -11000 -452 -10960
rect -852 -11320 -812 -11000
rect -492 -11320 -452 -11000
rect -852 -11360 -452 -11320
rect 160 -11000 560 -10960
rect 160 -11320 200 -11000
rect 520 -11320 560 -11000
rect 160 -11360 560 -11320
rect 1172 -11000 1572 -10960
rect 1172 -11320 1212 -11000
rect 1532 -11320 1572 -11000
rect 1172 -11360 1572 -11320
rect 2184 -11000 2584 -10960
rect 2184 -11320 2224 -11000
rect 2544 -11320 2584 -11000
rect 2184 -11360 2584 -11320
rect 3196 -11000 3596 -10960
rect 3196 -11320 3236 -11000
rect 3556 -11320 3596 -11000
rect 3196 -11360 3596 -11320
rect 4208 -11000 4608 -10960
rect 4208 -11320 4248 -11000
rect 4568 -11320 4608 -11000
rect 4208 -11360 4608 -11320
rect 5220 -11000 5620 -10960
rect 5220 -11320 5260 -11000
rect 5580 -11320 5620 -11000
rect 5220 -11360 5620 -11320
rect 6232 -11000 6632 -10960
rect 6232 -11320 6272 -11000
rect 6592 -11320 6632 -11000
rect 6232 -11360 6632 -11320
rect 7244 -11000 7644 -10960
rect 7244 -11320 7284 -11000
rect 7604 -11320 7644 -11000
rect 7244 -11360 7644 -11320
rect 8256 -11000 8656 -10960
rect 8256 -11320 8296 -11000
rect 8616 -11320 8656 -11000
rect 8256 -11360 8656 -11320
rect 9268 -11000 9668 -10960
rect 9268 -11320 9308 -11000
rect 9628 -11320 9668 -11000
rect 9268 -11360 9668 -11320
rect 10280 -11000 10680 -10960
rect 10280 -11320 10320 -11000
rect 10640 -11320 10680 -11000
rect 10280 -11360 10680 -11320
rect 11292 -11000 11692 -10960
rect 11292 -11320 11332 -11000
rect 11652 -11320 11692 -11000
rect 11292 -11360 11692 -11320
rect 12304 -11000 12704 -10960
rect 12304 -11320 12344 -11000
rect 12664 -11320 12704 -11000
rect 12304 -11360 12704 -11320
rect 13316 -11000 13716 -10960
rect 13316 -11320 13356 -11000
rect 13676 -11320 13716 -11000
rect 13316 -11360 13716 -11320
rect 14328 -11000 14728 -10960
rect 14328 -11320 14368 -11000
rect 14688 -11320 14728 -11000
rect 14328 -11360 14728 -11320
rect 15340 -11000 15740 -10960
rect 15340 -11320 15380 -11000
rect 15700 -11320 15740 -11000
rect 15340 -11360 15740 -11320
rect 16352 -11000 16752 -10960
rect 16352 -11320 16392 -11000
rect 16712 -11320 16752 -11000
rect 16352 -11360 16752 -11320
<< mimcapcontact >>
rect -17004 11000 -16684 11320
rect -15992 11000 -15672 11320
rect -14980 11000 -14660 11320
rect -13968 11000 -13648 11320
rect -12956 11000 -12636 11320
rect -11944 11000 -11624 11320
rect -10932 11000 -10612 11320
rect -9920 11000 -9600 11320
rect -8908 11000 -8588 11320
rect -7896 11000 -7576 11320
rect -6884 11000 -6564 11320
rect -5872 11000 -5552 11320
rect -4860 11000 -4540 11320
rect -3848 11000 -3528 11320
rect -2836 11000 -2516 11320
rect -1824 11000 -1504 11320
rect -812 11000 -492 11320
rect 200 11000 520 11320
rect 1212 11000 1532 11320
rect 2224 11000 2544 11320
rect 3236 11000 3556 11320
rect 4248 11000 4568 11320
rect 5260 11000 5580 11320
rect 6272 11000 6592 11320
rect 7284 11000 7604 11320
rect 8296 11000 8616 11320
rect 9308 11000 9628 11320
rect 10320 11000 10640 11320
rect 11332 11000 11652 11320
rect 12344 11000 12664 11320
rect 13356 11000 13676 11320
rect 14368 11000 14688 11320
rect 15380 11000 15700 11320
rect 16392 11000 16712 11320
rect -17004 10280 -16684 10600
rect -15992 10280 -15672 10600
rect -14980 10280 -14660 10600
rect -13968 10280 -13648 10600
rect -12956 10280 -12636 10600
rect -11944 10280 -11624 10600
rect -10932 10280 -10612 10600
rect -9920 10280 -9600 10600
rect -8908 10280 -8588 10600
rect -7896 10280 -7576 10600
rect -6884 10280 -6564 10600
rect -5872 10280 -5552 10600
rect -4860 10280 -4540 10600
rect -3848 10280 -3528 10600
rect -2836 10280 -2516 10600
rect -1824 10280 -1504 10600
rect -812 10280 -492 10600
rect 200 10280 520 10600
rect 1212 10280 1532 10600
rect 2224 10280 2544 10600
rect 3236 10280 3556 10600
rect 4248 10280 4568 10600
rect 5260 10280 5580 10600
rect 6272 10280 6592 10600
rect 7284 10280 7604 10600
rect 8296 10280 8616 10600
rect 9308 10280 9628 10600
rect 10320 10280 10640 10600
rect 11332 10280 11652 10600
rect 12344 10280 12664 10600
rect 13356 10280 13676 10600
rect 14368 10280 14688 10600
rect 15380 10280 15700 10600
rect 16392 10280 16712 10600
rect -17004 9560 -16684 9880
rect -15992 9560 -15672 9880
rect -14980 9560 -14660 9880
rect -13968 9560 -13648 9880
rect -12956 9560 -12636 9880
rect -11944 9560 -11624 9880
rect -10932 9560 -10612 9880
rect -9920 9560 -9600 9880
rect -8908 9560 -8588 9880
rect -7896 9560 -7576 9880
rect -6884 9560 -6564 9880
rect -5872 9560 -5552 9880
rect -4860 9560 -4540 9880
rect -3848 9560 -3528 9880
rect -2836 9560 -2516 9880
rect -1824 9560 -1504 9880
rect -812 9560 -492 9880
rect 200 9560 520 9880
rect 1212 9560 1532 9880
rect 2224 9560 2544 9880
rect 3236 9560 3556 9880
rect 4248 9560 4568 9880
rect 5260 9560 5580 9880
rect 6272 9560 6592 9880
rect 7284 9560 7604 9880
rect 8296 9560 8616 9880
rect 9308 9560 9628 9880
rect 10320 9560 10640 9880
rect 11332 9560 11652 9880
rect 12344 9560 12664 9880
rect 13356 9560 13676 9880
rect 14368 9560 14688 9880
rect 15380 9560 15700 9880
rect 16392 9560 16712 9880
rect -17004 8840 -16684 9160
rect -15992 8840 -15672 9160
rect -14980 8840 -14660 9160
rect -13968 8840 -13648 9160
rect -12956 8840 -12636 9160
rect -11944 8840 -11624 9160
rect -10932 8840 -10612 9160
rect -9920 8840 -9600 9160
rect -8908 8840 -8588 9160
rect -7896 8840 -7576 9160
rect -6884 8840 -6564 9160
rect -5872 8840 -5552 9160
rect -4860 8840 -4540 9160
rect -3848 8840 -3528 9160
rect -2836 8840 -2516 9160
rect -1824 8840 -1504 9160
rect -812 8840 -492 9160
rect 200 8840 520 9160
rect 1212 8840 1532 9160
rect 2224 8840 2544 9160
rect 3236 8840 3556 9160
rect 4248 8840 4568 9160
rect 5260 8840 5580 9160
rect 6272 8840 6592 9160
rect 7284 8840 7604 9160
rect 8296 8840 8616 9160
rect 9308 8840 9628 9160
rect 10320 8840 10640 9160
rect 11332 8840 11652 9160
rect 12344 8840 12664 9160
rect 13356 8840 13676 9160
rect 14368 8840 14688 9160
rect 15380 8840 15700 9160
rect 16392 8840 16712 9160
rect -17004 8120 -16684 8440
rect -15992 8120 -15672 8440
rect -14980 8120 -14660 8440
rect -13968 8120 -13648 8440
rect -12956 8120 -12636 8440
rect -11944 8120 -11624 8440
rect -10932 8120 -10612 8440
rect -9920 8120 -9600 8440
rect -8908 8120 -8588 8440
rect -7896 8120 -7576 8440
rect -6884 8120 -6564 8440
rect -5872 8120 -5552 8440
rect -4860 8120 -4540 8440
rect -3848 8120 -3528 8440
rect -2836 8120 -2516 8440
rect -1824 8120 -1504 8440
rect -812 8120 -492 8440
rect 200 8120 520 8440
rect 1212 8120 1532 8440
rect 2224 8120 2544 8440
rect 3236 8120 3556 8440
rect 4248 8120 4568 8440
rect 5260 8120 5580 8440
rect 6272 8120 6592 8440
rect 7284 8120 7604 8440
rect 8296 8120 8616 8440
rect 9308 8120 9628 8440
rect 10320 8120 10640 8440
rect 11332 8120 11652 8440
rect 12344 8120 12664 8440
rect 13356 8120 13676 8440
rect 14368 8120 14688 8440
rect 15380 8120 15700 8440
rect 16392 8120 16712 8440
rect -17004 7400 -16684 7720
rect -15992 7400 -15672 7720
rect -14980 7400 -14660 7720
rect -13968 7400 -13648 7720
rect -12956 7400 -12636 7720
rect -11944 7400 -11624 7720
rect -10932 7400 -10612 7720
rect -9920 7400 -9600 7720
rect -8908 7400 -8588 7720
rect -7896 7400 -7576 7720
rect -6884 7400 -6564 7720
rect -5872 7400 -5552 7720
rect -4860 7400 -4540 7720
rect -3848 7400 -3528 7720
rect -2836 7400 -2516 7720
rect -1824 7400 -1504 7720
rect -812 7400 -492 7720
rect 200 7400 520 7720
rect 1212 7400 1532 7720
rect 2224 7400 2544 7720
rect 3236 7400 3556 7720
rect 4248 7400 4568 7720
rect 5260 7400 5580 7720
rect 6272 7400 6592 7720
rect 7284 7400 7604 7720
rect 8296 7400 8616 7720
rect 9308 7400 9628 7720
rect 10320 7400 10640 7720
rect 11332 7400 11652 7720
rect 12344 7400 12664 7720
rect 13356 7400 13676 7720
rect 14368 7400 14688 7720
rect 15380 7400 15700 7720
rect 16392 7400 16712 7720
rect -17004 6680 -16684 7000
rect -15992 6680 -15672 7000
rect -14980 6680 -14660 7000
rect -13968 6680 -13648 7000
rect -12956 6680 -12636 7000
rect -11944 6680 -11624 7000
rect -10932 6680 -10612 7000
rect -9920 6680 -9600 7000
rect -8908 6680 -8588 7000
rect -7896 6680 -7576 7000
rect -6884 6680 -6564 7000
rect -5872 6680 -5552 7000
rect -4860 6680 -4540 7000
rect -3848 6680 -3528 7000
rect -2836 6680 -2516 7000
rect -1824 6680 -1504 7000
rect -812 6680 -492 7000
rect 200 6680 520 7000
rect 1212 6680 1532 7000
rect 2224 6680 2544 7000
rect 3236 6680 3556 7000
rect 4248 6680 4568 7000
rect 5260 6680 5580 7000
rect 6272 6680 6592 7000
rect 7284 6680 7604 7000
rect 8296 6680 8616 7000
rect 9308 6680 9628 7000
rect 10320 6680 10640 7000
rect 11332 6680 11652 7000
rect 12344 6680 12664 7000
rect 13356 6680 13676 7000
rect 14368 6680 14688 7000
rect 15380 6680 15700 7000
rect 16392 6680 16712 7000
rect -17004 5960 -16684 6280
rect -15992 5960 -15672 6280
rect -14980 5960 -14660 6280
rect -13968 5960 -13648 6280
rect -12956 5960 -12636 6280
rect -11944 5960 -11624 6280
rect -10932 5960 -10612 6280
rect -9920 5960 -9600 6280
rect -8908 5960 -8588 6280
rect -7896 5960 -7576 6280
rect -6884 5960 -6564 6280
rect -5872 5960 -5552 6280
rect -4860 5960 -4540 6280
rect -3848 5960 -3528 6280
rect -2836 5960 -2516 6280
rect -1824 5960 -1504 6280
rect -812 5960 -492 6280
rect 200 5960 520 6280
rect 1212 5960 1532 6280
rect 2224 5960 2544 6280
rect 3236 5960 3556 6280
rect 4248 5960 4568 6280
rect 5260 5960 5580 6280
rect 6272 5960 6592 6280
rect 7284 5960 7604 6280
rect 8296 5960 8616 6280
rect 9308 5960 9628 6280
rect 10320 5960 10640 6280
rect 11332 5960 11652 6280
rect 12344 5960 12664 6280
rect 13356 5960 13676 6280
rect 14368 5960 14688 6280
rect 15380 5960 15700 6280
rect 16392 5960 16712 6280
rect -17004 5240 -16684 5560
rect -15992 5240 -15672 5560
rect -14980 5240 -14660 5560
rect -13968 5240 -13648 5560
rect -12956 5240 -12636 5560
rect -11944 5240 -11624 5560
rect -10932 5240 -10612 5560
rect -9920 5240 -9600 5560
rect -8908 5240 -8588 5560
rect -7896 5240 -7576 5560
rect -6884 5240 -6564 5560
rect -5872 5240 -5552 5560
rect -4860 5240 -4540 5560
rect -3848 5240 -3528 5560
rect -2836 5240 -2516 5560
rect -1824 5240 -1504 5560
rect -812 5240 -492 5560
rect 200 5240 520 5560
rect 1212 5240 1532 5560
rect 2224 5240 2544 5560
rect 3236 5240 3556 5560
rect 4248 5240 4568 5560
rect 5260 5240 5580 5560
rect 6272 5240 6592 5560
rect 7284 5240 7604 5560
rect 8296 5240 8616 5560
rect 9308 5240 9628 5560
rect 10320 5240 10640 5560
rect 11332 5240 11652 5560
rect 12344 5240 12664 5560
rect 13356 5240 13676 5560
rect 14368 5240 14688 5560
rect 15380 5240 15700 5560
rect 16392 5240 16712 5560
rect -17004 4520 -16684 4840
rect -15992 4520 -15672 4840
rect -14980 4520 -14660 4840
rect -13968 4520 -13648 4840
rect -12956 4520 -12636 4840
rect -11944 4520 -11624 4840
rect -10932 4520 -10612 4840
rect -9920 4520 -9600 4840
rect -8908 4520 -8588 4840
rect -7896 4520 -7576 4840
rect -6884 4520 -6564 4840
rect -5872 4520 -5552 4840
rect -4860 4520 -4540 4840
rect -3848 4520 -3528 4840
rect -2836 4520 -2516 4840
rect -1824 4520 -1504 4840
rect -812 4520 -492 4840
rect 200 4520 520 4840
rect 1212 4520 1532 4840
rect 2224 4520 2544 4840
rect 3236 4520 3556 4840
rect 4248 4520 4568 4840
rect 5260 4520 5580 4840
rect 6272 4520 6592 4840
rect 7284 4520 7604 4840
rect 8296 4520 8616 4840
rect 9308 4520 9628 4840
rect 10320 4520 10640 4840
rect 11332 4520 11652 4840
rect 12344 4520 12664 4840
rect 13356 4520 13676 4840
rect 14368 4520 14688 4840
rect 15380 4520 15700 4840
rect 16392 4520 16712 4840
rect -17004 3800 -16684 4120
rect -15992 3800 -15672 4120
rect -14980 3800 -14660 4120
rect -13968 3800 -13648 4120
rect -12956 3800 -12636 4120
rect -11944 3800 -11624 4120
rect -10932 3800 -10612 4120
rect -9920 3800 -9600 4120
rect -8908 3800 -8588 4120
rect -7896 3800 -7576 4120
rect -6884 3800 -6564 4120
rect -5872 3800 -5552 4120
rect -4860 3800 -4540 4120
rect -3848 3800 -3528 4120
rect -2836 3800 -2516 4120
rect -1824 3800 -1504 4120
rect -812 3800 -492 4120
rect 200 3800 520 4120
rect 1212 3800 1532 4120
rect 2224 3800 2544 4120
rect 3236 3800 3556 4120
rect 4248 3800 4568 4120
rect 5260 3800 5580 4120
rect 6272 3800 6592 4120
rect 7284 3800 7604 4120
rect 8296 3800 8616 4120
rect 9308 3800 9628 4120
rect 10320 3800 10640 4120
rect 11332 3800 11652 4120
rect 12344 3800 12664 4120
rect 13356 3800 13676 4120
rect 14368 3800 14688 4120
rect 15380 3800 15700 4120
rect 16392 3800 16712 4120
rect -17004 3080 -16684 3400
rect -15992 3080 -15672 3400
rect -14980 3080 -14660 3400
rect -13968 3080 -13648 3400
rect -12956 3080 -12636 3400
rect -11944 3080 -11624 3400
rect -10932 3080 -10612 3400
rect -9920 3080 -9600 3400
rect -8908 3080 -8588 3400
rect -7896 3080 -7576 3400
rect -6884 3080 -6564 3400
rect -5872 3080 -5552 3400
rect -4860 3080 -4540 3400
rect -3848 3080 -3528 3400
rect -2836 3080 -2516 3400
rect -1824 3080 -1504 3400
rect -812 3080 -492 3400
rect 200 3080 520 3400
rect 1212 3080 1532 3400
rect 2224 3080 2544 3400
rect 3236 3080 3556 3400
rect 4248 3080 4568 3400
rect 5260 3080 5580 3400
rect 6272 3080 6592 3400
rect 7284 3080 7604 3400
rect 8296 3080 8616 3400
rect 9308 3080 9628 3400
rect 10320 3080 10640 3400
rect 11332 3080 11652 3400
rect 12344 3080 12664 3400
rect 13356 3080 13676 3400
rect 14368 3080 14688 3400
rect 15380 3080 15700 3400
rect 16392 3080 16712 3400
rect -17004 2360 -16684 2680
rect -15992 2360 -15672 2680
rect -14980 2360 -14660 2680
rect -13968 2360 -13648 2680
rect -12956 2360 -12636 2680
rect -11944 2360 -11624 2680
rect -10932 2360 -10612 2680
rect -9920 2360 -9600 2680
rect -8908 2360 -8588 2680
rect -7896 2360 -7576 2680
rect -6884 2360 -6564 2680
rect -5872 2360 -5552 2680
rect -4860 2360 -4540 2680
rect -3848 2360 -3528 2680
rect -2836 2360 -2516 2680
rect -1824 2360 -1504 2680
rect -812 2360 -492 2680
rect 200 2360 520 2680
rect 1212 2360 1532 2680
rect 2224 2360 2544 2680
rect 3236 2360 3556 2680
rect 4248 2360 4568 2680
rect 5260 2360 5580 2680
rect 6272 2360 6592 2680
rect 7284 2360 7604 2680
rect 8296 2360 8616 2680
rect 9308 2360 9628 2680
rect 10320 2360 10640 2680
rect 11332 2360 11652 2680
rect 12344 2360 12664 2680
rect 13356 2360 13676 2680
rect 14368 2360 14688 2680
rect 15380 2360 15700 2680
rect 16392 2360 16712 2680
rect -17004 1640 -16684 1960
rect -15992 1640 -15672 1960
rect -14980 1640 -14660 1960
rect -13968 1640 -13648 1960
rect -12956 1640 -12636 1960
rect -11944 1640 -11624 1960
rect -10932 1640 -10612 1960
rect -9920 1640 -9600 1960
rect -8908 1640 -8588 1960
rect -7896 1640 -7576 1960
rect -6884 1640 -6564 1960
rect -5872 1640 -5552 1960
rect -4860 1640 -4540 1960
rect -3848 1640 -3528 1960
rect -2836 1640 -2516 1960
rect -1824 1640 -1504 1960
rect -812 1640 -492 1960
rect 200 1640 520 1960
rect 1212 1640 1532 1960
rect 2224 1640 2544 1960
rect 3236 1640 3556 1960
rect 4248 1640 4568 1960
rect 5260 1640 5580 1960
rect 6272 1640 6592 1960
rect 7284 1640 7604 1960
rect 8296 1640 8616 1960
rect 9308 1640 9628 1960
rect 10320 1640 10640 1960
rect 11332 1640 11652 1960
rect 12344 1640 12664 1960
rect 13356 1640 13676 1960
rect 14368 1640 14688 1960
rect 15380 1640 15700 1960
rect 16392 1640 16712 1960
rect -17004 920 -16684 1240
rect -15992 920 -15672 1240
rect -14980 920 -14660 1240
rect -13968 920 -13648 1240
rect -12956 920 -12636 1240
rect -11944 920 -11624 1240
rect -10932 920 -10612 1240
rect -9920 920 -9600 1240
rect -8908 920 -8588 1240
rect -7896 920 -7576 1240
rect -6884 920 -6564 1240
rect -5872 920 -5552 1240
rect -4860 920 -4540 1240
rect -3848 920 -3528 1240
rect -2836 920 -2516 1240
rect -1824 920 -1504 1240
rect -812 920 -492 1240
rect 200 920 520 1240
rect 1212 920 1532 1240
rect 2224 920 2544 1240
rect 3236 920 3556 1240
rect 4248 920 4568 1240
rect 5260 920 5580 1240
rect 6272 920 6592 1240
rect 7284 920 7604 1240
rect 8296 920 8616 1240
rect 9308 920 9628 1240
rect 10320 920 10640 1240
rect 11332 920 11652 1240
rect 12344 920 12664 1240
rect 13356 920 13676 1240
rect 14368 920 14688 1240
rect 15380 920 15700 1240
rect 16392 920 16712 1240
rect -17004 200 -16684 520
rect -15992 200 -15672 520
rect -14980 200 -14660 520
rect -13968 200 -13648 520
rect -12956 200 -12636 520
rect -11944 200 -11624 520
rect -10932 200 -10612 520
rect -9920 200 -9600 520
rect -8908 200 -8588 520
rect -7896 200 -7576 520
rect -6884 200 -6564 520
rect -5872 200 -5552 520
rect -4860 200 -4540 520
rect -3848 200 -3528 520
rect -2836 200 -2516 520
rect -1824 200 -1504 520
rect -812 200 -492 520
rect 200 200 520 520
rect 1212 200 1532 520
rect 2224 200 2544 520
rect 3236 200 3556 520
rect 4248 200 4568 520
rect 5260 200 5580 520
rect 6272 200 6592 520
rect 7284 200 7604 520
rect 8296 200 8616 520
rect 9308 200 9628 520
rect 10320 200 10640 520
rect 11332 200 11652 520
rect 12344 200 12664 520
rect 13356 200 13676 520
rect 14368 200 14688 520
rect 15380 200 15700 520
rect 16392 200 16712 520
rect -17004 -520 -16684 -200
rect -15992 -520 -15672 -200
rect -14980 -520 -14660 -200
rect -13968 -520 -13648 -200
rect -12956 -520 -12636 -200
rect -11944 -520 -11624 -200
rect -10932 -520 -10612 -200
rect -9920 -520 -9600 -200
rect -8908 -520 -8588 -200
rect -7896 -520 -7576 -200
rect -6884 -520 -6564 -200
rect -5872 -520 -5552 -200
rect -4860 -520 -4540 -200
rect -3848 -520 -3528 -200
rect -2836 -520 -2516 -200
rect -1824 -520 -1504 -200
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect 1212 -520 1532 -200
rect 2224 -520 2544 -200
rect 3236 -520 3556 -200
rect 4248 -520 4568 -200
rect 5260 -520 5580 -200
rect 6272 -520 6592 -200
rect 7284 -520 7604 -200
rect 8296 -520 8616 -200
rect 9308 -520 9628 -200
rect 10320 -520 10640 -200
rect 11332 -520 11652 -200
rect 12344 -520 12664 -200
rect 13356 -520 13676 -200
rect 14368 -520 14688 -200
rect 15380 -520 15700 -200
rect 16392 -520 16712 -200
rect -17004 -1240 -16684 -920
rect -15992 -1240 -15672 -920
rect -14980 -1240 -14660 -920
rect -13968 -1240 -13648 -920
rect -12956 -1240 -12636 -920
rect -11944 -1240 -11624 -920
rect -10932 -1240 -10612 -920
rect -9920 -1240 -9600 -920
rect -8908 -1240 -8588 -920
rect -7896 -1240 -7576 -920
rect -6884 -1240 -6564 -920
rect -5872 -1240 -5552 -920
rect -4860 -1240 -4540 -920
rect -3848 -1240 -3528 -920
rect -2836 -1240 -2516 -920
rect -1824 -1240 -1504 -920
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect 1212 -1240 1532 -920
rect 2224 -1240 2544 -920
rect 3236 -1240 3556 -920
rect 4248 -1240 4568 -920
rect 5260 -1240 5580 -920
rect 6272 -1240 6592 -920
rect 7284 -1240 7604 -920
rect 8296 -1240 8616 -920
rect 9308 -1240 9628 -920
rect 10320 -1240 10640 -920
rect 11332 -1240 11652 -920
rect 12344 -1240 12664 -920
rect 13356 -1240 13676 -920
rect 14368 -1240 14688 -920
rect 15380 -1240 15700 -920
rect 16392 -1240 16712 -920
rect -17004 -1960 -16684 -1640
rect -15992 -1960 -15672 -1640
rect -14980 -1960 -14660 -1640
rect -13968 -1960 -13648 -1640
rect -12956 -1960 -12636 -1640
rect -11944 -1960 -11624 -1640
rect -10932 -1960 -10612 -1640
rect -9920 -1960 -9600 -1640
rect -8908 -1960 -8588 -1640
rect -7896 -1960 -7576 -1640
rect -6884 -1960 -6564 -1640
rect -5872 -1960 -5552 -1640
rect -4860 -1960 -4540 -1640
rect -3848 -1960 -3528 -1640
rect -2836 -1960 -2516 -1640
rect -1824 -1960 -1504 -1640
rect -812 -1960 -492 -1640
rect 200 -1960 520 -1640
rect 1212 -1960 1532 -1640
rect 2224 -1960 2544 -1640
rect 3236 -1960 3556 -1640
rect 4248 -1960 4568 -1640
rect 5260 -1960 5580 -1640
rect 6272 -1960 6592 -1640
rect 7284 -1960 7604 -1640
rect 8296 -1960 8616 -1640
rect 9308 -1960 9628 -1640
rect 10320 -1960 10640 -1640
rect 11332 -1960 11652 -1640
rect 12344 -1960 12664 -1640
rect 13356 -1960 13676 -1640
rect 14368 -1960 14688 -1640
rect 15380 -1960 15700 -1640
rect 16392 -1960 16712 -1640
rect -17004 -2680 -16684 -2360
rect -15992 -2680 -15672 -2360
rect -14980 -2680 -14660 -2360
rect -13968 -2680 -13648 -2360
rect -12956 -2680 -12636 -2360
rect -11944 -2680 -11624 -2360
rect -10932 -2680 -10612 -2360
rect -9920 -2680 -9600 -2360
rect -8908 -2680 -8588 -2360
rect -7896 -2680 -7576 -2360
rect -6884 -2680 -6564 -2360
rect -5872 -2680 -5552 -2360
rect -4860 -2680 -4540 -2360
rect -3848 -2680 -3528 -2360
rect -2836 -2680 -2516 -2360
rect -1824 -2680 -1504 -2360
rect -812 -2680 -492 -2360
rect 200 -2680 520 -2360
rect 1212 -2680 1532 -2360
rect 2224 -2680 2544 -2360
rect 3236 -2680 3556 -2360
rect 4248 -2680 4568 -2360
rect 5260 -2680 5580 -2360
rect 6272 -2680 6592 -2360
rect 7284 -2680 7604 -2360
rect 8296 -2680 8616 -2360
rect 9308 -2680 9628 -2360
rect 10320 -2680 10640 -2360
rect 11332 -2680 11652 -2360
rect 12344 -2680 12664 -2360
rect 13356 -2680 13676 -2360
rect 14368 -2680 14688 -2360
rect 15380 -2680 15700 -2360
rect 16392 -2680 16712 -2360
rect -17004 -3400 -16684 -3080
rect -15992 -3400 -15672 -3080
rect -14980 -3400 -14660 -3080
rect -13968 -3400 -13648 -3080
rect -12956 -3400 -12636 -3080
rect -11944 -3400 -11624 -3080
rect -10932 -3400 -10612 -3080
rect -9920 -3400 -9600 -3080
rect -8908 -3400 -8588 -3080
rect -7896 -3400 -7576 -3080
rect -6884 -3400 -6564 -3080
rect -5872 -3400 -5552 -3080
rect -4860 -3400 -4540 -3080
rect -3848 -3400 -3528 -3080
rect -2836 -3400 -2516 -3080
rect -1824 -3400 -1504 -3080
rect -812 -3400 -492 -3080
rect 200 -3400 520 -3080
rect 1212 -3400 1532 -3080
rect 2224 -3400 2544 -3080
rect 3236 -3400 3556 -3080
rect 4248 -3400 4568 -3080
rect 5260 -3400 5580 -3080
rect 6272 -3400 6592 -3080
rect 7284 -3400 7604 -3080
rect 8296 -3400 8616 -3080
rect 9308 -3400 9628 -3080
rect 10320 -3400 10640 -3080
rect 11332 -3400 11652 -3080
rect 12344 -3400 12664 -3080
rect 13356 -3400 13676 -3080
rect 14368 -3400 14688 -3080
rect 15380 -3400 15700 -3080
rect 16392 -3400 16712 -3080
rect -17004 -4120 -16684 -3800
rect -15992 -4120 -15672 -3800
rect -14980 -4120 -14660 -3800
rect -13968 -4120 -13648 -3800
rect -12956 -4120 -12636 -3800
rect -11944 -4120 -11624 -3800
rect -10932 -4120 -10612 -3800
rect -9920 -4120 -9600 -3800
rect -8908 -4120 -8588 -3800
rect -7896 -4120 -7576 -3800
rect -6884 -4120 -6564 -3800
rect -5872 -4120 -5552 -3800
rect -4860 -4120 -4540 -3800
rect -3848 -4120 -3528 -3800
rect -2836 -4120 -2516 -3800
rect -1824 -4120 -1504 -3800
rect -812 -4120 -492 -3800
rect 200 -4120 520 -3800
rect 1212 -4120 1532 -3800
rect 2224 -4120 2544 -3800
rect 3236 -4120 3556 -3800
rect 4248 -4120 4568 -3800
rect 5260 -4120 5580 -3800
rect 6272 -4120 6592 -3800
rect 7284 -4120 7604 -3800
rect 8296 -4120 8616 -3800
rect 9308 -4120 9628 -3800
rect 10320 -4120 10640 -3800
rect 11332 -4120 11652 -3800
rect 12344 -4120 12664 -3800
rect 13356 -4120 13676 -3800
rect 14368 -4120 14688 -3800
rect 15380 -4120 15700 -3800
rect 16392 -4120 16712 -3800
rect -17004 -4840 -16684 -4520
rect -15992 -4840 -15672 -4520
rect -14980 -4840 -14660 -4520
rect -13968 -4840 -13648 -4520
rect -12956 -4840 -12636 -4520
rect -11944 -4840 -11624 -4520
rect -10932 -4840 -10612 -4520
rect -9920 -4840 -9600 -4520
rect -8908 -4840 -8588 -4520
rect -7896 -4840 -7576 -4520
rect -6884 -4840 -6564 -4520
rect -5872 -4840 -5552 -4520
rect -4860 -4840 -4540 -4520
rect -3848 -4840 -3528 -4520
rect -2836 -4840 -2516 -4520
rect -1824 -4840 -1504 -4520
rect -812 -4840 -492 -4520
rect 200 -4840 520 -4520
rect 1212 -4840 1532 -4520
rect 2224 -4840 2544 -4520
rect 3236 -4840 3556 -4520
rect 4248 -4840 4568 -4520
rect 5260 -4840 5580 -4520
rect 6272 -4840 6592 -4520
rect 7284 -4840 7604 -4520
rect 8296 -4840 8616 -4520
rect 9308 -4840 9628 -4520
rect 10320 -4840 10640 -4520
rect 11332 -4840 11652 -4520
rect 12344 -4840 12664 -4520
rect 13356 -4840 13676 -4520
rect 14368 -4840 14688 -4520
rect 15380 -4840 15700 -4520
rect 16392 -4840 16712 -4520
rect -17004 -5560 -16684 -5240
rect -15992 -5560 -15672 -5240
rect -14980 -5560 -14660 -5240
rect -13968 -5560 -13648 -5240
rect -12956 -5560 -12636 -5240
rect -11944 -5560 -11624 -5240
rect -10932 -5560 -10612 -5240
rect -9920 -5560 -9600 -5240
rect -8908 -5560 -8588 -5240
rect -7896 -5560 -7576 -5240
rect -6884 -5560 -6564 -5240
rect -5872 -5560 -5552 -5240
rect -4860 -5560 -4540 -5240
rect -3848 -5560 -3528 -5240
rect -2836 -5560 -2516 -5240
rect -1824 -5560 -1504 -5240
rect -812 -5560 -492 -5240
rect 200 -5560 520 -5240
rect 1212 -5560 1532 -5240
rect 2224 -5560 2544 -5240
rect 3236 -5560 3556 -5240
rect 4248 -5560 4568 -5240
rect 5260 -5560 5580 -5240
rect 6272 -5560 6592 -5240
rect 7284 -5560 7604 -5240
rect 8296 -5560 8616 -5240
rect 9308 -5560 9628 -5240
rect 10320 -5560 10640 -5240
rect 11332 -5560 11652 -5240
rect 12344 -5560 12664 -5240
rect 13356 -5560 13676 -5240
rect 14368 -5560 14688 -5240
rect 15380 -5560 15700 -5240
rect 16392 -5560 16712 -5240
rect -17004 -6280 -16684 -5960
rect -15992 -6280 -15672 -5960
rect -14980 -6280 -14660 -5960
rect -13968 -6280 -13648 -5960
rect -12956 -6280 -12636 -5960
rect -11944 -6280 -11624 -5960
rect -10932 -6280 -10612 -5960
rect -9920 -6280 -9600 -5960
rect -8908 -6280 -8588 -5960
rect -7896 -6280 -7576 -5960
rect -6884 -6280 -6564 -5960
rect -5872 -6280 -5552 -5960
rect -4860 -6280 -4540 -5960
rect -3848 -6280 -3528 -5960
rect -2836 -6280 -2516 -5960
rect -1824 -6280 -1504 -5960
rect -812 -6280 -492 -5960
rect 200 -6280 520 -5960
rect 1212 -6280 1532 -5960
rect 2224 -6280 2544 -5960
rect 3236 -6280 3556 -5960
rect 4248 -6280 4568 -5960
rect 5260 -6280 5580 -5960
rect 6272 -6280 6592 -5960
rect 7284 -6280 7604 -5960
rect 8296 -6280 8616 -5960
rect 9308 -6280 9628 -5960
rect 10320 -6280 10640 -5960
rect 11332 -6280 11652 -5960
rect 12344 -6280 12664 -5960
rect 13356 -6280 13676 -5960
rect 14368 -6280 14688 -5960
rect 15380 -6280 15700 -5960
rect 16392 -6280 16712 -5960
rect -17004 -7000 -16684 -6680
rect -15992 -7000 -15672 -6680
rect -14980 -7000 -14660 -6680
rect -13968 -7000 -13648 -6680
rect -12956 -7000 -12636 -6680
rect -11944 -7000 -11624 -6680
rect -10932 -7000 -10612 -6680
rect -9920 -7000 -9600 -6680
rect -8908 -7000 -8588 -6680
rect -7896 -7000 -7576 -6680
rect -6884 -7000 -6564 -6680
rect -5872 -7000 -5552 -6680
rect -4860 -7000 -4540 -6680
rect -3848 -7000 -3528 -6680
rect -2836 -7000 -2516 -6680
rect -1824 -7000 -1504 -6680
rect -812 -7000 -492 -6680
rect 200 -7000 520 -6680
rect 1212 -7000 1532 -6680
rect 2224 -7000 2544 -6680
rect 3236 -7000 3556 -6680
rect 4248 -7000 4568 -6680
rect 5260 -7000 5580 -6680
rect 6272 -7000 6592 -6680
rect 7284 -7000 7604 -6680
rect 8296 -7000 8616 -6680
rect 9308 -7000 9628 -6680
rect 10320 -7000 10640 -6680
rect 11332 -7000 11652 -6680
rect 12344 -7000 12664 -6680
rect 13356 -7000 13676 -6680
rect 14368 -7000 14688 -6680
rect 15380 -7000 15700 -6680
rect 16392 -7000 16712 -6680
rect -17004 -7720 -16684 -7400
rect -15992 -7720 -15672 -7400
rect -14980 -7720 -14660 -7400
rect -13968 -7720 -13648 -7400
rect -12956 -7720 -12636 -7400
rect -11944 -7720 -11624 -7400
rect -10932 -7720 -10612 -7400
rect -9920 -7720 -9600 -7400
rect -8908 -7720 -8588 -7400
rect -7896 -7720 -7576 -7400
rect -6884 -7720 -6564 -7400
rect -5872 -7720 -5552 -7400
rect -4860 -7720 -4540 -7400
rect -3848 -7720 -3528 -7400
rect -2836 -7720 -2516 -7400
rect -1824 -7720 -1504 -7400
rect -812 -7720 -492 -7400
rect 200 -7720 520 -7400
rect 1212 -7720 1532 -7400
rect 2224 -7720 2544 -7400
rect 3236 -7720 3556 -7400
rect 4248 -7720 4568 -7400
rect 5260 -7720 5580 -7400
rect 6272 -7720 6592 -7400
rect 7284 -7720 7604 -7400
rect 8296 -7720 8616 -7400
rect 9308 -7720 9628 -7400
rect 10320 -7720 10640 -7400
rect 11332 -7720 11652 -7400
rect 12344 -7720 12664 -7400
rect 13356 -7720 13676 -7400
rect 14368 -7720 14688 -7400
rect 15380 -7720 15700 -7400
rect 16392 -7720 16712 -7400
rect -17004 -8440 -16684 -8120
rect -15992 -8440 -15672 -8120
rect -14980 -8440 -14660 -8120
rect -13968 -8440 -13648 -8120
rect -12956 -8440 -12636 -8120
rect -11944 -8440 -11624 -8120
rect -10932 -8440 -10612 -8120
rect -9920 -8440 -9600 -8120
rect -8908 -8440 -8588 -8120
rect -7896 -8440 -7576 -8120
rect -6884 -8440 -6564 -8120
rect -5872 -8440 -5552 -8120
rect -4860 -8440 -4540 -8120
rect -3848 -8440 -3528 -8120
rect -2836 -8440 -2516 -8120
rect -1824 -8440 -1504 -8120
rect -812 -8440 -492 -8120
rect 200 -8440 520 -8120
rect 1212 -8440 1532 -8120
rect 2224 -8440 2544 -8120
rect 3236 -8440 3556 -8120
rect 4248 -8440 4568 -8120
rect 5260 -8440 5580 -8120
rect 6272 -8440 6592 -8120
rect 7284 -8440 7604 -8120
rect 8296 -8440 8616 -8120
rect 9308 -8440 9628 -8120
rect 10320 -8440 10640 -8120
rect 11332 -8440 11652 -8120
rect 12344 -8440 12664 -8120
rect 13356 -8440 13676 -8120
rect 14368 -8440 14688 -8120
rect 15380 -8440 15700 -8120
rect 16392 -8440 16712 -8120
rect -17004 -9160 -16684 -8840
rect -15992 -9160 -15672 -8840
rect -14980 -9160 -14660 -8840
rect -13968 -9160 -13648 -8840
rect -12956 -9160 -12636 -8840
rect -11944 -9160 -11624 -8840
rect -10932 -9160 -10612 -8840
rect -9920 -9160 -9600 -8840
rect -8908 -9160 -8588 -8840
rect -7896 -9160 -7576 -8840
rect -6884 -9160 -6564 -8840
rect -5872 -9160 -5552 -8840
rect -4860 -9160 -4540 -8840
rect -3848 -9160 -3528 -8840
rect -2836 -9160 -2516 -8840
rect -1824 -9160 -1504 -8840
rect -812 -9160 -492 -8840
rect 200 -9160 520 -8840
rect 1212 -9160 1532 -8840
rect 2224 -9160 2544 -8840
rect 3236 -9160 3556 -8840
rect 4248 -9160 4568 -8840
rect 5260 -9160 5580 -8840
rect 6272 -9160 6592 -8840
rect 7284 -9160 7604 -8840
rect 8296 -9160 8616 -8840
rect 9308 -9160 9628 -8840
rect 10320 -9160 10640 -8840
rect 11332 -9160 11652 -8840
rect 12344 -9160 12664 -8840
rect 13356 -9160 13676 -8840
rect 14368 -9160 14688 -8840
rect 15380 -9160 15700 -8840
rect 16392 -9160 16712 -8840
rect -17004 -9880 -16684 -9560
rect -15992 -9880 -15672 -9560
rect -14980 -9880 -14660 -9560
rect -13968 -9880 -13648 -9560
rect -12956 -9880 -12636 -9560
rect -11944 -9880 -11624 -9560
rect -10932 -9880 -10612 -9560
rect -9920 -9880 -9600 -9560
rect -8908 -9880 -8588 -9560
rect -7896 -9880 -7576 -9560
rect -6884 -9880 -6564 -9560
rect -5872 -9880 -5552 -9560
rect -4860 -9880 -4540 -9560
rect -3848 -9880 -3528 -9560
rect -2836 -9880 -2516 -9560
rect -1824 -9880 -1504 -9560
rect -812 -9880 -492 -9560
rect 200 -9880 520 -9560
rect 1212 -9880 1532 -9560
rect 2224 -9880 2544 -9560
rect 3236 -9880 3556 -9560
rect 4248 -9880 4568 -9560
rect 5260 -9880 5580 -9560
rect 6272 -9880 6592 -9560
rect 7284 -9880 7604 -9560
rect 8296 -9880 8616 -9560
rect 9308 -9880 9628 -9560
rect 10320 -9880 10640 -9560
rect 11332 -9880 11652 -9560
rect 12344 -9880 12664 -9560
rect 13356 -9880 13676 -9560
rect 14368 -9880 14688 -9560
rect 15380 -9880 15700 -9560
rect 16392 -9880 16712 -9560
rect -17004 -10600 -16684 -10280
rect -15992 -10600 -15672 -10280
rect -14980 -10600 -14660 -10280
rect -13968 -10600 -13648 -10280
rect -12956 -10600 -12636 -10280
rect -11944 -10600 -11624 -10280
rect -10932 -10600 -10612 -10280
rect -9920 -10600 -9600 -10280
rect -8908 -10600 -8588 -10280
rect -7896 -10600 -7576 -10280
rect -6884 -10600 -6564 -10280
rect -5872 -10600 -5552 -10280
rect -4860 -10600 -4540 -10280
rect -3848 -10600 -3528 -10280
rect -2836 -10600 -2516 -10280
rect -1824 -10600 -1504 -10280
rect -812 -10600 -492 -10280
rect 200 -10600 520 -10280
rect 1212 -10600 1532 -10280
rect 2224 -10600 2544 -10280
rect 3236 -10600 3556 -10280
rect 4248 -10600 4568 -10280
rect 5260 -10600 5580 -10280
rect 6272 -10600 6592 -10280
rect 7284 -10600 7604 -10280
rect 8296 -10600 8616 -10280
rect 9308 -10600 9628 -10280
rect 10320 -10600 10640 -10280
rect 11332 -10600 11652 -10280
rect 12344 -10600 12664 -10280
rect 13356 -10600 13676 -10280
rect 14368 -10600 14688 -10280
rect 15380 -10600 15700 -10280
rect 16392 -10600 16712 -10280
rect -17004 -11320 -16684 -11000
rect -15992 -11320 -15672 -11000
rect -14980 -11320 -14660 -11000
rect -13968 -11320 -13648 -11000
rect -12956 -11320 -12636 -11000
rect -11944 -11320 -11624 -11000
rect -10932 -11320 -10612 -11000
rect -9920 -11320 -9600 -11000
rect -8908 -11320 -8588 -11000
rect -7896 -11320 -7576 -11000
rect -6884 -11320 -6564 -11000
rect -5872 -11320 -5552 -11000
rect -4860 -11320 -4540 -11000
rect -3848 -11320 -3528 -11000
rect -2836 -11320 -2516 -11000
rect -1824 -11320 -1504 -11000
rect -812 -11320 -492 -11000
rect 200 -11320 520 -11000
rect 1212 -11320 1532 -11000
rect 2224 -11320 2544 -11000
rect 3236 -11320 3556 -11000
rect 4248 -11320 4568 -11000
rect 5260 -11320 5580 -11000
rect 6272 -11320 6592 -11000
rect 7284 -11320 7604 -11000
rect 8296 -11320 8616 -11000
rect 9308 -11320 9628 -11000
rect 10320 -11320 10640 -11000
rect 11332 -11320 11652 -11000
rect 12344 -11320 12664 -11000
rect 13356 -11320 13676 -11000
rect 14368 -11320 14688 -11000
rect 15380 -11320 15700 -11000
rect 16392 -11320 16712 -11000
<< metal4 >>
rect -16412 11372 -16316 11388
rect -17005 11320 -16683 11321
rect -17005 11000 -17004 11320
rect -16684 11000 -16683 11320
rect -17005 10999 -16683 11000
rect -16412 10948 -16396 11372
rect -16332 10948 -16316 11372
rect -15400 11372 -15304 11388
rect -15993 11320 -15671 11321
rect -15993 11000 -15992 11320
rect -15672 11000 -15671 11320
rect -15993 10999 -15671 11000
rect -16412 10932 -16316 10948
rect -15400 10948 -15384 11372
rect -15320 10948 -15304 11372
rect -14388 11372 -14292 11388
rect -14981 11320 -14659 11321
rect -14981 11000 -14980 11320
rect -14660 11000 -14659 11320
rect -14981 10999 -14659 11000
rect -15400 10932 -15304 10948
rect -14388 10948 -14372 11372
rect -14308 10948 -14292 11372
rect -13376 11372 -13280 11388
rect -13969 11320 -13647 11321
rect -13969 11000 -13968 11320
rect -13648 11000 -13647 11320
rect -13969 10999 -13647 11000
rect -14388 10932 -14292 10948
rect -13376 10948 -13360 11372
rect -13296 10948 -13280 11372
rect -12364 11372 -12268 11388
rect -12957 11320 -12635 11321
rect -12957 11000 -12956 11320
rect -12636 11000 -12635 11320
rect -12957 10999 -12635 11000
rect -13376 10932 -13280 10948
rect -12364 10948 -12348 11372
rect -12284 10948 -12268 11372
rect -11352 11372 -11256 11388
rect -11945 11320 -11623 11321
rect -11945 11000 -11944 11320
rect -11624 11000 -11623 11320
rect -11945 10999 -11623 11000
rect -12364 10932 -12268 10948
rect -11352 10948 -11336 11372
rect -11272 10948 -11256 11372
rect -10340 11372 -10244 11388
rect -10933 11320 -10611 11321
rect -10933 11000 -10932 11320
rect -10612 11000 -10611 11320
rect -10933 10999 -10611 11000
rect -11352 10932 -11256 10948
rect -10340 10948 -10324 11372
rect -10260 10948 -10244 11372
rect -9328 11372 -9232 11388
rect -9921 11320 -9599 11321
rect -9921 11000 -9920 11320
rect -9600 11000 -9599 11320
rect -9921 10999 -9599 11000
rect -10340 10932 -10244 10948
rect -9328 10948 -9312 11372
rect -9248 10948 -9232 11372
rect -8316 11372 -8220 11388
rect -8909 11320 -8587 11321
rect -8909 11000 -8908 11320
rect -8588 11000 -8587 11320
rect -8909 10999 -8587 11000
rect -9328 10932 -9232 10948
rect -8316 10948 -8300 11372
rect -8236 10948 -8220 11372
rect -7304 11372 -7208 11388
rect -7897 11320 -7575 11321
rect -7897 11000 -7896 11320
rect -7576 11000 -7575 11320
rect -7897 10999 -7575 11000
rect -8316 10932 -8220 10948
rect -7304 10948 -7288 11372
rect -7224 10948 -7208 11372
rect -6292 11372 -6196 11388
rect -6885 11320 -6563 11321
rect -6885 11000 -6884 11320
rect -6564 11000 -6563 11320
rect -6885 10999 -6563 11000
rect -7304 10932 -7208 10948
rect -6292 10948 -6276 11372
rect -6212 10948 -6196 11372
rect -5280 11372 -5184 11388
rect -5873 11320 -5551 11321
rect -5873 11000 -5872 11320
rect -5552 11000 -5551 11320
rect -5873 10999 -5551 11000
rect -6292 10932 -6196 10948
rect -5280 10948 -5264 11372
rect -5200 10948 -5184 11372
rect -4268 11372 -4172 11388
rect -4861 11320 -4539 11321
rect -4861 11000 -4860 11320
rect -4540 11000 -4539 11320
rect -4861 10999 -4539 11000
rect -5280 10932 -5184 10948
rect -4268 10948 -4252 11372
rect -4188 10948 -4172 11372
rect -3256 11372 -3160 11388
rect -3849 11320 -3527 11321
rect -3849 11000 -3848 11320
rect -3528 11000 -3527 11320
rect -3849 10999 -3527 11000
rect -4268 10932 -4172 10948
rect -3256 10948 -3240 11372
rect -3176 10948 -3160 11372
rect -2244 11372 -2148 11388
rect -2837 11320 -2515 11321
rect -2837 11000 -2836 11320
rect -2516 11000 -2515 11320
rect -2837 10999 -2515 11000
rect -3256 10932 -3160 10948
rect -2244 10948 -2228 11372
rect -2164 10948 -2148 11372
rect -1232 11372 -1136 11388
rect -1825 11320 -1503 11321
rect -1825 11000 -1824 11320
rect -1504 11000 -1503 11320
rect -1825 10999 -1503 11000
rect -2244 10932 -2148 10948
rect -1232 10948 -1216 11372
rect -1152 10948 -1136 11372
rect -220 11372 -124 11388
rect -813 11320 -491 11321
rect -813 11000 -812 11320
rect -492 11000 -491 11320
rect -813 10999 -491 11000
rect -1232 10932 -1136 10948
rect -220 10948 -204 11372
rect -140 10948 -124 11372
rect 792 11372 888 11388
rect 199 11320 521 11321
rect 199 11000 200 11320
rect 520 11000 521 11320
rect 199 10999 521 11000
rect -220 10932 -124 10948
rect 792 10948 808 11372
rect 872 10948 888 11372
rect 1804 11372 1900 11388
rect 1211 11320 1533 11321
rect 1211 11000 1212 11320
rect 1532 11000 1533 11320
rect 1211 10999 1533 11000
rect 792 10932 888 10948
rect 1804 10948 1820 11372
rect 1884 10948 1900 11372
rect 2816 11372 2912 11388
rect 2223 11320 2545 11321
rect 2223 11000 2224 11320
rect 2544 11000 2545 11320
rect 2223 10999 2545 11000
rect 1804 10932 1900 10948
rect 2816 10948 2832 11372
rect 2896 10948 2912 11372
rect 3828 11372 3924 11388
rect 3235 11320 3557 11321
rect 3235 11000 3236 11320
rect 3556 11000 3557 11320
rect 3235 10999 3557 11000
rect 2816 10932 2912 10948
rect 3828 10948 3844 11372
rect 3908 10948 3924 11372
rect 4840 11372 4936 11388
rect 4247 11320 4569 11321
rect 4247 11000 4248 11320
rect 4568 11000 4569 11320
rect 4247 10999 4569 11000
rect 3828 10932 3924 10948
rect 4840 10948 4856 11372
rect 4920 10948 4936 11372
rect 5852 11372 5948 11388
rect 5259 11320 5581 11321
rect 5259 11000 5260 11320
rect 5580 11000 5581 11320
rect 5259 10999 5581 11000
rect 4840 10932 4936 10948
rect 5852 10948 5868 11372
rect 5932 10948 5948 11372
rect 6864 11372 6960 11388
rect 6271 11320 6593 11321
rect 6271 11000 6272 11320
rect 6592 11000 6593 11320
rect 6271 10999 6593 11000
rect 5852 10932 5948 10948
rect 6864 10948 6880 11372
rect 6944 10948 6960 11372
rect 7876 11372 7972 11388
rect 7283 11320 7605 11321
rect 7283 11000 7284 11320
rect 7604 11000 7605 11320
rect 7283 10999 7605 11000
rect 6864 10932 6960 10948
rect 7876 10948 7892 11372
rect 7956 10948 7972 11372
rect 8888 11372 8984 11388
rect 8295 11320 8617 11321
rect 8295 11000 8296 11320
rect 8616 11000 8617 11320
rect 8295 10999 8617 11000
rect 7876 10932 7972 10948
rect 8888 10948 8904 11372
rect 8968 10948 8984 11372
rect 9900 11372 9996 11388
rect 9307 11320 9629 11321
rect 9307 11000 9308 11320
rect 9628 11000 9629 11320
rect 9307 10999 9629 11000
rect 8888 10932 8984 10948
rect 9900 10948 9916 11372
rect 9980 10948 9996 11372
rect 10912 11372 11008 11388
rect 10319 11320 10641 11321
rect 10319 11000 10320 11320
rect 10640 11000 10641 11320
rect 10319 10999 10641 11000
rect 9900 10932 9996 10948
rect 10912 10948 10928 11372
rect 10992 10948 11008 11372
rect 11924 11372 12020 11388
rect 11331 11320 11653 11321
rect 11331 11000 11332 11320
rect 11652 11000 11653 11320
rect 11331 10999 11653 11000
rect 10912 10932 11008 10948
rect 11924 10948 11940 11372
rect 12004 10948 12020 11372
rect 12936 11372 13032 11388
rect 12343 11320 12665 11321
rect 12343 11000 12344 11320
rect 12664 11000 12665 11320
rect 12343 10999 12665 11000
rect 11924 10932 12020 10948
rect 12936 10948 12952 11372
rect 13016 10948 13032 11372
rect 13948 11372 14044 11388
rect 13355 11320 13677 11321
rect 13355 11000 13356 11320
rect 13676 11000 13677 11320
rect 13355 10999 13677 11000
rect 12936 10932 13032 10948
rect 13948 10948 13964 11372
rect 14028 10948 14044 11372
rect 14960 11372 15056 11388
rect 14367 11320 14689 11321
rect 14367 11000 14368 11320
rect 14688 11000 14689 11320
rect 14367 10999 14689 11000
rect 13948 10932 14044 10948
rect 14960 10948 14976 11372
rect 15040 10948 15056 11372
rect 15972 11372 16068 11388
rect 15379 11320 15701 11321
rect 15379 11000 15380 11320
rect 15700 11000 15701 11320
rect 15379 10999 15701 11000
rect 14960 10932 15056 10948
rect 15972 10948 15988 11372
rect 16052 10948 16068 11372
rect 16984 11372 17080 11388
rect 16391 11320 16713 11321
rect 16391 11000 16392 11320
rect 16712 11000 16713 11320
rect 16391 10999 16713 11000
rect 15972 10932 16068 10948
rect 16984 10948 17000 11372
rect 17064 10948 17080 11372
rect 16984 10932 17080 10948
rect -16412 10652 -16316 10668
rect -17005 10600 -16683 10601
rect -17005 10280 -17004 10600
rect -16684 10280 -16683 10600
rect -17005 10279 -16683 10280
rect -16412 10228 -16396 10652
rect -16332 10228 -16316 10652
rect -15400 10652 -15304 10668
rect -15993 10600 -15671 10601
rect -15993 10280 -15992 10600
rect -15672 10280 -15671 10600
rect -15993 10279 -15671 10280
rect -16412 10212 -16316 10228
rect -15400 10228 -15384 10652
rect -15320 10228 -15304 10652
rect -14388 10652 -14292 10668
rect -14981 10600 -14659 10601
rect -14981 10280 -14980 10600
rect -14660 10280 -14659 10600
rect -14981 10279 -14659 10280
rect -15400 10212 -15304 10228
rect -14388 10228 -14372 10652
rect -14308 10228 -14292 10652
rect -13376 10652 -13280 10668
rect -13969 10600 -13647 10601
rect -13969 10280 -13968 10600
rect -13648 10280 -13647 10600
rect -13969 10279 -13647 10280
rect -14388 10212 -14292 10228
rect -13376 10228 -13360 10652
rect -13296 10228 -13280 10652
rect -12364 10652 -12268 10668
rect -12957 10600 -12635 10601
rect -12957 10280 -12956 10600
rect -12636 10280 -12635 10600
rect -12957 10279 -12635 10280
rect -13376 10212 -13280 10228
rect -12364 10228 -12348 10652
rect -12284 10228 -12268 10652
rect -11352 10652 -11256 10668
rect -11945 10600 -11623 10601
rect -11945 10280 -11944 10600
rect -11624 10280 -11623 10600
rect -11945 10279 -11623 10280
rect -12364 10212 -12268 10228
rect -11352 10228 -11336 10652
rect -11272 10228 -11256 10652
rect -10340 10652 -10244 10668
rect -10933 10600 -10611 10601
rect -10933 10280 -10932 10600
rect -10612 10280 -10611 10600
rect -10933 10279 -10611 10280
rect -11352 10212 -11256 10228
rect -10340 10228 -10324 10652
rect -10260 10228 -10244 10652
rect -9328 10652 -9232 10668
rect -9921 10600 -9599 10601
rect -9921 10280 -9920 10600
rect -9600 10280 -9599 10600
rect -9921 10279 -9599 10280
rect -10340 10212 -10244 10228
rect -9328 10228 -9312 10652
rect -9248 10228 -9232 10652
rect -8316 10652 -8220 10668
rect -8909 10600 -8587 10601
rect -8909 10280 -8908 10600
rect -8588 10280 -8587 10600
rect -8909 10279 -8587 10280
rect -9328 10212 -9232 10228
rect -8316 10228 -8300 10652
rect -8236 10228 -8220 10652
rect -7304 10652 -7208 10668
rect -7897 10600 -7575 10601
rect -7897 10280 -7896 10600
rect -7576 10280 -7575 10600
rect -7897 10279 -7575 10280
rect -8316 10212 -8220 10228
rect -7304 10228 -7288 10652
rect -7224 10228 -7208 10652
rect -6292 10652 -6196 10668
rect -6885 10600 -6563 10601
rect -6885 10280 -6884 10600
rect -6564 10280 -6563 10600
rect -6885 10279 -6563 10280
rect -7304 10212 -7208 10228
rect -6292 10228 -6276 10652
rect -6212 10228 -6196 10652
rect -5280 10652 -5184 10668
rect -5873 10600 -5551 10601
rect -5873 10280 -5872 10600
rect -5552 10280 -5551 10600
rect -5873 10279 -5551 10280
rect -6292 10212 -6196 10228
rect -5280 10228 -5264 10652
rect -5200 10228 -5184 10652
rect -4268 10652 -4172 10668
rect -4861 10600 -4539 10601
rect -4861 10280 -4860 10600
rect -4540 10280 -4539 10600
rect -4861 10279 -4539 10280
rect -5280 10212 -5184 10228
rect -4268 10228 -4252 10652
rect -4188 10228 -4172 10652
rect -3256 10652 -3160 10668
rect -3849 10600 -3527 10601
rect -3849 10280 -3848 10600
rect -3528 10280 -3527 10600
rect -3849 10279 -3527 10280
rect -4268 10212 -4172 10228
rect -3256 10228 -3240 10652
rect -3176 10228 -3160 10652
rect -2244 10652 -2148 10668
rect -2837 10600 -2515 10601
rect -2837 10280 -2836 10600
rect -2516 10280 -2515 10600
rect -2837 10279 -2515 10280
rect -3256 10212 -3160 10228
rect -2244 10228 -2228 10652
rect -2164 10228 -2148 10652
rect -1232 10652 -1136 10668
rect -1825 10600 -1503 10601
rect -1825 10280 -1824 10600
rect -1504 10280 -1503 10600
rect -1825 10279 -1503 10280
rect -2244 10212 -2148 10228
rect -1232 10228 -1216 10652
rect -1152 10228 -1136 10652
rect -220 10652 -124 10668
rect -813 10600 -491 10601
rect -813 10280 -812 10600
rect -492 10280 -491 10600
rect -813 10279 -491 10280
rect -1232 10212 -1136 10228
rect -220 10228 -204 10652
rect -140 10228 -124 10652
rect 792 10652 888 10668
rect 199 10600 521 10601
rect 199 10280 200 10600
rect 520 10280 521 10600
rect 199 10279 521 10280
rect -220 10212 -124 10228
rect 792 10228 808 10652
rect 872 10228 888 10652
rect 1804 10652 1900 10668
rect 1211 10600 1533 10601
rect 1211 10280 1212 10600
rect 1532 10280 1533 10600
rect 1211 10279 1533 10280
rect 792 10212 888 10228
rect 1804 10228 1820 10652
rect 1884 10228 1900 10652
rect 2816 10652 2912 10668
rect 2223 10600 2545 10601
rect 2223 10280 2224 10600
rect 2544 10280 2545 10600
rect 2223 10279 2545 10280
rect 1804 10212 1900 10228
rect 2816 10228 2832 10652
rect 2896 10228 2912 10652
rect 3828 10652 3924 10668
rect 3235 10600 3557 10601
rect 3235 10280 3236 10600
rect 3556 10280 3557 10600
rect 3235 10279 3557 10280
rect 2816 10212 2912 10228
rect 3828 10228 3844 10652
rect 3908 10228 3924 10652
rect 4840 10652 4936 10668
rect 4247 10600 4569 10601
rect 4247 10280 4248 10600
rect 4568 10280 4569 10600
rect 4247 10279 4569 10280
rect 3828 10212 3924 10228
rect 4840 10228 4856 10652
rect 4920 10228 4936 10652
rect 5852 10652 5948 10668
rect 5259 10600 5581 10601
rect 5259 10280 5260 10600
rect 5580 10280 5581 10600
rect 5259 10279 5581 10280
rect 4840 10212 4936 10228
rect 5852 10228 5868 10652
rect 5932 10228 5948 10652
rect 6864 10652 6960 10668
rect 6271 10600 6593 10601
rect 6271 10280 6272 10600
rect 6592 10280 6593 10600
rect 6271 10279 6593 10280
rect 5852 10212 5948 10228
rect 6864 10228 6880 10652
rect 6944 10228 6960 10652
rect 7876 10652 7972 10668
rect 7283 10600 7605 10601
rect 7283 10280 7284 10600
rect 7604 10280 7605 10600
rect 7283 10279 7605 10280
rect 6864 10212 6960 10228
rect 7876 10228 7892 10652
rect 7956 10228 7972 10652
rect 8888 10652 8984 10668
rect 8295 10600 8617 10601
rect 8295 10280 8296 10600
rect 8616 10280 8617 10600
rect 8295 10279 8617 10280
rect 7876 10212 7972 10228
rect 8888 10228 8904 10652
rect 8968 10228 8984 10652
rect 9900 10652 9996 10668
rect 9307 10600 9629 10601
rect 9307 10280 9308 10600
rect 9628 10280 9629 10600
rect 9307 10279 9629 10280
rect 8888 10212 8984 10228
rect 9900 10228 9916 10652
rect 9980 10228 9996 10652
rect 10912 10652 11008 10668
rect 10319 10600 10641 10601
rect 10319 10280 10320 10600
rect 10640 10280 10641 10600
rect 10319 10279 10641 10280
rect 9900 10212 9996 10228
rect 10912 10228 10928 10652
rect 10992 10228 11008 10652
rect 11924 10652 12020 10668
rect 11331 10600 11653 10601
rect 11331 10280 11332 10600
rect 11652 10280 11653 10600
rect 11331 10279 11653 10280
rect 10912 10212 11008 10228
rect 11924 10228 11940 10652
rect 12004 10228 12020 10652
rect 12936 10652 13032 10668
rect 12343 10600 12665 10601
rect 12343 10280 12344 10600
rect 12664 10280 12665 10600
rect 12343 10279 12665 10280
rect 11924 10212 12020 10228
rect 12936 10228 12952 10652
rect 13016 10228 13032 10652
rect 13948 10652 14044 10668
rect 13355 10600 13677 10601
rect 13355 10280 13356 10600
rect 13676 10280 13677 10600
rect 13355 10279 13677 10280
rect 12936 10212 13032 10228
rect 13948 10228 13964 10652
rect 14028 10228 14044 10652
rect 14960 10652 15056 10668
rect 14367 10600 14689 10601
rect 14367 10280 14368 10600
rect 14688 10280 14689 10600
rect 14367 10279 14689 10280
rect 13948 10212 14044 10228
rect 14960 10228 14976 10652
rect 15040 10228 15056 10652
rect 15972 10652 16068 10668
rect 15379 10600 15701 10601
rect 15379 10280 15380 10600
rect 15700 10280 15701 10600
rect 15379 10279 15701 10280
rect 14960 10212 15056 10228
rect 15972 10228 15988 10652
rect 16052 10228 16068 10652
rect 16984 10652 17080 10668
rect 16391 10600 16713 10601
rect 16391 10280 16392 10600
rect 16712 10280 16713 10600
rect 16391 10279 16713 10280
rect 15972 10212 16068 10228
rect 16984 10228 17000 10652
rect 17064 10228 17080 10652
rect 16984 10212 17080 10228
rect -16412 9932 -16316 9948
rect -17005 9880 -16683 9881
rect -17005 9560 -17004 9880
rect -16684 9560 -16683 9880
rect -17005 9559 -16683 9560
rect -16412 9508 -16396 9932
rect -16332 9508 -16316 9932
rect -15400 9932 -15304 9948
rect -15993 9880 -15671 9881
rect -15993 9560 -15992 9880
rect -15672 9560 -15671 9880
rect -15993 9559 -15671 9560
rect -16412 9492 -16316 9508
rect -15400 9508 -15384 9932
rect -15320 9508 -15304 9932
rect -14388 9932 -14292 9948
rect -14981 9880 -14659 9881
rect -14981 9560 -14980 9880
rect -14660 9560 -14659 9880
rect -14981 9559 -14659 9560
rect -15400 9492 -15304 9508
rect -14388 9508 -14372 9932
rect -14308 9508 -14292 9932
rect -13376 9932 -13280 9948
rect -13969 9880 -13647 9881
rect -13969 9560 -13968 9880
rect -13648 9560 -13647 9880
rect -13969 9559 -13647 9560
rect -14388 9492 -14292 9508
rect -13376 9508 -13360 9932
rect -13296 9508 -13280 9932
rect -12364 9932 -12268 9948
rect -12957 9880 -12635 9881
rect -12957 9560 -12956 9880
rect -12636 9560 -12635 9880
rect -12957 9559 -12635 9560
rect -13376 9492 -13280 9508
rect -12364 9508 -12348 9932
rect -12284 9508 -12268 9932
rect -11352 9932 -11256 9948
rect -11945 9880 -11623 9881
rect -11945 9560 -11944 9880
rect -11624 9560 -11623 9880
rect -11945 9559 -11623 9560
rect -12364 9492 -12268 9508
rect -11352 9508 -11336 9932
rect -11272 9508 -11256 9932
rect -10340 9932 -10244 9948
rect -10933 9880 -10611 9881
rect -10933 9560 -10932 9880
rect -10612 9560 -10611 9880
rect -10933 9559 -10611 9560
rect -11352 9492 -11256 9508
rect -10340 9508 -10324 9932
rect -10260 9508 -10244 9932
rect -9328 9932 -9232 9948
rect -9921 9880 -9599 9881
rect -9921 9560 -9920 9880
rect -9600 9560 -9599 9880
rect -9921 9559 -9599 9560
rect -10340 9492 -10244 9508
rect -9328 9508 -9312 9932
rect -9248 9508 -9232 9932
rect -8316 9932 -8220 9948
rect -8909 9880 -8587 9881
rect -8909 9560 -8908 9880
rect -8588 9560 -8587 9880
rect -8909 9559 -8587 9560
rect -9328 9492 -9232 9508
rect -8316 9508 -8300 9932
rect -8236 9508 -8220 9932
rect -7304 9932 -7208 9948
rect -7897 9880 -7575 9881
rect -7897 9560 -7896 9880
rect -7576 9560 -7575 9880
rect -7897 9559 -7575 9560
rect -8316 9492 -8220 9508
rect -7304 9508 -7288 9932
rect -7224 9508 -7208 9932
rect -6292 9932 -6196 9948
rect -6885 9880 -6563 9881
rect -6885 9560 -6884 9880
rect -6564 9560 -6563 9880
rect -6885 9559 -6563 9560
rect -7304 9492 -7208 9508
rect -6292 9508 -6276 9932
rect -6212 9508 -6196 9932
rect -5280 9932 -5184 9948
rect -5873 9880 -5551 9881
rect -5873 9560 -5872 9880
rect -5552 9560 -5551 9880
rect -5873 9559 -5551 9560
rect -6292 9492 -6196 9508
rect -5280 9508 -5264 9932
rect -5200 9508 -5184 9932
rect -4268 9932 -4172 9948
rect -4861 9880 -4539 9881
rect -4861 9560 -4860 9880
rect -4540 9560 -4539 9880
rect -4861 9559 -4539 9560
rect -5280 9492 -5184 9508
rect -4268 9508 -4252 9932
rect -4188 9508 -4172 9932
rect -3256 9932 -3160 9948
rect -3849 9880 -3527 9881
rect -3849 9560 -3848 9880
rect -3528 9560 -3527 9880
rect -3849 9559 -3527 9560
rect -4268 9492 -4172 9508
rect -3256 9508 -3240 9932
rect -3176 9508 -3160 9932
rect -2244 9932 -2148 9948
rect -2837 9880 -2515 9881
rect -2837 9560 -2836 9880
rect -2516 9560 -2515 9880
rect -2837 9559 -2515 9560
rect -3256 9492 -3160 9508
rect -2244 9508 -2228 9932
rect -2164 9508 -2148 9932
rect -1232 9932 -1136 9948
rect -1825 9880 -1503 9881
rect -1825 9560 -1824 9880
rect -1504 9560 -1503 9880
rect -1825 9559 -1503 9560
rect -2244 9492 -2148 9508
rect -1232 9508 -1216 9932
rect -1152 9508 -1136 9932
rect -220 9932 -124 9948
rect -813 9880 -491 9881
rect -813 9560 -812 9880
rect -492 9560 -491 9880
rect -813 9559 -491 9560
rect -1232 9492 -1136 9508
rect -220 9508 -204 9932
rect -140 9508 -124 9932
rect 792 9932 888 9948
rect 199 9880 521 9881
rect 199 9560 200 9880
rect 520 9560 521 9880
rect 199 9559 521 9560
rect -220 9492 -124 9508
rect 792 9508 808 9932
rect 872 9508 888 9932
rect 1804 9932 1900 9948
rect 1211 9880 1533 9881
rect 1211 9560 1212 9880
rect 1532 9560 1533 9880
rect 1211 9559 1533 9560
rect 792 9492 888 9508
rect 1804 9508 1820 9932
rect 1884 9508 1900 9932
rect 2816 9932 2912 9948
rect 2223 9880 2545 9881
rect 2223 9560 2224 9880
rect 2544 9560 2545 9880
rect 2223 9559 2545 9560
rect 1804 9492 1900 9508
rect 2816 9508 2832 9932
rect 2896 9508 2912 9932
rect 3828 9932 3924 9948
rect 3235 9880 3557 9881
rect 3235 9560 3236 9880
rect 3556 9560 3557 9880
rect 3235 9559 3557 9560
rect 2816 9492 2912 9508
rect 3828 9508 3844 9932
rect 3908 9508 3924 9932
rect 4840 9932 4936 9948
rect 4247 9880 4569 9881
rect 4247 9560 4248 9880
rect 4568 9560 4569 9880
rect 4247 9559 4569 9560
rect 3828 9492 3924 9508
rect 4840 9508 4856 9932
rect 4920 9508 4936 9932
rect 5852 9932 5948 9948
rect 5259 9880 5581 9881
rect 5259 9560 5260 9880
rect 5580 9560 5581 9880
rect 5259 9559 5581 9560
rect 4840 9492 4936 9508
rect 5852 9508 5868 9932
rect 5932 9508 5948 9932
rect 6864 9932 6960 9948
rect 6271 9880 6593 9881
rect 6271 9560 6272 9880
rect 6592 9560 6593 9880
rect 6271 9559 6593 9560
rect 5852 9492 5948 9508
rect 6864 9508 6880 9932
rect 6944 9508 6960 9932
rect 7876 9932 7972 9948
rect 7283 9880 7605 9881
rect 7283 9560 7284 9880
rect 7604 9560 7605 9880
rect 7283 9559 7605 9560
rect 6864 9492 6960 9508
rect 7876 9508 7892 9932
rect 7956 9508 7972 9932
rect 8888 9932 8984 9948
rect 8295 9880 8617 9881
rect 8295 9560 8296 9880
rect 8616 9560 8617 9880
rect 8295 9559 8617 9560
rect 7876 9492 7972 9508
rect 8888 9508 8904 9932
rect 8968 9508 8984 9932
rect 9900 9932 9996 9948
rect 9307 9880 9629 9881
rect 9307 9560 9308 9880
rect 9628 9560 9629 9880
rect 9307 9559 9629 9560
rect 8888 9492 8984 9508
rect 9900 9508 9916 9932
rect 9980 9508 9996 9932
rect 10912 9932 11008 9948
rect 10319 9880 10641 9881
rect 10319 9560 10320 9880
rect 10640 9560 10641 9880
rect 10319 9559 10641 9560
rect 9900 9492 9996 9508
rect 10912 9508 10928 9932
rect 10992 9508 11008 9932
rect 11924 9932 12020 9948
rect 11331 9880 11653 9881
rect 11331 9560 11332 9880
rect 11652 9560 11653 9880
rect 11331 9559 11653 9560
rect 10912 9492 11008 9508
rect 11924 9508 11940 9932
rect 12004 9508 12020 9932
rect 12936 9932 13032 9948
rect 12343 9880 12665 9881
rect 12343 9560 12344 9880
rect 12664 9560 12665 9880
rect 12343 9559 12665 9560
rect 11924 9492 12020 9508
rect 12936 9508 12952 9932
rect 13016 9508 13032 9932
rect 13948 9932 14044 9948
rect 13355 9880 13677 9881
rect 13355 9560 13356 9880
rect 13676 9560 13677 9880
rect 13355 9559 13677 9560
rect 12936 9492 13032 9508
rect 13948 9508 13964 9932
rect 14028 9508 14044 9932
rect 14960 9932 15056 9948
rect 14367 9880 14689 9881
rect 14367 9560 14368 9880
rect 14688 9560 14689 9880
rect 14367 9559 14689 9560
rect 13948 9492 14044 9508
rect 14960 9508 14976 9932
rect 15040 9508 15056 9932
rect 15972 9932 16068 9948
rect 15379 9880 15701 9881
rect 15379 9560 15380 9880
rect 15700 9560 15701 9880
rect 15379 9559 15701 9560
rect 14960 9492 15056 9508
rect 15972 9508 15988 9932
rect 16052 9508 16068 9932
rect 16984 9932 17080 9948
rect 16391 9880 16713 9881
rect 16391 9560 16392 9880
rect 16712 9560 16713 9880
rect 16391 9559 16713 9560
rect 15972 9492 16068 9508
rect 16984 9508 17000 9932
rect 17064 9508 17080 9932
rect 16984 9492 17080 9508
rect -16412 9212 -16316 9228
rect -17005 9160 -16683 9161
rect -17005 8840 -17004 9160
rect -16684 8840 -16683 9160
rect -17005 8839 -16683 8840
rect -16412 8788 -16396 9212
rect -16332 8788 -16316 9212
rect -15400 9212 -15304 9228
rect -15993 9160 -15671 9161
rect -15993 8840 -15992 9160
rect -15672 8840 -15671 9160
rect -15993 8839 -15671 8840
rect -16412 8772 -16316 8788
rect -15400 8788 -15384 9212
rect -15320 8788 -15304 9212
rect -14388 9212 -14292 9228
rect -14981 9160 -14659 9161
rect -14981 8840 -14980 9160
rect -14660 8840 -14659 9160
rect -14981 8839 -14659 8840
rect -15400 8772 -15304 8788
rect -14388 8788 -14372 9212
rect -14308 8788 -14292 9212
rect -13376 9212 -13280 9228
rect -13969 9160 -13647 9161
rect -13969 8840 -13968 9160
rect -13648 8840 -13647 9160
rect -13969 8839 -13647 8840
rect -14388 8772 -14292 8788
rect -13376 8788 -13360 9212
rect -13296 8788 -13280 9212
rect -12364 9212 -12268 9228
rect -12957 9160 -12635 9161
rect -12957 8840 -12956 9160
rect -12636 8840 -12635 9160
rect -12957 8839 -12635 8840
rect -13376 8772 -13280 8788
rect -12364 8788 -12348 9212
rect -12284 8788 -12268 9212
rect -11352 9212 -11256 9228
rect -11945 9160 -11623 9161
rect -11945 8840 -11944 9160
rect -11624 8840 -11623 9160
rect -11945 8839 -11623 8840
rect -12364 8772 -12268 8788
rect -11352 8788 -11336 9212
rect -11272 8788 -11256 9212
rect -10340 9212 -10244 9228
rect -10933 9160 -10611 9161
rect -10933 8840 -10932 9160
rect -10612 8840 -10611 9160
rect -10933 8839 -10611 8840
rect -11352 8772 -11256 8788
rect -10340 8788 -10324 9212
rect -10260 8788 -10244 9212
rect -9328 9212 -9232 9228
rect -9921 9160 -9599 9161
rect -9921 8840 -9920 9160
rect -9600 8840 -9599 9160
rect -9921 8839 -9599 8840
rect -10340 8772 -10244 8788
rect -9328 8788 -9312 9212
rect -9248 8788 -9232 9212
rect -8316 9212 -8220 9228
rect -8909 9160 -8587 9161
rect -8909 8840 -8908 9160
rect -8588 8840 -8587 9160
rect -8909 8839 -8587 8840
rect -9328 8772 -9232 8788
rect -8316 8788 -8300 9212
rect -8236 8788 -8220 9212
rect -7304 9212 -7208 9228
rect -7897 9160 -7575 9161
rect -7897 8840 -7896 9160
rect -7576 8840 -7575 9160
rect -7897 8839 -7575 8840
rect -8316 8772 -8220 8788
rect -7304 8788 -7288 9212
rect -7224 8788 -7208 9212
rect -6292 9212 -6196 9228
rect -6885 9160 -6563 9161
rect -6885 8840 -6884 9160
rect -6564 8840 -6563 9160
rect -6885 8839 -6563 8840
rect -7304 8772 -7208 8788
rect -6292 8788 -6276 9212
rect -6212 8788 -6196 9212
rect -5280 9212 -5184 9228
rect -5873 9160 -5551 9161
rect -5873 8840 -5872 9160
rect -5552 8840 -5551 9160
rect -5873 8839 -5551 8840
rect -6292 8772 -6196 8788
rect -5280 8788 -5264 9212
rect -5200 8788 -5184 9212
rect -4268 9212 -4172 9228
rect -4861 9160 -4539 9161
rect -4861 8840 -4860 9160
rect -4540 8840 -4539 9160
rect -4861 8839 -4539 8840
rect -5280 8772 -5184 8788
rect -4268 8788 -4252 9212
rect -4188 8788 -4172 9212
rect -3256 9212 -3160 9228
rect -3849 9160 -3527 9161
rect -3849 8840 -3848 9160
rect -3528 8840 -3527 9160
rect -3849 8839 -3527 8840
rect -4268 8772 -4172 8788
rect -3256 8788 -3240 9212
rect -3176 8788 -3160 9212
rect -2244 9212 -2148 9228
rect -2837 9160 -2515 9161
rect -2837 8840 -2836 9160
rect -2516 8840 -2515 9160
rect -2837 8839 -2515 8840
rect -3256 8772 -3160 8788
rect -2244 8788 -2228 9212
rect -2164 8788 -2148 9212
rect -1232 9212 -1136 9228
rect -1825 9160 -1503 9161
rect -1825 8840 -1824 9160
rect -1504 8840 -1503 9160
rect -1825 8839 -1503 8840
rect -2244 8772 -2148 8788
rect -1232 8788 -1216 9212
rect -1152 8788 -1136 9212
rect -220 9212 -124 9228
rect -813 9160 -491 9161
rect -813 8840 -812 9160
rect -492 8840 -491 9160
rect -813 8839 -491 8840
rect -1232 8772 -1136 8788
rect -220 8788 -204 9212
rect -140 8788 -124 9212
rect 792 9212 888 9228
rect 199 9160 521 9161
rect 199 8840 200 9160
rect 520 8840 521 9160
rect 199 8839 521 8840
rect -220 8772 -124 8788
rect 792 8788 808 9212
rect 872 8788 888 9212
rect 1804 9212 1900 9228
rect 1211 9160 1533 9161
rect 1211 8840 1212 9160
rect 1532 8840 1533 9160
rect 1211 8839 1533 8840
rect 792 8772 888 8788
rect 1804 8788 1820 9212
rect 1884 8788 1900 9212
rect 2816 9212 2912 9228
rect 2223 9160 2545 9161
rect 2223 8840 2224 9160
rect 2544 8840 2545 9160
rect 2223 8839 2545 8840
rect 1804 8772 1900 8788
rect 2816 8788 2832 9212
rect 2896 8788 2912 9212
rect 3828 9212 3924 9228
rect 3235 9160 3557 9161
rect 3235 8840 3236 9160
rect 3556 8840 3557 9160
rect 3235 8839 3557 8840
rect 2816 8772 2912 8788
rect 3828 8788 3844 9212
rect 3908 8788 3924 9212
rect 4840 9212 4936 9228
rect 4247 9160 4569 9161
rect 4247 8840 4248 9160
rect 4568 8840 4569 9160
rect 4247 8839 4569 8840
rect 3828 8772 3924 8788
rect 4840 8788 4856 9212
rect 4920 8788 4936 9212
rect 5852 9212 5948 9228
rect 5259 9160 5581 9161
rect 5259 8840 5260 9160
rect 5580 8840 5581 9160
rect 5259 8839 5581 8840
rect 4840 8772 4936 8788
rect 5852 8788 5868 9212
rect 5932 8788 5948 9212
rect 6864 9212 6960 9228
rect 6271 9160 6593 9161
rect 6271 8840 6272 9160
rect 6592 8840 6593 9160
rect 6271 8839 6593 8840
rect 5852 8772 5948 8788
rect 6864 8788 6880 9212
rect 6944 8788 6960 9212
rect 7876 9212 7972 9228
rect 7283 9160 7605 9161
rect 7283 8840 7284 9160
rect 7604 8840 7605 9160
rect 7283 8839 7605 8840
rect 6864 8772 6960 8788
rect 7876 8788 7892 9212
rect 7956 8788 7972 9212
rect 8888 9212 8984 9228
rect 8295 9160 8617 9161
rect 8295 8840 8296 9160
rect 8616 8840 8617 9160
rect 8295 8839 8617 8840
rect 7876 8772 7972 8788
rect 8888 8788 8904 9212
rect 8968 8788 8984 9212
rect 9900 9212 9996 9228
rect 9307 9160 9629 9161
rect 9307 8840 9308 9160
rect 9628 8840 9629 9160
rect 9307 8839 9629 8840
rect 8888 8772 8984 8788
rect 9900 8788 9916 9212
rect 9980 8788 9996 9212
rect 10912 9212 11008 9228
rect 10319 9160 10641 9161
rect 10319 8840 10320 9160
rect 10640 8840 10641 9160
rect 10319 8839 10641 8840
rect 9900 8772 9996 8788
rect 10912 8788 10928 9212
rect 10992 8788 11008 9212
rect 11924 9212 12020 9228
rect 11331 9160 11653 9161
rect 11331 8840 11332 9160
rect 11652 8840 11653 9160
rect 11331 8839 11653 8840
rect 10912 8772 11008 8788
rect 11924 8788 11940 9212
rect 12004 8788 12020 9212
rect 12936 9212 13032 9228
rect 12343 9160 12665 9161
rect 12343 8840 12344 9160
rect 12664 8840 12665 9160
rect 12343 8839 12665 8840
rect 11924 8772 12020 8788
rect 12936 8788 12952 9212
rect 13016 8788 13032 9212
rect 13948 9212 14044 9228
rect 13355 9160 13677 9161
rect 13355 8840 13356 9160
rect 13676 8840 13677 9160
rect 13355 8839 13677 8840
rect 12936 8772 13032 8788
rect 13948 8788 13964 9212
rect 14028 8788 14044 9212
rect 14960 9212 15056 9228
rect 14367 9160 14689 9161
rect 14367 8840 14368 9160
rect 14688 8840 14689 9160
rect 14367 8839 14689 8840
rect 13948 8772 14044 8788
rect 14960 8788 14976 9212
rect 15040 8788 15056 9212
rect 15972 9212 16068 9228
rect 15379 9160 15701 9161
rect 15379 8840 15380 9160
rect 15700 8840 15701 9160
rect 15379 8839 15701 8840
rect 14960 8772 15056 8788
rect 15972 8788 15988 9212
rect 16052 8788 16068 9212
rect 16984 9212 17080 9228
rect 16391 9160 16713 9161
rect 16391 8840 16392 9160
rect 16712 8840 16713 9160
rect 16391 8839 16713 8840
rect 15972 8772 16068 8788
rect 16984 8788 17000 9212
rect 17064 8788 17080 9212
rect 16984 8772 17080 8788
rect -16412 8492 -16316 8508
rect -17005 8440 -16683 8441
rect -17005 8120 -17004 8440
rect -16684 8120 -16683 8440
rect -17005 8119 -16683 8120
rect -16412 8068 -16396 8492
rect -16332 8068 -16316 8492
rect -15400 8492 -15304 8508
rect -15993 8440 -15671 8441
rect -15993 8120 -15992 8440
rect -15672 8120 -15671 8440
rect -15993 8119 -15671 8120
rect -16412 8052 -16316 8068
rect -15400 8068 -15384 8492
rect -15320 8068 -15304 8492
rect -14388 8492 -14292 8508
rect -14981 8440 -14659 8441
rect -14981 8120 -14980 8440
rect -14660 8120 -14659 8440
rect -14981 8119 -14659 8120
rect -15400 8052 -15304 8068
rect -14388 8068 -14372 8492
rect -14308 8068 -14292 8492
rect -13376 8492 -13280 8508
rect -13969 8440 -13647 8441
rect -13969 8120 -13968 8440
rect -13648 8120 -13647 8440
rect -13969 8119 -13647 8120
rect -14388 8052 -14292 8068
rect -13376 8068 -13360 8492
rect -13296 8068 -13280 8492
rect -12364 8492 -12268 8508
rect -12957 8440 -12635 8441
rect -12957 8120 -12956 8440
rect -12636 8120 -12635 8440
rect -12957 8119 -12635 8120
rect -13376 8052 -13280 8068
rect -12364 8068 -12348 8492
rect -12284 8068 -12268 8492
rect -11352 8492 -11256 8508
rect -11945 8440 -11623 8441
rect -11945 8120 -11944 8440
rect -11624 8120 -11623 8440
rect -11945 8119 -11623 8120
rect -12364 8052 -12268 8068
rect -11352 8068 -11336 8492
rect -11272 8068 -11256 8492
rect -10340 8492 -10244 8508
rect -10933 8440 -10611 8441
rect -10933 8120 -10932 8440
rect -10612 8120 -10611 8440
rect -10933 8119 -10611 8120
rect -11352 8052 -11256 8068
rect -10340 8068 -10324 8492
rect -10260 8068 -10244 8492
rect -9328 8492 -9232 8508
rect -9921 8440 -9599 8441
rect -9921 8120 -9920 8440
rect -9600 8120 -9599 8440
rect -9921 8119 -9599 8120
rect -10340 8052 -10244 8068
rect -9328 8068 -9312 8492
rect -9248 8068 -9232 8492
rect -8316 8492 -8220 8508
rect -8909 8440 -8587 8441
rect -8909 8120 -8908 8440
rect -8588 8120 -8587 8440
rect -8909 8119 -8587 8120
rect -9328 8052 -9232 8068
rect -8316 8068 -8300 8492
rect -8236 8068 -8220 8492
rect -7304 8492 -7208 8508
rect -7897 8440 -7575 8441
rect -7897 8120 -7896 8440
rect -7576 8120 -7575 8440
rect -7897 8119 -7575 8120
rect -8316 8052 -8220 8068
rect -7304 8068 -7288 8492
rect -7224 8068 -7208 8492
rect -6292 8492 -6196 8508
rect -6885 8440 -6563 8441
rect -6885 8120 -6884 8440
rect -6564 8120 -6563 8440
rect -6885 8119 -6563 8120
rect -7304 8052 -7208 8068
rect -6292 8068 -6276 8492
rect -6212 8068 -6196 8492
rect -5280 8492 -5184 8508
rect -5873 8440 -5551 8441
rect -5873 8120 -5872 8440
rect -5552 8120 -5551 8440
rect -5873 8119 -5551 8120
rect -6292 8052 -6196 8068
rect -5280 8068 -5264 8492
rect -5200 8068 -5184 8492
rect -4268 8492 -4172 8508
rect -4861 8440 -4539 8441
rect -4861 8120 -4860 8440
rect -4540 8120 -4539 8440
rect -4861 8119 -4539 8120
rect -5280 8052 -5184 8068
rect -4268 8068 -4252 8492
rect -4188 8068 -4172 8492
rect -3256 8492 -3160 8508
rect -3849 8440 -3527 8441
rect -3849 8120 -3848 8440
rect -3528 8120 -3527 8440
rect -3849 8119 -3527 8120
rect -4268 8052 -4172 8068
rect -3256 8068 -3240 8492
rect -3176 8068 -3160 8492
rect -2244 8492 -2148 8508
rect -2837 8440 -2515 8441
rect -2837 8120 -2836 8440
rect -2516 8120 -2515 8440
rect -2837 8119 -2515 8120
rect -3256 8052 -3160 8068
rect -2244 8068 -2228 8492
rect -2164 8068 -2148 8492
rect -1232 8492 -1136 8508
rect -1825 8440 -1503 8441
rect -1825 8120 -1824 8440
rect -1504 8120 -1503 8440
rect -1825 8119 -1503 8120
rect -2244 8052 -2148 8068
rect -1232 8068 -1216 8492
rect -1152 8068 -1136 8492
rect -220 8492 -124 8508
rect -813 8440 -491 8441
rect -813 8120 -812 8440
rect -492 8120 -491 8440
rect -813 8119 -491 8120
rect -1232 8052 -1136 8068
rect -220 8068 -204 8492
rect -140 8068 -124 8492
rect 792 8492 888 8508
rect 199 8440 521 8441
rect 199 8120 200 8440
rect 520 8120 521 8440
rect 199 8119 521 8120
rect -220 8052 -124 8068
rect 792 8068 808 8492
rect 872 8068 888 8492
rect 1804 8492 1900 8508
rect 1211 8440 1533 8441
rect 1211 8120 1212 8440
rect 1532 8120 1533 8440
rect 1211 8119 1533 8120
rect 792 8052 888 8068
rect 1804 8068 1820 8492
rect 1884 8068 1900 8492
rect 2816 8492 2912 8508
rect 2223 8440 2545 8441
rect 2223 8120 2224 8440
rect 2544 8120 2545 8440
rect 2223 8119 2545 8120
rect 1804 8052 1900 8068
rect 2816 8068 2832 8492
rect 2896 8068 2912 8492
rect 3828 8492 3924 8508
rect 3235 8440 3557 8441
rect 3235 8120 3236 8440
rect 3556 8120 3557 8440
rect 3235 8119 3557 8120
rect 2816 8052 2912 8068
rect 3828 8068 3844 8492
rect 3908 8068 3924 8492
rect 4840 8492 4936 8508
rect 4247 8440 4569 8441
rect 4247 8120 4248 8440
rect 4568 8120 4569 8440
rect 4247 8119 4569 8120
rect 3828 8052 3924 8068
rect 4840 8068 4856 8492
rect 4920 8068 4936 8492
rect 5852 8492 5948 8508
rect 5259 8440 5581 8441
rect 5259 8120 5260 8440
rect 5580 8120 5581 8440
rect 5259 8119 5581 8120
rect 4840 8052 4936 8068
rect 5852 8068 5868 8492
rect 5932 8068 5948 8492
rect 6864 8492 6960 8508
rect 6271 8440 6593 8441
rect 6271 8120 6272 8440
rect 6592 8120 6593 8440
rect 6271 8119 6593 8120
rect 5852 8052 5948 8068
rect 6864 8068 6880 8492
rect 6944 8068 6960 8492
rect 7876 8492 7972 8508
rect 7283 8440 7605 8441
rect 7283 8120 7284 8440
rect 7604 8120 7605 8440
rect 7283 8119 7605 8120
rect 6864 8052 6960 8068
rect 7876 8068 7892 8492
rect 7956 8068 7972 8492
rect 8888 8492 8984 8508
rect 8295 8440 8617 8441
rect 8295 8120 8296 8440
rect 8616 8120 8617 8440
rect 8295 8119 8617 8120
rect 7876 8052 7972 8068
rect 8888 8068 8904 8492
rect 8968 8068 8984 8492
rect 9900 8492 9996 8508
rect 9307 8440 9629 8441
rect 9307 8120 9308 8440
rect 9628 8120 9629 8440
rect 9307 8119 9629 8120
rect 8888 8052 8984 8068
rect 9900 8068 9916 8492
rect 9980 8068 9996 8492
rect 10912 8492 11008 8508
rect 10319 8440 10641 8441
rect 10319 8120 10320 8440
rect 10640 8120 10641 8440
rect 10319 8119 10641 8120
rect 9900 8052 9996 8068
rect 10912 8068 10928 8492
rect 10992 8068 11008 8492
rect 11924 8492 12020 8508
rect 11331 8440 11653 8441
rect 11331 8120 11332 8440
rect 11652 8120 11653 8440
rect 11331 8119 11653 8120
rect 10912 8052 11008 8068
rect 11924 8068 11940 8492
rect 12004 8068 12020 8492
rect 12936 8492 13032 8508
rect 12343 8440 12665 8441
rect 12343 8120 12344 8440
rect 12664 8120 12665 8440
rect 12343 8119 12665 8120
rect 11924 8052 12020 8068
rect 12936 8068 12952 8492
rect 13016 8068 13032 8492
rect 13948 8492 14044 8508
rect 13355 8440 13677 8441
rect 13355 8120 13356 8440
rect 13676 8120 13677 8440
rect 13355 8119 13677 8120
rect 12936 8052 13032 8068
rect 13948 8068 13964 8492
rect 14028 8068 14044 8492
rect 14960 8492 15056 8508
rect 14367 8440 14689 8441
rect 14367 8120 14368 8440
rect 14688 8120 14689 8440
rect 14367 8119 14689 8120
rect 13948 8052 14044 8068
rect 14960 8068 14976 8492
rect 15040 8068 15056 8492
rect 15972 8492 16068 8508
rect 15379 8440 15701 8441
rect 15379 8120 15380 8440
rect 15700 8120 15701 8440
rect 15379 8119 15701 8120
rect 14960 8052 15056 8068
rect 15972 8068 15988 8492
rect 16052 8068 16068 8492
rect 16984 8492 17080 8508
rect 16391 8440 16713 8441
rect 16391 8120 16392 8440
rect 16712 8120 16713 8440
rect 16391 8119 16713 8120
rect 15972 8052 16068 8068
rect 16984 8068 17000 8492
rect 17064 8068 17080 8492
rect 16984 8052 17080 8068
rect -16412 7772 -16316 7788
rect -17005 7720 -16683 7721
rect -17005 7400 -17004 7720
rect -16684 7400 -16683 7720
rect -17005 7399 -16683 7400
rect -16412 7348 -16396 7772
rect -16332 7348 -16316 7772
rect -15400 7772 -15304 7788
rect -15993 7720 -15671 7721
rect -15993 7400 -15992 7720
rect -15672 7400 -15671 7720
rect -15993 7399 -15671 7400
rect -16412 7332 -16316 7348
rect -15400 7348 -15384 7772
rect -15320 7348 -15304 7772
rect -14388 7772 -14292 7788
rect -14981 7720 -14659 7721
rect -14981 7400 -14980 7720
rect -14660 7400 -14659 7720
rect -14981 7399 -14659 7400
rect -15400 7332 -15304 7348
rect -14388 7348 -14372 7772
rect -14308 7348 -14292 7772
rect -13376 7772 -13280 7788
rect -13969 7720 -13647 7721
rect -13969 7400 -13968 7720
rect -13648 7400 -13647 7720
rect -13969 7399 -13647 7400
rect -14388 7332 -14292 7348
rect -13376 7348 -13360 7772
rect -13296 7348 -13280 7772
rect -12364 7772 -12268 7788
rect -12957 7720 -12635 7721
rect -12957 7400 -12956 7720
rect -12636 7400 -12635 7720
rect -12957 7399 -12635 7400
rect -13376 7332 -13280 7348
rect -12364 7348 -12348 7772
rect -12284 7348 -12268 7772
rect -11352 7772 -11256 7788
rect -11945 7720 -11623 7721
rect -11945 7400 -11944 7720
rect -11624 7400 -11623 7720
rect -11945 7399 -11623 7400
rect -12364 7332 -12268 7348
rect -11352 7348 -11336 7772
rect -11272 7348 -11256 7772
rect -10340 7772 -10244 7788
rect -10933 7720 -10611 7721
rect -10933 7400 -10932 7720
rect -10612 7400 -10611 7720
rect -10933 7399 -10611 7400
rect -11352 7332 -11256 7348
rect -10340 7348 -10324 7772
rect -10260 7348 -10244 7772
rect -9328 7772 -9232 7788
rect -9921 7720 -9599 7721
rect -9921 7400 -9920 7720
rect -9600 7400 -9599 7720
rect -9921 7399 -9599 7400
rect -10340 7332 -10244 7348
rect -9328 7348 -9312 7772
rect -9248 7348 -9232 7772
rect -8316 7772 -8220 7788
rect -8909 7720 -8587 7721
rect -8909 7400 -8908 7720
rect -8588 7400 -8587 7720
rect -8909 7399 -8587 7400
rect -9328 7332 -9232 7348
rect -8316 7348 -8300 7772
rect -8236 7348 -8220 7772
rect -7304 7772 -7208 7788
rect -7897 7720 -7575 7721
rect -7897 7400 -7896 7720
rect -7576 7400 -7575 7720
rect -7897 7399 -7575 7400
rect -8316 7332 -8220 7348
rect -7304 7348 -7288 7772
rect -7224 7348 -7208 7772
rect -6292 7772 -6196 7788
rect -6885 7720 -6563 7721
rect -6885 7400 -6884 7720
rect -6564 7400 -6563 7720
rect -6885 7399 -6563 7400
rect -7304 7332 -7208 7348
rect -6292 7348 -6276 7772
rect -6212 7348 -6196 7772
rect -5280 7772 -5184 7788
rect -5873 7720 -5551 7721
rect -5873 7400 -5872 7720
rect -5552 7400 -5551 7720
rect -5873 7399 -5551 7400
rect -6292 7332 -6196 7348
rect -5280 7348 -5264 7772
rect -5200 7348 -5184 7772
rect -4268 7772 -4172 7788
rect -4861 7720 -4539 7721
rect -4861 7400 -4860 7720
rect -4540 7400 -4539 7720
rect -4861 7399 -4539 7400
rect -5280 7332 -5184 7348
rect -4268 7348 -4252 7772
rect -4188 7348 -4172 7772
rect -3256 7772 -3160 7788
rect -3849 7720 -3527 7721
rect -3849 7400 -3848 7720
rect -3528 7400 -3527 7720
rect -3849 7399 -3527 7400
rect -4268 7332 -4172 7348
rect -3256 7348 -3240 7772
rect -3176 7348 -3160 7772
rect -2244 7772 -2148 7788
rect -2837 7720 -2515 7721
rect -2837 7400 -2836 7720
rect -2516 7400 -2515 7720
rect -2837 7399 -2515 7400
rect -3256 7332 -3160 7348
rect -2244 7348 -2228 7772
rect -2164 7348 -2148 7772
rect -1232 7772 -1136 7788
rect -1825 7720 -1503 7721
rect -1825 7400 -1824 7720
rect -1504 7400 -1503 7720
rect -1825 7399 -1503 7400
rect -2244 7332 -2148 7348
rect -1232 7348 -1216 7772
rect -1152 7348 -1136 7772
rect -220 7772 -124 7788
rect -813 7720 -491 7721
rect -813 7400 -812 7720
rect -492 7400 -491 7720
rect -813 7399 -491 7400
rect -1232 7332 -1136 7348
rect -220 7348 -204 7772
rect -140 7348 -124 7772
rect 792 7772 888 7788
rect 199 7720 521 7721
rect 199 7400 200 7720
rect 520 7400 521 7720
rect 199 7399 521 7400
rect -220 7332 -124 7348
rect 792 7348 808 7772
rect 872 7348 888 7772
rect 1804 7772 1900 7788
rect 1211 7720 1533 7721
rect 1211 7400 1212 7720
rect 1532 7400 1533 7720
rect 1211 7399 1533 7400
rect 792 7332 888 7348
rect 1804 7348 1820 7772
rect 1884 7348 1900 7772
rect 2816 7772 2912 7788
rect 2223 7720 2545 7721
rect 2223 7400 2224 7720
rect 2544 7400 2545 7720
rect 2223 7399 2545 7400
rect 1804 7332 1900 7348
rect 2816 7348 2832 7772
rect 2896 7348 2912 7772
rect 3828 7772 3924 7788
rect 3235 7720 3557 7721
rect 3235 7400 3236 7720
rect 3556 7400 3557 7720
rect 3235 7399 3557 7400
rect 2816 7332 2912 7348
rect 3828 7348 3844 7772
rect 3908 7348 3924 7772
rect 4840 7772 4936 7788
rect 4247 7720 4569 7721
rect 4247 7400 4248 7720
rect 4568 7400 4569 7720
rect 4247 7399 4569 7400
rect 3828 7332 3924 7348
rect 4840 7348 4856 7772
rect 4920 7348 4936 7772
rect 5852 7772 5948 7788
rect 5259 7720 5581 7721
rect 5259 7400 5260 7720
rect 5580 7400 5581 7720
rect 5259 7399 5581 7400
rect 4840 7332 4936 7348
rect 5852 7348 5868 7772
rect 5932 7348 5948 7772
rect 6864 7772 6960 7788
rect 6271 7720 6593 7721
rect 6271 7400 6272 7720
rect 6592 7400 6593 7720
rect 6271 7399 6593 7400
rect 5852 7332 5948 7348
rect 6864 7348 6880 7772
rect 6944 7348 6960 7772
rect 7876 7772 7972 7788
rect 7283 7720 7605 7721
rect 7283 7400 7284 7720
rect 7604 7400 7605 7720
rect 7283 7399 7605 7400
rect 6864 7332 6960 7348
rect 7876 7348 7892 7772
rect 7956 7348 7972 7772
rect 8888 7772 8984 7788
rect 8295 7720 8617 7721
rect 8295 7400 8296 7720
rect 8616 7400 8617 7720
rect 8295 7399 8617 7400
rect 7876 7332 7972 7348
rect 8888 7348 8904 7772
rect 8968 7348 8984 7772
rect 9900 7772 9996 7788
rect 9307 7720 9629 7721
rect 9307 7400 9308 7720
rect 9628 7400 9629 7720
rect 9307 7399 9629 7400
rect 8888 7332 8984 7348
rect 9900 7348 9916 7772
rect 9980 7348 9996 7772
rect 10912 7772 11008 7788
rect 10319 7720 10641 7721
rect 10319 7400 10320 7720
rect 10640 7400 10641 7720
rect 10319 7399 10641 7400
rect 9900 7332 9996 7348
rect 10912 7348 10928 7772
rect 10992 7348 11008 7772
rect 11924 7772 12020 7788
rect 11331 7720 11653 7721
rect 11331 7400 11332 7720
rect 11652 7400 11653 7720
rect 11331 7399 11653 7400
rect 10912 7332 11008 7348
rect 11924 7348 11940 7772
rect 12004 7348 12020 7772
rect 12936 7772 13032 7788
rect 12343 7720 12665 7721
rect 12343 7400 12344 7720
rect 12664 7400 12665 7720
rect 12343 7399 12665 7400
rect 11924 7332 12020 7348
rect 12936 7348 12952 7772
rect 13016 7348 13032 7772
rect 13948 7772 14044 7788
rect 13355 7720 13677 7721
rect 13355 7400 13356 7720
rect 13676 7400 13677 7720
rect 13355 7399 13677 7400
rect 12936 7332 13032 7348
rect 13948 7348 13964 7772
rect 14028 7348 14044 7772
rect 14960 7772 15056 7788
rect 14367 7720 14689 7721
rect 14367 7400 14368 7720
rect 14688 7400 14689 7720
rect 14367 7399 14689 7400
rect 13948 7332 14044 7348
rect 14960 7348 14976 7772
rect 15040 7348 15056 7772
rect 15972 7772 16068 7788
rect 15379 7720 15701 7721
rect 15379 7400 15380 7720
rect 15700 7400 15701 7720
rect 15379 7399 15701 7400
rect 14960 7332 15056 7348
rect 15972 7348 15988 7772
rect 16052 7348 16068 7772
rect 16984 7772 17080 7788
rect 16391 7720 16713 7721
rect 16391 7400 16392 7720
rect 16712 7400 16713 7720
rect 16391 7399 16713 7400
rect 15972 7332 16068 7348
rect 16984 7348 17000 7772
rect 17064 7348 17080 7772
rect 16984 7332 17080 7348
rect -16412 7052 -16316 7068
rect -17005 7000 -16683 7001
rect -17005 6680 -17004 7000
rect -16684 6680 -16683 7000
rect -17005 6679 -16683 6680
rect -16412 6628 -16396 7052
rect -16332 6628 -16316 7052
rect -15400 7052 -15304 7068
rect -15993 7000 -15671 7001
rect -15993 6680 -15992 7000
rect -15672 6680 -15671 7000
rect -15993 6679 -15671 6680
rect -16412 6612 -16316 6628
rect -15400 6628 -15384 7052
rect -15320 6628 -15304 7052
rect -14388 7052 -14292 7068
rect -14981 7000 -14659 7001
rect -14981 6680 -14980 7000
rect -14660 6680 -14659 7000
rect -14981 6679 -14659 6680
rect -15400 6612 -15304 6628
rect -14388 6628 -14372 7052
rect -14308 6628 -14292 7052
rect -13376 7052 -13280 7068
rect -13969 7000 -13647 7001
rect -13969 6680 -13968 7000
rect -13648 6680 -13647 7000
rect -13969 6679 -13647 6680
rect -14388 6612 -14292 6628
rect -13376 6628 -13360 7052
rect -13296 6628 -13280 7052
rect -12364 7052 -12268 7068
rect -12957 7000 -12635 7001
rect -12957 6680 -12956 7000
rect -12636 6680 -12635 7000
rect -12957 6679 -12635 6680
rect -13376 6612 -13280 6628
rect -12364 6628 -12348 7052
rect -12284 6628 -12268 7052
rect -11352 7052 -11256 7068
rect -11945 7000 -11623 7001
rect -11945 6680 -11944 7000
rect -11624 6680 -11623 7000
rect -11945 6679 -11623 6680
rect -12364 6612 -12268 6628
rect -11352 6628 -11336 7052
rect -11272 6628 -11256 7052
rect -10340 7052 -10244 7068
rect -10933 7000 -10611 7001
rect -10933 6680 -10932 7000
rect -10612 6680 -10611 7000
rect -10933 6679 -10611 6680
rect -11352 6612 -11256 6628
rect -10340 6628 -10324 7052
rect -10260 6628 -10244 7052
rect -9328 7052 -9232 7068
rect -9921 7000 -9599 7001
rect -9921 6680 -9920 7000
rect -9600 6680 -9599 7000
rect -9921 6679 -9599 6680
rect -10340 6612 -10244 6628
rect -9328 6628 -9312 7052
rect -9248 6628 -9232 7052
rect -8316 7052 -8220 7068
rect -8909 7000 -8587 7001
rect -8909 6680 -8908 7000
rect -8588 6680 -8587 7000
rect -8909 6679 -8587 6680
rect -9328 6612 -9232 6628
rect -8316 6628 -8300 7052
rect -8236 6628 -8220 7052
rect -7304 7052 -7208 7068
rect -7897 7000 -7575 7001
rect -7897 6680 -7896 7000
rect -7576 6680 -7575 7000
rect -7897 6679 -7575 6680
rect -8316 6612 -8220 6628
rect -7304 6628 -7288 7052
rect -7224 6628 -7208 7052
rect -6292 7052 -6196 7068
rect -6885 7000 -6563 7001
rect -6885 6680 -6884 7000
rect -6564 6680 -6563 7000
rect -6885 6679 -6563 6680
rect -7304 6612 -7208 6628
rect -6292 6628 -6276 7052
rect -6212 6628 -6196 7052
rect -5280 7052 -5184 7068
rect -5873 7000 -5551 7001
rect -5873 6680 -5872 7000
rect -5552 6680 -5551 7000
rect -5873 6679 -5551 6680
rect -6292 6612 -6196 6628
rect -5280 6628 -5264 7052
rect -5200 6628 -5184 7052
rect -4268 7052 -4172 7068
rect -4861 7000 -4539 7001
rect -4861 6680 -4860 7000
rect -4540 6680 -4539 7000
rect -4861 6679 -4539 6680
rect -5280 6612 -5184 6628
rect -4268 6628 -4252 7052
rect -4188 6628 -4172 7052
rect -3256 7052 -3160 7068
rect -3849 7000 -3527 7001
rect -3849 6680 -3848 7000
rect -3528 6680 -3527 7000
rect -3849 6679 -3527 6680
rect -4268 6612 -4172 6628
rect -3256 6628 -3240 7052
rect -3176 6628 -3160 7052
rect -2244 7052 -2148 7068
rect -2837 7000 -2515 7001
rect -2837 6680 -2836 7000
rect -2516 6680 -2515 7000
rect -2837 6679 -2515 6680
rect -3256 6612 -3160 6628
rect -2244 6628 -2228 7052
rect -2164 6628 -2148 7052
rect -1232 7052 -1136 7068
rect -1825 7000 -1503 7001
rect -1825 6680 -1824 7000
rect -1504 6680 -1503 7000
rect -1825 6679 -1503 6680
rect -2244 6612 -2148 6628
rect -1232 6628 -1216 7052
rect -1152 6628 -1136 7052
rect -220 7052 -124 7068
rect -813 7000 -491 7001
rect -813 6680 -812 7000
rect -492 6680 -491 7000
rect -813 6679 -491 6680
rect -1232 6612 -1136 6628
rect -220 6628 -204 7052
rect -140 6628 -124 7052
rect 792 7052 888 7068
rect 199 7000 521 7001
rect 199 6680 200 7000
rect 520 6680 521 7000
rect 199 6679 521 6680
rect -220 6612 -124 6628
rect 792 6628 808 7052
rect 872 6628 888 7052
rect 1804 7052 1900 7068
rect 1211 7000 1533 7001
rect 1211 6680 1212 7000
rect 1532 6680 1533 7000
rect 1211 6679 1533 6680
rect 792 6612 888 6628
rect 1804 6628 1820 7052
rect 1884 6628 1900 7052
rect 2816 7052 2912 7068
rect 2223 7000 2545 7001
rect 2223 6680 2224 7000
rect 2544 6680 2545 7000
rect 2223 6679 2545 6680
rect 1804 6612 1900 6628
rect 2816 6628 2832 7052
rect 2896 6628 2912 7052
rect 3828 7052 3924 7068
rect 3235 7000 3557 7001
rect 3235 6680 3236 7000
rect 3556 6680 3557 7000
rect 3235 6679 3557 6680
rect 2816 6612 2912 6628
rect 3828 6628 3844 7052
rect 3908 6628 3924 7052
rect 4840 7052 4936 7068
rect 4247 7000 4569 7001
rect 4247 6680 4248 7000
rect 4568 6680 4569 7000
rect 4247 6679 4569 6680
rect 3828 6612 3924 6628
rect 4840 6628 4856 7052
rect 4920 6628 4936 7052
rect 5852 7052 5948 7068
rect 5259 7000 5581 7001
rect 5259 6680 5260 7000
rect 5580 6680 5581 7000
rect 5259 6679 5581 6680
rect 4840 6612 4936 6628
rect 5852 6628 5868 7052
rect 5932 6628 5948 7052
rect 6864 7052 6960 7068
rect 6271 7000 6593 7001
rect 6271 6680 6272 7000
rect 6592 6680 6593 7000
rect 6271 6679 6593 6680
rect 5852 6612 5948 6628
rect 6864 6628 6880 7052
rect 6944 6628 6960 7052
rect 7876 7052 7972 7068
rect 7283 7000 7605 7001
rect 7283 6680 7284 7000
rect 7604 6680 7605 7000
rect 7283 6679 7605 6680
rect 6864 6612 6960 6628
rect 7876 6628 7892 7052
rect 7956 6628 7972 7052
rect 8888 7052 8984 7068
rect 8295 7000 8617 7001
rect 8295 6680 8296 7000
rect 8616 6680 8617 7000
rect 8295 6679 8617 6680
rect 7876 6612 7972 6628
rect 8888 6628 8904 7052
rect 8968 6628 8984 7052
rect 9900 7052 9996 7068
rect 9307 7000 9629 7001
rect 9307 6680 9308 7000
rect 9628 6680 9629 7000
rect 9307 6679 9629 6680
rect 8888 6612 8984 6628
rect 9900 6628 9916 7052
rect 9980 6628 9996 7052
rect 10912 7052 11008 7068
rect 10319 7000 10641 7001
rect 10319 6680 10320 7000
rect 10640 6680 10641 7000
rect 10319 6679 10641 6680
rect 9900 6612 9996 6628
rect 10912 6628 10928 7052
rect 10992 6628 11008 7052
rect 11924 7052 12020 7068
rect 11331 7000 11653 7001
rect 11331 6680 11332 7000
rect 11652 6680 11653 7000
rect 11331 6679 11653 6680
rect 10912 6612 11008 6628
rect 11924 6628 11940 7052
rect 12004 6628 12020 7052
rect 12936 7052 13032 7068
rect 12343 7000 12665 7001
rect 12343 6680 12344 7000
rect 12664 6680 12665 7000
rect 12343 6679 12665 6680
rect 11924 6612 12020 6628
rect 12936 6628 12952 7052
rect 13016 6628 13032 7052
rect 13948 7052 14044 7068
rect 13355 7000 13677 7001
rect 13355 6680 13356 7000
rect 13676 6680 13677 7000
rect 13355 6679 13677 6680
rect 12936 6612 13032 6628
rect 13948 6628 13964 7052
rect 14028 6628 14044 7052
rect 14960 7052 15056 7068
rect 14367 7000 14689 7001
rect 14367 6680 14368 7000
rect 14688 6680 14689 7000
rect 14367 6679 14689 6680
rect 13948 6612 14044 6628
rect 14960 6628 14976 7052
rect 15040 6628 15056 7052
rect 15972 7052 16068 7068
rect 15379 7000 15701 7001
rect 15379 6680 15380 7000
rect 15700 6680 15701 7000
rect 15379 6679 15701 6680
rect 14960 6612 15056 6628
rect 15972 6628 15988 7052
rect 16052 6628 16068 7052
rect 16984 7052 17080 7068
rect 16391 7000 16713 7001
rect 16391 6680 16392 7000
rect 16712 6680 16713 7000
rect 16391 6679 16713 6680
rect 15972 6612 16068 6628
rect 16984 6628 17000 7052
rect 17064 6628 17080 7052
rect 16984 6612 17080 6628
rect -16412 6332 -16316 6348
rect -17005 6280 -16683 6281
rect -17005 5960 -17004 6280
rect -16684 5960 -16683 6280
rect -17005 5959 -16683 5960
rect -16412 5908 -16396 6332
rect -16332 5908 -16316 6332
rect -15400 6332 -15304 6348
rect -15993 6280 -15671 6281
rect -15993 5960 -15992 6280
rect -15672 5960 -15671 6280
rect -15993 5959 -15671 5960
rect -16412 5892 -16316 5908
rect -15400 5908 -15384 6332
rect -15320 5908 -15304 6332
rect -14388 6332 -14292 6348
rect -14981 6280 -14659 6281
rect -14981 5960 -14980 6280
rect -14660 5960 -14659 6280
rect -14981 5959 -14659 5960
rect -15400 5892 -15304 5908
rect -14388 5908 -14372 6332
rect -14308 5908 -14292 6332
rect -13376 6332 -13280 6348
rect -13969 6280 -13647 6281
rect -13969 5960 -13968 6280
rect -13648 5960 -13647 6280
rect -13969 5959 -13647 5960
rect -14388 5892 -14292 5908
rect -13376 5908 -13360 6332
rect -13296 5908 -13280 6332
rect -12364 6332 -12268 6348
rect -12957 6280 -12635 6281
rect -12957 5960 -12956 6280
rect -12636 5960 -12635 6280
rect -12957 5959 -12635 5960
rect -13376 5892 -13280 5908
rect -12364 5908 -12348 6332
rect -12284 5908 -12268 6332
rect -11352 6332 -11256 6348
rect -11945 6280 -11623 6281
rect -11945 5960 -11944 6280
rect -11624 5960 -11623 6280
rect -11945 5959 -11623 5960
rect -12364 5892 -12268 5908
rect -11352 5908 -11336 6332
rect -11272 5908 -11256 6332
rect -10340 6332 -10244 6348
rect -10933 6280 -10611 6281
rect -10933 5960 -10932 6280
rect -10612 5960 -10611 6280
rect -10933 5959 -10611 5960
rect -11352 5892 -11256 5908
rect -10340 5908 -10324 6332
rect -10260 5908 -10244 6332
rect -9328 6332 -9232 6348
rect -9921 6280 -9599 6281
rect -9921 5960 -9920 6280
rect -9600 5960 -9599 6280
rect -9921 5959 -9599 5960
rect -10340 5892 -10244 5908
rect -9328 5908 -9312 6332
rect -9248 5908 -9232 6332
rect -8316 6332 -8220 6348
rect -8909 6280 -8587 6281
rect -8909 5960 -8908 6280
rect -8588 5960 -8587 6280
rect -8909 5959 -8587 5960
rect -9328 5892 -9232 5908
rect -8316 5908 -8300 6332
rect -8236 5908 -8220 6332
rect -7304 6332 -7208 6348
rect -7897 6280 -7575 6281
rect -7897 5960 -7896 6280
rect -7576 5960 -7575 6280
rect -7897 5959 -7575 5960
rect -8316 5892 -8220 5908
rect -7304 5908 -7288 6332
rect -7224 5908 -7208 6332
rect -6292 6332 -6196 6348
rect -6885 6280 -6563 6281
rect -6885 5960 -6884 6280
rect -6564 5960 -6563 6280
rect -6885 5959 -6563 5960
rect -7304 5892 -7208 5908
rect -6292 5908 -6276 6332
rect -6212 5908 -6196 6332
rect -5280 6332 -5184 6348
rect -5873 6280 -5551 6281
rect -5873 5960 -5872 6280
rect -5552 5960 -5551 6280
rect -5873 5959 -5551 5960
rect -6292 5892 -6196 5908
rect -5280 5908 -5264 6332
rect -5200 5908 -5184 6332
rect -4268 6332 -4172 6348
rect -4861 6280 -4539 6281
rect -4861 5960 -4860 6280
rect -4540 5960 -4539 6280
rect -4861 5959 -4539 5960
rect -5280 5892 -5184 5908
rect -4268 5908 -4252 6332
rect -4188 5908 -4172 6332
rect -3256 6332 -3160 6348
rect -3849 6280 -3527 6281
rect -3849 5960 -3848 6280
rect -3528 5960 -3527 6280
rect -3849 5959 -3527 5960
rect -4268 5892 -4172 5908
rect -3256 5908 -3240 6332
rect -3176 5908 -3160 6332
rect -2244 6332 -2148 6348
rect -2837 6280 -2515 6281
rect -2837 5960 -2836 6280
rect -2516 5960 -2515 6280
rect -2837 5959 -2515 5960
rect -3256 5892 -3160 5908
rect -2244 5908 -2228 6332
rect -2164 5908 -2148 6332
rect -1232 6332 -1136 6348
rect -1825 6280 -1503 6281
rect -1825 5960 -1824 6280
rect -1504 5960 -1503 6280
rect -1825 5959 -1503 5960
rect -2244 5892 -2148 5908
rect -1232 5908 -1216 6332
rect -1152 5908 -1136 6332
rect -220 6332 -124 6348
rect -813 6280 -491 6281
rect -813 5960 -812 6280
rect -492 5960 -491 6280
rect -813 5959 -491 5960
rect -1232 5892 -1136 5908
rect -220 5908 -204 6332
rect -140 5908 -124 6332
rect 792 6332 888 6348
rect 199 6280 521 6281
rect 199 5960 200 6280
rect 520 5960 521 6280
rect 199 5959 521 5960
rect -220 5892 -124 5908
rect 792 5908 808 6332
rect 872 5908 888 6332
rect 1804 6332 1900 6348
rect 1211 6280 1533 6281
rect 1211 5960 1212 6280
rect 1532 5960 1533 6280
rect 1211 5959 1533 5960
rect 792 5892 888 5908
rect 1804 5908 1820 6332
rect 1884 5908 1900 6332
rect 2816 6332 2912 6348
rect 2223 6280 2545 6281
rect 2223 5960 2224 6280
rect 2544 5960 2545 6280
rect 2223 5959 2545 5960
rect 1804 5892 1900 5908
rect 2816 5908 2832 6332
rect 2896 5908 2912 6332
rect 3828 6332 3924 6348
rect 3235 6280 3557 6281
rect 3235 5960 3236 6280
rect 3556 5960 3557 6280
rect 3235 5959 3557 5960
rect 2816 5892 2912 5908
rect 3828 5908 3844 6332
rect 3908 5908 3924 6332
rect 4840 6332 4936 6348
rect 4247 6280 4569 6281
rect 4247 5960 4248 6280
rect 4568 5960 4569 6280
rect 4247 5959 4569 5960
rect 3828 5892 3924 5908
rect 4840 5908 4856 6332
rect 4920 5908 4936 6332
rect 5852 6332 5948 6348
rect 5259 6280 5581 6281
rect 5259 5960 5260 6280
rect 5580 5960 5581 6280
rect 5259 5959 5581 5960
rect 4840 5892 4936 5908
rect 5852 5908 5868 6332
rect 5932 5908 5948 6332
rect 6864 6332 6960 6348
rect 6271 6280 6593 6281
rect 6271 5960 6272 6280
rect 6592 5960 6593 6280
rect 6271 5959 6593 5960
rect 5852 5892 5948 5908
rect 6864 5908 6880 6332
rect 6944 5908 6960 6332
rect 7876 6332 7972 6348
rect 7283 6280 7605 6281
rect 7283 5960 7284 6280
rect 7604 5960 7605 6280
rect 7283 5959 7605 5960
rect 6864 5892 6960 5908
rect 7876 5908 7892 6332
rect 7956 5908 7972 6332
rect 8888 6332 8984 6348
rect 8295 6280 8617 6281
rect 8295 5960 8296 6280
rect 8616 5960 8617 6280
rect 8295 5959 8617 5960
rect 7876 5892 7972 5908
rect 8888 5908 8904 6332
rect 8968 5908 8984 6332
rect 9900 6332 9996 6348
rect 9307 6280 9629 6281
rect 9307 5960 9308 6280
rect 9628 5960 9629 6280
rect 9307 5959 9629 5960
rect 8888 5892 8984 5908
rect 9900 5908 9916 6332
rect 9980 5908 9996 6332
rect 10912 6332 11008 6348
rect 10319 6280 10641 6281
rect 10319 5960 10320 6280
rect 10640 5960 10641 6280
rect 10319 5959 10641 5960
rect 9900 5892 9996 5908
rect 10912 5908 10928 6332
rect 10992 5908 11008 6332
rect 11924 6332 12020 6348
rect 11331 6280 11653 6281
rect 11331 5960 11332 6280
rect 11652 5960 11653 6280
rect 11331 5959 11653 5960
rect 10912 5892 11008 5908
rect 11924 5908 11940 6332
rect 12004 5908 12020 6332
rect 12936 6332 13032 6348
rect 12343 6280 12665 6281
rect 12343 5960 12344 6280
rect 12664 5960 12665 6280
rect 12343 5959 12665 5960
rect 11924 5892 12020 5908
rect 12936 5908 12952 6332
rect 13016 5908 13032 6332
rect 13948 6332 14044 6348
rect 13355 6280 13677 6281
rect 13355 5960 13356 6280
rect 13676 5960 13677 6280
rect 13355 5959 13677 5960
rect 12936 5892 13032 5908
rect 13948 5908 13964 6332
rect 14028 5908 14044 6332
rect 14960 6332 15056 6348
rect 14367 6280 14689 6281
rect 14367 5960 14368 6280
rect 14688 5960 14689 6280
rect 14367 5959 14689 5960
rect 13948 5892 14044 5908
rect 14960 5908 14976 6332
rect 15040 5908 15056 6332
rect 15972 6332 16068 6348
rect 15379 6280 15701 6281
rect 15379 5960 15380 6280
rect 15700 5960 15701 6280
rect 15379 5959 15701 5960
rect 14960 5892 15056 5908
rect 15972 5908 15988 6332
rect 16052 5908 16068 6332
rect 16984 6332 17080 6348
rect 16391 6280 16713 6281
rect 16391 5960 16392 6280
rect 16712 5960 16713 6280
rect 16391 5959 16713 5960
rect 15972 5892 16068 5908
rect 16984 5908 17000 6332
rect 17064 5908 17080 6332
rect 16984 5892 17080 5908
rect -16412 5612 -16316 5628
rect -17005 5560 -16683 5561
rect -17005 5240 -17004 5560
rect -16684 5240 -16683 5560
rect -17005 5239 -16683 5240
rect -16412 5188 -16396 5612
rect -16332 5188 -16316 5612
rect -15400 5612 -15304 5628
rect -15993 5560 -15671 5561
rect -15993 5240 -15992 5560
rect -15672 5240 -15671 5560
rect -15993 5239 -15671 5240
rect -16412 5172 -16316 5188
rect -15400 5188 -15384 5612
rect -15320 5188 -15304 5612
rect -14388 5612 -14292 5628
rect -14981 5560 -14659 5561
rect -14981 5240 -14980 5560
rect -14660 5240 -14659 5560
rect -14981 5239 -14659 5240
rect -15400 5172 -15304 5188
rect -14388 5188 -14372 5612
rect -14308 5188 -14292 5612
rect -13376 5612 -13280 5628
rect -13969 5560 -13647 5561
rect -13969 5240 -13968 5560
rect -13648 5240 -13647 5560
rect -13969 5239 -13647 5240
rect -14388 5172 -14292 5188
rect -13376 5188 -13360 5612
rect -13296 5188 -13280 5612
rect -12364 5612 -12268 5628
rect -12957 5560 -12635 5561
rect -12957 5240 -12956 5560
rect -12636 5240 -12635 5560
rect -12957 5239 -12635 5240
rect -13376 5172 -13280 5188
rect -12364 5188 -12348 5612
rect -12284 5188 -12268 5612
rect -11352 5612 -11256 5628
rect -11945 5560 -11623 5561
rect -11945 5240 -11944 5560
rect -11624 5240 -11623 5560
rect -11945 5239 -11623 5240
rect -12364 5172 -12268 5188
rect -11352 5188 -11336 5612
rect -11272 5188 -11256 5612
rect -10340 5612 -10244 5628
rect -10933 5560 -10611 5561
rect -10933 5240 -10932 5560
rect -10612 5240 -10611 5560
rect -10933 5239 -10611 5240
rect -11352 5172 -11256 5188
rect -10340 5188 -10324 5612
rect -10260 5188 -10244 5612
rect -9328 5612 -9232 5628
rect -9921 5560 -9599 5561
rect -9921 5240 -9920 5560
rect -9600 5240 -9599 5560
rect -9921 5239 -9599 5240
rect -10340 5172 -10244 5188
rect -9328 5188 -9312 5612
rect -9248 5188 -9232 5612
rect -8316 5612 -8220 5628
rect -8909 5560 -8587 5561
rect -8909 5240 -8908 5560
rect -8588 5240 -8587 5560
rect -8909 5239 -8587 5240
rect -9328 5172 -9232 5188
rect -8316 5188 -8300 5612
rect -8236 5188 -8220 5612
rect -7304 5612 -7208 5628
rect -7897 5560 -7575 5561
rect -7897 5240 -7896 5560
rect -7576 5240 -7575 5560
rect -7897 5239 -7575 5240
rect -8316 5172 -8220 5188
rect -7304 5188 -7288 5612
rect -7224 5188 -7208 5612
rect -6292 5612 -6196 5628
rect -6885 5560 -6563 5561
rect -6885 5240 -6884 5560
rect -6564 5240 -6563 5560
rect -6885 5239 -6563 5240
rect -7304 5172 -7208 5188
rect -6292 5188 -6276 5612
rect -6212 5188 -6196 5612
rect -5280 5612 -5184 5628
rect -5873 5560 -5551 5561
rect -5873 5240 -5872 5560
rect -5552 5240 -5551 5560
rect -5873 5239 -5551 5240
rect -6292 5172 -6196 5188
rect -5280 5188 -5264 5612
rect -5200 5188 -5184 5612
rect -4268 5612 -4172 5628
rect -4861 5560 -4539 5561
rect -4861 5240 -4860 5560
rect -4540 5240 -4539 5560
rect -4861 5239 -4539 5240
rect -5280 5172 -5184 5188
rect -4268 5188 -4252 5612
rect -4188 5188 -4172 5612
rect -3256 5612 -3160 5628
rect -3849 5560 -3527 5561
rect -3849 5240 -3848 5560
rect -3528 5240 -3527 5560
rect -3849 5239 -3527 5240
rect -4268 5172 -4172 5188
rect -3256 5188 -3240 5612
rect -3176 5188 -3160 5612
rect -2244 5612 -2148 5628
rect -2837 5560 -2515 5561
rect -2837 5240 -2836 5560
rect -2516 5240 -2515 5560
rect -2837 5239 -2515 5240
rect -3256 5172 -3160 5188
rect -2244 5188 -2228 5612
rect -2164 5188 -2148 5612
rect -1232 5612 -1136 5628
rect -1825 5560 -1503 5561
rect -1825 5240 -1824 5560
rect -1504 5240 -1503 5560
rect -1825 5239 -1503 5240
rect -2244 5172 -2148 5188
rect -1232 5188 -1216 5612
rect -1152 5188 -1136 5612
rect -220 5612 -124 5628
rect -813 5560 -491 5561
rect -813 5240 -812 5560
rect -492 5240 -491 5560
rect -813 5239 -491 5240
rect -1232 5172 -1136 5188
rect -220 5188 -204 5612
rect -140 5188 -124 5612
rect 792 5612 888 5628
rect 199 5560 521 5561
rect 199 5240 200 5560
rect 520 5240 521 5560
rect 199 5239 521 5240
rect -220 5172 -124 5188
rect 792 5188 808 5612
rect 872 5188 888 5612
rect 1804 5612 1900 5628
rect 1211 5560 1533 5561
rect 1211 5240 1212 5560
rect 1532 5240 1533 5560
rect 1211 5239 1533 5240
rect 792 5172 888 5188
rect 1804 5188 1820 5612
rect 1884 5188 1900 5612
rect 2816 5612 2912 5628
rect 2223 5560 2545 5561
rect 2223 5240 2224 5560
rect 2544 5240 2545 5560
rect 2223 5239 2545 5240
rect 1804 5172 1900 5188
rect 2816 5188 2832 5612
rect 2896 5188 2912 5612
rect 3828 5612 3924 5628
rect 3235 5560 3557 5561
rect 3235 5240 3236 5560
rect 3556 5240 3557 5560
rect 3235 5239 3557 5240
rect 2816 5172 2912 5188
rect 3828 5188 3844 5612
rect 3908 5188 3924 5612
rect 4840 5612 4936 5628
rect 4247 5560 4569 5561
rect 4247 5240 4248 5560
rect 4568 5240 4569 5560
rect 4247 5239 4569 5240
rect 3828 5172 3924 5188
rect 4840 5188 4856 5612
rect 4920 5188 4936 5612
rect 5852 5612 5948 5628
rect 5259 5560 5581 5561
rect 5259 5240 5260 5560
rect 5580 5240 5581 5560
rect 5259 5239 5581 5240
rect 4840 5172 4936 5188
rect 5852 5188 5868 5612
rect 5932 5188 5948 5612
rect 6864 5612 6960 5628
rect 6271 5560 6593 5561
rect 6271 5240 6272 5560
rect 6592 5240 6593 5560
rect 6271 5239 6593 5240
rect 5852 5172 5948 5188
rect 6864 5188 6880 5612
rect 6944 5188 6960 5612
rect 7876 5612 7972 5628
rect 7283 5560 7605 5561
rect 7283 5240 7284 5560
rect 7604 5240 7605 5560
rect 7283 5239 7605 5240
rect 6864 5172 6960 5188
rect 7876 5188 7892 5612
rect 7956 5188 7972 5612
rect 8888 5612 8984 5628
rect 8295 5560 8617 5561
rect 8295 5240 8296 5560
rect 8616 5240 8617 5560
rect 8295 5239 8617 5240
rect 7876 5172 7972 5188
rect 8888 5188 8904 5612
rect 8968 5188 8984 5612
rect 9900 5612 9996 5628
rect 9307 5560 9629 5561
rect 9307 5240 9308 5560
rect 9628 5240 9629 5560
rect 9307 5239 9629 5240
rect 8888 5172 8984 5188
rect 9900 5188 9916 5612
rect 9980 5188 9996 5612
rect 10912 5612 11008 5628
rect 10319 5560 10641 5561
rect 10319 5240 10320 5560
rect 10640 5240 10641 5560
rect 10319 5239 10641 5240
rect 9900 5172 9996 5188
rect 10912 5188 10928 5612
rect 10992 5188 11008 5612
rect 11924 5612 12020 5628
rect 11331 5560 11653 5561
rect 11331 5240 11332 5560
rect 11652 5240 11653 5560
rect 11331 5239 11653 5240
rect 10912 5172 11008 5188
rect 11924 5188 11940 5612
rect 12004 5188 12020 5612
rect 12936 5612 13032 5628
rect 12343 5560 12665 5561
rect 12343 5240 12344 5560
rect 12664 5240 12665 5560
rect 12343 5239 12665 5240
rect 11924 5172 12020 5188
rect 12936 5188 12952 5612
rect 13016 5188 13032 5612
rect 13948 5612 14044 5628
rect 13355 5560 13677 5561
rect 13355 5240 13356 5560
rect 13676 5240 13677 5560
rect 13355 5239 13677 5240
rect 12936 5172 13032 5188
rect 13948 5188 13964 5612
rect 14028 5188 14044 5612
rect 14960 5612 15056 5628
rect 14367 5560 14689 5561
rect 14367 5240 14368 5560
rect 14688 5240 14689 5560
rect 14367 5239 14689 5240
rect 13948 5172 14044 5188
rect 14960 5188 14976 5612
rect 15040 5188 15056 5612
rect 15972 5612 16068 5628
rect 15379 5560 15701 5561
rect 15379 5240 15380 5560
rect 15700 5240 15701 5560
rect 15379 5239 15701 5240
rect 14960 5172 15056 5188
rect 15972 5188 15988 5612
rect 16052 5188 16068 5612
rect 16984 5612 17080 5628
rect 16391 5560 16713 5561
rect 16391 5240 16392 5560
rect 16712 5240 16713 5560
rect 16391 5239 16713 5240
rect 15972 5172 16068 5188
rect 16984 5188 17000 5612
rect 17064 5188 17080 5612
rect 16984 5172 17080 5188
rect -16412 4892 -16316 4908
rect -17005 4840 -16683 4841
rect -17005 4520 -17004 4840
rect -16684 4520 -16683 4840
rect -17005 4519 -16683 4520
rect -16412 4468 -16396 4892
rect -16332 4468 -16316 4892
rect -15400 4892 -15304 4908
rect -15993 4840 -15671 4841
rect -15993 4520 -15992 4840
rect -15672 4520 -15671 4840
rect -15993 4519 -15671 4520
rect -16412 4452 -16316 4468
rect -15400 4468 -15384 4892
rect -15320 4468 -15304 4892
rect -14388 4892 -14292 4908
rect -14981 4840 -14659 4841
rect -14981 4520 -14980 4840
rect -14660 4520 -14659 4840
rect -14981 4519 -14659 4520
rect -15400 4452 -15304 4468
rect -14388 4468 -14372 4892
rect -14308 4468 -14292 4892
rect -13376 4892 -13280 4908
rect -13969 4840 -13647 4841
rect -13969 4520 -13968 4840
rect -13648 4520 -13647 4840
rect -13969 4519 -13647 4520
rect -14388 4452 -14292 4468
rect -13376 4468 -13360 4892
rect -13296 4468 -13280 4892
rect -12364 4892 -12268 4908
rect -12957 4840 -12635 4841
rect -12957 4520 -12956 4840
rect -12636 4520 -12635 4840
rect -12957 4519 -12635 4520
rect -13376 4452 -13280 4468
rect -12364 4468 -12348 4892
rect -12284 4468 -12268 4892
rect -11352 4892 -11256 4908
rect -11945 4840 -11623 4841
rect -11945 4520 -11944 4840
rect -11624 4520 -11623 4840
rect -11945 4519 -11623 4520
rect -12364 4452 -12268 4468
rect -11352 4468 -11336 4892
rect -11272 4468 -11256 4892
rect -10340 4892 -10244 4908
rect -10933 4840 -10611 4841
rect -10933 4520 -10932 4840
rect -10612 4520 -10611 4840
rect -10933 4519 -10611 4520
rect -11352 4452 -11256 4468
rect -10340 4468 -10324 4892
rect -10260 4468 -10244 4892
rect -9328 4892 -9232 4908
rect -9921 4840 -9599 4841
rect -9921 4520 -9920 4840
rect -9600 4520 -9599 4840
rect -9921 4519 -9599 4520
rect -10340 4452 -10244 4468
rect -9328 4468 -9312 4892
rect -9248 4468 -9232 4892
rect -8316 4892 -8220 4908
rect -8909 4840 -8587 4841
rect -8909 4520 -8908 4840
rect -8588 4520 -8587 4840
rect -8909 4519 -8587 4520
rect -9328 4452 -9232 4468
rect -8316 4468 -8300 4892
rect -8236 4468 -8220 4892
rect -7304 4892 -7208 4908
rect -7897 4840 -7575 4841
rect -7897 4520 -7896 4840
rect -7576 4520 -7575 4840
rect -7897 4519 -7575 4520
rect -8316 4452 -8220 4468
rect -7304 4468 -7288 4892
rect -7224 4468 -7208 4892
rect -6292 4892 -6196 4908
rect -6885 4840 -6563 4841
rect -6885 4520 -6884 4840
rect -6564 4520 -6563 4840
rect -6885 4519 -6563 4520
rect -7304 4452 -7208 4468
rect -6292 4468 -6276 4892
rect -6212 4468 -6196 4892
rect -5280 4892 -5184 4908
rect -5873 4840 -5551 4841
rect -5873 4520 -5872 4840
rect -5552 4520 -5551 4840
rect -5873 4519 -5551 4520
rect -6292 4452 -6196 4468
rect -5280 4468 -5264 4892
rect -5200 4468 -5184 4892
rect -4268 4892 -4172 4908
rect -4861 4840 -4539 4841
rect -4861 4520 -4860 4840
rect -4540 4520 -4539 4840
rect -4861 4519 -4539 4520
rect -5280 4452 -5184 4468
rect -4268 4468 -4252 4892
rect -4188 4468 -4172 4892
rect -3256 4892 -3160 4908
rect -3849 4840 -3527 4841
rect -3849 4520 -3848 4840
rect -3528 4520 -3527 4840
rect -3849 4519 -3527 4520
rect -4268 4452 -4172 4468
rect -3256 4468 -3240 4892
rect -3176 4468 -3160 4892
rect -2244 4892 -2148 4908
rect -2837 4840 -2515 4841
rect -2837 4520 -2836 4840
rect -2516 4520 -2515 4840
rect -2837 4519 -2515 4520
rect -3256 4452 -3160 4468
rect -2244 4468 -2228 4892
rect -2164 4468 -2148 4892
rect -1232 4892 -1136 4908
rect -1825 4840 -1503 4841
rect -1825 4520 -1824 4840
rect -1504 4520 -1503 4840
rect -1825 4519 -1503 4520
rect -2244 4452 -2148 4468
rect -1232 4468 -1216 4892
rect -1152 4468 -1136 4892
rect -220 4892 -124 4908
rect -813 4840 -491 4841
rect -813 4520 -812 4840
rect -492 4520 -491 4840
rect -813 4519 -491 4520
rect -1232 4452 -1136 4468
rect -220 4468 -204 4892
rect -140 4468 -124 4892
rect 792 4892 888 4908
rect 199 4840 521 4841
rect 199 4520 200 4840
rect 520 4520 521 4840
rect 199 4519 521 4520
rect -220 4452 -124 4468
rect 792 4468 808 4892
rect 872 4468 888 4892
rect 1804 4892 1900 4908
rect 1211 4840 1533 4841
rect 1211 4520 1212 4840
rect 1532 4520 1533 4840
rect 1211 4519 1533 4520
rect 792 4452 888 4468
rect 1804 4468 1820 4892
rect 1884 4468 1900 4892
rect 2816 4892 2912 4908
rect 2223 4840 2545 4841
rect 2223 4520 2224 4840
rect 2544 4520 2545 4840
rect 2223 4519 2545 4520
rect 1804 4452 1900 4468
rect 2816 4468 2832 4892
rect 2896 4468 2912 4892
rect 3828 4892 3924 4908
rect 3235 4840 3557 4841
rect 3235 4520 3236 4840
rect 3556 4520 3557 4840
rect 3235 4519 3557 4520
rect 2816 4452 2912 4468
rect 3828 4468 3844 4892
rect 3908 4468 3924 4892
rect 4840 4892 4936 4908
rect 4247 4840 4569 4841
rect 4247 4520 4248 4840
rect 4568 4520 4569 4840
rect 4247 4519 4569 4520
rect 3828 4452 3924 4468
rect 4840 4468 4856 4892
rect 4920 4468 4936 4892
rect 5852 4892 5948 4908
rect 5259 4840 5581 4841
rect 5259 4520 5260 4840
rect 5580 4520 5581 4840
rect 5259 4519 5581 4520
rect 4840 4452 4936 4468
rect 5852 4468 5868 4892
rect 5932 4468 5948 4892
rect 6864 4892 6960 4908
rect 6271 4840 6593 4841
rect 6271 4520 6272 4840
rect 6592 4520 6593 4840
rect 6271 4519 6593 4520
rect 5852 4452 5948 4468
rect 6864 4468 6880 4892
rect 6944 4468 6960 4892
rect 7876 4892 7972 4908
rect 7283 4840 7605 4841
rect 7283 4520 7284 4840
rect 7604 4520 7605 4840
rect 7283 4519 7605 4520
rect 6864 4452 6960 4468
rect 7876 4468 7892 4892
rect 7956 4468 7972 4892
rect 8888 4892 8984 4908
rect 8295 4840 8617 4841
rect 8295 4520 8296 4840
rect 8616 4520 8617 4840
rect 8295 4519 8617 4520
rect 7876 4452 7972 4468
rect 8888 4468 8904 4892
rect 8968 4468 8984 4892
rect 9900 4892 9996 4908
rect 9307 4840 9629 4841
rect 9307 4520 9308 4840
rect 9628 4520 9629 4840
rect 9307 4519 9629 4520
rect 8888 4452 8984 4468
rect 9900 4468 9916 4892
rect 9980 4468 9996 4892
rect 10912 4892 11008 4908
rect 10319 4840 10641 4841
rect 10319 4520 10320 4840
rect 10640 4520 10641 4840
rect 10319 4519 10641 4520
rect 9900 4452 9996 4468
rect 10912 4468 10928 4892
rect 10992 4468 11008 4892
rect 11924 4892 12020 4908
rect 11331 4840 11653 4841
rect 11331 4520 11332 4840
rect 11652 4520 11653 4840
rect 11331 4519 11653 4520
rect 10912 4452 11008 4468
rect 11924 4468 11940 4892
rect 12004 4468 12020 4892
rect 12936 4892 13032 4908
rect 12343 4840 12665 4841
rect 12343 4520 12344 4840
rect 12664 4520 12665 4840
rect 12343 4519 12665 4520
rect 11924 4452 12020 4468
rect 12936 4468 12952 4892
rect 13016 4468 13032 4892
rect 13948 4892 14044 4908
rect 13355 4840 13677 4841
rect 13355 4520 13356 4840
rect 13676 4520 13677 4840
rect 13355 4519 13677 4520
rect 12936 4452 13032 4468
rect 13948 4468 13964 4892
rect 14028 4468 14044 4892
rect 14960 4892 15056 4908
rect 14367 4840 14689 4841
rect 14367 4520 14368 4840
rect 14688 4520 14689 4840
rect 14367 4519 14689 4520
rect 13948 4452 14044 4468
rect 14960 4468 14976 4892
rect 15040 4468 15056 4892
rect 15972 4892 16068 4908
rect 15379 4840 15701 4841
rect 15379 4520 15380 4840
rect 15700 4520 15701 4840
rect 15379 4519 15701 4520
rect 14960 4452 15056 4468
rect 15972 4468 15988 4892
rect 16052 4468 16068 4892
rect 16984 4892 17080 4908
rect 16391 4840 16713 4841
rect 16391 4520 16392 4840
rect 16712 4520 16713 4840
rect 16391 4519 16713 4520
rect 15972 4452 16068 4468
rect 16984 4468 17000 4892
rect 17064 4468 17080 4892
rect 16984 4452 17080 4468
rect -16412 4172 -16316 4188
rect -17005 4120 -16683 4121
rect -17005 3800 -17004 4120
rect -16684 3800 -16683 4120
rect -17005 3799 -16683 3800
rect -16412 3748 -16396 4172
rect -16332 3748 -16316 4172
rect -15400 4172 -15304 4188
rect -15993 4120 -15671 4121
rect -15993 3800 -15992 4120
rect -15672 3800 -15671 4120
rect -15993 3799 -15671 3800
rect -16412 3732 -16316 3748
rect -15400 3748 -15384 4172
rect -15320 3748 -15304 4172
rect -14388 4172 -14292 4188
rect -14981 4120 -14659 4121
rect -14981 3800 -14980 4120
rect -14660 3800 -14659 4120
rect -14981 3799 -14659 3800
rect -15400 3732 -15304 3748
rect -14388 3748 -14372 4172
rect -14308 3748 -14292 4172
rect -13376 4172 -13280 4188
rect -13969 4120 -13647 4121
rect -13969 3800 -13968 4120
rect -13648 3800 -13647 4120
rect -13969 3799 -13647 3800
rect -14388 3732 -14292 3748
rect -13376 3748 -13360 4172
rect -13296 3748 -13280 4172
rect -12364 4172 -12268 4188
rect -12957 4120 -12635 4121
rect -12957 3800 -12956 4120
rect -12636 3800 -12635 4120
rect -12957 3799 -12635 3800
rect -13376 3732 -13280 3748
rect -12364 3748 -12348 4172
rect -12284 3748 -12268 4172
rect -11352 4172 -11256 4188
rect -11945 4120 -11623 4121
rect -11945 3800 -11944 4120
rect -11624 3800 -11623 4120
rect -11945 3799 -11623 3800
rect -12364 3732 -12268 3748
rect -11352 3748 -11336 4172
rect -11272 3748 -11256 4172
rect -10340 4172 -10244 4188
rect -10933 4120 -10611 4121
rect -10933 3800 -10932 4120
rect -10612 3800 -10611 4120
rect -10933 3799 -10611 3800
rect -11352 3732 -11256 3748
rect -10340 3748 -10324 4172
rect -10260 3748 -10244 4172
rect -9328 4172 -9232 4188
rect -9921 4120 -9599 4121
rect -9921 3800 -9920 4120
rect -9600 3800 -9599 4120
rect -9921 3799 -9599 3800
rect -10340 3732 -10244 3748
rect -9328 3748 -9312 4172
rect -9248 3748 -9232 4172
rect -8316 4172 -8220 4188
rect -8909 4120 -8587 4121
rect -8909 3800 -8908 4120
rect -8588 3800 -8587 4120
rect -8909 3799 -8587 3800
rect -9328 3732 -9232 3748
rect -8316 3748 -8300 4172
rect -8236 3748 -8220 4172
rect -7304 4172 -7208 4188
rect -7897 4120 -7575 4121
rect -7897 3800 -7896 4120
rect -7576 3800 -7575 4120
rect -7897 3799 -7575 3800
rect -8316 3732 -8220 3748
rect -7304 3748 -7288 4172
rect -7224 3748 -7208 4172
rect -6292 4172 -6196 4188
rect -6885 4120 -6563 4121
rect -6885 3800 -6884 4120
rect -6564 3800 -6563 4120
rect -6885 3799 -6563 3800
rect -7304 3732 -7208 3748
rect -6292 3748 -6276 4172
rect -6212 3748 -6196 4172
rect -5280 4172 -5184 4188
rect -5873 4120 -5551 4121
rect -5873 3800 -5872 4120
rect -5552 3800 -5551 4120
rect -5873 3799 -5551 3800
rect -6292 3732 -6196 3748
rect -5280 3748 -5264 4172
rect -5200 3748 -5184 4172
rect -4268 4172 -4172 4188
rect -4861 4120 -4539 4121
rect -4861 3800 -4860 4120
rect -4540 3800 -4539 4120
rect -4861 3799 -4539 3800
rect -5280 3732 -5184 3748
rect -4268 3748 -4252 4172
rect -4188 3748 -4172 4172
rect -3256 4172 -3160 4188
rect -3849 4120 -3527 4121
rect -3849 3800 -3848 4120
rect -3528 3800 -3527 4120
rect -3849 3799 -3527 3800
rect -4268 3732 -4172 3748
rect -3256 3748 -3240 4172
rect -3176 3748 -3160 4172
rect -2244 4172 -2148 4188
rect -2837 4120 -2515 4121
rect -2837 3800 -2836 4120
rect -2516 3800 -2515 4120
rect -2837 3799 -2515 3800
rect -3256 3732 -3160 3748
rect -2244 3748 -2228 4172
rect -2164 3748 -2148 4172
rect -1232 4172 -1136 4188
rect -1825 4120 -1503 4121
rect -1825 3800 -1824 4120
rect -1504 3800 -1503 4120
rect -1825 3799 -1503 3800
rect -2244 3732 -2148 3748
rect -1232 3748 -1216 4172
rect -1152 3748 -1136 4172
rect -220 4172 -124 4188
rect -813 4120 -491 4121
rect -813 3800 -812 4120
rect -492 3800 -491 4120
rect -813 3799 -491 3800
rect -1232 3732 -1136 3748
rect -220 3748 -204 4172
rect -140 3748 -124 4172
rect 792 4172 888 4188
rect 199 4120 521 4121
rect 199 3800 200 4120
rect 520 3800 521 4120
rect 199 3799 521 3800
rect -220 3732 -124 3748
rect 792 3748 808 4172
rect 872 3748 888 4172
rect 1804 4172 1900 4188
rect 1211 4120 1533 4121
rect 1211 3800 1212 4120
rect 1532 3800 1533 4120
rect 1211 3799 1533 3800
rect 792 3732 888 3748
rect 1804 3748 1820 4172
rect 1884 3748 1900 4172
rect 2816 4172 2912 4188
rect 2223 4120 2545 4121
rect 2223 3800 2224 4120
rect 2544 3800 2545 4120
rect 2223 3799 2545 3800
rect 1804 3732 1900 3748
rect 2816 3748 2832 4172
rect 2896 3748 2912 4172
rect 3828 4172 3924 4188
rect 3235 4120 3557 4121
rect 3235 3800 3236 4120
rect 3556 3800 3557 4120
rect 3235 3799 3557 3800
rect 2816 3732 2912 3748
rect 3828 3748 3844 4172
rect 3908 3748 3924 4172
rect 4840 4172 4936 4188
rect 4247 4120 4569 4121
rect 4247 3800 4248 4120
rect 4568 3800 4569 4120
rect 4247 3799 4569 3800
rect 3828 3732 3924 3748
rect 4840 3748 4856 4172
rect 4920 3748 4936 4172
rect 5852 4172 5948 4188
rect 5259 4120 5581 4121
rect 5259 3800 5260 4120
rect 5580 3800 5581 4120
rect 5259 3799 5581 3800
rect 4840 3732 4936 3748
rect 5852 3748 5868 4172
rect 5932 3748 5948 4172
rect 6864 4172 6960 4188
rect 6271 4120 6593 4121
rect 6271 3800 6272 4120
rect 6592 3800 6593 4120
rect 6271 3799 6593 3800
rect 5852 3732 5948 3748
rect 6864 3748 6880 4172
rect 6944 3748 6960 4172
rect 7876 4172 7972 4188
rect 7283 4120 7605 4121
rect 7283 3800 7284 4120
rect 7604 3800 7605 4120
rect 7283 3799 7605 3800
rect 6864 3732 6960 3748
rect 7876 3748 7892 4172
rect 7956 3748 7972 4172
rect 8888 4172 8984 4188
rect 8295 4120 8617 4121
rect 8295 3800 8296 4120
rect 8616 3800 8617 4120
rect 8295 3799 8617 3800
rect 7876 3732 7972 3748
rect 8888 3748 8904 4172
rect 8968 3748 8984 4172
rect 9900 4172 9996 4188
rect 9307 4120 9629 4121
rect 9307 3800 9308 4120
rect 9628 3800 9629 4120
rect 9307 3799 9629 3800
rect 8888 3732 8984 3748
rect 9900 3748 9916 4172
rect 9980 3748 9996 4172
rect 10912 4172 11008 4188
rect 10319 4120 10641 4121
rect 10319 3800 10320 4120
rect 10640 3800 10641 4120
rect 10319 3799 10641 3800
rect 9900 3732 9996 3748
rect 10912 3748 10928 4172
rect 10992 3748 11008 4172
rect 11924 4172 12020 4188
rect 11331 4120 11653 4121
rect 11331 3800 11332 4120
rect 11652 3800 11653 4120
rect 11331 3799 11653 3800
rect 10912 3732 11008 3748
rect 11924 3748 11940 4172
rect 12004 3748 12020 4172
rect 12936 4172 13032 4188
rect 12343 4120 12665 4121
rect 12343 3800 12344 4120
rect 12664 3800 12665 4120
rect 12343 3799 12665 3800
rect 11924 3732 12020 3748
rect 12936 3748 12952 4172
rect 13016 3748 13032 4172
rect 13948 4172 14044 4188
rect 13355 4120 13677 4121
rect 13355 3800 13356 4120
rect 13676 3800 13677 4120
rect 13355 3799 13677 3800
rect 12936 3732 13032 3748
rect 13948 3748 13964 4172
rect 14028 3748 14044 4172
rect 14960 4172 15056 4188
rect 14367 4120 14689 4121
rect 14367 3800 14368 4120
rect 14688 3800 14689 4120
rect 14367 3799 14689 3800
rect 13948 3732 14044 3748
rect 14960 3748 14976 4172
rect 15040 3748 15056 4172
rect 15972 4172 16068 4188
rect 15379 4120 15701 4121
rect 15379 3800 15380 4120
rect 15700 3800 15701 4120
rect 15379 3799 15701 3800
rect 14960 3732 15056 3748
rect 15972 3748 15988 4172
rect 16052 3748 16068 4172
rect 16984 4172 17080 4188
rect 16391 4120 16713 4121
rect 16391 3800 16392 4120
rect 16712 3800 16713 4120
rect 16391 3799 16713 3800
rect 15972 3732 16068 3748
rect 16984 3748 17000 4172
rect 17064 3748 17080 4172
rect 16984 3732 17080 3748
rect -16412 3452 -16316 3468
rect -17005 3400 -16683 3401
rect -17005 3080 -17004 3400
rect -16684 3080 -16683 3400
rect -17005 3079 -16683 3080
rect -16412 3028 -16396 3452
rect -16332 3028 -16316 3452
rect -15400 3452 -15304 3468
rect -15993 3400 -15671 3401
rect -15993 3080 -15992 3400
rect -15672 3080 -15671 3400
rect -15993 3079 -15671 3080
rect -16412 3012 -16316 3028
rect -15400 3028 -15384 3452
rect -15320 3028 -15304 3452
rect -14388 3452 -14292 3468
rect -14981 3400 -14659 3401
rect -14981 3080 -14980 3400
rect -14660 3080 -14659 3400
rect -14981 3079 -14659 3080
rect -15400 3012 -15304 3028
rect -14388 3028 -14372 3452
rect -14308 3028 -14292 3452
rect -13376 3452 -13280 3468
rect -13969 3400 -13647 3401
rect -13969 3080 -13968 3400
rect -13648 3080 -13647 3400
rect -13969 3079 -13647 3080
rect -14388 3012 -14292 3028
rect -13376 3028 -13360 3452
rect -13296 3028 -13280 3452
rect -12364 3452 -12268 3468
rect -12957 3400 -12635 3401
rect -12957 3080 -12956 3400
rect -12636 3080 -12635 3400
rect -12957 3079 -12635 3080
rect -13376 3012 -13280 3028
rect -12364 3028 -12348 3452
rect -12284 3028 -12268 3452
rect -11352 3452 -11256 3468
rect -11945 3400 -11623 3401
rect -11945 3080 -11944 3400
rect -11624 3080 -11623 3400
rect -11945 3079 -11623 3080
rect -12364 3012 -12268 3028
rect -11352 3028 -11336 3452
rect -11272 3028 -11256 3452
rect -10340 3452 -10244 3468
rect -10933 3400 -10611 3401
rect -10933 3080 -10932 3400
rect -10612 3080 -10611 3400
rect -10933 3079 -10611 3080
rect -11352 3012 -11256 3028
rect -10340 3028 -10324 3452
rect -10260 3028 -10244 3452
rect -9328 3452 -9232 3468
rect -9921 3400 -9599 3401
rect -9921 3080 -9920 3400
rect -9600 3080 -9599 3400
rect -9921 3079 -9599 3080
rect -10340 3012 -10244 3028
rect -9328 3028 -9312 3452
rect -9248 3028 -9232 3452
rect -8316 3452 -8220 3468
rect -8909 3400 -8587 3401
rect -8909 3080 -8908 3400
rect -8588 3080 -8587 3400
rect -8909 3079 -8587 3080
rect -9328 3012 -9232 3028
rect -8316 3028 -8300 3452
rect -8236 3028 -8220 3452
rect -7304 3452 -7208 3468
rect -7897 3400 -7575 3401
rect -7897 3080 -7896 3400
rect -7576 3080 -7575 3400
rect -7897 3079 -7575 3080
rect -8316 3012 -8220 3028
rect -7304 3028 -7288 3452
rect -7224 3028 -7208 3452
rect -6292 3452 -6196 3468
rect -6885 3400 -6563 3401
rect -6885 3080 -6884 3400
rect -6564 3080 -6563 3400
rect -6885 3079 -6563 3080
rect -7304 3012 -7208 3028
rect -6292 3028 -6276 3452
rect -6212 3028 -6196 3452
rect -5280 3452 -5184 3468
rect -5873 3400 -5551 3401
rect -5873 3080 -5872 3400
rect -5552 3080 -5551 3400
rect -5873 3079 -5551 3080
rect -6292 3012 -6196 3028
rect -5280 3028 -5264 3452
rect -5200 3028 -5184 3452
rect -4268 3452 -4172 3468
rect -4861 3400 -4539 3401
rect -4861 3080 -4860 3400
rect -4540 3080 -4539 3400
rect -4861 3079 -4539 3080
rect -5280 3012 -5184 3028
rect -4268 3028 -4252 3452
rect -4188 3028 -4172 3452
rect -3256 3452 -3160 3468
rect -3849 3400 -3527 3401
rect -3849 3080 -3848 3400
rect -3528 3080 -3527 3400
rect -3849 3079 -3527 3080
rect -4268 3012 -4172 3028
rect -3256 3028 -3240 3452
rect -3176 3028 -3160 3452
rect -2244 3452 -2148 3468
rect -2837 3400 -2515 3401
rect -2837 3080 -2836 3400
rect -2516 3080 -2515 3400
rect -2837 3079 -2515 3080
rect -3256 3012 -3160 3028
rect -2244 3028 -2228 3452
rect -2164 3028 -2148 3452
rect -1232 3452 -1136 3468
rect -1825 3400 -1503 3401
rect -1825 3080 -1824 3400
rect -1504 3080 -1503 3400
rect -1825 3079 -1503 3080
rect -2244 3012 -2148 3028
rect -1232 3028 -1216 3452
rect -1152 3028 -1136 3452
rect -220 3452 -124 3468
rect -813 3400 -491 3401
rect -813 3080 -812 3400
rect -492 3080 -491 3400
rect -813 3079 -491 3080
rect -1232 3012 -1136 3028
rect -220 3028 -204 3452
rect -140 3028 -124 3452
rect 792 3452 888 3468
rect 199 3400 521 3401
rect 199 3080 200 3400
rect 520 3080 521 3400
rect 199 3079 521 3080
rect -220 3012 -124 3028
rect 792 3028 808 3452
rect 872 3028 888 3452
rect 1804 3452 1900 3468
rect 1211 3400 1533 3401
rect 1211 3080 1212 3400
rect 1532 3080 1533 3400
rect 1211 3079 1533 3080
rect 792 3012 888 3028
rect 1804 3028 1820 3452
rect 1884 3028 1900 3452
rect 2816 3452 2912 3468
rect 2223 3400 2545 3401
rect 2223 3080 2224 3400
rect 2544 3080 2545 3400
rect 2223 3079 2545 3080
rect 1804 3012 1900 3028
rect 2816 3028 2832 3452
rect 2896 3028 2912 3452
rect 3828 3452 3924 3468
rect 3235 3400 3557 3401
rect 3235 3080 3236 3400
rect 3556 3080 3557 3400
rect 3235 3079 3557 3080
rect 2816 3012 2912 3028
rect 3828 3028 3844 3452
rect 3908 3028 3924 3452
rect 4840 3452 4936 3468
rect 4247 3400 4569 3401
rect 4247 3080 4248 3400
rect 4568 3080 4569 3400
rect 4247 3079 4569 3080
rect 3828 3012 3924 3028
rect 4840 3028 4856 3452
rect 4920 3028 4936 3452
rect 5852 3452 5948 3468
rect 5259 3400 5581 3401
rect 5259 3080 5260 3400
rect 5580 3080 5581 3400
rect 5259 3079 5581 3080
rect 4840 3012 4936 3028
rect 5852 3028 5868 3452
rect 5932 3028 5948 3452
rect 6864 3452 6960 3468
rect 6271 3400 6593 3401
rect 6271 3080 6272 3400
rect 6592 3080 6593 3400
rect 6271 3079 6593 3080
rect 5852 3012 5948 3028
rect 6864 3028 6880 3452
rect 6944 3028 6960 3452
rect 7876 3452 7972 3468
rect 7283 3400 7605 3401
rect 7283 3080 7284 3400
rect 7604 3080 7605 3400
rect 7283 3079 7605 3080
rect 6864 3012 6960 3028
rect 7876 3028 7892 3452
rect 7956 3028 7972 3452
rect 8888 3452 8984 3468
rect 8295 3400 8617 3401
rect 8295 3080 8296 3400
rect 8616 3080 8617 3400
rect 8295 3079 8617 3080
rect 7876 3012 7972 3028
rect 8888 3028 8904 3452
rect 8968 3028 8984 3452
rect 9900 3452 9996 3468
rect 9307 3400 9629 3401
rect 9307 3080 9308 3400
rect 9628 3080 9629 3400
rect 9307 3079 9629 3080
rect 8888 3012 8984 3028
rect 9900 3028 9916 3452
rect 9980 3028 9996 3452
rect 10912 3452 11008 3468
rect 10319 3400 10641 3401
rect 10319 3080 10320 3400
rect 10640 3080 10641 3400
rect 10319 3079 10641 3080
rect 9900 3012 9996 3028
rect 10912 3028 10928 3452
rect 10992 3028 11008 3452
rect 11924 3452 12020 3468
rect 11331 3400 11653 3401
rect 11331 3080 11332 3400
rect 11652 3080 11653 3400
rect 11331 3079 11653 3080
rect 10912 3012 11008 3028
rect 11924 3028 11940 3452
rect 12004 3028 12020 3452
rect 12936 3452 13032 3468
rect 12343 3400 12665 3401
rect 12343 3080 12344 3400
rect 12664 3080 12665 3400
rect 12343 3079 12665 3080
rect 11924 3012 12020 3028
rect 12936 3028 12952 3452
rect 13016 3028 13032 3452
rect 13948 3452 14044 3468
rect 13355 3400 13677 3401
rect 13355 3080 13356 3400
rect 13676 3080 13677 3400
rect 13355 3079 13677 3080
rect 12936 3012 13032 3028
rect 13948 3028 13964 3452
rect 14028 3028 14044 3452
rect 14960 3452 15056 3468
rect 14367 3400 14689 3401
rect 14367 3080 14368 3400
rect 14688 3080 14689 3400
rect 14367 3079 14689 3080
rect 13948 3012 14044 3028
rect 14960 3028 14976 3452
rect 15040 3028 15056 3452
rect 15972 3452 16068 3468
rect 15379 3400 15701 3401
rect 15379 3080 15380 3400
rect 15700 3080 15701 3400
rect 15379 3079 15701 3080
rect 14960 3012 15056 3028
rect 15972 3028 15988 3452
rect 16052 3028 16068 3452
rect 16984 3452 17080 3468
rect 16391 3400 16713 3401
rect 16391 3080 16392 3400
rect 16712 3080 16713 3400
rect 16391 3079 16713 3080
rect 15972 3012 16068 3028
rect 16984 3028 17000 3452
rect 17064 3028 17080 3452
rect 16984 3012 17080 3028
rect -16412 2732 -16316 2748
rect -17005 2680 -16683 2681
rect -17005 2360 -17004 2680
rect -16684 2360 -16683 2680
rect -17005 2359 -16683 2360
rect -16412 2308 -16396 2732
rect -16332 2308 -16316 2732
rect -15400 2732 -15304 2748
rect -15993 2680 -15671 2681
rect -15993 2360 -15992 2680
rect -15672 2360 -15671 2680
rect -15993 2359 -15671 2360
rect -16412 2292 -16316 2308
rect -15400 2308 -15384 2732
rect -15320 2308 -15304 2732
rect -14388 2732 -14292 2748
rect -14981 2680 -14659 2681
rect -14981 2360 -14980 2680
rect -14660 2360 -14659 2680
rect -14981 2359 -14659 2360
rect -15400 2292 -15304 2308
rect -14388 2308 -14372 2732
rect -14308 2308 -14292 2732
rect -13376 2732 -13280 2748
rect -13969 2680 -13647 2681
rect -13969 2360 -13968 2680
rect -13648 2360 -13647 2680
rect -13969 2359 -13647 2360
rect -14388 2292 -14292 2308
rect -13376 2308 -13360 2732
rect -13296 2308 -13280 2732
rect -12364 2732 -12268 2748
rect -12957 2680 -12635 2681
rect -12957 2360 -12956 2680
rect -12636 2360 -12635 2680
rect -12957 2359 -12635 2360
rect -13376 2292 -13280 2308
rect -12364 2308 -12348 2732
rect -12284 2308 -12268 2732
rect -11352 2732 -11256 2748
rect -11945 2680 -11623 2681
rect -11945 2360 -11944 2680
rect -11624 2360 -11623 2680
rect -11945 2359 -11623 2360
rect -12364 2292 -12268 2308
rect -11352 2308 -11336 2732
rect -11272 2308 -11256 2732
rect -10340 2732 -10244 2748
rect -10933 2680 -10611 2681
rect -10933 2360 -10932 2680
rect -10612 2360 -10611 2680
rect -10933 2359 -10611 2360
rect -11352 2292 -11256 2308
rect -10340 2308 -10324 2732
rect -10260 2308 -10244 2732
rect -9328 2732 -9232 2748
rect -9921 2680 -9599 2681
rect -9921 2360 -9920 2680
rect -9600 2360 -9599 2680
rect -9921 2359 -9599 2360
rect -10340 2292 -10244 2308
rect -9328 2308 -9312 2732
rect -9248 2308 -9232 2732
rect -8316 2732 -8220 2748
rect -8909 2680 -8587 2681
rect -8909 2360 -8908 2680
rect -8588 2360 -8587 2680
rect -8909 2359 -8587 2360
rect -9328 2292 -9232 2308
rect -8316 2308 -8300 2732
rect -8236 2308 -8220 2732
rect -7304 2732 -7208 2748
rect -7897 2680 -7575 2681
rect -7897 2360 -7896 2680
rect -7576 2360 -7575 2680
rect -7897 2359 -7575 2360
rect -8316 2292 -8220 2308
rect -7304 2308 -7288 2732
rect -7224 2308 -7208 2732
rect -6292 2732 -6196 2748
rect -6885 2680 -6563 2681
rect -6885 2360 -6884 2680
rect -6564 2360 -6563 2680
rect -6885 2359 -6563 2360
rect -7304 2292 -7208 2308
rect -6292 2308 -6276 2732
rect -6212 2308 -6196 2732
rect -5280 2732 -5184 2748
rect -5873 2680 -5551 2681
rect -5873 2360 -5872 2680
rect -5552 2360 -5551 2680
rect -5873 2359 -5551 2360
rect -6292 2292 -6196 2308
rect -5280 2308 -5264 2732
rect -5200 2308 -5184 2732
rect -4268 2732 -4172 2748
rect -4861 2680 -4539 2681
rect -4861 2360 -4860 2680
rect -4540 2360 -4539 2680
rect -4861 2359 -4539 2360
rect -5280 2292 -5184 2308
rect -4268 2308 -4252 2732
rect -4188 2308 -4172 2732
rect -3256 2732 -3160 2748
rect -3849 2680 -3527 2681
rect -3849 2360 -3848 2680
rect -3528 2360 -3527 2680
rect -3849 2359 -3527 2360
rect -4268 2292 -4172 2308
rect -3256 2308 -3240 2732
rect -3176 2308 -3160 2732
rect -2244 2732 -2148 2748
rect -2837 2680 -2515 2681
rect -2837 2360 -2836 2680
rect -2516 2360 -2515 2680
rect -2837 2359 -2515 2360
rect -3256 2292 -3160 2308
rect -2244 2308 -2228 2732
rect -2164 2308 -2148 2732
rect -1232 2732 -1136 2748
rect -1825 2680 -1503 2681
rect -1825 2360 -1824 2680
rect -1504 2360 -1503 2680
rect -1825 2359 -1503 2360
rect -2244 2292 -2148 2308
rect -1232 2308 -1216 2732
rect -1152 2308 -1136 2732
rect -220 2732 -124 2748
rect -813 2680 -491 2681
rect -813 2360 -812 2680
rect -492 2360 -491 2680
rect -813 2359 -491 2360
rect -1232 2292 -1136 2308
rect -220 2308 -204 2732
rect -140 2308 -124 2732
rect 792 2732 888 2748
rect 199 2680 521 2681
rect 199 2360 200 2680
rect 520 2360 521 2680
rect 199 2359 521 2360
rect -220 2292 -124 2308
rect 792 2308 808 2732
rect 872 2308 888 2732
rect 1804 2732 1900 2748
rect 1211 2680 1533 2681
rect 1211 2360 1212 2680
rect 1532 2360 1533 2680
rect 1211 2359 1533 2360
rect 792 2292 888 2308
rect 1804 2308 1820 2732
rect 1884 2308 1900 2732
rect 2816 2732 2912 2748
rect 2223 2680 2545 2681
rect 2223 2360 2224 2680
rect 2544 2360 2545 2680
rect 2223 2359 2545 2360
rect 1804 2292 1900 2308
rect 2816 2308 2832 2732
rect 2896 2308 2912 2732
rect 3828 2732 3924 2748
rect 3235 2680 3557 2681
rect 3235 2360 3236 2680
rect 3556 2360 3557 2680
rect 3235 2359 3557 2360
rect 2816 2292 2912 2308
rect 3828 2308 3844 2732
rect 3908 2308 3924 2732
rect 4840 2732 4936 2748
rect 4247 2680 4569 2681
rect 4247 2360 4248 2680
rect 4568 2360 4569 2680
rect 4247 2359 4569 2360
rect 3828 2292 3924 2308
rect 4840 2308 4856 2732
rect 4920 2308 4936 2732
rect 5852 2732 5948 2748
rect 5259 2680 5581 2681
rect 5259 2360 5260 2680
rect 5580 2360 5581 2680
rect 5259 2359 5581 2360
rect 4840 2292 4936 2308
rect 5852 2308 5868 2732
rect 5932 2308 5948 2732
rect 6864 2732 6960 2748
rect 6271 2680 6593 2681
rect 6271 2360 6272 2680
rect 6592 2360 6593 2680
rect 6271 2359 6593 2360
rect 5852 2292 5948 2308
rect 6864 2308 6880 2732
rect 6944 2308 6960 2732
rect 7876 2732 7972 2748
rect 7283 2680 7605 2681
rect 7283 2360 7284 2680
rect 7604 2360 7605 2680
rect 7283 2359 7605 2360
rect 6864 2292 6960 2308
rect 7876 2308 7892 2732
rect 7956 2308 7972 2732
rect 8888 2732 8984 2748
rect 8295 2680 8617 2681
rect 8295 2360 8296 2680
rect 8616 2360 8617 2680
rect 8295 2359 8617 2360
rect 7876 2292 7972 2308
rect 8888 2308 8904 2732
rect 8968 2308 8984 2732
rect 9900 2732 9996 2748
rect 9307 2680 9629 2681
rect 9307 2360 9308 2680
rect 9628 2360 9629 2680
rect 9307 2359 9629 2360
rect 8888 2292 8984 2308
rect 9900 2308 9916 2732
rect 9980 2308 9996 2732
rect 10912 2732 11008 2748
rect 10319 2680 10641 2681
rect 10319 2360 10320 2680
rect 10640 2360 10641 2680
rect 10319 2359 10641 2360
rect 9900 2292 9996 2308
rect 10912 2308 10928 2732
rect 10992 2308 11008 2732
rect 11924 2732 12020 2748
rect 11331 2680 11653 2681
rect 11331 2360 11332 2680
rect 11652 2360 11653 2680
rect 11331 2359 11653 2360
rect 10912 2292 11008 2308
rect 11924 2308 11940 2732
rect 12004 2308 12020 2732
rect 12936 2732 13032 2748
rect 12343 2680 12665 2681
rect 12343 2360 12344 2680
rect 12664 2360 12665 2680
rect 12343 2359 12665 2360
rect 11924 2292 12020 2308
rect 12936 2308 12952 2732
rect 13016 2308 13032 2732
rect 13948 2732 14044 2748
rect 13355 2680 13677 2681
rect 13355 2360 13356 2680
rect 13676 2360 13677 2680
rect 13355 2359 13677 2360
rect 12936 2292 13032 2308
rect 13948 2308 13964 2732
rect 14028 2308 14044 2732
rect 14960 2732 15056 2748
rect 14367 2680 14689 2681
rect 14367 2360 14368 2680
rect 14688 2360 14689 2680
rect 14367 2359 14689 2360
rect 13948 2292 14044 2308
rect 14960 2308 14976 2732
rect 15040 2308 15056 2732
rect 15972 2732 16068 2748
rect 15379 2680 15701 2681
rect 15379 2360 15380 2680
rect 15700 2360 15701 2680
rect 15379 2359 15701 2360
rect 14960 2292 15056 2308
rect 15972 2308 15988 2732
rect 16052 2308 16068 2732
rect 16984 2732 17080 2748
rect 16391 2680 16713 2681
rect 16391 2360 16392 2680
rect 16712 2360 16713 2680
rect 16391 2359 16713 2360
rect 15972 2292 16068 2308
rect 16984 2308 17000 2732
rect 17064 2308 17080 2732
rect 16984 2292 17080 2308
rect -16412 2012 -16316 2028
rect -17005 1960 -16683 1961
rect -17005 1640 -17004 1960
rect -16684 1640 -16683 1960
rect -17005 1639 -16683 1640
rect -16412 1588 -16396 2012
rect -16332 1588 -16316 2012
rect -15400 2012 -15304 2028
rect -15993 1960 -15671 1961
rect -15993 1640 -15992 1960
rect -15672 1640 -15671 1960
rect -15993 1639 -15671 1640
rect -16412 1572 -16316 1588
rect -15400 1588 -15384 2012
rect -15320 1588 -15304 2012
rect -14388 2012 -14292 2028
rect -14981 1960 -14659 1961
rect -14981 1640 -14980 1960
rect -14660 1640 -14659 1960
rect -14981 1639 -14659 1640
rect -15400 1572 -15304 1588
rect -14388 1588 -14372 2012
rect -14308 1588 -14292 2012
rect -13376 2012 -13280 2028
rect -13969 1960 -13647 1961
rect -13969 1640 -13968 1960
rect -13648 1640 -13647 1960
rect -13969 1639 -13647 1640
rect -14388 1572 -14292 1588
rect -13376 1588 -13360 2012
rect -13296 1588 -13280 2012
rect -12364 2012 -12268 2028
rect -12957 1960 -12635 1961
rect -12957 1640 -12956 1960
rect -12636 1640 -12635 1960
rect -12957 1639 -12635 1640
rect -13376 1572 -13280 1588
rect -12364 1588 -12348 2012
rect -12284 1588 -12268 2012
rect -11352 2012 -11256 2028
rect -11945 1960 -11623 1961
rect -11945 1640 -11944 1960
rect -11624 1640 -11623 1960
rect -11945 1639 -11623 1640
rect -12364 1572 -12268 1588
rect -11352 1588 -11336 2012
rect -11272 1588 -11256 2012
rect -10340 2012 -10244 2028
rect -10933 1960 -10611 1961
rect -10933 1640 -10932 1960
rect -10612 1640 -10611 1960
rect -10933 1639 -10611 1640
rect -11352 1572 -11256 1588
rect -10340 1588 -10324 2012
rect -10260 1588 -10244 2012
rect -9328 2012 -9232 2028
rect -9921 1960 -9599 1961
rect -9921 1640 -9920 1960
rect -9600 1640 -9599 1960
rect -9921 1639 -9599 1640
rect -10340 1572 -10244 1588
rect -9328 1588 -9312 2012
rect -9248 1588 -9232 2012
rect -8316 2012 -8220 2028
rect -8909 1960 -8587 1961
rect -8909 1640 -8908 1960
rect -8588 1640 -8587 1960
rect -8909 1639 -8587 1640
rect -9328 1572 -9232 1588
rect -8316 1588 -8300 2012
rect -8236 1588 -8220 2012
rect -7304 2012 -7208 2028
rect -7897 1960 -7575 1961
rect -7897 1640 -7896 1960
rect -7576 1640 -7575 1960
rect -7897 1639 -7575 1640
rect -8316 1572 -8220 1588
rect -7304 1588 -7288 2012
rect -7224 1588 -7208 2012
rect -6292 2012 -6196 2028
rect -6885 1960 -6563 1961
rect -6885 1640 -6884 1960
rect -6564 1640 -6563 1960
rect -6885 1639 -6563 1640
rect -7304 1572 -7208 1588
rect -6292 1588 -6276 2012
rect -6212 1588 -6196 2012
rect -5280 2012 -5184 2028
rect -5873 1960 -5551 1961
rect -5873 1640 -5872 1960
rect -5552 1640 -5551 1960
rect -5873 1639 -5551 1640
rect -6292 1572 -6196 1588
rect -5280 1588 -5264 2012
rect -5200 1588 -5184 2012
rect -4268 2012 -4172 2028
rect -4861 1960 -4539 1961
rect -4861 1640 -4860 1960
rect -4540 1640 -4539 1960
rect -4861 1639 -4539 1640
rect -5280 1572 -5184 1588
rect -4268 1588 -4252 2012
rect -4188 1588 -4172 2012
rect -3256 2012 -3160 2028
rect -3849 1960 -3527 1961
rect -3849 1640 -3848 1960
rect -3528 1640 -3527 1960
rect -3849 1639 -3527 1640
rect -4268 1572 -4172 1588
rect -3256 1588 -3240 2012
rect -3176 1588 -3160 2012
rect -2244 2012 -2148 2028
rect -2837 1960 -2515 1961
rect -2837 1640 -2836 1960
rect -2516 1640 -2515 1960
rect -2837 1639 -2515 1640
rect -3256 1572 -3160 1588
rect -2244 1588 -2228 2012
rect -2164 1588 -2148 2012
rect -1232 2012 -1136 2028
rect -1825 1960 -1503 1961
rect -1825 1640 -1824 1960
rect -1504 1640 -1503 1960
rect -1825 1639 -1503 1640
rect -2244 1572 -2148 1588
rect -1232 1588 -1216 2012
rect -1152 1588 -1136 2012
rect -220 2012 -124 2028
rect -813 1960 -491 1961
rect -813 1640 -812 1960
rect -492 1640 -491 1960
rect -813 1639 -491 1640
rect -1232 1572 -1136 1588
rect -220 1588 -204 2012
rect -140 1588 -124 2012
rect 792 2012 888 2028
rect 199 1960 521 1961
rect 199 1640 200 1960
rect 520 1640 521 1960
rect 199 1639 521 1640
rect -220 1572 -124 1588
rect 792 1588 808 2012
rect 872 1588 888 2012
rect 1804 2012 1900 2028
rect 1211 1960 1533 1961
rect 1211 1640 1212 1960
rect 1532 1640 1533 1960
rect 1211 1639 1533 1640
rect 792 1572 888 1588
rect 1804 1588 1820 2012
rect 1884 1588 1900 2012
rect 2816 2012 2912 2028
rect 2223 1960 2545 1961
rect 2223 1640 2224 1960
rect 2544 1640 2545 1960
rect 2223 1639 2545 1640
rect 1804 1572 1900 1588
rect 2816 1588 2832 2012
rect 2896 1588 2912 2012
rect 3828 2012 3924 2028
rect 3235 1960 3557 1961
rect 3235 1640 3236 1960
rect 3556 1640 3557 1960
rect 3235 1639 3557 1640
rect 2816 1572 2912 1588
rect 3828 1588 3844 2012
rect 3908 1588 3924 2012
rect 4840 2012 4936 2028
rect 4247 1960 4569 1961
rect 4247 1640 4248 1960
rect 4568 1640 4569 1960
rect 4247 1639 4569 1640
rect 3828 1572 3924 1588
rect 4840 1588 4856 2012
rect 4920 1588 4936 2012
rect 5852 2012 5948 2028
rect 5259 1960 5581 1961
rect 5259 1640 5260 1960
rect 5580 1640 5581 1960
rect 5259 1639 5581 1640
rect 4840 1572 4936 1588
rect 5852 1588 5868 2012
rect 5932 1588 5948 2012
rect 6864 2012 6960 2028
rect 6271 1960 6593 1961
rect 6271 1640 6272 1960
rect 6592 1640 6593 1960
rect 6271 1639 6593 1640
rect 5852 1572 5948 1588
rect 6864 1588 6880 2012
rect 6944 1588 6960 2012
rect 7876 2012 7972 2028
rect 7283 1960 7605 1961
rect 7283 1640 7284 1960
rect 7604 1640 7605 1960
rect 7283 1639 7605 1640
rect 6864 1572 6960 1588
rect 7876 1588 7892 2012
rect 7956 1588 7972 2012
rect 8888 2012 8984 2028
rect 8295 1960 8617 1961
rect 8295 1640 8296 1960
rect 8616 1640 8617 1960
rect 8295 1639 8617 1640
rect 7876 1572 7972 1588
rect 8888 1588 8904 2012
rect 8968 1588 8984 2012
rect 9900 2012 9996 2028
rect 9307 1960 9629 1961
rect 9307 1640 9308 1960
rect 9628 1640 9629 1960
rect 9307 1639 9629 1640
rect 8888 1572 8984 1588
rect 9900 1588 9916 2012
rect 9980 1588 9996 2012
rect 10912 2012 11008 2028
rect 10319 1960 10641 1961
rect 10319 1640 10320 1960
rect 10640 1640 10641 1960
rect 10319 1639 10641 1640
rect 9900 1572 9996 1588
rect 10912 1588 10928 2012
rect 10992 1588 11008 2012
rect 11924 2012 12020 2028
rect 11331 1960 11653 1961
rect 11331 1640 11332 1960
rect 11652 1640 11653 1960
rect 11331 1639 11653 1640
rect 10912 1572 11008 1588
rect 11924 1588 11940 2012
rect 12004 1588 12020 2012
rect 12936 2012 13032 2028
rect 12343 1960 12665 1961
rect 12343 1640 12344 1960
rect 12664 1640 12665 1960
rect 12343 1639 12665 1640
rect 11924 1572 12020 1588
rect 12936 1588 12952 2012
rect 13016 1588 13032 2012
rect 13948 2012 14044 2028
rect 13355 1960 13677 1961
rect 13355 1640 13356 1960
rect 13676 1640 13677 1960
rect 13355 1639 13677 1640
rect 12936 1572 13032 1588
rect 13948 1588 13964 2012
rect 14028 1588 14044 2012
rect 14960 2012 15056 2028
rect 14367 1960 14689 1961
rect 14367 1640 14368 1960
rect 14688 1640 14689 1960
rect 14367 1639 14689 1640
rect 13948 1572 14044 1588
rect 14960 1588 14976 2012
rect 15040 1588 15056 2012
rect 15972 2012 16068 2028
rect 15379 1960 15701 1961
rect 15379 1640 15380 1960
rect 15700 1640 15701 1960
rect 15379 1639 15701 1640
rect 14960 1572 15056 1588
rect 15972 1588 15988 2012
rect 16052 1588 16068 2012
rect 16984 2012 17080 2028
rect 16391 1960 16713 1961
rect 16391 1640 16392 1960
rect 16712 1640 16713 1960
rect 16391 1639 16713 1640
rect 15972 1572 16068 1588
rect 16984 1588 17000 2012
rect 17064 1588 17080 2012
rect 16984 1572 17080 1588
rect -16412 1292 -16316 1308
rect -17005 1240 -16683 1241
rect -17005 920 -17004 1240
rect -16684 920 -16683 1240
rect -17005 919 -16683 920
rect -16412 868 -16396 1292
rect -16332 868 -16316 1292
rect -15400 1292 -15304 1308
rect -15993 1240 -15671 1241
rect -15993 920 -15992 1240
rect -15672 920 -15671 1240
rect -15993 919 -15671 920
rect -16412 852 -16316 868
rect -15400 868 -15384 1292
rect -15320 868 -15304 1292
rect -14388 1292 -14292 1308
rect -14981 1240 -14659 1241
rect -14981 920 -14980 1240
rect -14660 920 -14659 1240
rect -14981 919 -14659 920
rect -15400 852 -15304 868
rect -14388 868 -14372 1292
rect -14308 868 -14292 1292
rect -13376 1292 -13280 1308
rect -13969 1240 -13647 1241
rect -13969 920 -13968 1240
rect -13648 920 -13647 1240
rect -13969 919 -13647 920
rect -14388 852 -14292 868
rect -13376 868 -13360 1292
rect -13296 868 -13280 1292
rect -12364 1292 -12268 1308
rect -12957 1240 -12635 1241
rect -12957 920 -12956 1240
rect -12636 920 -12635 1240
rect -12957 919 -12635 920
rect -13376 852 -13280 868
rect -12364 868 -12348 1292
rect -12284 868 -12268 1292
rect -11352 1292 -11256 1308
rect -11945 1240 -11623 1241
rect -11945 920 -11944 1240
rect -11624 920 -11623 1240
rect -11945 919 -11623 920
rect -12364 852 -12268 868
rect -11352 868 -11336 1292
rect -11272 868 -11256 1292
rect -10340 1292 -10244 1308
rect -10933 1240 -10611 1241
rect -10933 920 -10932 1240
rect -10612 920 -10611 1240
rect -10933 919 -10611 920
rect -11352 852 -11256 868
rect -10340 868 -10324 1292
rect -10260 868 -10244 1292
rect -9328 1292 -9232 1308
rect -9921 1240 -9599 1241
rect -9921 920 -9920 1240
rect -9600 920 -9599 1240
rect -9921 919 -9599 920
rect -10340 852 -10244 868
rect -9328 868 -9312 1292
rect -9248 868 -9232 1292
rect -8316 1292 -8220 1308
rect -8909 1240 -8587 1241
rect -8909 920 -8908 1240
rect -8588 920 -8587 1240
rect -8909 919 -8587 920
rect -9328 852 -9232 868
rect -8316 868 -8300 1292
rect -8236 868 -8220 1292
rect -7304 1292 -7208 1308
rect -7897 1240 -7575 1241
rect -7897 920 -7896 1240
rect -7576 920 -7575 1240
rect -7897 919 -7575 920
rect -8316 852 -8220 868
rect -7304 868 -7288 1292
rect -7224 868 -7208 1292
rect -6292 1292 -6196 1308
rect -6885 1240 -6563 1241
rect -6885 920 -6884 1240
rect -6564 920 -6563 1240
rect -6885 919 -6563 920
rect -7304 852 -7208 868
rect -6292 868 -6276 1292
rect -6212 868 -6196 1292
rect -5280 1292 -5184 1308
rect -5873 1240 -5551 1241
rect -5873 920 -5872 1240
rect -5552 920 -5551 1240
rect -5873 919 -5551 920
rect -6292 852 -6196 868
rect -5280 868 -5264 1292
rect -5200 868 -5184 1292
rect -4268 1292 -4172 1308
rect -4861 1240 -4539 1241
rect -4861 920 -4860 1240
rect -4540 920 -4539 1240
rect -4861 919 -4539 920
rect -5280 852 -5184 868
rect -4268 868 -4252 1292
rect -4188 868 -4172 1292
rect -3256 1292 -3160 1308
rect -3849 1240 -3527 1241
rect -3849 920 -3848 1240
rect -3528 920 -3527 1240
rect -3849 919 -3527 920
rect -4268 852 -4172 868
rect -3256 868 -3240 1292
rect -3176 868 -3160 1292
rect -2244 1292 -2148 1308
rect -2837 1240 -2515 1241
rect -2837 920 -2836 1240
rect -2516 920 -2515 1240
rect -2837 919 -2515 920
rect -3256 852 -3160 868
rect -2244 868 -2228 1292
rect -2164 868 -2148 1292
rect -1232 1292 -1136 1308
rect -1825 1240 -1503 1241
rect -1825 920 -1824 1240
rect -1504 920 -1503 1240
rect -1825 919 -1503 920
rect -2244 852 -2148 868
rect -1232 868 -1216 1292
rect -1152 868 -1136 1292
rect -220 1292 -124 1308
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -1232 852 -1136 868
rect -220 868 -204 1292
rect -140 868 -124 1292
rect 792 1292 888 1308
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -220 852 -124 868
rect 792 868 808 1292
rect 872 868 888 1292
rect 1804 1292 1900 1308
rect 1211 1240 1533 1241
rect 1211 920 1212 1240
rect 1532 920 1533 1240
rect 1211 919 1533 920
rect 792 852 888 868
rect 1804 868 1820 1292
rect 1884 868 1900 1292
rect 2816 1292 2912 1308
rect 2223 1240 2545 1241
rect 2223 920 2224 1240
rect 2544 920 2545 1240
rect 2223 919 2545 920
rect 1804 852 1900 868
rect 2816 868 2832 1292
rect 2896 868 2912 1292
rect 3828 1292 3924 1308
rect 3235 1240 3557 1241
rect 3235 920 3236 1240
rect 3556 920 3557 1240
rect 3235 919 3557 920
rect 2816 852 2912 868
rect 3828 868 3844 1292
rect 3908 868 3924 1292
rect 4840 1292 4936 1308
rect 4247 1240 4569 1241
rect 4247 920 4248 1240
rect 4568 920 4569 1240
rect 4247 919 4569 920
rect 3828 852 3924 868
rect 4840 868 4856 1292
rect 4920 868 4936 1292
rect 5852 1292 5948 1308
rect 5259 1240 5581 1241
rect 5259 920 5260 1240
rect 5580 920 5581 1240
rect 5259 919 5581 920
rect 4840 852 4936 868
rect 5852 868 5868 1292
rect 5932 868 5948 1292
rect 6864 1292 6960 1308
rect 6271 1240 6593 1241
rect 6271 920 6272 1240
rect 6592 920 6593 1240
rect 6271 919 6593 920
rect 5852 852 5948 868
rect 6864 868 6880 1292
rect 6944 868 6960 1292
rect 7876 1292 7972 1308
rect 7283 1240 7605 1241
rect 7283 920 7284 1240
rect 7604 920 7605 1240
rect 7283 919 7605 920
rect 6864 852 6960 868
rect 7876 868 7892 1292
rect 7956 868 7972 1292
rect 8888 1292 8984 1308
rect 8295 1240 8617 1241
rect 8295 920 8296 1240
rect 8616 920 8617 1240
rect 8295 919 8617 920
rect 7876 852 7972 868
rect 8888 868 8904 1292
rect 8968 868 8984 1292
rect 9900 1292 9996 1308
rect 9307 1240 9629 1241
rect 9307 920 9308 1240
rect 9628 920 9629 1240
rect 9307 919 9629 920
rect 8888 852 8984 868
rect 9900 868 9916 1292
rect 9980 868 9996 1292
rect 10912 1292 11008 1308
rect 10319 1240 10641 1241
rect 10319 920 10320 1240
rect 10640 920 10641 1240
rect 10319 919 10641 920
rect 9900 852 9996 868
rect 10912 868 10928 1292
rect 10992 868 11008 1292
rect 11924 1292 12020 1308
rect 11331 1240 11653 1241
rect 11331 920 11332 1240
rect 11652 920 11653 1240
rect 11331 919 11653 920
rect 10912 852 11008 868
rect 11924 868 11940 1292
rect 12004 868 12020 1292
rect 12936 1292 13032 1308
rect 12343 1240 12665 1241
rect 12343 920 12344 1240
rect 12664 920 12665 1240
rect 12343 919 12665 920
rect 11924 852 12020 868
rect 12936 868 12952 1292
rect 13016 868 13032 1292
rect 13948 1292 14044 1308
rect 13355 1240 13677 1241
rect 13355 920 13356 1240
rect 13676 920 13677 1240
rect 13355 919 13677 920
rect 12936 852 13032 868
rect 13948 868 13964 1292
rect 14028 868 14044 1292
rect 14960 1292 15056 1308
rect 14367 1240 14689 1241
rect 14367 920 14368 1240
rect 14688 920 14689 1240
rect 14367 919 14689 920
rect 13948 852 14044 868
rect 14960 868 14976 1292
rect 15040 868 15056 1292
rect 15972 1292 16068 1308
rect 15379 1240 15701 1241
rect 15379 920 15380 1240
rect 15700 920 15701 1240
rect 15379 919 15701 920
rect 14960 852 15056 868
rect 15972 868 15988 1292
rect 16052 868 16068 1292
rect 16984 1292 17080 1308
rect 16391 1240 16713 1241
rect 16391 920 16392 1240
rect 16712 920 16713 1240
rect 16391 919 16713 920
rect 15972 852 16068 868
rect 16984 868 17000 1292
rect 17064 868 17080 1292
rect 16984 852 17080 868
rect -16412 572 -16316 588
rect -17005 520 -16683 521
rect -17005 200 -17004 520
rect -16684 200 -16683 520
rect -17005 199 -16683 200
rect -16412 148 -16396 572
rect -16332 148 -16316 572
rect -15400 572 -15304 588
rect -15993 520 -15671 521
rect -15993 200 -15992 520
rect -15672 200 -15671 520
rect -15993 199 -15671 200
rect -16412 132 -16316 148
rect -15400 148 -15384 572
rect -15320 148 -15304 572
rect -14388 572 -14292 588
rect -14981 520 -14659 521
rect -14981 200 -14980 520
rect -14660 200 -14659 520
rect -14981 199 -14659 200
rect -15400 132 -15304 148
rect -14388 148 -14372 572
rect -14308 148 -14292 572
rect -13376 572 -13280 588
rect -13969 520 -13647 521
rect -13969 200 -13968 520
rect -13648 200 -13647 520
rect -13969 199 -13647 200
rect -14388 132 -14292 148
rect -13376 148 -13360 572
rect -13296 148 -13280 572
rect -12364 572 -12268 588
rect -12957 520 -12635 521
rect -12957 200 -12956 520
rect -12636 200 -12635 520
rect -12957 199 -12635 200
rect -13376 132 -13280 148
rect -12364 148 -12348 572
rect -12284 148 -12268 572
rect -11352 572 -11256 588
rect -11945 520 -11623 521
rect -11945 200 -11944 520
rect -11624 200 -11623 520
rect -11945 199 -11623 200
rect -12364 132 -12268 148
rect -11352 148 -11336 572
rect -11272 148 -11256 572
rect -10340 572 -10244 588
rect -10933 520 -10611 521
rect -10933 200 -10932 520
rect -10612 200 -10611 520
rect -10933 199 -10611 200
rect -11352 132 -11256 148
rect -10340 148 -10324 572
rect -10260 148 -10244 572
rect -9328 572 -9232 588
rect -9921 520 -9599 521
rect -9921 200 -9920 520
rect -9600 200 -9599 520
rect -9921 199 -9599 200
rect -10340 132 -10244 148
rect -9328 148 -9312 572
rect -9248 148 -9232 572
rect -8316 572 -8220 588
rect -8909 520 -8587 521
rect -8909 200 -8908 520
rect -8588 200 -8587 520
rect -8909 199 -8587 200
rect -9328 132 -9232 148
rect -8316 148 -8300 572
rect -8236 148 -8220 572
rect -7304 572 -7208 588
rect -7897 520 -7575 521
rect -7897 200 -7896 520
rect -7576 200 -7575 520
rect -7897 199 -7575 200
rect -8316 132 -8220 148
rect -7304 148 -7288 572
rect -7224 148 -7208 572
rect -6292 572 -6196 588
rect -6885 520 -6563 521
rect -6885 200 -6884 520
rect -6564 200 -6563 520
rect -6885 199 -6563 200
rect -7304 132 -7208 148
rect -6292 148 -6276 572
rect -6212 148 -6196 572
rect -5280 572 -5184 588
rect -5873 520 -5551 521
rect -5873 200 -5872 520
rect -5552 200 -5551 520
rect -5873 199 -5551 200
rect -6292 132 -6196 148
rect -5280 148 -5264 572
rect -5200 148 -5184 572
rect -4268 572 -4172 588
rect -4861 520 -4539 521
rect -4861 200 -4860 520
rect -4540 200 -4539 520
rect -4861 199 -4539 200
rect -5280 132 -5184 148
rect -4268 148 -4252 572
rect -4188 148 -4172 572
rect -3256 572 -3160 588
rect -3849 520 -3527 521
rect -3849 200 -3848 520
rect -3528 200 -3527 520
rect -3849 199 -3527 200
rect -4268 132 -4172 148
rect -3256 148 -3240 572
rect -3176 148 -3160 572
rect -2244 572 -2148 588
rect -2837 520 -2515 521
rect -2837 200 -2836 520
rect -2516 200 -2515 520
rect -2837 199 -2515 200
rect -3256 132 -3160 148
rect -2244 148 -2228 572
rect -2164 148 -2148 572
rect -1232 572 -1136 588
rect -1825 520 -1503 521
rect -1825 200 -1824 520
rect -1504 200 -1503 520
rect -1825 199 -1503 200
rect -2244 132 -2148 148
rect -1232 148 -1216 572
rect -1152 148 -1136 572
rect -220 572 -124 588
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -1232 132 -1136 148
rect -220 148 -204 572
rect -140 148 -124 572
rect 792 572 888 588
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -220 132 -124 148
rect 792 148 808 572
rect 872 148 888 572
rect 1804 572 1900 588
rect 1211 520 1533 521
rect 1211 200 1212 520
rect 1532 200 1533 520
rect 1211 199 1533 200
rect 792 132 888 148
rect 1804 148 1820 572
rect 1884 148 1900 572
rect 2816 572 2912 588
rect 2223 520 2545 521
rect 2223 200 2224 520
rect 2544 200 2545 520
rect 2223 199 2545 200
rect 1804 132 1900 148
rect 2816 148 2832 572
rect 2896 148 2912 572
rect 3828 572 3924 588
rect 3235 520 3557 521
rect 3235 200 3236 520
rect 3556 200 3557 520
rect 3235 199 3557 200
rect 2816 132 2912 148
rect 3828 148 3844 572
rect 3908 148 3924 572
rect 4840 572 4936 588
rect 4247 520 4569 521
rect 4247 200 4248 520
rect 4568 200 4569 520
rect 4247 199 4569 200
rect 3828 132 3924 148
rect 4840 148 4856 572
rect 4920 148 4936 572
rect 5852 572 5948 588
rect 5259 520 5581 521
rect 5259 200 5260 520
rect 5580 200 5581 520
rect 5259 199 5581 200
rect 4840 132 4936 148
rect 5852 148 5868 572
rect 5932 148 5948 572
rect 6864 572 6960 588
rect 6271 520 6593 521
rect 6271 200 6272 520
rect 6592 200 6593 520
rect 6271 199 6593 200
rect 5852 132 5948 148
rect 6864 148 6880 572
rect 6944 148 6960 572
rect 7876 572 7972 588
rect 7283 520 7605 521
rect 7283 200 7284 520
rect 7604 200 7605 520
rect 7283 199 7605 200
rect 6864 132 6960 148
rect 7876 148 7892 572
rect 7956 148 7972 572
rect 8888 572 8984 588
rect 8295 520 8617 521
rect 8295 200 8296 520
rect 8616 200 8617 520
rect 8295 199 8617 200
rect 7876 132 7972 148
rect 8888 148 8904 572
rect 8968 148 8984 572
rect 9900 572 9996 588
rect 9307 520 9629 521
rect 9307 200 9308 520
rect 9628 200 9629 520
rect 9307 199 9629 200
rect 8888 132 8984 148
rect 9900 148 9916 572
rect 9980 148 9996 572
rect 10912 572 11008 588
rect 10319 520 10641 521
rect 10319 200 10320 520
rect 10640 200 10641 520
rect 10319 199 10641 200
rect 9900 132 9996 148
rect 10912 148 10928 572
rect 10992 148 11008 572
rect 11924 572 12020 588
rect 11331 520 11653 521
rect 11331 200 11332 520
rect 11652 200 11653 520
rect 11331 199 11653 200
rect 10912 132 11008 148
rect 11924 148 11940 572
rect 12004 148 12020 572
rect 12936 572 13032 588
rect 12343 520 12665 521
rect 12343 200 12344 520
rect 12664 200 12665 520
rect 12343 199 12665 200
rect 11924 132 12020 148
rect 12936 148 12952 572
rect 13016 148 13032 572
rect 13948 572 14044 588
rect 13355 520 13677 521
rect 13355 200 13356 520
rect 13676 200 13677 520
rect 13355 199 13677 200
rect 12936 132 13032 148
rect 13948 148 13964 572
rect 14028 148 14044 572
rect 14960 572 15056 588
rect 14367 520 14689 521
rect 14367 200 14368 520
rect 14688 200 14689 520
rect 14367 199 14689 200
rect 13948 132 14044 148
rect 14960 148 14976 572
rect 15040 148 15056 572
rect 15972 572 16068 588
rect 15379 520 15701 521
rect 15379 200 15380 520
rect 15700 200 15701 520
rect 15379 199 15701 200
rect 14960 132 15056 148
rect 15972 148 15988 572
rect 16052 148 16068 572
rect 16984 572 17080 588
rect 16391 520 16713 521
rect 16391 200 16392 520
rect 16712 200 16713 520
rect 16391 199 16713 200
rect 15972 132 16068 148
rect 16984 148 17000 572
rect 17064 148 17080 572
rect 16984 132 17080 148
rect -16412 -148 -16316 -132
rect -17005 -200 -16683 -199
rect -17005 -520 -17004 -200
rect -16684 -520 -16683 -200
rect -17005 -521 -16683 -520
rect -16412 -572 -16396 -148
rect -16332 -572 -16316 -148
rect -15400 -148 -15304 -132
rect -15993 -200 -15671 -199
rect -15993 -520 -15992 -200
rect -15672 -520 -15671 -200
rect -15993 -521 -15671 -520
rect -16412 -588 -16316 -572
rect -15400 -572 -15384 -148
rect -15320 -572 -15304 -148
rect -14388 -148 -14292 -132
rect -14981 -200 -14659 -199
rect -14981 -520 -14980 -200
rect -14660 -520 -14659 -200
rect -14981 -521 -14659 -520
rect -15400 -588 -15304 -572
rect -14388 -572 -14372 -148
rect -14308 -572 -14292 -148
rect -13376 -148 -13280 -132
rect -13969 -200 -13647 -199
rect -13969 -520 -13968 -200
rect -13648 -520 -13647 -200
rect -13969 -521 -13647 -520
rect -14388 -588 -14292 -572
rect -13376 -572 -13360 -148
rect -13296 -572 -13280 -148
rect -12364 -148 -12268 -132
rect -12957 -200 -12635 -199
rect -12957 -520 -12956 -200
rect -12636 -520 -12635 -200
rect -12957 -521 -12635 -520
rect -13376 -588 -13280 -572
rect -12364 -572 -12348 -148
rect -12284 -572 -12268 -148
rect -11352 -148 -11256 -132
rect -11945 -200 -11623 -199
rect -11945 -520 -11944 -200
rect -11624 -520 -11623 -200
rect -11945 -521 -11623 -520
rect -12364 -588 -12268 -572
rect -11352 -572 -11336 -148
rect -11272 -572 -11256 -148
rect -10340 -148 -10244 -132
rect -10933 -200 -10611 -199
rect -10933 -520 -10932 -200
rect -10612 -520 -10611 -200
rect -10933 -521 -10611 -520
rect -11352 -588 -11256 -572
rect -10340 -572 -10324 -148
rect -10260 -572 -10244 -148
rect -9328 -148 -9232 -132
rect -9921 -200 -9599 -199
rect -9921 -520 -9920 -200
rect -9600 -520 -9599 -200
rect -9921 -521 -9599 -520
rect -10340 -588 -10244 -572
rect -9328 -572 -9312 -148
rect -9248 -572 -9232 -148
rect -8316 -148 -8220 -132
rect -8909 -200 -8587 -199
rect -8909 -520 -8908 -200
rect -8588 -520 -8587 -200
rect -8909 -521 -8587 -520
rect -9328 -588 -9232 -572
rect -8316 -572 -8300 -148
rect -8236 -572 -8220 -148
rect -7304 -148 -7208 -132
rect -7897 -200 -7575 -199
rect -7897 -520 -7896 -200
rect -7576 -520 -7575 -200
rect -7897 -521 -7575 -520
rect -8316 -588 -8220 -572
rect -7304 -572 -7288 -148
rect -7224 -572 -7208 -148
rect -6292 -148 -6196 -132
rect -6885 -200 -6563 -199
rect -6885 -520 -6884 -200
rect -6564 -520 -6563 -200
rect -6885 -521 -6563 -520
rect -7304 -588 -7208 -572
rect -6292 -572 -6276 -148
rect -6212 -572 -6196 -148
rect -5280 -148 -5184 -132
rect -5873 -200 -5551 -199
rect -5873 -520 -5872 -200
rect -5552 -520 -5551 -200
rect -5873 -521 -5551 -520
rect -6292 -588 -6196 -572
rect -5280 -572 -5264 -148
rect -5200 -572 -5184 -148
rect -4268 -148 -4172 -132
rect -4861 -200 -4539 -199
rect -4861 -520 -4860 -200
rect -4540 -520 -4539 -200
rect -4861 -521 -4539 -520
rect -5280 -588 -5184 -572
rect -4268 -572 -4252 -148
rect -4188 -572 -4172 -148
rect -3256 -148 -3160 -132
rect -3849 -200 -3527 -199
rect -3849 -520 -3848 -200
rect -3528 -520 -3527 -200
rect -3849 -521 -3527 -520
rect -4268 -588 -4172 -572
rect -3256 -572 -3240 -148
rect -3176 -572 -3160 -148
rect -2244 -148 -2148 -132
rect -2837 -200 -2515 -199
rect -2837 -520 -2836 -200
rect -2516 -520 -2515 -200
rect -2837 -521 -2515 -520
rect -3256 -588 -3160 -572
rect -2244 -572 -2228 -148
rect -2164 -572 -2148 -148
rect -1232 -148 -1136 -132
rect -1825 -200 -1503 -199
rect -1825 -520 -1824 -200
rect -1504 -520 -1503 -200
rect -1825 -521 -1503 -520
rect -2244 -588 -2148 -572
rect -1232 -572 -1216 -148
rect -1152 -572 -1136 -148
rect -220 -148 -124 -132
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -1232 -588 -1136 -572
rect -220 -572 -204 -148
rect -140 -572 -124 -148
rect 792 -148 888 -132
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -220 -588 -124 -572
rect 792 -572 808 -148
rect 872 -572 888 -148
rect 1804 -148 1900 -132
rect 1211 -200 1533 -199
rect 1211 -520 1212 -200
rect 1532 -520 1533 -200
rect 1211 -521 1533 -520
rect 792 -588 888 -572
rect 1804 -572 1820 -148
rect 1884 -572 1900 -148
rect 2816 -148 2912 -132
rect 2223 -200 2545 -199
rect 2223 -520 2224 -200
rect 2544 -520 2545 -200
rect 2223 -521 2545 -520
rect 1804 -588 1900 -572
rect 2816 -572 2832 -148
rect 2896 -572 2912 -148
rect 3828 -148 3924 -132
rect 3235 -200 3557 -199
rect 3235 -520 3236 -200
rect 3556 -520 3557 -200
rect 3235 -521 3557 -520
rect 2816 -588 2912 -572
rect 3828 -572 3844 -148
rect 3908 -572 3924 -148
rect 4840 -148 4936 -132
rect 4247 -200 4569 -199
rect 4247 -520 4248 -200
rect 4568 -520 4569 -200
rect 4247 -521 4569 -520
rect 3828 -588 3924 -572
rect 4840 -572 4856 -148
rect 4920 -572 4936 -148
rect 5852 -148 5948 -132
rect 5259 -200 5581 -199
rect 5259 -520 5260 -200
rect 5580 -520 5581 -200
rect 5259 -521 5581 -520
rect 4840 -588 4936 -572
rect 5852 -572 5868 -148
rect 5932 -572 5948 -148
rect 6864 -148 6960 -132
rect 6271 -200 6593 -199
rect 6271 -520 6272 -200
rect 6592 -520 6593 -200
rect 6271 -521 6593 -520
rect 5852 -588 5948 -572
rect 6864 -572 6880 -148
rect 6944 -572 6960 -148
rect 7876 -148 7972 -132
rect 7283 -200 7605 -199
rect 7283 -520 7284 -200
rect 7604 -520 7605 -200
rect 7283 -521 7605 -520
rect 6864 -588 6960 -572
rect 7876 -572 7892 -148
rect 7956 -572 7972 -148
rect 8888 -148 8984 -132
rect 8295 -200 8617 -199
rect 8295 -520 8296 -200
rect 8616 -520 8617 -200
rect 8295 -521 8617 -520
rect 7876 -588 7972 -572
rect 8888 -572 8904 -148
rect 8968 -572 8984 -148
rect 9900 -148 9996 -132
rect 9307 -200 9629 -199
rect 9307 -520 9308 -200
rect 9628 -520 9629 -200
rect 9307 -521 9629 -520
rect 8888 -588 8984 -572
rect 9900 -572 9916 -148
rect 9980 -572 9996 -148
rect 10912 -148 11008 -132
rect 10319 -200 10641 -199
rect 10319 -520 10320 -200
rect 10640 -520 10641 -200
rect 10319 -521 10641 -520
rect 9900 -588 9996 -572
rect 10912 -572 10928 -148
rect 10992 -572 11008 -148
rect 11924 -148 12020 -132
rect 11331 -200 11653 -199
rect 11331 -520 11332 -200
rect 11652 -520 11653 -200
rect 11331 -521 11653 -520
rect 10912 -588 11008 -572
rect 11924 -572 11940 -148
rect 12004 -572 12020 -148
rect 12936 -148 13032 -132
rect 12343 -200 12665 -199
rect 12343 -520 12344 -200
rect 12664 -520 12665 -200
rect 12343 -521 12665 -520
rect 11924 -588 12020 -572
rect 12936 -572 12952 -148
rect 13016 -572 13032 -148
rect 13948 -148 14044 -132
rect 13355 -200 13677 -199
rect 13355 -520 13356 -200
rect 13676 -520 13677 -200
rect 13355 -521 13677 -520
rect 12936 -588 13032 -572
rect 13948 -572 13964 -148
rect 14028 -572 14044 -148
rect 14960 -148 15056 -132
rect 14367 -200 14689 -199
rect 14367 -520 14368 -200
rect 14688 -520 14689 -200
rect 14367 -521 14689 -520
rect 13948 -588 14044 -572
rect 14960 -572 14976 -148
rect 15040 -572 15056 -148
rect 15972 -148 16068 -132
rect 15379 -200 15701 -199
rect 15379 -520 15380 -200
rect 15700 -520 15701 -200
rect 15379 -521 15701 -520
rect 14960 -588 15056 -572
rect 15972 -572 15988 -148
rect 16052 -572 16068 -148
rect 16984 -148 17080 -132
rect 16391 -200 16713 -199
rect 16391 -520 16392 -200
rect 16712 -520 16713 -200
rect 16391 -521 16713 -520
rect 15972 -588 16068 -572
rect 16984 -572 17000 -148
rect 17064 -572 17080 -148
rect 16984 -588 17080 -572
rect -16412 -868 -16316 -852
rect -17005 -920 -16683 -919
rect -17005 -1240 -17004 -920
rect -16684 -1240 -16683 -920
rect -17005 -1241 -16683 -1240
rect -16412 -1292 -16396 -868
rect -16332 -1292 -16316 -868
rect -15400 -868 -15304 -852
rect -15993 -920 -15671 -919
rect -15993 -1240 -15992 -920
rect -15672 -1240 -15671 -920
rect -15993 -1241 -15671 -1240
rect -16412 -1308 -16316 -1292
rect -15400 -1292 -15384 -868
rect -15320 -1292 -15304 -868
rect -14388 -868 -14292 -852
rect -14981 -920 -14659 -919
rect -14981 -1240 -14980 -920
rect -14660 -1240 -14659 -920
rect -14981 -1241 -14659 -1240
rect -15400 -1308 -15304 -1292
rect -14388 -1292 -14372 -868
rect -14308 -1292 -14292 -868
rect -13376 -868 -13280 -852
rect -13969 -920 -13647 -919
rect -13969 -1240 -13968 -920
rect -13648 -1240 -13647 -920
rect -13969 -1241 -13647 -1240
rect -14388 -1308 -14292 -1292
rect -13376 -1292 -13360 -868
rect -13296 -1292 -13280 -868
rect -12364 -868 -12268 -852
rect -12957 -920 -12635 -919
rect -12957 -1240 -12956 -920
rect -12636 -1240 -12635 -920
rect -12957 -1241 -12635 -1240
rect -13376 -1308 -13280 -1292
rect -12364 -1292 -12348 -868
rect -12284 -1292 -12268 -868
rect -11352 -868 -11256 -852
rect -11945 -920 -11623 -919
rect -11945 -1240 -11944 -920
rect -11624 -1240 -11623 -920
rect -11945 -1241 -11623 -1240
rect -12364 -1308 -12268 -1292
rect -11352 -1292 -11336 -868
rect -11272 -1292 -11256 -868
rect -10340 -868 -10244 -852
rect -10933 -920 -10611 -919
rect -10933 -1240 -10932 -920
rect -10612 -1240 -10611 -920
rect -10933 -1241 -10611 -1240
rect -11352 -1308 -11256 -1292
rect -10340 -1292 -10324 -868
rect -10260 -1292 -10244 -868
rect -9328 -868 -9232 -852
rect -9921 -920 -9599 -919
rect -9921 -1240 -9920 -920
rect -9600 -1240 -9599 -920
rect -9921 -1241 -9599 -1240
rect -10340 -1308 -10244 -1292
rect -9328 -1292 -9312 -868
rect -9248 -1292 -9232 -868
rect -8316 -868 -8220 -852
rect -8909 -920 -8587 -919
rect -8909 -1240 -8908 -920
rect -8588 -1240 -8587 -920
rect -8909 -1241 -8587 -1240
rect -9328 -1308 -9232 -1292
rect -8316 -1292 -8300 -868
rect -8236 -1292 -8220 -868
rect -7304 -868 -7208 -852
rect -7897 -920 -7575 -919
rect -7897 -1240 -7896 -920
rect -7576 -1240 -7575 -920
rect -7897 -1241 -7575 -1240
rect -8316 -1308 -8220 -1292
rect -7304 -1292 -7288 -868
rect -7224 -1292 -7208 -868
rect -6292 -868 -6196 -852
rect -6885 -920 -6563 -919
rect -6885 -1240 -6884 -920
rect -6564 -1240 -6563 -920
rect -6885 -1241 -6563 -1240
rect -7304 -1308 -7208 -1292
rect -6292 -1292 -6276 -868
rect -6212 -1292 -6196 -868
rect -5280 -868 -5184 -852
rect -5873 -920 -5551 -919
rect -5873 -1240 -5872 -920
rect -5552 -1240 -5551 -920
rect -5873 -1241 -5551 -1240
rect -6292 -1308 -6196 -1292
rect -5280 -1292 -5264 -868
rect -5200 -1292 -5184 -868
rect -4268 -868 -4172 -852
rect -4861 -920 -4539 -919
rect -4861 -1240 -4860 -920
rect -4540 -1240 -4539 -920
rect -4861 -1241 -4539 -1240
rect -5280 -1308 -5184 -1292
rect -4268 -1292 -4252 -868
rect -4188 -1292 -4172 -868
rect -3256 -868 -3160 -852
rect -3849 -920 -3527 -919
rect -3849 -1240 -3848 -920
rect -3528 -1240 -3527 -920
rect -3849 -1241 -3527 -1240
rect -4268 -1308 -4172 -1292
rect -3256 -1292 -3240 -868
rect -3176 -1292 -3160 -868
rect -2244 -868 -2148 -852
rect -2837 -920 -2515 -919
rect -2837 -1240 -2836 -920
rect -2516 -1240 -2515 -920
rect -2837 -1241 -2515 -1240
rect -3256 -1308 -3160 -1292
rect -2244 -1292 -2228 -868
rect -2164 -1292 -2148 -868
rect -1232 -868 -1136 -852
rect -1825 -920 -1503 -919
rect -1825 -1240 -1824 -920
rect -1504 -1240 -1503 -920
rect -1825 -1241 -1503 -1240
rect -2244 -1308 -2148 -1292
rect -1232 -1292 -1216 -868
rect -1152 -1292 -1136 -868
rect -220 -868 -124 -852
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -1232 -1308 -1136 -1292
rect -220 -1292 -204 -868
rect -140 -1292 -124 -868
rect 792 -868 888 -852
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -220 -1308 -124 -1292
rect 792 -1292 808 -868
rect 872 -1292 888 -868
rect 1804 -868 1900 -852
rect 1211 -920 1533 -919
rect 1211 -1240 1212 -920
rect 1532 -1240 1533 -920
rect 1211 -1241 1533 -1240
rect 792 -1308 888 -1292
rect 1804 -1292 1820 -868
rect 1884 -1292 1900 -868
rect 2816 -868 2912 -852
rect 2223 -920 2545 -919
rect 2223 -1240 2224 -920
rect 2544 -1240 2545 -920
rect 2223 -1241 2545 -1240
rect 1804 -1308 1900 -1292
rect 2816 -1292 2832 -868
rect 2896 -1292 2912 -868
rect 3828 -868 3924 -852
rect 3235 -920 3557 -919
rect 3235 -1240 3236 -920
rect 3556 -1240 3557 -920
rect 3235 -1241 3557 -1240
rect 2816 -1308 2912 -1292
rect 3828 -1292 3844 -868
rect 3908 -1292 3924 -868
rect 4840 -868 4936 -852
rect 4247 -920 4569 -919
rect 4247 -1240 4248 -920
rect 4568 -1240 4569 -920
rect 4247 -1241 4569 -1240
rect 3828 -1308 3924 -1292
rect 4840 -1292 4856 -868
rect 4920 -1292 4936 -868
rect 5852 -868 5948 -852
rect 5259 -920 5581 -919
rect 5259 -1240 5260 -920
rect 5580 -1240 5581 -920
rect 5259 -1241 5581 -1240
rect 4840 -1308 4936 -1292
rect 5852 -1292 5868 -868
rect 5932 -1292 5948 -868
rect 6864 -868 6960 -852
rect 6271 -920 6593 -919
rect 6271 -1240 6272 -920
rect 6592 -1240 6593 -920
rect 6271 -1241 6593 -1240
rect 5852 -1308 5948 -1292
rect 6864 -1292 6880 -868
rect 6944 -1292 6960 -868
rect 7876 -868 7972 -852
rect 7283 -920 7605 -919
rect 7283 -1240 7284 -920
rect 7604 -1240 7605 -920
rect 7283 -1241 7605 -1240
rect 6864 -1308 6960 -1292
rect 7876 -1292 7892 -868
rect 7956 -1292 7972 -868
rect 8888 -868 8984 -852
rect 8295 -920 8617 -919
rect 8295 -1240 8296 -920
rect 8616 -1240 8617 -920
rect 8295 -1241 8617 -1240
rect 7876 -1308 7972 -1292
rect 8888 -1292 8904 -868
rect 8968 -1292 8984 -868
rect 9900 -868 9996 -852
rect 9307 -920 9629 -919
rect 9307 -1240 9308 -920
rect 9628 -1240 9629 -920
rect 9307 -1241 9629 -1240
rect 8888 -1308 8984 -1292
rect 9900 -1292 9916 -868
rect 9980 -1292 9996 -868
rect 10912 -868 11008 -852
rect 10319 -920 10641 -919
rect 10319 -1240 10320 -920
rect 10640 -1240 10641 -920
rect 10319 -1241 10641 -1240
rect 9900 -1308 9996 -1292
rect 10912 -1292 10928 -868
rect 10992 -1292 11008 -868
rect 11924 -868 12020 -852
rect 11331 -920 11653 -919
rect 11331 -1240 11332 -920
rect 11652 -1240 11653 -920
rect 11331 -1241 11653 -1240
rect 10912 -1308 11008 -1292
rect 11924 -1292 11940 -868
rect 12004 -1292 12020 -868
rect 12936 -868 13032 -852
rect 12343 -920 12665 -919
rect 12343 -1240 12344 -920
rect 12664 -1240 12665 -920
rect 12343 -1241 12665 -1240
rect 11924 -1308 12020 -1292
rect 12936 -1292 12952 -868
rect 13016 -1292 13032 -868
rect 13948 -868 14044 -852
rect 13355 -920 13677 -919
rect 13355 -1240 13356 -920
rect 13676 -1240 13677 -920
rect 13355 -1241 13677 -1240
rect 12936 -1308 13032 -1292
rect 13948 -1292 13964 -868
rect 14028 -1292 14044 -868
rect 14960 -868 15056 -852
rect 14367 -920 14689 -919
rect 14367 -1240 14368 -920
rect 14688 -1240 14689 -920
rect 14367 -1241 14689 -1240
rect 13948 -1308 14044 -1292
rect 14960 -1292 14976 -868
rect 15040 -1292 15056 -868
rect 15972 -868 16068 -852
rect 15379 -920 15701 -919
rect 15379 -1240 15380 -920
rect 15700 -1240 15701 -920
rect 15379 -1241 15701 -1240
rect 14960 -1308 15056 -1292
rect 15972 -1292 15988 -868
rect 16052 -1292 16068 -868
rect 16984 -868 17080 -852
rect 16391 -920 16713 -919
rect 16391 -1240 16392 -920
rect 16712 -1240 16713 -920
rect 16391 -1241 16713 -1240
rect 15972 -1308 16068 -1292
rect 16984 -1292 17000 -868
rect 17064 -1292 17080 -868
rect 16984 -1308 17080 -1292
rect -16412 -1588 -16316 -1572
rect -17005 -1640 -16683 -1639
rect -17005 -1960 -17004 -1640
rect -16684 -1960 -16683 -1640
rect -17005 -1961 -16683 -1960
rect -16412 -2012 -16396 -1588
rect -16332 -2012 -16316 -1588
rect -15400 -1588 -15304 -1572
rect -15993 -1640 -15671 -1639
rect -15993 -1960 -15992 -1640
rect -15672 -1960 -15671 -1640
rect -15993 -1961 -15671 -1960
rect -16412 -2028 -16316 -2012
rect -15400 -2012 -15384 -1588
rect -15320 -2012 -15304 -1588
rect -14388 -1588 -14292 -1572
rect -14981 -1640 -14659 -1639
rect -14981 -1960 -14980 -1640
rect -14660 -1960 -14659 -1640
rect -14981 -1961 -14659 -1960
rect -15400 -2028 -15304 -2012
rect -14388 -2012 -14372 -1588
rect -14308 -2012 -14292 -1588
rect -13376 -1588 -13280 -1572
rect -13969 -1640 -13647 -1639
rect -13969 -1960 -13968 -1640
rect -13648 -1960 -13647 -1640
rect -13969 -1961 -13647 -1960
rect -14388 -2028 -14292 -2012
rect -13376 -2012 -13360 -1588
rect -13296 -2012 -13280 -1588
rect -12364 -1588 -12268 -1572
rect -12957 -1640 -12635 -1639
rect -12957 -1960 -12956 -1640
rect -12636 -1960 -12635 -1640
rect -12957 -1961 -12635 -1960
rect -13376 -2028 -13280 -2012
rect -12364 -2012 -12348 -1588
rect -12284 -2012 -12268 -1588
rect -11352 -1588 -11256 -1572
rect -11945 -1640 -11623 -1639
rect -11945 -1960 -11944 -1640
rect -11624 -1960 -11623 -1640
rect -11945 -1961 -11623 -1960
rect -12364 -2028 -12268 -2012
rect -11352 -2012 -11336 -1588
rect -11272 -2012 -11256 -1588
rect -10340 -1588 -10244 -1572
rect -10933 -1640 -10611 -1639
rect -10933 -1960 -10932 -1640
rect -10612 -1960 -10611 -1640
rect -10933 -1961 -10611 -1960
rect -11352 -2028 -11256 -2012
rect -10340 -2012 -10324 -1588
rect -10260 -2012 -10244 -1588
rect -9328 -1588 -9232 -1572
rect -9921 -1640 -9599 -1639
rect -9921 -1960 -9920 -1640
rect -9600 -1960 -9599 -1640
rect -9921 -1961 -9599 -1960
rect -10340 -2028 -10244 -2012
rect -9328 -2012 -9312 -1588
rect -9248 -2012 -9232 -1588
rect -8316 -1588 -8220 -1572
rect -8909 -1640 -8587 -1639
rect -8909 -1960 -8908 -1640
rect -8588 -1960 -8587 -1640
rect -8909 -1961 -8587 -1960
rect -9328 -2028 -9232 -2012
rect -8316 -2012 -8300 -1588
rect -8236 -2012 -8220 -1588
rect -7304 -1588 -7208 -1572
rect -7897 -1640 -7575 -1639
rect -7897 -1960 -7896 -1640
rect -7576 -1960 -7575 -1640
rect -7897 -1961 -7575 -1960
rect -8316 -2028 -8220 -2012
rect -7304 -2012 -7288 -1588
rect -7224 -2012 -7208 -1588
rect -6292 -1588 -6196 -1572
rect -6885 -1640 -6563 -1639
rect -6885 -1960 -6884 -1640
rect -6564 -1960 -6563 -1640
rect -6885 -1961 -6563 -1960
rect -7304 -2028 -7208 -2012
rect -6292 -2012 -6276 -1588
rect -6212 -2012 -6196 -1588
rect -5280 -1588 -5184 -1572
rect -5873 -1640 -5551 -1639
rect -5873 -1960 -5872 -1640
rect -5552 -1960 -5551 -1640
rect -5873 -1961 -5551 -1960
rect -6292 -2028 -6196 -2012
rect -5280 -2012 -5264 -1588
rect -5200 -2012 -5184 -1588
rect -4268 -1588 -4172 -1572
rect -4861 -1640 -4539 -1639
rect -4861 -1960 -4860 -1640
rect -4540 -1960 -4539 -1640
rect -4861 -1961 -4539 -1960
rect -5280 -2028 -5184 -2012
rect -4268 -2012 -4252 -1588
rect -4188 -2012 -4172 -1588
rect -3256 -1588 -3160 -1572
rect -3849 -1640 -3527 -1639
rect -3849 -1960 -3848 -1640
rect -3528 -1960 -3527 -1640
rect -3849 -1961 -3527 -1960
rect -4268 -2028 -4172 -2012
rect -3256 -2012 -3240 -1588
rect -3176 -2012 -3160 -1588
rect -2244 -1588 -2148 -1572
rect -2837 -1640 -2515 -1639
rect -2837 -1960 -2836 -1640
rect -2516 -1960 -2515 -1640
rect -2837 -1961 -2515 -1960
rect -3256 -2028 -3160 -2012
rect -2244 -2012 -2228 -1588
rect -2164 -2012 -2148 -1588
rect -1232 -1588 -1136 -1572
rect -1825 -1640 -1503 -1639
rect -1825 -1960 -1824 -1640
rect -1504 -1960 -1503 -1640
rect -1825 -1961 -1503 -1960
rect -2244 -2028 -2148 -2012
rect -1232 -2012 -1216 -1588
rect -1152 -2012 -1136 -1588
rect -220 -1588 -124 -1572
rect -813 -1640 -491 -1639
rect -813 -1960 -812 -1640
rect -492 -1960 -491 -1640
rect -813 -1961 -491 -1960
rect -1232 -2028 -1136 -2012
rect -220 -2012 -204 -1588
rect -140 -2012 -124 -1588
rect 792 -1588 888 -1572
rect 199 -1640 521 -1639
rect 199 -1960 200 -1640
rect 520 -1960 521 -1640
rect 199 -1961 521 -1960
rect -220 -2028 -124 -2012
rect 792 -2012 808 -1588
rect 872 -2012 888 -1588
rect 1804 -1588 1900 -1572
rect 1211 -1640 1533 -1639
rect 1211 -1960 1212 -1640
rect 1532 -1960 1533 -1640
rect 1211 -1961 1533 -1960
rect 792 -2028 888 -2012
rect 1804 -2012 1820 -1588
rect 1884 -2012 1900 -1588
rect 2816 -1588 2912 -1572
rect 2223 -1640 2545 -1639
rect 2223 -1960 2224 -1640
rect 2544 -1960 2545 -1640
rect 2223 -1961 2545 -1960
rect 1804 -2028 1900 -2012
rect 2816 -2012 2832 -1588
rect 2896 -2012 2912 -1588
rect 3828 -1588 3924 -1572
rect 3235 -1640 3557 -1639
rect 3235 -1960 3236 -1640
rect 3556 -1960 3557 -1640
rect 3235 -1961 3557 -1960
rect 2816 -2028 2912 -2012
rect 3828 -2012 3844 -1588
rect 3908 -2012 3924 -1588
rect 4840 -1588 4936 -1572
rect 4247 -1640 4569 -1639
rect 4247 -1960 4248 -1640
rect 4568 -1960 4569 -1640
rect 4247 -1961 4569 -1960
rect 3828 -2028 3924 -2012
rect 4840 -2012 4856 -1588
rect 4920 -2012 4936 -1588
rect 5852 -1588 5948 -1572
rect 5259 -1640 5581 -1639
rect 5259 -1960 5260 -1640
rect 5580 -1960 5581 -1640
rect 5259 -1961 5581 -1960
rect 4840 -2028 4936 -2012
rect 5852 -2012 5868 -1588
rect 5932 -2012 5948 -1588
rect 6864 -1588 6960 -1572
rect 6271 -1640 6593 -1639
rect 6271 -1960 6272 -1640
rect 6592 -1960 6593 -1640
rect 6271 -1961 6593 -1960
rect 5852 -2028 5948 -2012
rect 6864 -2012 6880 -1588
rect 6944 -2012 6960 -1588
rect 7876 -1588 7972 -1572
rect 7283 -1640 7605 -1639
rect 7283 -1960 7284 -1640
rect 7604 -1960 7605 -1640
rect 7283 -1961 7605 -1960
rect 6864 -2028 6960 -2012
rect 7876 -2012 7892 -1588
rect 7956 -2012 7972 -1588
rect 8888 -1588 8984 -1572
rect 8295 -1640 8617 -1639
rect 8295 -1960 8296 -1640
rect 8616 -1960 8617 -1640
rect 8295 -1961 8617 -1960
rect 7876 -2028 7972 -2012
rect 8888 -2012 8904 -1588
rect 8968 -2012 8984 -1588
rect 9900 -1588 9996 -1572
rect 9307 -1640 9629 -1639
rect 9307 -1960 9308 -1640
rect 9628 -1960 9629 -1640
rect 9307 -1961 9629 -1960
rect 8888 -2028 8984 -2012
rect 9900 -2012 9916 -1588
rect 9980 -2012 9996 -1588
rect 10912 -1588 11008 -1572
rect 10319 -1640 10641 -1639
rect 10319 -1960 10320 -1640
rect 10640 -1960 10641 -1640
rect 10319 -1961 10641 -1960
rect 9900 -2028 9996 -2012
rect 10912 -2012 10928 -1588
rect 10992 -2012 11008 -1588
rect 11924 -1588 12020 -1572
rect 11331 -1640 11653 -1639
rect 11331 -1960 11332 -1640
rect 11652 -1960 11653 -1640
rect 11331 -1961 11653 -1960
rect 10912 -2028 11008 -2012
rect 11924 -2012 11940 -1588
rect 12004 -2012 12020 -1588
rect 12936 -1588 13032 -1572
rect 12343 -1640 12665 -1639
rect 12343 -1960 12344 -1640
rect 12664 -1960 12665 -1640
rect 12343 -1961 12665 -1960
rect 11924 -2028 12020 -2012
rect 12936 -2012 12952 -1588
rect 13016 -2012 13032 -1588
rect 13948 -1588 14044 -1572
rect 13355 -1640 13677 -1639
rect 13355 -1960 13356 -1640
rect 13676 -1960 13677 -1640
rect 13355 -1961 13677 -1960
rect 12936 -2028 13032 -2012
rect 13948 -2012 13964 -1588
rect 14028 -2012 14044 -1588
rect 14960 -1588 15056 -1572
rect 14367 -1640 14689 -1639
rect 14367 -1960 14368 -1640
rect 14688 -1960 14689 -1640
rect 14367 -1961 14689 -1960
rect 13948 -2028 14044 -2012
rect 14960 -2012 14976 -1588
rect 15040 -2012 15056 -1588
rect 15972 -1588 16068 -1572
rect 15379 -1640 15701 -1639
rect 15379 -1960 15380 -1640
rect 15700 -1960 15701 -1640
rect 15379 -1961 15701 -1960
rect 14960 -2028 15056 -2012
rect 15972 -2012 15988 -1588
rect 16052 -2012 16068 -1588
rect 16984 -1588 17080 -1572
rect 16391 -1640 16713 -1639
rect 16391 -1960 16392 -1640
rect 16712 -1960 16713 -1640
rect 16391 -1961 16713 -1960
rect 15972 -2028 16068 -2012
rect 16984 -2012 17000 -1588
rect 17064 -2012 17080 -1588
rect 16984 -2028 17080 -2012
rect -16412 -2308 -16316 -2292
rect -17005 -2360 -16683 -2359
rect -17005 -2680 -17004 -2360
rect -16684 -2680 -16683 -2360
rect -17005 -2681 -16683 -2680
rect -16412 -2732 -16396 -2308
rect -16332 -2732 -16316 -2308
rect -15400 -2308 -15304 -2292
rect -15993 -2360 -15671 -2359
rect -15993 -2680 -15992 -2360
rect -15672 -2680 -15671 -2360
rect -15993 -2681 -15671 -2680
rect -16412 -2748 -16316 -2732
rect -15400 -2732 -15384 -2308
rect -15320 -2732 -15304 -2308
rect -14388 -2308 -14292 -2292
rect -14981 -2360 -14659 -2359
rect -14981 -2680 -14980 -2360
rect -14660 -2680 -14659 -2360
rect -14981 -2681 -14659 -2680
rect -15400 -2748 -15304 -2732
rect -14388 -2732 -14372 -2308
rect -14308 -2732 -14292 -2308
rect -13376 -2308 -13280 -2292
rect -13969 -2360 -13647 -2359
rect -13969 -2680 -13968 -2360
rect -13648 -2680 -13647 -2360
rect -13969 -2681 -13647 -2680
rect -14388 -2748 -14292 -2732
rect -13376 -2732 -13360 -2308
rect -13296 -2732 -13280 -2308
rect -12364 -2308 -12268 -2292
rect -12957 -2360 -12635 -2359
rect -12957 -2680 -12956 -2360
rect -12636 -2680 -12635 -2360
rect -12957 -2681 -12635 -2680
rect -13376 -2748 -13280 -2732
rect -12364 -2732 -12348 -2308
rect -12284 -2732 -12268 -2308
rect -11352 -2308 -11256 -2292
rect -11945 -2360 -11623 -2359
rect -11945 -2680 -11944 -2360
rect -11624 -2680 -11623 -2360
rect -11945 -2681 -11623 -2680
rect -12364 -2748 -12268 -2732
rect -11352 -2732 -11336 -2308
rect -11272 -2732 -11256 -2308
rect -10340 -2308 -10244 -2292
rect -10933 -2360 -10611 -2359
rect -10933 -2680 -10932 -2360
rect -10612 -2680 -10611 -2360
rect -10933 -2681 -10611 -2680
rect -11352 -2748 -11256 -2732
rect -10340 -2732 -10324 -2308
rect -10260 -2732 -10244 -2308
rect -9328 -2308 -9232 -2292
rect -9921 -2360 -9599 -2359
rect -9921 -2680 -9920 -2360
rect -9600 -2680 -9599 -2360
rect -9921 -2681 -9599 -2680
rect -10340 -2748 -10244 -2732
rect -9328 -2732 -9312 -2308
rect -9248 -2732 -9232 -2308
rect -8316 -2308 -8220 -2292
rect -8909 -2360 -8587 -2359
rect -8909 -2680 -8908 -2360
rect -8588 -2680 -8587 -2360
rect -8909 -2681 -8587 -2680
rect -9328 -2748 -9232 -2732
rect -8316 -2732 -8300 -2308
rect -8236 -2732 -8220 -2308
rect -7304 -2308 -7208 -2292
rect -7897 -2360 -7575 -2359
rect -7897 -2680 -7896 -2360
rect -7576 -2680 -7575 -2360
rect -7897 -2681 -7575 -2680
rect -8316 -2748 -8220 -2732
rect -7304 -2732 -7288 -2308
rect -7224 -2732 -7208 -2308
rect -6292 -2308 -6196 -2292
rect -6885 -2360 -6563 -2359
rect -6885 -2680 -6884 -2360
rect -6564 -2680 -6563 -2360
rect -6885 -2681 -6563 -2680
rect -7304 -2748 -7208 -2732
rect -6292 -2732 -6276 -2308
rect -6212 -2732 -6196 -2308
rect -5280 -2308 -5184 -2292
rect -5873 -2360 -5551 -2359
rect -5873 -2680 -5872 -2360
rect -5552 -2680 -5551 -2360
rect -5873 -2681 -5551 -2680
rect -6292 -2748 -6196 -2732
rect -5280 -2732 -5264 -2308
rect -5200 -2732 -5184 -2308
rect -4268 -2308 -4172 -2292
rect -4861 -2360 -4539 -2359
rect -4861 -2680 -4860 -2360
rect -4540 -2680 -4539 -2360
rect -4861 -2681 -4539 -2680
rect -5280 -2748 -5184 -2732
rect -4268 -2732 -4252 -2308
rect -4188 -2732 -4172 -2308
rect -3256 -2308 -3160 -2292
rect -3849 -2360 -3527 -2359
rect -3849 -2680 -3848 -2360
rect -3528 -2680 -3527 -2360
rect -3849 -2681 -3527 -2680
rect -4268 -2748 -4172 -2732
rect -3256 -2732 -3240 -2308
rect -3176 -2732 -3160 -2308
rect -2244 -2308 -2148 -2292
rect -2837 -2360 -2515 -2359
rect -2837 -2680 -2836 -2360
rect -2516 -2680 -2515 -2360
rect -2837 -2681 -2515 -2680
rect -3256 -2748 -3160 -2732
rect -2244 -2732 -2228 -2308
rect -2164 -2732 -2148 -2308
rect -1232 -2308 -1136 -2292
rect -1825 -2360 -1503 -2359
rect -1825 -2680 -1824 -2360
rect -1504 -2680 -1503 -2360
rect -1825 -2681 -1503 -2680
rect -2244 -2748 -2148 -2732
rect -1232 -2732 -1216 -2308
rect -1152 -2732 -1136 -2308
rect -220 -2308 -124 -2292
rect -813 -2360 -491 -2359
rect -813 -2680 -812 -2360
rect -492 -2680 -491 -2360
rect -813 -2681 -491 -2680
rect -1232 -2748 -1136 -2732
rect -220 -2732 -204 -2308
rect -140 -2732 -124 -2308
rect 792 -2308 888 -2292
rect 199 -2360 521 -2359
rect 199 -2680 200 -2360
rect 520 -2680 521 -2360
rect 199 -2681 521 -2680
rect -220 -2748 -124 -2732
rect 792 -2732 808 -2308
rect 872 -2732 888 -2308
rect 1804 -2308 1900 -2292
rect 1211 -2360 1533 -2359
rect 1211 -2680 1212 -2360
rect 1532 -2680 1533 -2360
rect 1211 -2681 1533 -2680
rect 792 -2748 888 -2732
rect 1804 -2732 1820 -2308
rect 1884 -2732 1900 -2308
rect 2816 -2308 2912 -2292
rect 2223 -2360 2545 -2359
rect 2223 -2680 2224 -2360
rect 2544 -2680 2545 -2360
rect 2223 -2681 2545 -2680
rect 1804 -2748 1900 -2732
rect 2816 -2732 2832 -2308
rect 2896 -2732 2912 -2308
rect 3828 -2308 3924 -2292
rect 3235 -2360 3557 -2359
rect 3235 -2680 3236 -2360
rect 3556 -2680 3557 -2360
rect 3235 -2681 3557 -2680
rect 2816 -2748 2912 -2732
rect 3828 -2732 3844 -2308
rect 3908 -2732 3924 -2308
rect 4840 -2308 4936 -2292
rect 4247 -2360 4569 -2359
rect 4247 -2680 4248 -2360
rect 4568 -2680 4569 -2360
rect 4247 -2681 4569 -2680
rect 3828 -2748 3924 -2732
rect 4840 -2732 4856 -2308
rect 4920 -2732 4936 -2308
rect 5852 -2308 5948 -2292
rect 5259 -2360 5581 -2359
rect 5259 -2680 5260 -2360
rect 5580 -2680 5581 -2360
rect 5259 -2681 5581 -2680
rect 4840 -2748 4936 -2732
rect 5852 -2732 5868 -2308
rect 5932 -2732 5948 -2308
rect 6864 -2308 6960 -2292
rect 6271 -2360 6593 -2359
rect 6271 -2680 6272 -2360
rect 6592 -2680 6593 -2360
rect 6271 -2681 6593 -2680
rect 5852 -2748 5948 -2732
rect 6864 -2732 6880 -2308
rect 6944 -2732 6960 -2308
rect 7876 -2308 7972 -2292
rect 7283 -2360 7605 -2359
rect 7283 -2680 7284 -2360
rect 7604 -2680 7605 -2360
rect 7283 -2681 7605 -2680
rect 6864 -2748 6960 -2732
rect 7876 -2732 7892 -2308
rect 7956 -2732 7972 -2308
rect 8888 -2308 8984 -2292
rect 8295 -2360 8617 -2359
rect 8295 -2680 8296 -2360
rect 8616 -2680 8617 -2360
rect 8295 -2681 8617 -2680
rect 7876 -2748 7972 -2732
rect 8888 -2732 8904 -2308
rect 8968 -2732 8984 -2308
rect 9900 -2308 9996 -2292
rect 9307 -2360 9629 -2359
rect 9307 -2680 9308 -2360
rect 9628 -2680 9629 -2360
rect 9307 -2681 9629 -2680
rect 8888 -2748 8984 -2732
rect 9900 -2732 9916 -2308
rect 9980 -2732 9996 -2308
rect 10912 -2308 11008 -2292
rect 10319 -2360 10641 -2359
rect 10319 -2680 10320 -2360
rect 10640 -2680 10641 -2360
rect 10319 -2681 10641 -2680
rect 9900 -2748 9996 -2732
rect 10912 -2732 10928 -2308
rect 10992 -2732 11008 -2308
rect 11924 -2308 12020 -2292
rect 11331 -2360 11653 -2359
rect 11331 -2680 11332 -2360
rect 11652 -2680 11653 -2360
rect 11331 -2681 11653 -2680
rect 10912 -2748 11008 -2732
rect 11924 -2732 11940 -2308
rect 12004 -2732 12020 -2308
rect 12936 -2308 13032 -2292
rect 12343 -2360 12665 -2359
rect 12343 -2680 12344 -2360
rect 12664 -2680 12665 -2360
rect 12343 -2681 12665 -2680
rect 11924 -2748 12020 -2732
rect 12936 -2732 12952 -2308
rect 13016 -2732 13032 -2308
rect 13948 -2308 14044 -2292
rect 13355 -2360 13677 -2359
rect 13355 -2680 13356 -2360
rect 13676 -2680 13677 -2360
rect 13355 -2681 13677 -2680
rect 12936 -2748 13032 -2732
rect 13948 -2732 13964 -2308
rect 14028 -2732 14044 -2308
rect 14960 -2308 15056 -2292
rect 14367 -2360 14689 -2359
rect 14367 -2680 14368 -2360
rect 14688 -2680 14689 -2360
rect 14367 -2681 14689 -2680
rect 13948 -2748 14044 -2732
rect 14960 -2732 14976 -2308
rect 15040 -2732 15056 -2308
rect 15972 -2308 16068 -2292
rect 15379 -2360 15701 -2359
rect 15379 -2680 15380 -2360
rect 15700 -2680 15701 -2360
rect 15379 -2681 15701 -2680
rect 14960 -2748 15056 -2732
rect 15972 -2732 15988 -2308
rect 16052 -2732 16068 -2308
rect 16984 -2308 17080 -2292
rect 16391 -2360 16713 -2359
rect 16391 -2680 16392 -2360
rect 16712 -2680 16713 -2360
rect 16391 -2681 16713 -2680
rect 15972 -2748 16068 -2732
rect 16984 -2732 17000 -2308
rect 17064 -2732 17080 -2308
rect 16984 -2748 17080 -2732
rect -16412 -3028 -16316 -3012
rect -17005 -3080 -16683 -3079
rect -17005 -3400 -17004 -3080
rect -16684 -3400 -16683 -3080
rect -17005 -3401 -16683 -3400
rect -16412 -3452 -16396 -3028
rect -16332 -3452 -16316 -3028
rect -15400 -3028 -15304 -3012
rect -15993 -3080 -15671 -3079
rect -15993 -3400 -15992 -3080
rect -15672 -3400 -15671 -3080
rect -15993 -3401 -15671 -3400
rect -16412 -3468 -16316 -3452
rect -15400 -3452 -15384 -3028
rect -15320 -3452 -15304 -3028
rect -14388 -3028 -14292 -3012
rect -14981 -3080 -14659 -3079
rect -14981 -3400 -14980 -3080
rect -14660 -3400 -14659 -3080
rect -14981 -3401 -14659 -3400
rect -15400 -3468 -15304 -3452
rect -14388 -3452 -14372 -3028
rect -14308 -3452 -14292 -3028
rect -13376 -3028 -13280 -3012
rect -13969 -3080 -13647 -3079
rect -13969 -3400 -13968 -3080
rect -13648 -3400 -13647 -3080
rect -13969 -3401 -13647 -3400
rect -14388 -3468 -14292 -3452
rect -13376 -3452 -13360 -3028
rect -13296 -3452 -13280 -3028
rect -12364 -3028 -12268 -3012
rect -12957 -3080 -12635 -3079
rect -12957 -3400 -12956 -3080
rect -12636 -3400 -12635 -3080
rect -12957 -3401 -12635 -3400
rect -13376 -3468 -13280 -3452
rect -12364 -3452 -12348 -3028
rect -12284 -3452 -12268 -3028
rect -11352 -3028 -11256 -3012
rect -11945 -3080 -11623 -3079
rect -11945 -3400 -11944 -3080
rect -11624 -3400 -11623 -3080
rect -11945 -3401 -11623 -3400
rect -12364 -3468 -12268 -3452
rect -11352 -3452 -11336 -3028
rect -11272 -3452 -11256 -3028
rect -10340 -3028 -10244 -3012
rect -10933 -3080 -10611 -3079
rect -10933 -3400 -10932 -3080
rect -10612 -3400 -10611 -3080
rect -10933 -3401 -10611 -3400
rect -11352 -3468 -11256 -3452
rect -10340 -3452 -10324 -3028
rect -10260 -3452 -10244 -3028
rect -9328 -3028 -9232 -3012
rect -9921 -3080 -9599 -3079
rect -9921 -3400 -9920 -3080
rect -9600 -3400 -9599 -3080
rect -9921 -3401 -9599 -3400
rect -10340 -3468 -10244 -3452
rect -9328 -3452 -9312 -3028
rect -9248 -3452 -9232 -3028
rect -8316 -3028 -8220 -3012
rect -8909 -3080 -8587 -3079
rect -8909 -3400 -8908 -3080
rect -8588 -3400 -8587 -3080
rect -8909 -3401 -8587 -3400
rect -9328 -3468 -9232 -3452
rect -8316 -3452 -8300 -3028
rect -8236 -3452 -8220 -3028
rect -7304 -3028 -7208 -3012
rect -7897 -3080 -7575 -3079
rect -7897 -3400 -7896 -3080
rect -7576 -3400 -7575 -3080
rect -7897 -3401 -7575 -3400
rect -8316 -3468 -8220 -3452
rect -7304 -3452 -7288 -3028
rect -7224 -3452 -7208 -3028
rect -6292 -3028 -6196 -3012
rect -6885 -3080 -6563 -3079
rect -6885 -3400 -6884 -3080
rect -6564 -3400 -6563 -3080
rect -6885 -3401 -6563 -3400
rect -7304 -3468 -7208 -3452
rect -6292 -3452 -6276 -3028
rect -6212 -3452 -6196 -3028
rect -5280 -3028 -5184 -3012
rect -5873 -3080 -5551 -3079
rect -5873 -3400 -5872 -3080
rect -5552 -3400 -5551 -3080
rect -5873 -3401 -5551 -3400
rect -6292 -3468 -6196 -3452
rect -5280 -3452 -5264 -3028
rect -5200 -3452 -5184 -3028
rect -4268 -3028 -4172 -3012
rect -4861 -3080 -4539 -3079
rect -4861 -3400 -4860 -3080
rect -4540 -3400 -4539 -3080
rect -4861 -3401 -4539 -3400
rect -5280 -3468 -5184 -3452
rect -4268 -3452 -4252 -3028
rect -4188 -3452 -4172 -3028
rect -3256 -3028 -3160 -3012
rect -3849 -3080 -3527 -3079
rect -3849 -3400 -3848 -3080
rect -3528 -3400 -3527 -3080
rect -3849 -3401 -3527 -3400
rect -4268 -3468 -4172 -3452
rect -3256 -3452 -3240 -3028
rect -3176 -3452 -3160 -3028
rect -2244 -3028 -2148 -3012
rect -2837 -3080 -2515 -3079
rect -2837 -3400 -2836 -3080
rect -2516 -3400 -2515 -3080
rect -2837 -3401 -2515 -3400
rect -3256 -3468 -3160 -3452
rect -2244 -3452 -2228 -3028
rect -2164 -3452 -2148 -3028
rect -1232 -3028 -1136 -3012
rect -1825 -3080 -1503 -3079
rect -1825 -3400 -1824 -3080
rect -1504 -3400 -1503 -3080
rect -1825 -3401 -1503 -3400
rect -2244 -3468 -2148 -3452
rect -1232 -3452 -1216 -3028
rect -1152 -3452 -1136 -3028
rect -220 -3028 -124 -3012
rect -813 -3080 -491 -3079
rect -813 -3400 -812 -3080
rect -492 -3400 -491 -3080
rect -813 -3401 -491 -3400
rect -1232 -3468 -1136 -3452
rect -220 -3452 -204 -3028
rect -140 -3452 -124 -3028
rect 792 -3028 888 -3012
rect 199 -3080 521 -3079
rect 199 -3400 200 -3080
rect 520 -3400 521 -3080
rect 199 -3401 521 -3400
rect -220 -3468 -124 -3452
rect 792 -3452 808 -3028
rect 872 -3452 888 -3028
rect 1804 -3028 1900 -3012
rect 1211 -3080 1533 -3079
rect 1211 -3400 1212 -3080
rect 1532 -3400 1533 -3080
rect 1211 -3401 1533 -3400
rect 792 -3468 888 -3452
rect 1804 -3452 1820 -3028
rect 1884 -3452 1900 -3028
rect 2816 -3028 2912 -3012
rect 2223 -3080 2545 -3079
rect 2223 -3400 2224 -3080
rect 2544 -3400 2545 -3080
rect 2223 -3401 2545 -3400
rect 1804 -3468 1900 -3452
rect 2816 -3452 2832 -3028
rect 2896 -3452 2912 -3028
rect 3828 -3028 3924 -3012
rect 3235 -3080 3557 -3079
rect 3235 -3400 3236 -3080
rect 3556 -3400 3557 -3080
rect 3235 -3401 3557 -3400
rect 2816 -3468 2912 -3452
rect 3828 -3452 3844 -3028
rect 3908 -3452 3924 -3028
rect 4840 -3028 4936 -3012
rect 4247 -3080 4569 -3079
rect 4247 -3400 4248 -3080
rect 4568 -3400 4569 -3080
rect 4247 -3401 4569 -3400
rect 3828 -3468 3924 -3452
rect 4840 -3452 4856 -3028
rect 4920 -3452 4936 -3028
rect 5852 -3028 5948 -3012
rect 5259 -3080 5581 -3079
rect 5259 -3400 5260 -3080
rect 5580 -3400 5581 -3080
rect 5259 -3401 5581 -3400
rect 4840 -3468 4936 -3452
rect 5852 -3452 5868 -3028
rect 5932 -3452 5948 -3028
rect 6864 -3028 6960 -3012
rect 6271 -3080 6593 -3079
rect 6271 -3400 6272 -3080
rect 6592 -3400 6593 -3080
rect 6271 -3401 6593 -3400
rect 5852 -3468 5948 -3452
rect 6864 -3452 6880 -3028
rect 6944 -3452 6960 -3028
rect 7876 -3028 7972 -3012
rect 7283 -3080 7605 -3079
rect 7283 -3400 7284 -3080
rect 7604 -3400 7605 -3080
rect 7283 -3401 7605 -3400
rect 6864 -3468 6960 -3452
rect 7876 -3452 7892 -3028
rect 7956 -3452 7972 -3028
rect 8888 -3028 8984 -3012
rect 8295 -3080 8617 -3079
rect 8295 -3400 8296 -3080
rect 8616 -3400 8617 -3080
rect 8295 -3401 8617 -3400
rect 7876 -3468 7972 -3452
rect 8888 -3452 8904 -3028
rect 8968 -3452 8984 -3028
rect 9900 -3028 9996 -3012
rect 9307 -3080 9629 -3079
rect 9307 -3400 9308 -3080
rect 9628 -3400 9629 -3080
rect 9307 -3401 9629 -3400
rect 8888 -3468 8984 -3452
rect 9900 -3452 9916 -3028
rect 9980 -3452 9996 -3028
rect 10912 -3028 11008 -3012
rect 10319 -3080 10641 -3079
rect 10319 -3400 10320 -3080
rect 10640 -3400 10641 -3080
rect 10319 -3401 10641 -3400
rect 9900 -3468 9996 -3452
rect 10912 -3452 10928 -3028
rect 10992 -3452 11008 -3028
rect 11924 -3028 12020 -3012
rect 11331 -3080 11653 -3079
rect 11331 -3400 11332 -3080
rect 11652 -3400 11653 -3080
rect 11331 -3401 11653 -3400
rect 10912 -3468 11008 -3452
rect 11924 -3452 11940 -3028
rect 12004 -3452 12020 -3028
rect 12936 -3028 13032 -3012
rect 12343 -3080 12665 -3079
rect 12343 -3400 12344 -3080
rect 12664 -3400 12665 -3080
rect 12343 -3401 12665 -3400
rect 11924 -3468 12020 -3452
rect 12936 -3452 12952 -3028
rect 13016 -3452 13032 -3028
rect 13948 -3028 14044 -3012
rect 13355 -3080 13677 -3079
rect 13355 -3400 13356 -3080
rect 13676 -3400 13677 -3080
rect 13355 -3401 13677 -3400
rect 12936 -3468 13032 -3452
rect 13948 -3452 13964 -3028
rect 14028 -3452 14044 -3028
rect 14960 -3028 15056 -3012
rect 14367 -3080 14689 -3079
rect 14367 -3400 14368 -3080
rect 14688 -3400 14689 -3080
rect 14367 -3401 14689 -3400
rect 13948 -3468 14044 -3452
rect 14960 -3452 14976 -3028
rect 15040 -3452 15056 -3028
rect 15972 -3028 16068 -3012
rect 15379 -3080 15701 -3079
rect 15379 -3400 15380 -3080
rect 15700 -3400 15701 -3080
rect 15379 -3401 15701 -3400
rect 14960 -3468 15056 -3452
rect 15972 -3452 15988 -3028
rect 16052 -3452 16068 -3028
rect 16984 -3028 17080 -3012
rect 16391 -3080 16713 -3079
rect 16391 -3400 16392 -3080
rect 16712 -3400 16713 -3080
rect 16391 -3401 16713 -3400
rect 15972 -3468 16068 -3452
rect 16984 -3452 17000 -3028
rect 17064 -3452 17080 -3028
rect 16984 -3468 17080 -3452
rect -16412 -3748 -16316 -3732
rect -17005 -3800 -16683 -3799
rect -17005 -4120 -17004 -3800
rect -16684 -4120 -16683 -3800
rect -17005 -4121 -16683 -4120
rect -16412 -4172 -16396 -3748
rect -16332 -4172 -16316 -3748
rect -15400 -3748 -15304 -3732
rect -15993 -3800 -15671 -3799
rect -15993 -4120 -15992 -3800
rect -15672 -4120 -15671 -3800
rect -15993 -4121 -15671 -4120
rect -16412 -4188 -16316 -4172
rect -15400 -4172 -15384 -3748
rect -15320 -4172 -15304 -3748
rect -14388 -3748 -14292 -3732
rect -14981 -3800 -14659 -3799
rect -14981 -4120 -14980 -3800
rect -14660 -4120 -14659 -3800
rect -14981 -4121 -14659 -4120
rect -15400 -4188 -15304 -4172
rect -14388 -4172 -14372 -3748
rect -14308 -4172 -14292 -3748
rect -13376 -3748 -13280 -3732
rect -13969 -3800 -13647 -3799
rect -13969 -4120 -13968 -3800
rect -13648 -4120 -13647 -3800
rect -13969 -4121 -13647 -4120
rect -14388 -4188 -14292 -4172
rect -13376 -4172 -13360 -3748
rect -13296 -4172 -13280 -3748
rect -12364 -3748 -12268 -3732
rect -12957 -3800 -12635 -3799
rect -12957 -4120 -12956 -3800
rect -12636 -4120 -12635 -3800
rect -12957 -4121 -12635 -4120
rect -13376 -4188 -13280 -4172
rect -12364 -4172 -12348 -3748
rect -12284 -4172 -12268 -3748
rect -11352 -3748 -11256 -3732
rect -11945 -3800 -11623 -3799
rect -11945 -4120 -11944 -3800
rect -11624 -4120 -11623 -3800
rect -11945 -4121 -11623 -4120
rect -12364 -4188 -12268 -4172
rect -11352 -4172 -11336 -3748
rect -11272 -4172 -11256 -3748
rect -10340 -3748 -10244 -3732
rect -10933 -3800 -10611 -3799
rect -10933 -4120 -10932 -3800
rect -10612 -4120 -10611 -3800
rect -10933 -4121 -10611 -4120
rect -11352 -4188 -11256 -4172
rect -10340 -4172 -10324 -3748
rect -10260 -4172 -10244 -3748
rect -9328 -3748 -9232 -3732
rect -9921 -3800 -9599 -3799
rect -9921 -4120 -9920 -3800
rect -9600 -4120 -9599 -3800
rect -9921 -4121 -9599 -4120
rect -10340 -4188 -10244 -4172
rect -9328 -4172 -9312 -3748
rect -9248 -4172 -9232 -3748
rect -8316 -3748 -8220 -3732
rect -8909 -3800 -8587 -3799
rect -8909 -4120 -8908 -3800
rect -8588 -4120 -8587 -3800
rect -8909 -4121 -8587 -4120
rect -9328 -4188 -9232 -4172
rect -8316 -4172 -8300 -3748
rect -8236 -4172 -8220 -3748
rect -7304 -3748 -7208 -3732
rect -7897 -3800 -7575 -3799
rect -7897 -4120 -7896 -3800
rect -7576 -4120 -7575 -3800
rect -7897 -4121 -7575 -4120
rect -8316 -4188 -8220 -4172
rect -7304 -4172 -7288 -3748
rect -7224 -4172 -7208 -3748
rect -6292 -3748 -6196 -3732
rect -6885 -3800 -6563 -3799
rect -6885 -4120 -6884 -3800
rect -6564 -4120 -6563 -3800
rect -6885 -4121 -6563 -4120
rect -7304 -4188 -7208 -4172
rect -6292 -4172 -6276 -3748
rect -6212 -4172 -6196 -3748
rect -5280 -3748 -5184 -3732
rect -5873 -3800 -5551 -3799
rect -5873 -4120 -5872 -3800
rect -5552 -4120 -5551 -3800
rect -5873 -4121 -5551 -4120
rect -6292 -4188 -6196 -4172
rect -5280 -4172 -5264 -3748
rect -5200 -4172 -5184 -3748
rect -4268 -3748 -4172 -3732
rect -4861 -3800 -4539 -3799
rect -4861 -4120 -4860 -3800
rect -4540 -4120 -4539 -3800
rect -4861 -4121 -4539 -4120
rect -5280 -4188 -5184 -4172
rect -4268 -4172 -4252 -3748
rect -4188 -4172 -4172 -3748
rect -3256 -3748 -3160 -3732
rect -3849 -3800 -3527 -3799
rect -3849 -4120 -3848 -3800
rect -3528 -4120 -3527 -3800
rect -3849 -4121 -3527 -4120
rect -4268 -4188 -4172 -4172
rect -3256 -4172 -3240 -3748
rect -3176 -4172 -3160 -3748
rect -2244 -3748 -2148 -3732
rect -2837 -3800 -2515 -3799
rect -2837 -4120 -2836 -3800
rect -2516 -4120 -2515 -3800
rect -2837 -4121 -2515 -4120
rect -3256 -4188 -3160 -4172
rect -2244 -4172 -2228 -3748
rect -2164 -4172 -2148 -3748
rect -1232 -3748 -1136 -3732
rect -1825 -3800 -1503 -3799
rect -1825 -4120 -1824 -3800
rect -1504 -4120 -1503 -3800
rect -1825 -4121 -1503 -4120
rect -2244 -4188 -2148 -4172
rect -1232 -4172 -1216 -3748
rect -1152 -4172 -1136 -3748
rect -220 -3748 -124 -3732
rect -813 -3800 -491 -3799
rect -813 -4120 -812 -3800
rect -492 -4120 -491 -3800
rect -813 -4121 -491 -4120
rect -1232 -4188 -1136 -4172
rect -220 -4172 -204 -3748
rect -140 -4172 -124 -3748
rect 792 -3748 888 -3732
rect 199 -3800 521 -3799
rect 199 -4120 200 -3800
rect 520 -4120 521 -3800
rect 199 -4121 521 -4120
rect -220 -4188 -124 -4172
rect 792 -4172 808 -3748
rect 872 -4172 888 -3748
rect 1804 -3748 1900 -3732
rect 1211 -3800 1533 -3799
rect 1211 -4120 1212 -3800
rect 1532 -4120 1533 -3800
rect 1211 -4121 1533 -4120
rect 792 -4188 888 -4172
rect 1804 -4172 1820 -3748
rect 1884 -4172 1900 -3748
rect 2816 -3748 2912 -3732
rect 2223 -3800 2545 -3799
rect 2223 -4120 2224 -3800
rect 2544 -4120 2545 -3800
rect 2223 -4121 2545 -4120
rect 1804 -4188 1900 -4172
rect 2816 -4172 2832 -3748
rect 2896 -4172 2912 -3748
rect 3828 -3748 3924 -3732
rect 3235 -3800 3557 -3799
rect 3235 -4120 3236 -3800
rect 3556 -4120 3557 -3800
rect 3235 -4121 3557 -4120
rect 2816 -4188 2912 -4172
rect 3828 -4172 3844 -3748
rect 3908 -4172 3924 -3748
rect 4840 -3748 4936 -3732
rect 4247 -3800 4569 -3799
rect 4247 -4120 4248 -3800
rect 4568 -4120 4569 -3800
rect 4247 -4121 4569 -4120
rect 3828 -4188 3924 -4172
rect 4840 -4172 4856 -3748
rect 4920 -4172 4936 -3748
rect 5852 -3748 5948 -3732
rect 5259 -3800 5581 -3799
rect 5259 -4120 5260 -3800
rect 5580 -4120 5581 -3800
rect 5259 -4121 5581 -4120
rect 4840 -4188 4936 -4172
rect 5852 -4172 5868 -3748
rect 5932 -4172 5948 -3748
rect 6864 -3748 6960 -3732
rect 6271 -3800 6593 -3799
rect 6271 -4120 6272 -3800
rect 6592 -4120 6593 -3800
rect 6271 -4121 6593 -4120
rect 5852 -4188 5948 -4172
rect 6864 -4172 6880 -3748
rect 6944 -4172 6960 -3748
rect 7876 -3748 7972 -3732
rect 7283 -3800 7605 -3799
rect 7283 -4120 7284 -3800
rect 7604 -4120 7605 -3800
rect 7283 -4121 7605 -4120
rect 6864 -4188 6960 -4172
rect 7876 -4172 7892 -3748
rect 7956 -4172 7972 -3748
rect 8888 -3748 8984 -3732
rect 8295 -3800 8617 -3799
rect 8295 -4120 8296 -3800
rect 8616 -4120 8617 -3800
rect 8295 -4121 8617 -4120
rect 7876 -4188 7972 -4172
rect 8888 -4172 8904 -3748
rect 8968 -4172 8984 -3748
rect 9900 -3748 9996 -3732
rect 9307 -3800 9629 -3799
rect 9307 -4120 9308 -3800
rect 9628 -4120 9629 -3800
rect 9307 -4121 9629 -4120
rect 8888 -4188 8984 -4172
rect 9900 -4172 9916 -3748
rect 9980 -4172 9996 -3748
rect 10912 -3748 11008 -3732
rect 10319 -3800 10641 -3799
rect 10319 -4120 10320 -3800
rect 10640 -4120 10641 -3800
rect 10319 -4121 10641 -4120
rect 9900 -4188 9996 -4172
rect 10912 -4172 10928 -3748
rect 10992 -4172 11008 -3748
rect 11924 -3748 12020 -3732
rect 11331 -3800 11653 -3799
rect 11331 -4120 11332 -3800
rect 11652 -4120 11653 -3800
rect 11331 -4121 11653 -4120
rect 10912 -4188 11008 -4172
rect 11924 -4172 11940 -3748
rect 12004 -4172 12020 -3748
rect 12936 -3748 13032 -3732
rect 12343 -3800 12665 -3799
rect 12343 -4120 12344 -3800
rect 12664 -4120 12665 -3800
rect 12343 -4121 12665 -4120
rect 11924 -4188 12020 -4172
rect 12936 -4172 12952 -3748
rect 13016 -4172 13032 -3748
rect 13948 -3748 14044 -3732
rect 13355 -3800 13677 -3799
rect 13355 -4120 13356 -3800
rect 13676 -4120 13677 -3800
rect 13355 -4121 13677 -4120
rect 12936 -4188 13032 -4172
rect 13948 -4172 13964 -3748
rect 14028 -4172 14044 -3748
rect 14960 -3748 15056 -3732
rect 14367 -3800 14689 -3799
rect 14367 -4120 14368 -3800
rect 14688 -4120 14689 -3800
rect 14367 -4121 14689 -4120
rect 13948 -4188 14044 -4172
rect 14960 -4172 14976 -3748
rect 15040 -4172 15056 -3748
rect 15972 -3748 16068 -3732
rect 15379 -3800 15701 -3799
rect 15379 -4120 15380 -3800
rect 15700 -4120 15701 -3800
rect 15379 -4121 15701 -4120
rect 14960 -4188 15056 -4172
rect 15972 -4172 15988 -3748
rect 16052 -4172 16068 -3748
rect 16984 -3748 17080 -3732
rect 16391 -3800 16713 -3799
rect 16391 -4120 16392 -3800
rect 16712 -4120 16713 -3800
rect 16391 -4121 16713 -4120
rect 15972 -4188 16068 -4172
rect 16984 -4172 17000 -3748
rect 17064 -4172 17080 -3748
rect 16984 -4188 17080 -4172
rect -16412 -4468 -16316 -4452
rect -17005 -4520 -16683 -4519
rect -17005 -4840 -17004 -4520
rect -16684 -4840 -16683 -4520
rect -17005 -4841 -16683 -4840
rect -16412 -4892 -16396 -4468
rect -16332 -4892 -16316 -4468
rect -15400 -4468 -15304 -4452
rect -15993 -4520 -15671 -4519
rect -15993 -4840 -15992 -4520
rect -15672 -4840 -15671 -4520
rect -15993 -4841 -15671 -4840
rect -16412 -4908 -16316 -4892
rect -15400 -4892 -15384 -4468
rect -15320 -4892 -15304 -4468
rect -14388 -4468 -14292 -4452
rect -14981 -4520 -14659 -4519
rect -14981 -4840 -14980 -4520
rect -14660 -4840 -14659 -4520
rect -14981 -4841 -14659 -4840
rect -15400 -4908 -15304 -4892
rect -14388 -4892 -14372 -4468
rect -14308 -4892 -14292 -4468
rect -13376 -4468 -13280 -4452
rect -13969 -4520 -13647 -4519
rect -13969 -4840 -13968 -4520
rect -13648 -4840 -13647 -4520
rect -13969 -4841 -13647 -4840
rect -14388 -4908 -14292 -4892
rect -13376 -4892 -13360 -4468
rect -13296 -4892 -13280 -4468
rect -12364 -4468 -12268 -4452
rect -12957 -4520 -12635 -4519
rect -12957 -4840 -12956 -4520
rect -12636 -4840 -12635 -4520
rect -12957 -4841 -12635 -4840
rect -13376 -4908 -13280 -4892
rect -12364 -4892 -12348 -4468
rect -12284 -4892 -12268 -4468
rect -11352 -4468 -11256 -4452
rect -11945 -4520 -11623 -4519
rect -11945 -4840 -11944 -4520
rect -11624 -4840 -11623 -4520
rect -11945 -4841 -11623 -4840
rect -12364 -4908 -12268 -4892
rect -11352 -4892 -11336 -4468
rect -11272 -4892 -11256 -4468
rect -10340 -4468 -10244 -4452
rect -10933 -4520 -10611 -4519
rect -10933 -4840 -10932 -4520
rect -10612 -4840 -10611 -4520
rect -10933 -4841 -10611 -4840
rect -11352 -4908 -11256 -4892
rect -10340 -4892 -10324 -4468
rect -10260 -4892 -10244 -4468
rect -9328 -4468 -9232 -4452
rect -9921 -4520 -9599 -4519
rect -9921 -4840 -9920 -4520
rect -9600 -4840 -9599 -4520
rect -9921 -4841 -9599 -4840
rect -10340 -4908 -10244 -4892
rect -9328 -4892 -9312 -4468
rect -9248 -4892 -9232 -4468
rect -8316 -4468 -8220 -4452
rect -8909 -4520 -8587 -4519
rect -8909 -4840 -8908 -4520
rect -8588 -4840 -8587 -4520
rect -8909 -4841 -8587 -4840
rect -9328 -4908 -9232 -4892
rect -8316 -4892 -8300 -4468
rect -8236 -4892 -8220 -4468
rect -7304 -4468 -7208 -4452
rect -7897 -4520 -7575 -4519
rect -7897 -4840 -7896 -4520
rect -7576 -4840 -7575 -4520
rect -7897 -4841 -7575 -4840
rect -8316 -4908 -8220 -4892
rect -7304 -4892 -7288 -4468
rect -7224 -4892 -7208 -4468
rect -6292 -4468 -6196 -4452
rect -6885 -4520 -6563 -4519
rect -6885 -4840 -6884 -4520
rect -6564 -4840 -6563 -4520
rect -6885 -4841 -6563 -4840
rect -7304 -4908 -7208 -4892
rect -6292 -4892 -6276 -4468
rect -6212 -4892 -6196 -4468
rect -5280 -4468 -5184 -4452
rect -5873 -4520 -5551 -4519
rect -5873 -4840 -5872 -4520
rect -5552 -4840 -5551 -4520
rect -5873 -4841 -5551 -4840
rect -6292 -4908 -6196 -4892
rect -5280 -4892 -5264 -4468
rect -5200 -4892 -5184 -4468
rect -4268 -4468 -4172 -4452
rect -4861 -4520 -4539 -4519
rect -4861 -4840 -4860 -4520
rect -4540 -4840 -4539 -4520
rect -4861 -4841 -4539 -4840
rect -5280 -4908 -5184 -4892
rect -4268 -4892 -4252 -4468
rect -4188 -4892 -4172 -4468
rect -3256 -4468 -3160 -4452
rect -3849 -4520 -3527 -4519
rect -3849 -4840 -3848 -4520
rect -3528 -4840 -3527 -4520
rect -3849 -4841 -3527 -4840
rect -4268 -4908 -4172 -4892
rect -3256 -4892 -3240 -4468
rect -3176 -4892 -3160 -4468
rect -2244 -4468 -2148 -4452
rect -2837 -4520 -2515 -4519
rect -2837 -4840 -2836 -4520
rect -2516 -4840 -2515 -4520
rect -2837 -4841 -2515 -4840
rect -3256 -4908 -3160 -4892
rect -2244 -4892 -2228 -4468
rect -2164 -4892 -2148 -4468
rect -1232 -4468 -1136 -4452
rect -1825 -4520 -1503 -4519
rect -1825 -4840 -1824 -4520
rect -1504 -4840 -1503 -4520
rect -1825 -4841 -1503 -4840
rect -2244 -4908 -2148 -4892
rect -1232 -4892 -1216 -4468
rect -1152 -4892 -1136 -4468
rect -220 -4468 -124 -4452
rect -813 -4520 -491 -4519
rect -813 -4840 -812 -4520
rect -492 -4840 -491 -4520
rect -813 -4841 -491 -4840
rect -1232 -4908 -1136 -4892
rect -220 -4892 -204 -4468
rect -140 -4892 -124 -4468
rect 792 -4468 888 -4452
rect 199 -4520 521 -4519
rect 199 -4840 200 -4520
rect 520 -4840 521 -4520
rect 199 -4841 521 -4840
rect -220 -4908 -124 -4892
rect 792 -4892 808 -4468
rect 872 -4892 888 -4468
rect 1804 -4468 1900 -4452
rect 1211 -4520 1533 -4519
rect 1211 -4840 1212 -4520
rect 1532 -4840 1533 -4520
rect 1211 -4841 1533 -4840
rect 792 -4908 888 -4892
rect 1804 -4892 1820 -4468
rect 1884 -4892 1900 -4468
rect 2816 -4468 2912 -4452
rect 2223 -4520 2545 -4519
rect 2223 -4840 2224 -4520
rect 2544 -4840 2545 -4520
rect 2223 -4841 2545 -4840
rect 1804 -4908 1900 -4892
rect 2816 -4892 2832 -4468
rect 2896 -4892 2912 -4468
rect 3828 -4468 3924 -4452
rect 3235 -4520 3557 -4519
rect 3235 -4840 3236 -4520
rect 3556 -4840 3557 -4520
rect 3235 -4841 3557 -4840
rect 2816 -4908 2912 -4892
rect 3828 -4892 3844 -4468
rect 3908 -4892 3924 -4468
rect 4840 -4468 4936 -4452
rect 4247 -4520 4569 -4519
rect 4247 -4840 4248 -4520
rect 4568 -4840 4569 -4520
rect 4247 -4841 4569 -4840
rect 3828 -4908 3924 -4892
rect 4840 -4892 4856 -4468
rect 4920 -4892 4936 -4468
rect 5852 -4468 5948 -4452
rect 5259 -4520 5581 -4519
rect 5259 -4840 5260 -4520
rect 5580 -4840 5581 -4520
rect 5259 -4841 5581 -4840
rect 4840 -4908 4936 -4892
rect 5852 -4892 5868 -4468
rect 5932 -4892 5948 -4468
rect 6864 -4468 6960 -4452
rect 6271 -4520 6593 -4519
rect 6271 -4840 6272 -4520
rect 6592 -4840 6593 -4520
rect 6271 -4841 6593 -4840
rect 5852 -4908 5948 -4892
rect 6864 -4892 6880 -4468
rect 6944 -4892 6960 -4468
rect 7876 -4468 7972 -4452
rect 7283 -4520 7605 -4519
rect 7283 -4840 7284 -4520
rect 7604 -4840 7605 -4520
rect 7283 -4841 7605 -4840
rect 6864 -4908 6960 -4892
rect 7876 -4892 7892 -4468
rect 7956 -4892 7972 -4468
rect 8888 -4468 8984 -4452
rect 8295 -4520 8617 -4519
rect 8295 -4840 8296 -4520
rect 8616 -4840 8617 -4520
rect 8295 -4841 8617 -4840
rect 7876 -4908 7972 -4892
rect 8888 -4892 8904 -4468
rect 8968 -4892 8984 -4468
rect 9900 -4468 9996 -4452
rect 9307 -4520 9629 -4519
rect 9307 -4840 9308 -4520
rect 9628 -4840 9629 -4520
rect 9307 -4841 9629 -4840
rect 8888 -4908 8984 -4892
rect 9900 -4892 9916 -4468
rect 9980 -4892 9996 -4468
rect 10912 -4468 11008 -4452
rect 10319 -4520 10641 -4519
rect 10319 -4840 10320 -4520
rect 10640 -4840 10641 -4520
rect 10319 -4841 10641 -4840
rect 9900 -4908 9996 -4892
rect 10912 -4892 10928 -4468
rect 10992 -4892 11008 -4468
rect 11924 -4468 12020 -4452
rect 11331 -4520 11653 -4519
rect 11331 -4840 11332 -4520
rect 11652 -4840 11653 -4520
rect 11331 -4841 11653 -4840
rect 10912 -4908 11008 -4892
rect 11924 -4892 11940 -4468
rect 12004 -4892 12020 -4468
rect 12936 -4468 13032 -4452
rect 12343 -4520 12665 -4519
rect 12343 -4840 12344 -4520
rect 12664 -4840 12665 -4520
rect 12343 -4841 12665 -4840
rect 11924 -4908 12020 -4892
rect 12936 -4892 12952 -4468
rect 13016 -4892 13032 -4468
rect 13948 -4468 14044 -4452
rect 13355 -4520 13677 -4519
rect 13355 -4840 13356 -4520
rect 13676 -4840 13677 -4520
rect 13355 -4841 13677 -4840
rect 12936 -4908 13032 -4892
rect 13948 -4892 13964 -4468
rect 14028 -4892 14044 -4468
rect 14960 -4468 15056 -4452
rect 14367 -4520 14689 -4519
rect 14367 -4840 14368 -4520
rect 14688 -4840 14689 -4520
rect 14367 -4841 14689 -4840
rect 13948 -4908 14044 -4892
rect 14960 -4892 14976 -4468
rect 15040 -4892 15056 -4468
rect 15972 -4468 16068 -4452
rect 15379 -4520 15701 -4519
rect 15379 -4840 15380 -4520
rect 15700 -4840 15701 -4520
rect 15379 -4841 15701 -4840
rect 14960 -4908 15056 -4892
rect 15972 -4892 15988 -4468
rect 16052 -4892 16068 -4468
rect 16984 -4468 17080 -4452
rect 16391 -4520 16713 -4519
rect 16391 -4840 16392 -4520
rect 16712 -4840 16713 -4520
rect 16391 -4841 16713 -4840
rect 15972 -4908 16068 -4892
rect 16984 -4892 17000 -4468
rect 17064 -4892 17080 -4468
rect 16984 -4908 17080 -4892
rect -16412 -5188 -16316 -5172
rect -17005 -5240 -16683 -5239
rect -17005 -5560 -17004 -5240
rect -16684 -5560 -16683 -5240
rect -17005 -5561 -16683 -5560
rect -16412 -5612 -16396 -5188
rect -16332 -5612 -16316 -5188
rect -15400 -5188 -15304 -5172
rect -15993 -5240 -15671 -5239
rect -15993 -5560 -15992 -5240
rect -15672 -5560 -15671 -5240
rect -15993 -5561 -15671 -5560
rect -16412 -5628 -16316 -5612
rect -15400 -5612 -15384 -5188
rect -15320 -5612 -15304 -5188
rect -14388 -5188 -14292 -5172
rect -14981 -5240 -14659 -5239
rect -14981 -5560 -14980 -5240
rect -14660 -5560 -14659 -5240
rect -14981 -5561 -14659 -5560
rect -15400 -5628 -15304 -5612
rect -14388 -5612 -14372 -5188
rect -14308 -5612 -14292 -5188
rect -13376 -5188 -13280 -5172
rect -13969 -5240 -13647 -5239
rect -13969 -5560 -13968 -5240
rect -13648 -5560 -13647 -5240
rect -13969 -5561 -13647 -5560
rect -14388 -5628 -14292 -5612
rect -13376 -5612 -13360 -5188
rect -13296 -5612 -13280 -5188
rect -12364 -5188 -12268 -5172
rect -12957 -5240 -12635 -5239
rect -12957 -5560 -12956 -5240
rect -12636 -5560 -12635 -5240
rect -12957 -5561 -12635 -5560
rect -13376 -5628 -13280 -5612
rect -12364 -5612 -12348 -5188
rect -12284 -5612 -12268 -5188
rect -11352 -5188 -11256 -5172
rect -11945 -5240 -11623 -5239
rect -11945 -5560 -11944 -5240
rect -11624 -5560 -11623 -5240
rect -11945 -5561 -11623 -5560
rect -12364 -5628 -12268 -5612
rect -11352 -5612 -11336 -5188
rect -11272 -5612 -11256 -5188
rect -10340 -5188 -10244 -5172
rect -10933 -5240 -10611 -5239
rect -10933 -5560 -10932 -5240
rect -10612 -5560 -10611 -5240
rect -10933 -5561 -10611 -5560
rect -11352 -5628 -11256 -5612
rect -10340 -5612 -10324 -5188
rect -10260 -5612 -10244 -5188
rect -9328 -5188 -9232 -5172
rect -9921 -5240 -9599 -5239
rect -9921 -5560 -9920 -5240
rect -9600 -5560 -9599 -5240
rect -9921 -5561 -9599 -5560
rect -10340 -5628 -10244 -5612
rect -9328 -5612 -9312 -5188
rect -9248 -5612 -9232 -5188
rect -8316 -5188 -8220 -5172
rect -8909 -5240 -8587 -5239
rect -8909 -5560 -8908 -5240
rect -8588 -5560 -8587 -5240
rect -8909 -5561 -8587 -5560
rect -9328 -5628 -9232 -5612
rect -8316 -5612 -8300 -5188
rect -8236 -5612 -8220 -5188
rect -7304 -5188 -7208 -5172
rect -7897 -5240 -7575 -5239
rect -7897 -5560 -7896 -5240
rect -7576 -5560 -7575 -5240
rect -7897 -5561 -7575 -5560
rect -8316 -5628 -8220 -5612
rect -7304 -5612 -7288 -5188
rect -7224 -5612 -7208 -5188
rect -6292 -5188 -6196 -5172
rect -6885 -5240 -6563 -5239
rect -6885 -5560 -6884 -5240
rect -6564 -5560 -6563 -5240
rect -6885 -5561 -6563 -5560
rect -7304 -5628 -7208 -5612
rect -6292 -5612 -6276 -5188
rect -6212 -5612 -6196 -5188
rect -5280 -5188 -5184 -5172
rect -5873 -5240 -5551 -5239
rect -5873 -5560 -5872 -5240
rect -5552 -5560 -5551 -5240
rect -5873 -5561 -5551 -5560
rect -6292 -5628 -6196 -5612
rect -5280 -5612 -5264 -5188
rect -5200 -5612 -5184 -5188
rect -4268 -5188 -4172 -5172
rect -4861 -5240 -4539 -5239
rect -4861 -5560 -4860 -5240
rect -4540 -5560 -4539 -5240
rect -4861 -5561 -4539 -5560
rect -5280 -5628 -5184 -5612
rect -4268 -5612 -4252 -5188
rect -4188 -5612 -4172 -5188
rect -3256 -5188 -3160 -5172
rect -3849 -5240 -3527 -5239
rect -3849 -5560 -3848 -5240
rect -3528 -5560 -3527 -5240
rect -3849 -5561 -3527 -5560
rect -4268 -5628 -4172 -5612
rect -3256 -5612 -3240 -5188
rect -3176 -5612 -3160 -5188
rect -2244 -5188 -2148 -5172
rect -2837 -5240 -2515 -5239
rect -2837 -5560 -2836 -5240
rect -2516 -5560 -2515 -5240
rect -2837 -5561 -2515 -5560
rect -3256 -5628 -3160 -5612
rect -2244 -5612 -2228 -5188
rect -2164 -5612 -2148 -5188
rect -1232 -5188 -1136 -5172
rect -1825 -5240 -1503 -5239
rect -1825 -5560 -1824 -5240
rect -1504 -5560 -1503 -5240
rect -1825 -5561 -1503 -5560
rect -2244 -5628 -2148 -5612
rect -1232 -5612 -1216 -5188
rect -1152 -5612 -1136 -5188
rect -220 -5188 -124 -5172
rect -813 -5240 -491 -5239
rect -813 -5560 -812 -5240
rect -492 -5560 -491 -5240
rect -813 -5561 -491 -5560
rect -1232 -5628 -1136 -5612
rect -220 -5612 -204 -5188
rect -140 -5612 -124 -5188
rect 792 -5188 888 -5172
rect 199 -5240 521 -5239
rect 199 -5560 200 -5240
rect 520 -5560 521 -5240
rect 199 -5561 521 -5560
rect -220 -5628 -124 -5612
rect 792 -5612 808 -5188
rect 872 -5612 888 -5188
rect 1804 -5188 1900 -5172
rect 1211 -5240 1533 -5239
rect 1211 -5560 1212 -5240
rect 1532 -5560 1533 -5240
rect 1211 -5561 1533 -5560
rect 792 -5628 888 -5612
rect 1804 -5612 1820 -5188
rect 1884 -5612 1900 -5188
rect 2816 -5188 2912 -5172
rect 2223 -5240 2545 -5239
rect 2223 -5560 2224 -5240
rect 2544 -5560 2545 -5240
rect 2223 -5561 2545 -5560
rect 1804 -5628 1900 -5612
rect 2816 -5612 2832 -5188
rect 2896 -5612 2912 -5188
rect 3828 -5188 3924 -5172
rect 3235 -5240 3557 -5239
rect 3235 -5560 3236 -5240
rect 3556 -5560 3557 -5240
rect 3235 -5561 3557 -5560
rect 2816 -5628 2912 -5612
rect 3828 -5612 3844 -5188
rect 3908 -5612 3924 -5188
rect 4840 -5188 4936 -5172
rect 4247 -5240 4569 -5239
rect 4247 -5560 4248 -5240
rect 4568 -5560 4569 -5240
rect 4247 -5561 4569 -5560
rect 3828 -5628 3924 -5612
rect 4840 -5612 4856 -5188
rect 4920 -5612 4936 -5188
rect 5852 -5188 5948 -5172
rect 5259 -5240 5581 -5239
rect 5259 -5560 5260 -5240
rect 5580 -5560 5581 -5240
rect 5259 -5561 5581 -5560
rect 4840 -5628 4936 -5612
rect 5852 -5612 5868 -5188
rect 5932 -5612 5948 -5188
rect 6864 -5188 6960 -5172
rect 6271 -5240 6593 -5239
rect 6271 -5560 6272 -5240
rect 6592 -5560 6593 -5240
rect 6271 -5561 6593 -5560
rect 5852 -5628 5948 -5612
rect 6864 -5612 6880 -5188
rect 6944 -5612 6960 -5188
rect 7876 -5188 7972 -5172
rect 7283 -5240 7605 -5239
rect 7283 -5560 7284 -5240
rect 7604 -5560 7605 -5240
rect 7283 -5561 7605 -5560
rect 6864 -5628 6960 -5612
rect 7876 -5612 7892 -5188
rect 7956 -5612 7972 -5188
rect 8888 -5188 8984 -5172
rect 8295 -5240 8617 -5239
rect 8295 -5560 8296 -5240
rect 8616 -5560 8617 -5240
rect 8295 -5561 8617 -5560
rect 7876 -5628 7972 -5612
rect 8888 -5612 8904 -5188
rect 8968 -5612 8984 -5188
rect 9900 -5188 9996 -5172
rect 9307 -5240 9629 -5239
rect 9307 -5560 9308 -5240
rect 9628 -5560 9629 -5240
rect 9307 -5561 9629 -5560
rect 8888 -5628 8984 -5612
rect 9900 -5612 9916 -5188
rect 9980 -5612 9996 -5188
rect 10912 -5188 11008 -5172
rect 10319 -5240 10641 -5239
rect 10319 -5560 10320 -5240
rect 10640 -5560 10641 -5240
rect 10319 -5561 10641 -5560
rect 9900 -5628 9996 -5612
rect 10912 -5612 10928 -5188
rect 10992 -5612 11008 -5188
rect 11924 -5188 12020 -5172
rect 11331 -5240 11653 -5239
rect 11331 -5560 11332 -5240
rect 11652 -5560 11653 -5240
rect 11331 -5561 11653 -5560
rect 10912 -5628 11008 -5612
rect 11924 -5612 11940 -5188
rect 12004 -5612 12020 -5188
rect 12936 -5188 13032 -5172
rect 12343 -5240 12665 -5239
rect 12343 -5560 12344 -5240
rect 12664 -5560 12665 -5240
rect 12343 -5561 12665 -5560
rect 11924 -5628 12020 -5612
rect 12936 -5612 12952 -5188
rect 13016 -5612 13032 -5188
rect 13948 -5188 14044 -5172
rect 13355 -5240 13677 -5239
rect 13355 -5560 13356 -5240
rect 13676 -5560 13677 -5240
rect 13355 -5561 13677 -5560
rect 12936 -5628 13032 -5612
rect 13948 -5612 13964 -5188
rect 14028 -5612 14044 -5188
rect 14960 -5188 15056 -5172
rect 14367 -5240 14689 -5239
rect 14367 -5560 14368 -5240
rect 14688 -5560 14689 -5240
rect 14367 -5561 14689 -5560
rect 13948 -5628 14044 -5612
rect 14960 -5612 14976 -5188
rect 15040 -5612 15056 -5188
rect 15972 -5188 16068 -5172
rect 15379 -5240 15701 -5239
rect 15379 -5560 15380 -5240
rect 15700 -5560 15701 -5240
rect 15379 -5561 15701 -5560
rect 14960 -5628 15056 -5612
rect 15972 -5612 15988 -5188
rect 16052 -5612 16068 -5188
rect 16984 -5188 17080 -5172
rect 16391 -5240 16713 -5239
rect 16391 -5560 16392 -5240
rect 16712 -5560 16713 -5240
rect 16391 -5561 16713 -5560
rect 15972 -5628 16068 -5612
rect 16984 -5612 17000 -5188
rect 17064 -5612 17080 -5188
rect 16984 -5628 17080 -5612
rect -16412 -5908 -16316 -5892
rect -17005 -5960 -16683 -5959
rect -17005 -6280 -17004 -5960
rect -16684 -6280 -16683 -5960
rect -17005 -6281 -16683 -6280
rect -16412 -6332 -16396 -5908
rect -16332 -6332 -16316 -5908
rect -15400 -5908 -15304 -5892
rect -15993 -5960 -15671 -5959
rect -15993 -6280 -15992 -5960
rect -15672 -6280 -15671 -5960
rect -15993 -6281 -15671 -6280
rect -16412 -6348 -16316 -6332
rect -15400 -6332 -15384 -5908
rect -15320 -6332 -15304 -5908
rect -14388 -5908 -14292 -5892
rect -14981 -5960 -14659 -5959
rect -14981 -6280 -14980 -5960
rect -14660 -6280 -14659 -5960
rect -14981 -6281 -14659 -6280
rect -15400 -6348 -15304 -6332
rect -14388 -6332 -14372 -5908
rect -14308 -6332 -14292 -5908
rect -13376 -5908 -13280 -5892
rect -13969 -5960 -13647 -5959
rect -13969 -6280 -13968 -5960
rect -13648 -6280 -13647 -5960
rect -13969 -6281 -13647 -6280
rect -14388 -6348 -14292 -6332
rect -13376 -6332 -13360 -5908
rect -13296 -6332 -13280 -5908
rect -12364 -5908 -12268 -5892
rect -12957 -5960 -12635 -5959
rect -12957 -6280 -12956 -5960
rect -12636 -6280 -12635 -5960
rect -12957 -6281 -12635 -6280
rect -13376 -6348 -13280 -6332
rect -12364 -6332 -12348 -5908
rect -12284 -6332 -12268 -5908
rect -11352 -5908 -11256 -5892
rect -11945 -5960 -11623 -5959
rect -11945 -6280 -11944 -5960
rect -11624 -6280 -11623 -5960
rect -11945 -6281 -11623 -6280
rect -12364 -6348 -12268 -6332
rect -11352 -6332 -11336 -5908
rect -11272 -6332 -11256 -5908
rect -10340 -5908 -10244 -5892
rect -10933 -5960 -10611 -5959
rect -10933 -6280 -10932 -5960
rect -10612 -6280 -10611 -5960
rect -10933 -6281 -10611 -6280
rect -11352 -6348 -11256 -6332
rect -10340 -6332 -10324 -5908
rect -10260 -6332 -10244 -5908
rect -9328 -5908 -9232 -5892
rect -9921 -5960 -9599 -5959
rect -9921 -6280 -9920 -5960
rect -9600 -6280 -9599 -5960
rect -9921 -6281 -9599 -6280
rect -10340 -6348 -10244 -6332
rect -9328 -6332 -9312 -5908
rect -9248 -6332 -9232 -5908
rect -8316 -5908 -8220 -5892
rect -8909 -5960 -8587 -5959
rect -8909 -6280 -8908 -5960
rect -8588 -6280 -8587 -5960
rect -8909 -6281 -8587 -6280
rect -9328 -6348 -9232 -6332
rect -8316 -6332 -8300 -5908
rect -8236 -6332 -8220 -5908
rect -7304 -5908 -7208 -5892
rect -7897 -5960 -7575 -5959
rect -7897 -6280 -7896 -5960
rect -7576 -6280 -7575 -5960
rect -7897 -6281 -7575 -6280
rect -8316 -6348 -8220 -6332
rect -7304 -6332 -7288 -5908
rect -7224 -6332 -7208 -5908
rect -6292 -5908 -6196 -5892
rect -6885 -5960 -6563 -5959
rect -6885 -6280 -6884 -5960
rect -6564 -6280 -6563 -5960
rect -6885 -6281 -6563 -6280
rect -7304 -6348 -7208 -6332
rect -6292 -6332 -6276 -5908
rect -6212 -6332 -6196 -5908
rect -5280 -5908 -5184 -5892
rect -5873 -5960 -5551 -5959
rect -5873 -6280 -5872 -5960
rect -5552 -6280 -5551 -5960
rect -5873 -6281 -5551 -6280
rect -6292 -6348 -6196 -6332
rect -5280 -6332 -5264 -5908
rect -5200 -6332 -5184 -5908
rect -4268 -5908 -4172 -5892
rect -4861 -5960 -4539 -5959
rect -4861 -6280 -4860 -5960
rect -4540 -6280 -4539 -5960
rect -4861 -6281 -4539 -6280
rect -5280 -6348 -5184 -6332
rect -4268 -6332 -4252 -5908
rect -4188 -6332 -4172 -5908
rect -3256 -5908 -3160 -5892
rect -3849 -5960 -3527 -5959
rect -3849 -6280 -3848 -5960
rect -3528 -6280 -3527 -5960
rect -3849 -6281 -3527 -6280
rect -4268 -6348 -4172 -6332
rect -3256 -6332 -3240 -5908
rect -3176 -6332 -3160 -5908
rect -2244 -5908 -2148 -5892
rect -2837 -5960 -2515 -5959
rect -2837 -6280 -2836 -5960
rect -2516 -6280 -2515 -5960
rect -2837 -6281 -2515 -6280
rect -3256 -6348 -3160 -6332
rect -2244 -6332 -2228 -5908
rect -2164 -6332 -2148 -5908
rect -1232 -5908 -1136 -5892
rect -1825 -5960 -1503 -5959
rect -1825 -6280 -1824 -5960
rect -1504 -6280 -1503 -5960
rect -1825 -6281 -1503 -6280
rect -2244 -6348 -2148 -6332
rect -1232 -6332 -1216 -5908
rect -1152 -6332 -1136 -5908
rect -220 -5908 -124 -5892
rect -813 -5960 -491 -5959
rect -813 -6280 -812 -5960
rect -492 -6280 -491 -5960
rect -813 -6281 -491 -6280
rect -1232 -6348 -1136 -6332
rect -220 -6332 -204 -5908
rect -140 -6332 -124 -5908
rect 792 -5908 888 -5892
rect 199 -5960 521 -5959
rect 199 -6280 200 -5960
rect 520 -6280 521 -5960
rect 199 -6281 521 -6280
rect -220 -6348 -124 -6332
rect 792 -6332 808 -5908
rect 872 -6332 888 -5908
rect 1804 -5908 1900 -5892
rect 1211 -5960 1533 -5959
rect 1211 -6280 1212 -5960
rect 1532 -6280 1533 -5960
rect 1211 -6281 1533 -6280
rect 792 -6348 888 -6332
rect 1804 -6332 1820 -5908
rect 1884 -6332 1900 -5908
rect 2816 -5908 2912 -5892
rect 2223 -5960 2545 -5959
rect 2223 -6280 2224 -5960
rect 2544 -6280 2545 -5960
rect 2223 -6281 2545 -6280
rect 1804 -6348 1900 -6332
rect 2816 -6332 2832 -5908
rect 2896 -6332 2912 -5908
rect 3828 -5908 3924 -5892
rect 3235 -5960 3557 -5959
rect 3235 -6280 3236 -5960
rect 3556 -6280 3557 -5960
rect 3235 -6281 3557 -6280
rect 2816 -6348 2912 -6332
rect 3828 -6332 3844 -5908
rect 3908 -6332 3924 -5908
rect 4840 -5908 4936 -5892
rect 4247 -5960 4569 -5959
rect 4247 -6280 4248 -5960
rect 4568 -6280 4569 -5960
rect 4247 -6281 4569 -6280
rect 3828 -6348 3924 -6332
rect 4840 -6332 4856 -5908
rect 4920 -6332 4936 -5908
rect 5852 -5908 5948 -5892
rect 5259 -5960 5581 -5959
rect 5259 -6280 5260 -5960
rect 5580 -6280 5581 -5960
rect 5259 -6281 5581 -6280
rect 4840 -6348 4936 -6332
rect 5852 -6332 5868 -5908
rect 5932 -6332 5948 -5908
rect 6864 -5908 6960 -5892
rect 6271 -5960 6593 -5959
rect 6271 -6280 6272 -5960
rect 6592 -6280 6593 -5960
rect 6271 -6281 6593 -6280
rect 5852 -6348 5948 -6332
rect 6864 -6332 6880 -5908
rect 6944 -6332 6960 -5908
rect 7876 -5908 7972 -5892
rect 7283 -5960 7605 -5959
rect 7283 -6280 7284 -5960
rect 7604 -6280 7605 -5960
rect 7283 -6281 7605 -6280
rect 6864 -6348 6960 -6332
rect 7876 -6332 7892 -5908
rect 7956 -6332 7972 -5908
rect 8888 -5908 8984 -5892
rect 8295 -5960 8617 -5959
rect 8295 -6280 8296 -5960
rect 8616 -6280 8617 -5960
rect 8295 -6281 8617 -6280
rect 7876 -6348 7972 -6332
rect 8888 -6332 8904 -5908
rect 8968 -6332 8984 -5908
rect 9900 -5908 9996 -5892
rect 9307 -5960 9629 -5959
rect 9307 -6280 9308 -5960
rect 9628 -6280 9629 -5960
rect 9307 -6281 9629 -6280
rect 8888 -6348 8984 -6332
rect 9900 -6332 9916 -5908
rect 9980 -6332 9996 -5908
rect 10912 -5908 11008 -5892
rect 10319 -5960 10641 -5959
rect 10319 -6280 10320 -5960
rect 10640 -6280 10641 -5960
rect 10319 -6281 10641 -6280
rect 9900 -6348 9996 -6332
rect 10912 -6332 10928 -5908
rect 10992 -6332 11008 -5908
rect 11924 -5908 12020 -5892
rect 11331 -5960 11653 -5959
rect 11331 -6280 11332 -5960
rect 11652 -6280 11653 -5960
rect 11331 -6281 11653 -6280
rect 10912 -6348 11008 -6332
rect 11924 -6332 11940 -5908
rect 12004 -6332 12020 -5908
rect 12936 -5908 13032 -5892
rect 12343 -5960 12665 -5959
rect 12343 -6280 12344 -5960
rect 12664 -6280 12665 -5960
rect 12343 -6281 12665 -6280
rect 11924 -6348 12020 -6332
rect 12936 -6332 12952 -5908
rect 13016 -6332 13032 -5908
rect 13948 -5908 14044 -5892
rect 13355 -5960 13677 -5959
rect 13355 -6280 13356 -5960
rect 13676 -6280 13677 -5960
rect 13355 -6281 13677 -6280
rect 12936 -6348 13032 -6332
rect 13948 -6332 13964 -5908
rect 14028 -6332 14044 -5908
rect 14960 -5908 15056 -5892
rect 14367 -5960 14689 -5959
rect 14367 -6280 14368 -5960
rect 14688 -6280 14689 -5960
rect 14367 -6281 14689 -6280
rect 13948 -6348 14044 -6332
rect 14960 -6332 14976 -5908
rect 15040 -6332 15056 -5908
rect 15972 -5908 16068 -5892
rect 15379 -5960 15701 -5959
rect 15379 -6280 15380 -5960
rect 15700 -6280 15701 -5960
rect 15379 -6281 15701 -6280
rect 14960 -6348 15056 -6332
rect 15972 -6332 15988 -5908
rect 16052 -6332 16068 -5908
rect 16984 -5908 17080 -5892
rect 16391 -5960 16713 -5959
rect 16391 -6280 16392 -5960
rect 16712 -6280 16713 -5960
rect 16391 -6281 16713 -6280
rect 15972 -6348 16068 -6332
rect 16984 -6332 17000 -5908
rect 17064 -6332 17080 -5908
rect 16984 -6348 17080 -6332
rect -16412 -6628 -16316 -6612
rect -17005 -6680 -16683 -6679
rect -17005 -7000 -17004 -6680
rect -16684 -7000 -16683 -6680
rect -17005 -7001 -16683 -7000
rect -16412 -7052 -16396 -6628
rect -16332 -7052 -16316 -6628
rect -15400 -6628 -15304 -6612
rect -15993 -6680 -15671 -6679
rect -15993 -7000 -15992 -6680
rect -15672 -7000 -15671 -6680
rect -15993 -7001 -15671 -7000
rect -16412 -7068 -16316 -7052
rect -15400 -7052 -15384 -6628
rect -15320 -7052 -15304 -6628
rect -14388 -6628 -14292 -6612
rect -14981 -6680 -14659 -6679
rect -14981 -7000 -14980 -6680
rect -14660 -7000 -14659 -6680
rect -14981 -7001 -14659 -7000
rect -15400 -7068 -15304 -7052
rect -14388 -7052 -14372 -6628
rect -14308 -7052 -14292 -6628
rect -13376 -6628 -13280 -6612
rect -13969 -6680 -13647 -6679
rect -13969 -7000 -13968 -6680
rect -13648 -7000 -13647 -6680
rect -13969 -7001 -13647 -7000
rect -14388 -7068 -14292 -7052
rect -13376 -7052 -13360 -6628
rect -13296 -7052 -13280 -6628
rect -12364 -6628 -12268 -6612
rect -12957 -6680 -12635 -6679
rect -12957 -7000 -12956 -6680
rect -12636 -7000 -12635 -6680
rect -12957 -7001 -12635 -7000
rect -13376 -7068 -13280 -7052
rect -12364 -7052 -12348 -6628
rect -12284 -7052 -12268 -6628
rect -11352 -6628 -11256 -6612
rect -11945 -6680 -11623 -6679
rect -11945 -7000 -11944 -6680
rect -11624 -7000 -11623 -6680
rect -11945 -7001 -11623 -7000
rect -12364 -7068 -12268 -7052
rect -11352 -7052 -11336 -6628
rect -11272 -7052 -11256 -6628
rect -10340 -6628 -10244 -6612
rect -10933 -6680 -10611 -6679
rect -10933 -7000 -10932 -6680
rect -10612 -7000 -10611 -6680
rect -10933 -7001 -10611 -7000
rect -11352 -7068 -11256 -7052
rect -10340 -7052 -10324 -6628
rect -10260 -7052 -10244 -6628
rect -9328 -6628 -9232 -6612
rect -9921 -6680 -9599 -6679
rect -9921 -7000 -9920 -6680
rect -9600 -7000 -9599 -6680
rect -9921 -7001 -9599 -7000
rect -10340 -7068 -10244 -7052
rect -9328 -7052 -9312 -6628
rect -9248 -7052 -9232 -6628
rect -8316 -6628 -8220 -6612
rect -8909 -6680 -8587 -6679
rect -8909 -7000 -8908 -6680
rect -8588 -7000 -8587 -6680
rect -8909 -7001 -8587 -7000
rect -9328 -7068 -9232 -7052
rect -8316 -7052 -8300 -6628
rect -8236 -7052 -8220 -6628
rect -7304 -6628 -7208 -6612
rect -7897 -6680 -7575 -6679
rect -7897 -7000 -7896 -6680
rect -7576 -7000 -7575 -6680
rect -7897 -7001 -7575 -7000
rect -8316 -7068 -8220 -7052
rect -7304 -7052 -7288 -6628
rect -7224 -7052 -7208 -6628
rect -6292 -6628 -6196 -6612
rect -6885 -6680 -6563 -6679
rect -6885 -7000 -6884 -6680
rect -6564 -7000 -6563 -6680
rect -6885 -7001 -6563 -7000
rect -7304 -7068 -7208 -7052
rect -6292 -7052 -6276 -6628
rect -6212 -7052 -6196 -6628
rect -5280 -6628 -5184 -6612
rect -5873 -6680 -5551 -6679
rect -5873 -7000 -5872 -6680
rect -5552 -7000 -5551 -6680
rect -5873 -7001 -5551 -7000
rect -6292 -7068 -6196 -7052
rect -5280 -7052 -5264 -6628
rect -5200 -7052 -5184 -6628
rect -4268 -6628 -4172 -6612
rect -4861 -6680 -4539 -6679
rect -4861 -7000 -4860 -6680
rect -4540 -7000 -4539 -6680
rect -4861 -7001 -4539 -7000
rect -5280 -7068 -5184 -7052
rect -4268 -7052 -4252 -6628
rect -4188 -7052 -4172 -6628
rect -3256 -6628 -3160 -6612
rect -3849 -6680 -3527 -6679
rect -3849 -7000 -3848 -6680
rect -3528 -7000 -3527 -6680
rect -3849 -7001 -3527 -7000
rect -4268 -7068 -4172 -7052
rect -3256 -7052 -3240 -6628
rect -3176 -7052 -3160 -6628
rect -2244 -6628 -2148 -6612
rect -2837 -6680 -2515 -6679
rect -2837 -7000 -2836 -6680
rect -2516 -7000 -2515 -6680
rect -2837 -7001 -2515 -7000
rect -3256 -7068 -3160 -7052
rect -2244 -7052 -2228 -6628
rect -2164 -7052 -2148 -6628
rect -1232 -6628 -1136 -6612
rect -1825 -6680 -1503 -6679
rect -1825 -7000 -1824 -6680
rect -1504 -7000 -1503 -6680
rect -1825 -7001 -1503 -7000
rect -2244 -7068 -2148 -7052
rect -1232 -7052 -1216 -6628
rect -1152 -7052 -1136 -6628
rect -220 -6628 -124 -6612
rect -813 -6680 -491 -6679
rect -813 -7000 -812 -6680
rect -492 -7000 -491 -6680
rect -813 -7001 -491 -7000
rect -1232 -7068 -1136 -7052
rect -220 -7052 -204 -6628
rect -140 -7052 -124 -6628
rect 792 -6628 888 -6612
rect 199 -6680 521 -6679
rect 199 -7000 200 -6680
rect 520 -7000 521 -6680
rect 199 -7001 521 -7000
rect -220 -7068 -124 -7052
rect 792 -7052 808 -6628
rect 872 -7052 888 -6628
rect 1804 -6628 1900 -6612
rect 1211 -6680 1533 -6679
rect 1211 -7000 1212 -6680
rect 1532 -7000 1533 -6680
rect 1211 -7001 1533 -7000
rect 792 -7068 888 -7052
rect 1804 -7052 1820 -6628
rect 1884 -7052 1900 -6628
rect 2816 -6628 2912 -6612
rect 2223 -6680 2545 -6679
rect 2223 -7000 2224 -6680
rect 2544 -7000 2545 -6680
rect 2223 -7001 2545 -7000
rect 1804 -7068 1900 -7052
rect 2816 -7052 2832 -6628
rect 2896 -7052 2912 -6628
rect 3828 -6628 3924 -6612
rect 3235 -6680 3557 -6679
rect 3235 -7000 3236 -6680
rect 3556 -7000 3557 -6680
rect 3235 -7001 3557 -7000
rect 2816 -7068 2912 -7052
rect 3828 -7052 3844 -6628
rect 3908 -7052 3924 -6628
rect 4840 -6628 4936 -6612
rect 4247 -6680 4569 -6679
rect 4247 -7000 4248 -6680
rect 4568 -7000 4569 -6680
rect 4247 -7001 4569 -7000
rect 3828 -7068 3924 -7052
rect 4840 -7052 4856 -6628
rect 4920 -7052 4936 -6628
rect 5852 -6628 5948 -6612
rect 5259 -6680 5581 -6679
rect 5259 -7000 5260 -6680
rect 5580 -7000 5581 -6680
rect 5259 -7001 5581 -7000
rect 4840 -7068 4936 -7052
rect 5852 -7052 5868 -6628
rect 5932 -7052 5948 -6628
rect 6864 -6628 6960 -6612
rect 6271 -6680 6593 -6679
rect 6271 -7000 6272 -6680
rect 6592 -7000 6593 -6680
rect 6271 -7001 6593 -7000
rect 5852 -7068 5948 -7052
rect 6864 -7052 6880 -6628
rect 6944 -7052 6960 -6628
rect 7876 -6628 7972 -6612
rect 7283 -6680 7605 -6679
rect 7283 -7000 7284 -6680
rect 7604 -7000 7605 -6680
rect 7283 -7001 7605 -7000
rect 6864 -7068 6960 -7052
rect 7876 -7052 7892 -6628
rect 7956 -7052 7972 -6628
rect 8888 -6628 8984 -6612
rect 8295 -6680 8617 -6679
rect 8295 -7000 8296 -6680
rect 8616 -7000 8617 -6680
rect 8295 -7001 8617 -7000
rect 7876 -7068 7972 -7052
rect 8888 -7052 8904 -6628
rect 8968 -7052 8984 -6628
rect 9900 -6628 9996 -6612
rect 9307 -6680 9629 -6679
rect 9307 -7000 9308 -6680
rect 9628 -7000 9629 -6680
rect 9307 -7001 9629 -7000
rect 8888 -7068 8984 -7052
rect 9900 -7052 9916 -6628
rect 9980 -7052 9996 -6628
rect 10912 -6628 11008 -6612
rect 10319 -6680 10641 -6679
rect 10319 -7000 10320 -6680
rect 10640 -7000 10641 -6680
rect 10319 -7001 10641 -7000
rect 9900 -7068 9996 -7052
rect 10912 -7052 10928 -6628
rect 10992 -7052 11008 -6628
rect 11924 -6628 12020 -6612
rect 11331 -6680 11653 -6679
rect 11331 -7000 11332 -6680
rect 11652 -7000 11653 -6680
rect 11331 -7001 11653 -7000
rect 10912 -7068 11008 -7052
rect 11924 -7052 11940 -6628
rect 12004 -7052 12020 -6628
rect 12936 -6628 13032 -6612
rect 12343 -6680 12665 -6679
rect 12343 -7000 12344 -6680
rect 12664 -7000 12665 -6680
rect 12343 -7001 12665 -7000
rect 11924 -7068 12020 -7052
rect 12936 -7052 12952 -6628
rect 13016 -7052 13032 -6628
rect 13948 -6628 14044 -6612
rect 13355 -6680 13677 -6679
rect 13355 -7000 13356 -6680
rect 13676 -7000 13677 -6680
rect 13355 -7001 13677 -7000
rect 12936 -7068 13032 -7052
rect 13948 -7052 13964 -6628
rect 14028 -7052 14044 -6628
rect 14960 -6628 15056 -6612
rect 14367 -6680 14689 -6679
rect 14367 -7000 14368 -6680
rect 14688 -7000 14689 -6680
rect 14367 -7001 14689 -7000
rect 13948 -7068 14044 -7052
rect 14960 -7052 14976 -6628
rect 15040 -7052 15056 -6628
rect 15972 -6628 16068 -6612
rect 15379 -6680 15701 -6679
rect 15379 -7000 15380 -6680
rect 15700 -7000 15701 -6680
rect 15379 -7001 15701 -7000
rect 14960 -7068 15056 -7052
rect 15972 -7052 15988 -6628
rect 16052 -7052 16068 -6628
rect 16984 -6628 17080 -6612
rect 16391 -6680 16713 -6679
rect 16391 -7000 16392 -6680
rect 16712 -7000 16713 -6680
rect 16391 -7001 16713 -7000
rect 15972 -7068 16068 -7052
rect 16984 -7052 17000 -6628
rect 17064 -7052 17080 -6628
rect 16984 -7068 17080 -7052
rect -16412 -7348 -16316 -7332
rect -17005 -7400 -16683 -7399
rect -17005 -7720 -17004 -7400
rect -16684 -7720 -16683 -7400
rect -17005 -7721 -16683 -7720
rect -16412 -7772 -16396 -7348
rect -16332 -7772 -16316 -7348
rect -15400 -7348 -15304 -7332
rect -15993 -7400 -15671 -7399
rect -15993 -7720 -15992 -7400
rect -15672 -7720 -15671 -7400
rect -15993 -7721 -15671 -7720
rect -16412 -7788 -16316 -7772
rect -15400 -7772 -15384 -7348
rect -15320 -7772 -15304 -7348
rect -14388 -7348 -14292 -7332
rect -14981 -7400 -14659 -7399
rect -14981 -7720 -14980 -7400
rect -14660 -7720 -14659 -7400
rect -14981 -7721 -14659 -7720
rect -15400 -7788 -15304 -7772
rect -14388 -7772 -14372 -7348
rect -14308 -7772 -14292 -7348
rect -13376 -7348 -13280 -7332
rect -13969 -7400 -13647 -7399
rect -13969 -7720 -13968 -7400
rect -13648 -7720 -13647 -7400
rect -13969 -7721 -13647 -7720
rect -14388 -7788 -14292 -7772
rect -13376 -7772 -13360 -7348
rect -13296 -7772 -13280 -7348
rect -12364 -7348 -12268 -7332
rect -12957 -7400 -12635 -7399
rect -12957 -7720 -12956 -7400
rect -12636 -7720 -12635 -7400
rect -12957 -7721 -12635 -7720
rect -13376 -7788 -13280 -7772
rect -12364 -7772 -12348 -7348
rect -12284 -7772 -12268 -7348
rect -11352 -7348 -11256 -7332
rect -11945 -7400 -11623 -7399
rect -11945 -7720 -11944 -7400
rect -11624 -7720 -11623 -7400
rect -11945 -7721 -11623 -7720
rect -12364 -7788 -12268 -7772
rect -11352 -7772 -11336 -7348
rect -11272 -7772 -11256 -7348
rect -10340 -7348 -10244 -7332
rect -10933 -7400 -10611 -7399
rect -10933 -7720 -10932 -7400
rect -10612 -7720 -10611 -7400
rect -10933 -7721 -10611 -7720
rect -11352 -7788 -11256 -7772
rect -10340 -7772 -10324 -7348
rect -10260 -7772 -10244 -7348
rect -9328 -7348 -9232 -7332
rect -9921 -7400 -9599 -7399
rect -9921 -7720 -9920 -7400
rect -9600 -7720 -9599 -7400
rect -9921 -7721 -9599 -7720
rect -10340 -7788 -10244 -7772
rect -9328 -7772 -9312 -7348
rect -9248 -7772 -9232 -7348
rect -8316 -7348 -8220 -7332
rect -8909 -7400 -8587 -7399
rect -8909 -7720 -8908 -7400
rect -8588 -7720 -8587 -7400
rect -8909 -7721 -8587 -7720
rect -9328 -7788 -9232 -7772
rect -8316 -7772 -8300 -7348
rect -8236 -7772 -8220 -7348
rect -7304 -7348 -7208 -7332
rect -7897 -7400 -7575 -7399
rect -7897 -7720 -7896 -7400
rect -7576 -7720 -7575 -7400
rect -7897 -7721 -7575 -7720
rect -8316 -7788 -8220 -7772
rect -7304 -7772 -7288 -7348
rect -7224 -7772 -7208 -7348
rect -6292 -7348 -6196 -7332
rect -6885 -7400 -6563 -7399
rect -6885 -7720 -6884 -7400
rect -6564 -7720 -6563 -7400
rect -6885 -7721 -6563 -7720
rect -7304 -7788 -7208 -7772
rect -6292 -7772 -6276 -7348
rect -6212 -7772 -6196 -7348
rect -5280 -7348 -5184 -7332
rect -5873 -7400 -5551 -7399
rect -5873 -7720 -5872 -7400
rect -5552 -7720 -5551 -7400
rect -5873 -7721 -5551 -7720
rect -6292 -7788 -6196 -7772
rect -5280 -7772 -5264 -7348
rect -5200 -7772 -5184 -7348
rect -4268 -7348 -4172 -7332
rect -4861 -7400 -4539 -7399
rect -4861 -7720 -4860 -7400
rect -4540 -7720 -4539 -7400
rect -4861 -7721 -4539 -7720
rect -5280 -7788 -5184 -7772
rect -4268 -7772 -4252 -7348
rect -4188 -7772 -4172 -7348
rect -3256 -7348 -3160 -7332
rect -3849 -7400 -3527 -7399
rect -3849 -7720 -3848 -7400
rect -3528 -7720 -3527 -7400
rect -3849 -7721 -3527 -7720
rect -4268 -7788 -4172 -7772
rect -3256 -7772 -3240 -7348
rect -3176 -7772 -3160 -7348
rect -2244 -7348 -2148 -7332
rect -2837 -7400 -2515 -7399
rect -2837 -7720 -2836 -7400
rect -2516 -7720 -2515 -7400
rect -2837 -7721 -2515 -7720
rect -3256 -7788 -3160 -7772
rect -2244 -7772 -2228 -7348
rect -2164 -7772 -2148 -7348
rect -1232 -7348 -1136 -7332
rect -1825 -7400 -1503 -7399
rect -1825 -7720 -1824 -7400
rect -1504 -7720 -1503 -7400
rect -1825 -7721 -1503 -7720
rect -2244 -7788 -2148 -7772
rect -1232 -7772 -1216 -7348
rect -1152 -7772 -1136 -7348
rect -220 -7348 -124 -7332
rect -813 -7400 -491 -7399
rect -813 -7720 -812 -7400
rect -492 -7720 -491 -7400
rect -813 -7721 -491 -7720
rect -1232 -7788 -1136 -7772
rect -220 -7772 -204 -7348
rect -140 -7772 -124 -7348
rect 792 -7348 888 -7332
rect 199 -7400 521 -7399
rect 199 -7720 200 -7400
rect 520 -7720 521 -7400
rect 199 -7721 521 -7720
rect -220 -7788 -124 -7772
rect 792 -7772 808 -7348
rect 872 -7772 888 -7348
rect 1804 -7348 1900 -7332
rect 1211 -7400 1533 -7399
rect 1211 -7720 1212 -7400
rect 1532 -7720 1533 -7400
rect 1211 -7721 1533 -7720
rect 792 -7788 888 -7772
rect 1804 -7772 1820 -7348
rect 1884 -7772 1900 -7348
rect 2816 -7348 2912 -7332
rect 2223 -7400 2545 -7399
rect 2223 -7720 2224 -7400
rect 2544 -7720 2545 -7400
rect 2223 -7721 2545 -7720
rect 1804 -7788 1900 -7772
rect 2816 -7772 2832 -7348
rect 2896 -7772 2912 -7348
rect 3828 -7348 3924 -7332
rect 3235 -7400 3557 -7399
rect 3235 -7720 3236 -7400
rect 3556 -7720 3557 -7400
rect 3235 -7721 3557 -7720
rect 2816 -7788 2912 -7772
rect 3828 -7772 3844 -7348
rect 3908 -7772 3924 -7348
rect 4840 -7348 4936 -7332
rect 4247 -7400 4569 -7399
rect 4247 -7720 4248 -7400
rect 4568 -7720 4569 -7400
rect 4247 -7721 4569 -7720
rect 3828 -7788 3924 -7772
rect 4840 -7772 4856 -7348
rect 4920 -7772 4936 -7348
rect 5852 -7348 5948 -7332
rect 5259 -7400 5581 -7399
rect 5259 -7720 5260 -7400
rect 5580 -7720 5581 -7400
rect 5259 -7721 5581 -7720
rect 4840 -7788 4936 -7772
rect 5852 -7772 5868 -7348
rect 5932 -7772 5948 -7348
rect 6864 -7348 6960 -7332
rect 6271 -7400 6593 -7399
rect 6271 -7720 6272 -7400
rect 6592 -7720 6593 -7400
rect 6271 -7721 6593 -7720
rect 5852 -7788 5948 -7772
rect 6864 -7772 6880 -7348
rect 6944 -7772 6960 -7348
rect 7876 -7348 7972 -7332
rect 7283 -7400 7605 -7399
rect 7283 -7720 7284 -7400
rect 7604 -7720 7605 -7400
rect 7283 -7721 7605 -7720
rect 6864 -7788 6960 -7772
rect 7876 -7772 7892 -7348
rect 7956 -7772 7972 -7348
rect 8888 -7348 8984 -7332
rect 8295 -7400 8617 -7399
rect 8295 -7720 8296 -7400
rect 8616 -7720 8617 -7400
rect 8295 -7721 8617 -7720
rect 7876 -7788 7972 -7772
rect 8888 -7772 8904 -7348
rect 8968 -7772 8984 -7348
rect 9900 -7348 9996 -7332
rect 9307 -7400 9629 -7399
rect 9307 -7720 9308 -7400
rect 9628 -7720 9629 -7400
rect 9307 -7721 9629 -7720
rect 8888 -7788 8984 -7772
rect 9900 -7772 9916 -7348
rect 9980 -7772 9996 -7348
rect 10912 -7348 11008 -7332
rect 10319 -7400 10641 -7399
rect 10319 -7720 10320 -7400
rect 10640 -7720 10641 -7400
rect 10319 -7721 10641 -7720
rect 9900 -7788 9996 -7772
rect 10912 -7772 10928 -7348
rect 10992 -7772 11008 -7348
rect 11924 -7348 12020 -7332
rect 11331 -7400 11653 -7399
rect 11331 -7720 11332 -7400
rect 11652 -7720 11653 -7400
rect 11331 -7721 11653 -7720
rect 10912 -7788 11008 -7772
rect 11924 -7772 11940 -7348
rect 12004 -7772 12020 -7348
rect 12936 -7348 13032 -7332
rect 12343 -7400 12665 -7399
rect 12343 -7720 12344 -7400
rect 12664 -7720 12665 -7400
rect 12343 -7721 12665 -7720
rect 11924 -7788 12020 -7772
rect 12936 -7772 12952 -7348
rect 13016 -7772 13032 -7348
rect 13948 -7348 14044 -7332
rect 13355 -7400 13677 -7399
rect 13355 -7720 13356 -7400
rect 13676 -7720 13677 -7400
rect 13355 -7721 13677 -7720
rect 12936 -7788 13032 -7772
rect 13948 -7772 13964 -7348
rect 14028 -7772 14044 -7348
rect 14960 -7348 15056 -7332
rect 14367 -7400 14689 -7399
rect 14367 -7720 14368 -7400
rect 14688 -7720 14689 -7400
rect 14367 -7721 14689 -7720
rect 13948 -7788 14044 -7772
rect 14960 -7772 14976 -7348
rect 15040 -7772 15056 -7348
rect 15972 -7348 16068 -7332
rect 15379 -7400 15701 -7399
rect 15379 -7720 15380 -7400
rect 15700 -7720 15701 -7400
rect 15379 -7721 15701 -7720
rect 14960 -7788 15056 -7772
rect 15972 -7772 15988 -7348
rect 16052 -7772 16068 -7348
rect 16984 -7348 17080 -7332
rect 16391 -7400 16713 -7399
rect 16391 -7720 16392 -7400
rect 16712 -7720 16713 -7400
rect 16391 -7721 16713 -7720
rect 15972 -7788 16068 -7772
rect 16984 -7772 17000 -7348
rect 17064 -7772 17080 -7348
rect 16984 -7788 17080 -7772
rect -16412 -8068 -16316 -8052
rect -17005 -8120 -16683 -8119
rect -17005 -8440 -17004 -8120
rect -16684 -8440 -16683 -8120
rect -17005 -8441 -16683 -8440
rect -16412 -8492 -16396 -8068
rect -16332 -8492 -16316 -8068
rect -15400 -8068 -15304 -8052
rect -15993 -8120 -15671 -8119
rect -15993 -8440 -15992 -8120
rect -15672 -8440 -15671 -8120
rect -15993 -8441 -15671 -8440
rect -16412 -8508 -16316 -8492
rect -15400 -8492 -15384 -8068
rect -15320 -8492 -15304 -8068
rect -14388 -8068 -14292 -8052
rect -14981 -8120 -14659 -8119
rect -14981 -8440 -14980 -8120
rect -14660 -8440 -14659 -8120
rect -14981 -8441 -14659 -8440
rect -15400 -8508 -15304 -8492
rect -14388 -8492 -14372 -8068
rect -14308 -8492 -14292 -8068
rect -13376 -8068 -13280 -8052
rect -13969 -8120 -13647 -8119
rect -13969 -8440 -13968 -8120
rect -13648 -8440 -13647 -8120
rect -13969 -8441 -13647 -8440
rect -14388 -8508 -14292 -8492
rect -13376 -8492 -13360 -8068
rect -13296 -8492 -13280 -8068
rect -12364 -8068 -12268 -8052
rect -12957 -8120 -12635 -8119
rect -12957 -8440 -12956 -8120
rect -12636 -8440 -12635 -8120
rect -12957 -8441 -12635 -8440
rect -13376 -8508 -13280 -8492
rect -12364 -8492 -12348 -8068
rect -12284 -8492 -12268 -8068
rect -11352 -8068 -11256 -8052
rect -11945 -8120 -11623 -8119
rect -11945 -8440 -11944 -8120
rect -11624 -8440 -11623 -8120
rect -11945 -8441 -11623 -8440
rect -12364 -8508 -12268 -8492
rect -11352 -8492 -11336 -8068
rect -11272 -8492 -11256 -8068
rect -10340 -8068 -10244 -8052
rect -10933 -8120 -10611 -8119
rect -10933 -8440 -10932 -8120
rect -10612 -8440 -10611 -8120
rect -10933 -8441 -10611 -8440
rect -11352 -8508 -11256 -8492
rect -10340 -8492 -10324 -8068
rect -10260 -8492 -10244 -8068
rect -9328 -8068 -9232 -8052
rect -9921 -8120 -9599 -8119
rect -9921 -8440 -9920 -8120
rect -9600 -8440 -9599 -8120
rect -9921 -8441 -9599 -8440
rect -10340 -8508 -10244 -8492
rect -9328 -8492 -9312 -8068
rect -9248 -8492 -9232 -8068
rect -8316 -8068 -8220 -8052
rect -8909 -8120 -8587 -8119
rect -8909 -8440 -8908 -8120
rect -8588 -8440 -8587 -8120
rect -8909 -8441 -8587 -8440
rect -9328 -8508 -9232 -8492
rect -8316 -8492 -8300 -8068
rect -8236 -8492 -8220 -8068
rect -7304 -8068 -7208 -8052
rect -7897 -8120 -7575 -8119
rect -7897 -8440 -7896 -8120
rect -7576 -8440 -7575 -8120
rect -7897 -8441 -7575 -8440
rect -8316 -8508 -8220 -8492
rect -7304 -8492 -7288 -8068
rect -7224 -8492 -7208 -8068
rect -6292 -8068 -6196 -8052
rect -6885 -8120 -6563 -8119
rect -6885 -8440 -6884 -8120
rect -6564 -8440 -6563 -8120
rect -6885 -8441 -6563 -8440
rect -7304 -8508 -7208 -8492
rect -6292 -8492 -6276 -8068
rect -6212 -8492 -6196 -8068
rect -5280 -8068 -5184 -8052
rect -5873 -8120 -5551 -8119
rect -5873 -8440 -5872 -8120
rect -5552 -8440 -5551 -8120
rect -5873 -8441 -5551 -8440
rect -6292 -8508 -6196 -8492
rect -5280 -8492 -5264 -8068
rect -5200 -8492 -5184 -8068
rect -4268 -8068 -4172 -8052
rect -4861 -8120 -4539 -8119
rect -4861 -8440 -4860 -8120
rect -4540 -8440 -4539 -8120
rect -4861 -8441 -4539 -8440
rect -5280 -8508 -5184 -8492
rect -4268 -8492 -4252 -8068
rect -4188 -8492 -4172 -8068
rect -3256 -8068 -3160 -8052
rect -3849 -8120 -3527 -8119
rect -3849 -8440 -3848 -8120
rect -3528 -8440 -3527 -8120
rect -3849 -8441 -3527 -8440
rect -4268 -8508 -4172 -8492
rect -3256 -8492 -3240 -8068
rect -3176 -8492 -3160 -8068
rect -2244 -8068 -2148 -8052
rect -2837 -8120 -2515 -8119
rect -2837 -8440 -2836 -8120
rect -2516 -8440 -2515 -8120
rect -2837 -8441 -2515 -8440
rect -3256 -8508 -3160 -8492
rect -2244 -8492 -2228 -8068
rect -2164 -8492 -2148 -8068
rect -1232 -8068 -1136 -8052
rect -1825 -8120 -1503 -8119
rect -1825 -8440 -1824 -8120
rect -1504 -8440 -1503 -8120
rect -1825 -8441 -1503 -8440
rect -2244 -8508 -2148 -8492
rect -1232 -8492 -1216 -8068
rect -1152 -8492 -1136 -8068
rect -220 -8068 -124 -8052
rect -813 -8120 -491 -8119
rect -813 -8440 -812 -8120
rect -492 -8440 -491 -8120
rect -813 -8441 -491 -8440
rect -1232 -8508 -1136 -8492
rect -220 -8492 -204 -8068
rect -140 -8492 -124 -8068
rect 792 -8068 888 -8052
rect 199 -8120 521 -8119
rect 199 -8440 200 -8120
rect 520 -8440 521 -8120
rect 199 -8441 521 -8440
rect -220 -8508 -124 -8492
rect 792 -8492 808 -8068
rect 872 -8492 888 -8068
rect 1804 -8068 1900 -8052
rect 1211 -8120 1533 -8119
rect 1211 -8440 1212 -8120
rect 1532 -8440 1533 -8120
rect 1211 -8441 1533 -8440
rect 792 -8508 888 -8492
rect 1804 -8492 1820 -8068
rect 1884 -8492 1900 -8068
rect 2816 -8068 2912 -8052
rect 2223 -8120 2545 -8119
rect 2223 -8440 2224 -8120
rect 2544 -8440 2545 -8120
rect 2223 -8441 2545 -8440
rect 1804 -8508 1900 -8492
rect 2816 -8492 2832 -8068
rect 2896 -8492 2912 -8068
rect 3828 -8068 3924 -8052
rect 3235 -8120 3557 -8119
rect 3235 -8440 3236 -8120
rect 3556 -8440 3557 -8120
rect 3235 -8441 3557 -8440
rect 2816 -8508 2912 -8492
rect 3828 -8492 3844 -8068
rect 3908 -8492 3924 -8068
rect 4840 -8068 4936 -8052
rect 4247 -8120 4569 -8119
rect 4247 -8440 4248 -8120
rect 4568 -8440 4569 -8120
rect 4247 -8441 4569 -8440
rect 3828 -8508 3924 -8492
rect 4840 -8492 4856 -8068
rect 4920 -8492 4936 -8068
rect 5852 -8068 5948 -8052
rect 5259 -8120 5581 -8119
rect 5259 -8440 5260 -8120
rect 5580 -8440 5581 -8120
rect 5259 -8441 5581 -8440
rect 4840 -8508 4936 -8492
rect 5852 -8492 5868 -8068
rect 5932 -8492 5948 -8068
rect 6864 -8068 6960 -8052
rect 6271 -8120 6593 -8119
rect 6271 -8440 6272 -8120
rect 6592 -8440 6593 -8120
rect 6271 -8441 6593 -8440
rect 5852 -8508 5948 -8492
rect 6864 -8492 6880 -8068
rect 6944 -8492 6960 -8068
rect 7876 -8068 7972 -8052
rect 7283 -8120 7605 -8119
rect 7283 -8440 7284 -8120
rect 7604 -8440 7605 -8120
rect 7283 -8441 7605 -8440
rect 6864 -8508 6960 -8492
rect 7876 -8492 7892 -8068
rect 7956 -8492 7972 -8068
rect 8888 -8068 8984 -8052
rect 8295 -8120 8617 -8119
rect 8295 -8440 8296 -8120
rect 8616 -8440 8617 -8120
rect 8295 -8441 8617 -8440
rect 7876 -8508 7972 -8492
rect 8888 -8492 8904 -8068
rect 8968 -8492 8984 -8068
rect 9900 -8068 9996 -8052
rect 9307 -8120 9629 -8119
rect 9307 -8440 9308 -8120
rect 9628 -8440 9629 -8120
rect 9307 -8441 9629 -8440
rect 8888 -8508 8984 -8492
rect 9900 -8492 9916 -8068
rect 9980 -8492 9996 -8068
rect 10912 -8068 11008 -8052
rect 10319 -8120 10641 -8119
rect 10319 -8440 10320 -8120
rect 10640 -8440 10641 -8120
rect 10319 -8441 10641 -8440
rect 9900 -8508 9996 -8492
rect 10912 -8492 10928 -8068
rect 10992 -8492 11008 -8068
rect 11924 -8068 12020 -8052
rect 11331 -8120 11653 -8119
rect 11331 -8440 11332 -8120
rect 11652 -8440 11653 -8120
rect 11331 -8441 11653 -8440
rect 10912 -8508 11008 -8492
rect 11924 -8492 11940 -8068
rect 12004 -8492 12020 -8068
rect 12936 -8068 13032 -8052
rect 12343 -8120 12665 -8119
rect 12343 -8440 12344 -8120
rect 12664 -8440 12665 -8120
rect 12343 -8441 12665 -8440
rect 11924 -8508 12020 -8492
rect 12936 -8492 12952 -8068
rect 13016 -8492 13032 -8068
rect 13948 -8068 14044 -8052
rect 13355 -8120 13677 -8119
rect 13355 -8440 13356 -8120
rect 13676 -8440 13677 -8120
rect 13355 -8441 13677 -8440
rect 12936 -8508 13032 -8492
rect 13948 -8492 13964 -8068
rect 14028 -8492 14044 -8068
rect 14960 -8068 15056 -8052
rect 14367 -8120 14689 -8119
rect 14367 -8440 14368 -8120
rect 14688 -8440 14689 -8120
rect 14367 -8441 14689 -8440
rect 13948 -8508 14044 -8492
rect 14960 -8492 14976 -8068
rect 15040 -8492 15056 -8068
rect 15972 -8068 16068 -8052
rect 15379 -8120 15701 -8119
rect 15379 -8440 15380 -8120
rect 15700 -8440 15701 -8120
rect 15379 -8441 15701 -8440
rect 14960 -8508 15056 -8492
rect 15972 -8492 15988 -8068
rect 16052 -8492 16068 -8068
rect 16984 -8068 17080 -8052
rect 16391 -8120 16713 -8119
rect 16391 -8440 16392 -8120
rect 16712 -8440 16713 -8120
rect 16391 -8441 16713 -8440
rect 15972 -8508 16068 -8492
rect 16984 -8492 17000 -8068
rect 17064 -8492 17080 -8068
rect 16984 -8508 17080 -8492
rect -16412 -8788 -16316 -8772
rect -17005 -8840 -16683 -8839
rect -17005 -9160 -17004 -8840
rect -16684 -9160 -16683 -8840
rect -17005 -9161 -16683 -9160
rect -16412 -9212 -16396 -8788
rect -16332 -9212 -16316 -8788
rect -15400 -8788 -15304 -8772
rect -15993 -8840 -15671 -8839
rect -15993 -9160 -15992 -8840
rect -15672 -9160 -15671 -8840
rect -15993 -9161 -15671 -9160
rect -16412 -9228 -16316 -9212
rect -15400 -9212 -15384 -8788
rect -15320 -9212 -15304 -8788
rect -14388 -8788 -14292 -8772
rect -14981 -8840 -14659 -8839
rect -14981 -9160 -14980 -8840
rect -14660 -9160 -14659 -8840
rect -14981 -9161 -14659 -9160
rect -15400 -9228 -15304 -9212
rect -14388 -9212 -14372 -8788
rect -14308 -9212 -14292 -8788
rect -13376 -8788 -13280 -8772
rect -13969 -8840 -13647 -8839
rect -13969 -9160 -13968 -8840
rect -13648 -9160 -13647 -8840
rect -13969 -9161 -13647 -9160
rect -14388 -9228 -14292 -9212
rect -13376 -9212 -13360 -8788
rect -13296 -9212 -13280 -8788
rect -12364 -8788 -12268 -8772
rect -12957 -8840 -12635 -8839
rect -12957 -9160 -12956 -8840
rect -12636 -9160 -12635 -8840
rect -12957 -9161 -12635 -9160
rect -13376 -9228 -13280 -9212
rect -12364 -9212 -12348 -8788
rect -12284 -9212 -12268 -8788
rect -11352 -8788 -11256 -8772
rect -11945 -8840 -11623 -8839
rect -11945 -9160 -11944 -8840
rect -11624 -9160 -11623 -8840
rect -11945 -9161 -11623 -9160
rect -12364 -9228 -12268 -9212
rect -11352 -9212 -11336 -8788
rect -11272 -9212 -11256 -8788
rect -10340 -8788 -10244 -8772
rect -10933 -8840 -10611 -8839
rect -10933 -9160 -10932 -8840
rect -10612 -9160 -10611 -8840
rect -10933 -9161 -10611 -9160
rect -11352 -9228 -11256 -9212
rect -10340 -9212 -10324 -8788
rect -10260 -9212 -10244 -8788
rect -9328 -8788 -9232 -8772
rect -9921 -8840 -9599 -8839
rect -9921 -9160 -9920 -8840
rect -9600 -9160 -9599 -8840
rect -9921 -9161 -9599 -9160
rect -10340 -9228 -10244 -9212
rect -9328 -9212 -9312 -8788
rect -9248 -9212 -9232 -8788
rect -8316 -8788 -8220 -8772
rect -8909 -8840 -8587 -8839
rect -8909 -9160 -8908 -8840
rect -8588 -9160 -8587 -8840
rect -8909 -9161 -8587 -9160
rect -9328 -9228 -9232 -9212
rect -8316 -9212 -8300 -8788
rect -8236 -9212 -8220 -8788
rect -7304 -8788 -7208 -8772
rect -7897 -8840 -7575 -8839
rect -7897 -9160 -7896 -8840
rect -7576 -9160 -7575 -8840
rect -7897 -9161 -7575 -9160
rect -8316 -9228 -8220 -9212
rect -7304 -9212 -7288 -8788
rect -7224 -9212 -7208 -8788
rect -6292 -8788 -6196 -8772
rect -6885 -8840 -6563 -8839
rect -6885 -9160 -6884 -8840
rect -6564 -9160 -6563 -8840
rect -6885 -9161 -6563 -9160
rect -7304 -9228 -7208 -9212
rect -6292 -9212 -6276 -8788
rect -6212 -9212 -6196 -8788
rect -5280 -8788 -5184 -8772
rect -5873 -8840 -5551 -8839
rect -5873 -9160 -5872 -8840
rect -5552 -9160 -5551 -8840
rect -5873 -9161 -5551 -9160
rect -6292 -9228 -6196 -9212
rect -5280 -9212 -5264 -8788
rect -5200 -9212 -5184 -8788
rect -4268 -8788 -4172 -8772
rect -4861 -8840 -4539 -8839
rect -4861 -9160 -4860 -8840
rect -4540 -9160 -4539 -8840
rect -4861 -9161 -4539 -9160
rect -5280 -9228 -5184 -9212
rect -4268 -9212 -4252 -8788
rect -4188 -9212 -4172 -8788
rect -3256 -8788 -3160 -8772
rect -3849 -8840 -3527 -8839
rect -3849 -9160 -3848 -8840
rect -3528 -9160 -3527 -8840
rect -3849 -9161 -3527 -9160
rect -4268 -9228 -4172 -9212
rect -3256 -9212 -3240 -8788
rect -3176 -9212 -3160 -8788
rect -2244 -8788 -2148 -8772
rect -2837 -8840 -2515 -8839
rect -2837 -9160 -2836 -8840
rect -2516 -9160 -2515 -8840
rect -2837 -9161 -2515 -9160
rect -3256 -9228 -3160 -9212
rect -2244 -9212 -2228 -8788
rect -2164 -9212 -2148 -8788
rect -1232 -8788 -1136 -8772
rect -1825 -8840 -1503 -8839
rect -1825 -9160 -1824 -8840
rect -1504 -9160 -1503 -8840
rect -1825 -9161 -1503 -9160
rect -2244 -9228 -2148 -9212
rect -1232 -9212 -1216 -8788
rect -1152 -9212 -1136 -8788
rect -220 -8788 -124 -8772
rect -813 -8840 -491 -8839
rect -813 -9160 -812 -8840
rect -492 -9160 -491 -8840
rect -813 -9161 -491 -9160
rect -1232 -9228 -1136 -9212
rect -220 -9212 -204 -8788
rect -140 -9212 -124 -8788
rect 792 -8788 888 -8772
rect 199 -8840 521 -8839
rect 199 -9160 200 -8840
rect 520 -9160 521 -8840
rect 199 -9161 521 -9160
rect -220 -9228 -124 -9212
rect 792 -9212 808 -8788
rect 872 -9212 888 -8788
rect 1804 -8788 1900 -8772
rect 1211 -8840 1533 -8839
rect 1211 -9160 1212 -8840
rect 1532 -9160 1533 -8840
rect 1211 -9161 1533 -9160
rect 792 -9228 888 -9212
rect 1804 -9212 1820 -8788
rect 1884 -9212 1900 -8788
rect 2816 -8788 2912 -8772
rect 2223 -8840 2545 -8839
rect 2223 -9160 2224 -8840
rect 2544 -9160 2545 -8840
rect 2223 -9161 2545 -9160
rect 1804 -9228 1900 -9212
rect 2816 -9212 2832 -8788
rect 2896 -9212 2912 -8788
rect 3828 -8788 3924 -8772
rect 3235 -8840 3557 -8839
rect 3235 -9160 3236 -8840
rect 3556 -9160 3557 -8840
rect 3235 -9161 3557 -9160
rect 2816 -9228 2912 -9212
rect 3828 -9212 3844 -8788
rect 3908 -9212 3924 -8788
rect 4840 -8788 4936 -8772
rect 4247 -8840 4569 -8839
rect 4247 -9160 4248 -8840
rect 4568 -9160 4569 -8840
rect 4247 -9161 4569 -9160
rect 3828 -9228 3924 -9212
rect 4840 -9212 4856 -8788
rect 4920 -9212 4936 -8788
rect 5852 -8788 5948 -8772
rect 5259 -8840 5581 -8839
rect 5259 -9160 5260 -8840
rect 5580 -9160 5581 -8840
rect 5259 -9161 5581 -9160
rect 4840 -9228 4936 -9212
rect 5852 -9212 5868 -8788
rect 5932 -9212 5948 -8788
rect 6864 -8788 6960 -8772
rect 6271 -8840 6593 -8839
rect 6271 -9160 6272 -8840
rect 6592 -9160 6593 -8840
rect 6271 -9161 6593 -9160
rect 5852 -9228 5948 -9212
rect 6864 -9212 6880 -8788
rect 6944 -9212 6960 -8788
rect 7876 -8788 7972 -8772
rect 7283 -8840 7605 -8839
rect 7283 -9160 7284 -8840
rect 7604 -9160 7605 -8840
rect 7283 -9161 7605 -9160
rect 6864 -9228 6960 -9212
rect 7876 -9212 7892 -8788
rect 7956 -9212 7972 -8788
rect 8888 -8788 8984 -8772
rect 8295 -8840 8617 -8839
rect 8295 -9160 8296 -8840
rect 8616 -9160 8617 -8840
rect 8295 -9161 8617 -9160
rect 7876 -9228 7972 -9212
rect 8888 -9212 8904 -8788
rect 8968 -9212 8984 -8788
rect 9900 -8788 9996 -8772
rect 9307 -8840 9629 -8839
rect 9307 -9160 9308 -8840
rect 9628 -9160 9629 -8840
rect 9307 -9161 9629 -9160
rect 8888 -9228 8984 -9212
rect 9900 -9212 9916 -8788
rect 9980 -9212 9996 -8788
rect 10912 -8788 11008 -8772
rect 10319 -8840 10641 -8839
rect 10319 -9160 10320 -8840
rect 10640 -9160 10641 -8840
rect 10319 -9161 10641 -9160
rect 9900 -9228 9996 -9212
rect 10912 -9212 10928 -8788
rect 10992 -9212 11008 -8788
rect 11924 -8788 12020 -8772
rect 11331 -8840 11653 -8839
rect 11331 -9160 11332 -8840
rect 11652 -9160 11653 -8840
rect 11331 -9161 11653 -9160
rect 10912 -9228 11008 -9212
rect 11924 -9212 11940 -8788
rect 12004 -9212 12020 -8788
rect 12936 -8788 13032 -8772
rect 12343 -8840 12665 -8839
rect 12343 -9160 12344 -8840
rect 12664 -9160 12665 -8840
rect 12343 -9161 12665 -9160
rect 11924 -9228 12020 -9212
rect 12936 -9212 12952 -8788
rect 13016 -9212 13032 -8788
rect 13948 -8788 14044 -8772
rect 13355 -8840 13677 -8839
rect 13355 -9160 13356 -8840
rect 13676 -9160 13677 -8840
rect 13355 -9161 13677 -9160
rect 12936 -9228 13032 -9212
rect 13948 -9212 13964 -8788
rect 14028 -9212 14044 -8788
rect 14960 -8788 15056 -8772
rect 14367 -8840 14689 -8839
rect 14367 -9160 14368 -8840
rect 14688 -9160 14689 -8840
rect 14367 -9161 14689 -9160
rect 13948 -9228 14044 -9212
rect 14960 -9212 14976 -8788
rect 15040 -9212 15056 -8788
rect 15972 -8788 16068 -8772
rect 15379 -8840 15701 -8839
rect 15379 -9160 15380 -8840
rect 15700 -9160 15701 -8840
rect 15379 -9161 15701 -9160
rect 14960 -9228 15056 -9212
rect 15972 -9212 15988 -8788
rect 16052 -9212 16068 -8788
rect 16984 -8788 17080 -8772
rect 16391 -8840 16713 -8839
rect 16391 -9160 16392 -8840
rect 16712 -9160 16713 -8840
rect 16391 -9161 16713 -9160
rect 15972 -9228 16068 -9212
rect 16984 -9212 17000 -8788
rect 17064 -9212 17080 -8788
rect 16984 -9228 17080 -9212
rect -16412 -9508 -16316 -9492
rect -17005 -9560 -16683 -9559
rect -17005 -9880 -17004 -9560
rect -16684 -9880 -16683 -9560
rect -17005 -9881 -16683 -9880
rect -16412 -9932 -16396 -9508
rect -16332 -9932 -16316 -9508
rect -15400 -9508 -15304 -9492
rect -15993 -9560 -15671 -9559
rect -15993 -9880 -15992 -9560
rect -15672 -9880 -15671 -9560
rect -15993 -9881 -15671 -9880
rect -16412 -9948 -16316 -9932
rect -15400 -9932 -15384 -9508
rect -15320 -9932 -15304 -9508
rect -14388 -9508 -14292 -9492
rect -14981 -9560 -14659 -9559
rect -14981 -9880 -14980 -9560
rect -14660 -9880 -14659 -9560
rect -14981 -9881 -14659 -9880
rect -15400 -9948 -15304 -9932
rect -14388 -9932 -14372 -9508
rect -14308 -9932 -14292 -9508
rect -13376 -9508 -13280 -9492
rect -13969 -9560 -13647 -9559
rect -13969 -9880 -13968 -9560
rect -13648 -9880 -13647 -9560
rect -13969 -9881 -13647 -9880
rect -14388 -9948 -14292 -9932
rect -13376 -9932 -13360 -9508
rect -13296 -9932 -13280 -9508
rect -12364 -9508 -12268 -9492
rect -12957 -9560 -12635 -9559
rect -12957 -9880 -12956 -9560
rect -12636 -9880 -12635 -9560
rect -12957 -9881 -12635 -9880
rect -13376 -9948 -13280 -9932
rect -12364 -9932 -12348 -9508
rect -12284 -9932 -12268 -9508
rect -11352 -9508 -11256 -9492
rect -11945 -9560 -11623 -9559
rect -11945 -9880 -11944 -9560
rect -11624 -9880 -11623 -9560
rect -11945 -9881 -11623 -9880
rect -12364 -9948 -12268 -9932
rect -11352 -9932 -11336 -9508
rect -11272 -9932 -11256 -9508
rect -10340 -9508 -10244 -9492
rect -10933 -9560 -10611 -9559
rect -10933 -9880 -10932 -9560
rect -10612 -9880 -10611 -9560
rect -10933 -9881 -10611 -9880
rect -11352 -9948 -11256 -9932
rect -10340 -9932 -10324 -9508
rect -10260 -9932 -10244 -9508
rect -9328 -9508 -9232 -9492
rect -9921 -9560 -9599 -9559
rect -9921 -9880 -9920 -9560
rect -9600 -9880 -9599 -9560
rect -9921 -9881 -9599 -9880
rect -10340 -9948 -10244 -9932
rect -9328 -9932 -9312 -9508
rect -9248 -9932 -9232 -9508
rect -8316 -9508 -8220 -9492
rect -8909 -9560 -8587 -9559
rect -8909 -9880 -8908 -9560
rect -8588 -9880 -8587 -9560
rect -8909 -9881 -8587 -9880
rect -9328 -9948 -9232 -9932
rect -8316 -9932 -8300 -9508
rect -8236 -9932 -8220 -9508
rect -7304 -9508 -7208 -9492
rect -7897 -9560 -7575 -9559
rect -7897 -9880 -7896 -9560
rect -7576 -9880 -7575 -9560
rect -7897 -9881 -7575 -9880
rect -8316 -9948 -8220 -9932
rect -7304 -9932 -7288 -9508
rect -7224 -9932 -7208 -9508
rect -6292 -9508 -6196 -9492
rect -6885 -9560 -6563 -9559
rect -6885 -9880 -6884 -9560
rect -6564 -9880 -6563 -9560
rect -6885 -9881 -6563 -9880
rect -7304 -9948 -7208 -9932
rect -6292 -9932 -6276 -9508
rect -6212 -9932 -6196 -9508
rect -5280 -9508 -5184 -9492
rect -5873 -9560 -5551 -9559
rect -5873 -9880 -5872 -9560
rect -5552 -9880 -5551 -9560
rect -5873 -9881 -5551 -9880
rect -6292 -9948 -6196 -9932
rect -5280 -9932 -5264 -9508
rect -5200 -9932 -5184 -9508
rect -4268 -9508 -4172 -9492
rect -4861 -9560 -4539 -9559
rect -4861 -9880 -4860 -9560
rect -4540 -9880 -4539 -9560
rect -4861 -9881 -4539 -9880
rect -5280 -9948 -5184 -9932
rect -4268 -9932 -4252 -9508
rect -4188 -9932 -4172 -9508
rect -3256 -9508 -3160 -9492
rect -3849 -9560 -3527 -9559
rect -3849 -9880 -3848 -9560
rect -3528 -9880 -3527 -9560
rect -3849 -9881 -3527 -9880
rect -4268 -9948 -4172 -9932
rect -3256 -9932 -3240 -9508
rect -3176 -9932 -3160 -9508
rect -2244 -9508 -2148 -9492
rect -2837 -9560 -2515 -9559
rect -2837 -9880 -2836 -9560
rect -2516 -9880 -2515 -9560
rect -2837 -9881 -2515 -9880
rect -3256 -9948 -3160 -9932
rect -2244 -9932 -2228 -9508
rect -2164 -9932 -2148 -9508
rect -1232 -9508 -1136 -9492
rect -1825 -9560 -1503 -9559
rect -1825 -9880 -1824 -9560
rect -1504 -9880 -1503 -9560
rect -1825 -9881 -1503 -9880
rect -2244 -9948 -2148 -9932
rect -1232 -9932 -1216 -9508
rect -1152 -9932 -1136 -9508
rect -220 -9508 -124 -9492
rect -813 -9560 -491 -9559
rect -813 -9880 -812 -9560
rect -492 -9880 -491 -9560
rect -813 -9881 -491 -9880
rect -1232 -9948 -1136 -9932
rect -220 -9932 -204 -9508
rect -140 -9932 -124 -9508
rect 792 -9508 888 -9492
rect 199 -9560 521 -9559
rect 199 -9880 200 -9560
rect 520 -9880 521 -9560
rect 199 -9881 521 -9880
rect -220 -9948 -124 -9932
rect 792 -9932 808 -9508
rect 872 -9932 888 -9508
rect 1804 -9508 1900 -9492
rect 1211 -9560 1533 -9559
rect 1211 -9880 1212 -9560
rect 1532 -9880 1533 -9560
rect 1211 -9881 1533 -9880
rect 792 -9948 888 -9932
rect 1804 -9932 1820 -9508
rect 1884 -9932 1900 -9508
rect 2816 -9508 2912 -9492
rect 2223 -9560 2545 -9559
rect 2223 -9880 2224 -9560
rect 2544 -9880 2545 -9560
rect 2223 -9881 2545 -9880
rect 1804 -9948 1900 -9932
rect 2816 -9932 2832 -9508
rect 2896 -9932 2912 -9508
rect 3828 -9508 3924 -9492
rect 3235 -9560 3557 -9559
rect 3235 -9880 3236 -9560
rect 3556 -9880 3557 -9560
rect 3235 -9881 3557 -9880
rect 2816 -9948 2912 -9932
rect 3828 -9932 3844 -9508
rect 3908 -9932 3924 -9508
rect 4840 -9508 4936 -9492
rect 4247 -9560 4569 -9559
rect 4247 -9880 4248 -9560
rect 4568 -9880 4569 -9560
rect 4247 -9881 4569 -9880
rect 3828 -9948 3924 -9932
rect 4840 -9932 4856 -9508
rect 4920 -9932 4936 -9508
rect 5852 -9508 5948 -9492
rect 5259 -9560 5581 -9559
rect 5259 -9880 5260 -9560
rect 5580 -9880 5581 -9560
rect 5259 -9881 5581 -9880
rect 4840 -9948 4936 -9932
rect 5852 -9932 5868 -9508
rect 5932 -9932 5948 -9508
rect 6864 -9508 6960 -9492
rect 6271 -9560 6593 -9559
rect 6271 -9880 6272 -9560
rect 6592 -9880 6593 -9560
rect 6271 -9881 6593 -9880
rect 5852 -9948 5948 -9932
rect 6864 -9932 6880 -9508
rect 6944 -9932 6960 -9508
rect 7876 -9508 7972 -9492
rect 7283 -9560 7605 -9559
rect 7283 -9880 7284 -9560
rect 7604 -9880 7605 -9560
rect 7283 -9881 7605 -9880
rect 6864 -9948 6960 -9932
rect 7876 -9932 7892 -9508
rect 7956 -9932 7972 -9508
rect 8888 -9508 8984 -9492
rect 8295 -9560 8617 -9559
rect 8295 -9880 8296 -9560
rect 8616 -9880 8617 -9560
rect 8295 -9881 8617 -9880
rect 7876 -9948 7972 -9932
rect 8888 -9932 8904 -9508
rect 8968 -9932 8984 -9508
rect 9900 -9508 9996 -9492
rect 9307 -9560 9629 -9559
rect 9307 -9880 9308 -9560
rect 9628 -9880 9629 -9560
rect 9307 -9881 9629 -9880
rect 8888 -9948 8984 -9932
rect 9900 -9932 9916 -9508
rect 9980 -9932 9996 -9508
rect 10912 -9508 11008 -9492
rect 10319 -9560 10641 -9559
rect 10319 -9880 10320 -9560
rect 10640 -9880 10641 -9560
rect 10319 -9881 10641 -9880
rect 9900 -9948 9996 -9932
rect 10912 -9932 10928 -9508
rect 10992 -9932 11008 -9508
rect 11924 -9508 12020 -9492
rect 11331 -9560 11653 -9559
rect 11331 -9880 11332 -9560
rect 11652 -9880 11653 -9560
rect 11331 -9881 11653 -9880
rect 10912 -9948 11008 -9932
rect 11924 -9932 11940 -9508
rect 12004 -9932 12020 -9508
rect 12936 -9508 13032 -9492
rect 12343 -9560 12665 -9559
rect 12343 -9880 12344 -9560
rect 12664 -9880 12665 -9560
rect 12343 -9881 12665 -9880
rect 11924 -9948 12020 -9932
rect 12936 -9932 12952 -9508
rect 13016 -9932 13032 -9508
rect 13948 -9508 14044 -9492
rect 13355 -9560 13677 -9559
rect 13355 -9880 13356 -9560
rect 13676 -9880 13677 -9560
rect 13355 -9881 13677 -9880
rect 12936 -9948 13032 -9932
rect 13948 -9932 13964 -9508
rect 14028 -9932 14044 -9508
rect 14960 -9508 15056 -9492
rect 14367 -9560 14689 -9559
rect 14367 -9880 14368 -9560
rect 14688 -9880 14689 -9560
rect 14367 -9881 14689 -9880
rect 13948 -9948 14044 -9932
rect 14960 -9932 14976 -9508
rect 15040 -9932 15056 -9508
rect 15972 -9508 16068 -9492
rect 15379 -9560 15701 -9559
rect 15379 -9880 15380 -9560
rect 15700 -9880 15701 -9560
rect 15379 -9881 15701 -9880
rect 14960 -9948 15056 -9932
rect 15972 -9932 15988 -9508
rect 16052 -9932 16068 -9508
rect 16984 -9508 17080 -9492
rect 16391 -9560 16713 -9559
rect 16391 -9880 16392 -9560
rect 16712 -9880 16713 -9560
rect 16391 -9881 16713 -9880
rect 15972 -9948 16068 -9932
rect 16984 -9932 17000 -9508
rect 17064 -9932 17080 -9508
rect 16984 -9948 17080 -9932
rect -16412 -10228 -16316 -10212
rect -17005 -10280 -16683 -10279
rect -17005 -10600 -17004 -10280
rect -16684 -10600 -16683 -10280
rect -17005 -10601 -16683 -10600
rect -16412 -10652 -16396 -10228
rect -16332 -10652 -16316 -10228
rect -15400 -10228 -15304 -10212
rect -15993 -10280 -15671 -10279
rect -15993 -10600 -15992 -10280
rect -15672 -10600 -15671 -10280
rect -15993 -10601 -15671 -10600
rect -16412 -10668 -16316 -10652
rect -15400 -10652 -15384 -10228
rect -15320 -10652 -15304 -10228
rect -14388 -10228 -14292 -10212
rect -14981 -10280 -14659 -10279
rect -14981 -10600 -14980 -10280
rect -14660 -10600 -14659 -10280
rect -14981 -10601 -14659 -10600
rect -15400 -10668 -15304 -10652
rect -14388 -10652 -14372 -10228
rect -14308 -10652 -14292 -10228
rect -13376 -10228 -13280 -10212
rect -13969 -10280 -13647 -10279
rect -13969 -10600 -13968 -10280
rect -13648 -10600 -13647 -10280
rect -13969 -10601 -13647 -10600
rect -14388 -10668 -14292 -10652
rect -13376 -10652 -13360 -10228
rect -13296 -10652 -13280 -10228
rect -12364 -10228 -12268 -10212
rect -12957 -10280 -12635 -10279
rect -12957 -10600 -12956 -10280
rect -12636 -10600 -12635 -10280
rect -12957 -10601 -12635 -10600
rect -13376 -10668 -13280 -10652
rect -12364 -10652 -12348 -10228
rect -12284 -10652 -12268 -10228
rect -11352 -10228 -11256 -10212
rect -11945 -10280 -11623 -10279
rect -11945 -10600 -11944 -10280
rect -11624 -10600 -11623 -10280
rect -11945 -10601 -11623 -10600
rect -12364 -10668 -12268 -10652
rect -11352 -10652 -11336 -10228
rect -11272 -10652 -11256 -10228
rect -10340 -10228 -10244 -10212
rect -10933 -10280 -10611 -10279
rect -10933 -10600 -10932 -10280
rect -10612 -10600 -10611 -10280
rect -10933 -10601 -10611 -10600
rect -11352 -10668 -11256 -10652
rect -10340 -10652 -10324 -10228
rect -10260 -10652 -10244 -10228
rect -9328 -10228 -9232 -10212
rect -9921 -10280 -9599 -10279
rect -9921 -10600 -9920 -10280
rect -9600 -10600 -9599 -10280
rect -9921 -10601 -9599 -10600
rect -10340 -10668 -10244 -10652
rect -9328 -10652 -9312 -10228
rect -9248 -10652 -9232 -10228
rect -8316 -10228 -8220 -10212
rect -8909 -10280 -8587 -10279
rect -8909 -10600 -8908 -10280
rect -8588 -10600 -8587 -10280
rect -8909 -10601 -8587 -10600
rect -9328 -10668 -9232 -10652
rect -8316 -10652 -8300 -10228
rect -8236 -10652 -8220 -10228
rect -7304 -10228 -7208 -10212
rect -7897 -10280 -7575 -10279
rect -7897 -10600 -7896 -10280
rect -7576 -10600 -7575 -10280
rect -7897 -10601 -7575 -10600
rect -8316 -10668 -8220 -10652
rect -7304 -10652 -7288 -10228
rect -7224 -10652 -7208 -10228
rect -6292 -10228 -6196 -10212
rect -6885 -10280 -6563 -10279
rect -6885 -10600 -6884 -10280
rect -6564 -10600 -6563 -10280
rect -6885 -10601 -6563 -10600
rect -7304 -10668 -7208 -10652
rect -6292 -10652 -6276 -10228
rect -6212 -10652 -6196 -10228
rect -5280 -10228 -5184 -10212
rect -5873 -10280 -5551 -10279
rect -5873 -10600 -5872 -10280
rect -5552 -10600 -5551 -10280
rect -5873 -10601 -5551 -10600
rect -6292 -10668 -6196 -10652
rect -5280 -10652 -5264 -10228
rect -5200 -10652 -5184 -10228
rect -4268 -10228 -4172 -10212
rect -4861 -10280 -4539 -10279
rect -4861 -10600 -4860 -10280
rect -4540 -10600 -4539 -10280
rect -4861 -10601 -4539 -10600
rect -5280 -10668 -5184 -10652
rect -4268 -10652 -4252 -10228
rect -4188 -10652 -4172 -10228
rect -3256 -10228 -3160 -10212
rect -3849 -10280 -3527 -10279
rect -3849 -10600 -3848 -10280
rect -3528 -10600 -3527 -10280
rect -3849 -10601 -3527 -10600
rect -4268 -10668 -4172 -10652
rect -3256 -10652 -3240 -10228
rect -3176 -10652 -3160 -10228
rect -2244 -10228 -2148 -10212
rect -2837 -10280 -2515 -10279
rect -2837 -10600 -2836 -10280
rect -2516 -10600 -2515 -10280
rect -2837 -10601 -2515 -10600
rect -3256 -10668 -3160 -10652
rect -2244 -10652 -2228 -10228
rect -2164 -10652 -2148 -10228
rect -1232 -10228 -1136 -10212
rect -1825 -10280 -1503 -10279
rect -1825 -10600 -1824 -10280
rect -1504 -10600 -1503 -10280
rect -1825 -10601 -1503 -10600
rect -2244 -10668 -2148 -10652
rect -1232 -10652 -1216 -10228
rect -1152 -10652 -1136 -10228
rect -220 -10228 -124 -10212
rect -813 -10280 -491 -10279
rect -813 -10600 -812 -10280
rect -492 -10600 -491 -10280
rect -813 -10601 -491 -10600
rect -1232 -10668 -1136 -10652
rect -220 -10652 -204 -10228
rect -140 -10652 -124 -10228
rect 792 -10228 888 -10212
rect 199 -10280 521 -10279
rect 199 -10600 200 -10280
rect 520 -10600 521 -10280
rect 199 -10601 521 -10600
rect -220 -10668 -124 -10652
rect 792 -10652 808 -10228
rect 872 -10652 888 -10228
rect 1804 -10228 1900 -10212
rect 1211 -10280 1533 -10279
rect 1211 -10600 1212 -10280
rect 1532 -10600 1533 -10280
rect 1211 -10601 1533 -10600
rect 792 -10668 888 -10652
rect 1804 -10652 1820 -10228
rect 1884 -10652 1900 -10228
rect 2816 -10228 2912 -10212
rect 2223 -10280 2545 -10279
rect 2223 -10600 2224 -10280
rect 2544 -10600 2545 -10280
rect 2223 -10601 2545 -10600
rect 1804 -10668 1900 -10652
rect 2816 -10652 2832 -10228
rect 2896 -10652 2912 -10228
rect 3828 -10228 3924 -10212
rect 3235 -10280 3557 -10279
rect 3235 -10600 3236 -10280
rect 3556 -10600 3557 -10280
rect 3235 -10601 3557 -10600
rect 2816 -10668 2912 -10652
rect 3828 -10652 3844 -10228
rect 3908 -10652 3924 -10228
rect 4840 -10228 4936 -10212
rect 4247 -10280 4569 -10279
rect 4247 -10600 4248 -10280
rect 4568 -10600 4569 -10280
rect 4247 -10601 4569 -10600
rect 3828 -10668 3924 -10652
rect 4840 -10652 4856 -10228
rect 4920 -10652 4936 -10228
rect 5852 -10228 5948 -10212
rect 5259 -10280 5581 -10279
rect 5259 -10600 5260 -10280
rect 5580 -10600 5581 -10280
rect 5259 -10601 5581 -10600
rect 4840 -10668 4936 -10652
rect 5852 -10652 5868 -10228
rect 5932 -10652 5948 -10228
rect 6864 -10228 6960 -10212
rect 6271 -10280 6593 -10279
rect 6271 -10600 6272 -10280
rect 6592 -10600 6593 -10280
rect 6271 -10601 6593 -10600
rect 5852 -10668 5948 -10652
rect 6864 -10652 6880 -10228
rect 6944 -10652 6960 -10228
rect 7876 -10228 7972 -10212
rect 7283 -10280 7605 -10279
rect 7283 -10600 7284 -10280
rect 7604 -10600 7605 -10280
rect 7283 -10601 7605 -10600
rect 6864 -10668 6960 -10652
rect 7876 -10652 7892 -10228
rect 7956 -10652 7972 -10228
rect 8888 -10228 8984 -10212
rect 8295 -10280 8617 -10279
rect 8295 -10600 8296 -10280
rect 8616 -10600 8617 -10280
rect 8295 -10601 8617 -10600
rect 7876 -10668 7972 -10652
rect 8888 -10652 8904 -10228
rect 8968 -10652 8984 -10228
rect 9900 -10228 9996 -10212
rect 9307 -10280 9629 -10279
rect 9307 -10600 9308 -10280
rect 9628 -10600 9629 -10280
rect 9307 -10601 9629 -10600
rect 8888 -10668 8984 -10652
rect 9900 -10652 9916 -10228
rect 9980 -10652 9996 -10228
rect 10912 -10228 11008 -10212
rect 10319 -10280 10641 -10279
rect 10319 -10600 10320 -10280
rect 10640 -10600 10641 -10280
rect 10319 -10601 10641 -10600
rect 9900 -10668 9996 -10652
rect 10912 -10652 10928 -10228
rect 10992 -10652 11008 -10228
rect 11924 -10228 12020 -10212
rect 11331 -10280 11653 -10279
rect 11331 -10600 11332 -10280
rect 11652 -10600 11653 -10280
rect 11331 -10601 11653 -10600
rect 10912 -10668 11008 -10652
rect 11924 -10652 11940 -10228
rect 12004 -10652 12020 -10228
rect 12936 -10228 13032 -10212
rect 12343 -10280 12665 -10279
rect 12343 -10600 12344 -10280
rect 12664 -10600 12665 -10280
rect 12343 -10601 12665 -10600
rect 11924 -10668 12020 -10652
rect 12936 -10652 12952 -10228
rect 13016 -10652 13032 -10228
rect 13948 -10228 14044 -10212
rect 13355 -10280 13677 -10279
rect 13355 -10600 13356 -10280
rect 13676 -10600 13677 -10280
rect 13355 -10601 13677 -10600
rect 12936 -10668 13032 -10652
rect 13948 -10652 13964 -10228
rect 14028 -10652 14044 -10228
rect 14960 -10228 15056 -10212
rect 14367 -10280 14689 -10279
rect 14367 -10600 14368 -10280
rect 14688 -10600 14689 -10280
rect 14367 -10601 14689 -10600
rect 13948 -10668 14044 -10652
rect 14960 -10652 14976 -10228
rect 15040 -10652 15056 -10228
rect 15972 -10228 16068 -10212
rect 15379 -10280 15701 -10279
rect 15379 -10600 15380 -10280
rect 15700 -10600 15701 -10280
rect 15379 -10601 15701 -10600
rect 14960 -10668 15056 -10652
rect 15972 -10652 15988 -10228
rect 16052 -10652 16068 -10228
rect 16984 -10228 17080 -10212
rect 16391 -10280 16713 -10279
rect 16391 -10600 16392 -10280
rect 16712 -10600 16713 -10280
rect 16391 -10601 16713 -10600
rect 15972 -10668 16068 -10652
rect 16984 -10652 17000 -10228
rect 17064 -10652 17080 -10228
rect 16984 -10668 17080 -10652
rect -16412 -10948 -16316 -10932
rect -17005 -11000 -16683 -10999
rect -17005 -11320 -17004 -11000
rect -16684 -11320 -16683 -11000
rect -17005 -11321 -16683 -11320
rect -16412 -11372 -16396 -10948
rect -16332 -11372 -16316 -10948
rect -15400 -10948 -15304 -10932
rect -15993 -11000 -15671 -10999
rect -15993 -11320 -15992 -11000
rect -15672 -11320 -15671 -11000
rect -15993 -11321 -15671 -11320
rect -16412 -11388 -16316 -11372
rect -15400 -11372 -15384 -10948
rect -15320 -11372 -15304 -10948
rect -14388 -10948 -14292 -10932
rect -14981 -11000 -14659 -10999
rect -14981 -11320 -14980 -11000
rect -14660 -11320 -14659 -11000
rect -14981 -11321 -14659 -11320
rect -15400 -11388 -15304 -11372
rect -14388 -11372 -14372 -10948
rect -14308 -11372 -14292 -10948
rect -13376 -10948 -13280 -10932
rect -13969 -11000 -13647 -10999
rect -13969 -11320 -13968 -11000
rect -13648 -11320 -13647 -11000
rect -13969 -11321 -13647 -11320
rect -14388 -11388 -14292 -11372
rect -13376 -11372 -13360 -10948
rect -13296 -11372 -13280 -10948
rect -12364 -10948 -12268 -10932
rect -12957 -11000 -12635 -10999
rect -12957 -11320 -12956 -11000
rect -12636 -11320 -12635 -11000
rect -12957 -11321 -12635 -11320
rect -13376 -11388 -13280 -11372
rect -12364 -11372 -12348 -10948
rect -12284 -11372 -12268 -10948
rect -11352 -10948 -11256 -10932
rect -11945 -11000 -11623 -10999
rect -11945 -11320 -11944 -11000
rect -11624 -11320 -11623 -11000
rect -11945 -11321 -11623 -11320
rect -12364 -11388 -12268 -11372
rect -11352 -11372 -11336 -10948
rect -11272 -11372 -11256 -10948
rect -10340 -10948 -10244 -10932
rect -10933 -11000 -10611 -10999
rect -10933 -11320 -10932 -11000
rect -10612 -11320 -10611 -11000
rect -10933 -11321 -10611 -11320
rect -11352 -11388 -11256 -11372
rect -10340 -11372 -10324 -10948
rect -10260 -11372 -10244 -10948
rect -9328 -10948 -9232 -10932
rect -9921 -11000 -9599 -10999
rect -9921 -11320 -9920 -11000
rect -9600 -11320 -9599 -11000
rect -9921 -11321 -9599 -11320
rect -10340 -11388 -10244 -11372
rect -9328 -11372 -9312 -10948
rect -9248 -11372 -9232 -10948
rect -8316 -10948 -8220 -10932
rect -8909 -11000 -8587 -10999
rect -8909 -11320 -8908 -11000
rect -8588 -11320 -8587 -11000
rect -8909 -11321 -8587 -11320
rect -9328 -11388 -9232 -11372
rect -8316 -11372 -8300 -10948
rect -8236 -11372 -8220 -10948
rect -7304 -10948 -7208 -10932
rect -7897 -11000 -7575 -10999
rect -7897 -11320 -7896 -11000
rect -7576 -11320 -7575 -11000
rect -7897 -11321 -7575 -11320
rect -8316 -11388 -8220 -11372
rect -7304 -11372 -7288 -10948
rect -7224 -11372 -7208 -10948
rect -6292 -10948 -6196 -10932
rect -6885 -11000 -6563 -10999
rect -6885 -11320 -6884 -11000
rect -6564 -11320 -6563 -11000
rect -6885 -11321 -6563 -11320
rect -7304 -11388 -7208 -11372
rect -6292 -11372 -6276 -10948
rect -6212 -11372 -6196 -10948
rect -5280 -10948 -5184 -10932
rect -5873 -11000 -5551 -10999
rect -5873 -11320 -5872 -11000
rect -5552 -11320 -5551 -11000
rect -5873 -11321 -5551 -11320
rect -6292 -11388 -6196 -11372
rect -5280 -11372 -5264 -10948
rect -5200 -11372 -5184 -10948
rect -4268 -10948 -4172 -10932
rect -4861 -11000 -4539 -10999
rect -4861 -11320 -4860 -11000
rect -4540 -11320 -4539 -11000
rect -4861 -11321 -4539 -11320
rect -5280 -11388 -5184 -11372
rect -4268 -11372 -4252 -10948
rect -4188 -11372 -4172 -10948
rect -3256 -10948 -3160 -10932
rect -3849 -11000 -3527 -10999
rect -3849 -11320 -3848 -11000
rect -3528 -11320 -3527 -11000
rect -3849 -11321 -3527 -11320
rect -4268 -11388 -4172 -11372
rect -3256 -11372 -3240 -10948
rect -3176 -11372 -3160 -10948
rect -2244 -10948 -2148 -10932
rect -2837 -11000 -2515 -10999
rect -2837 -11320 -2836 -11000
rect -2516 -11320 -2515 -11000
rect -2837 -11321 -2515 -11320
rect -3256 -11388 -3160 -11372
rect -2244 -11372 -2228 -10948
rect -2164 -11372 -2148 -10948
rect -1232 -10948 -1136 -10932
rect -1825 -11000 -1503 -10999
rect -1825 -11320 -1824 -11000
rect -1504 -11320 -1503 -11000
rect -1825 -11321 -1503 -11320
rect -2244 -11388 -2148 -11372
rect -1232 -11372 -1216 -10948
rect -1152 -11372 -1136 -10948
rect -220 -10948 -124 -10932
rect -813 -11000 -491 -10999
rect -813 -11320 -812 -11000
rect -492 -11320 -491 -11000
rect -813 -11321 -491 -11320
rect -1232 -11388 -1136 -11372
rect -220 -11372 -204 -10948
rect -140 -11372 -124 -10948
rect 792 -10948 888 -10932
rect 199 -11000 521 -10999
rect 199 -11320 200 -11000
rect 520 -11320 521 -11000
rect 199 -11321 521 -11320
rect -220 -11388 -124 -11372
rect 792 -11372 808 -10948
rect 872 -11372 888 -10948
rect 1804 -10948 1900 -10932
rect 1211 -11000 1533 -10999
rect 1211 -11320 1212 -11000
rect 1532 -11320 1533 -11000
rect 1211 -11321 1533 -11320
rect 792 -11388 888 -11372
rect 1804 -11372 1820 -10948
rect 1884 -11372 1900 -10948
rect 2816 -10948 2912 -10932
rect 2223 -11000 2545 -10999
rect 2223 -11320 2224 -11000
rect 2544 -11320 2545 -11000
rect 2223 -11321 2545 -11320
rect 1804 -11388 1900 -11372
rect 2816 -11372 2832 -10948
rect 2896 -11372 2912 -10948
rect 3828 -10948 3924 -10932
rect 3235 -11000 3557 -10999
rect 3235 -11320 3236 -11000
rect 3556 -11320 3557 -11000
rect 3235 -11321 3557 -11320
rect 2816 -11388 2912 -11372
rect 3828 -11372 3844 -10948
rect 3908 -11372 3924 -10948
rect 4840 -10948 4936 -10932
rect 4247 -11000 4569 -10999
rect 4247 -11320 4248 -11000
rect 4568 -11320 4569 -11000
rect 4247 -11321 4569 -11320
rect 3828 -11388 3924 -11372
rect 4840 -11372 4856 -10948
rect 4920 -11372 4936 -10948
rect 5852 -10948 5948 -10932
rect 5259 -11000 5581 -10999
rect 5259 -11320 5260 -11000
rect 5580 -11320 5581 -11000
rect 5259 -11321 5581 -11320
rect 4840 -11388 4936 -11372
rect 5852 -11372 5868 -10948
rect 5932 -11372 5948 -10948
rect 6864 -10948 6960 -10932
rect 6271 -11000 6593 -10999
rect 6271 -11320 6272 -11000
rect 6592 -11320 6593 -11000
rect 6271 -11321 6593 -11320
rect 5852 -11388 5948 -11372
rect 6864 -11372 6880 -10948
rect 6944 -11372 6960 -10948
rect 7876 -10948 7972 -10932
rect 7283 -11000 7605 -10999
rect 7283 -11320 7284 -11000
rect 7604 -11320 7605 -11000
rect 7283 -11321 7605 -11320
rect 6864 -11388 6960 -11372
rect 7876 -11372 7892 -10948
rect 7956 -11372 7972 -10948
rect 8888 -10948 8984 -10932
rect 8295 -11000 8617 -10999
rect 8295 -11320 8296 -11000
rect 8616 -11320 8617 -11000
rect 8295 -11321 8617 -11320
rect 7876 -11388 7972 -11372
rect 8888 -11372 8904 -10948
rect 8968 -11372 8984 -10948
rect 9900 -10948 9996 -10932
rect 9307 -11000 9629 -10999
rect 9307 -11320 9308 -11000
rect 9628 -11320 9629 -11000
rect 9307 -11321 9629 -11320
rect 8888 -11388 8984 -11372
rect 9900 -11372 9916 -10948
rect 9980 -11372 9996 -10948
rect 10912 -10948 11008 -10932
rect 10319 -11000 10641 -10999
rect 10319 -11320 10320 -11000
rect 10640 -11320 10641 -11000
rect 10319 -11321 10641 -11320
rect 9900 -11388 9996 -11372
rect 10912 -11372 10928 -10948
rect 10992 -11372 11008 -10948
rect 11924 -10948 12020 -10932
rect 11331 -11000 11653 -10999
rect 11331 -11320 11332 -11000
rect 11652 -11320 11653 -11000
rect 11331 -11321 11653 -11320
rect 10912 -11388 11008 -11372
rect 11924 -11372 11940 -10948
rect 12004 -11372 12020 -10948
rect 12936 -10948 13032 -10932
rect 12343 -11000 12665 -10999
rect 12343 -11320 12344 -11000
rect 12664 -11320 12665 -11000
rect 12343 -11321 12665 -11320
rect 11924 -11388 12020 -11372
rect 12936 -11372 12952 -10948
rect 13016 -11372 13032 -10948
rect 13948 -10948 14044 -10932
rect 13355 -11000 13677 -10999
rect 13355 -11320 13356 -11000
rect 13676 -11320 13677 -11000
rect 13355 -11321 13677 -11320
rect 12936 -11388 13032 -11372
rect 13948 -11372 13964 -10948
rect 14028 -11372 14044 -10948
rect 14960 -10948 15056 -10932
rect 14367 -11000 14689 -10999
rect 14367 -11320 14368 -11000
rect 14688 -11320 14689 -11000
rect 14367 -11321 14689 -11320
rect 13948 -11388 14044 -11372
rect 14960 -11372 14976 -10948
rect 15040 -11372 15056 -10948
rect 15972 -10948 16068 -10932
rect 15379 -11000 15701 -10999
rect 15379 -11320 15380 -11000
rect 15700 -11320 15701 -11000
rect 15379 -11321 15701 -11320
rect 14960 -11388 15056 -11372
rect 15972 -11372 15988 -10948
rect 16052 -11372 16068 -10948
rect 16984 -10948 17080 -10932
rect 16391 -11000 16713 -10999
rect 16391 -11320 16392 -11000
rect 16712 -11320 16713 -11000
rect 16391 -11321 16713 -11320
rect 15972 -11388 16068 -11372
rect 16984 -11372 17000 -10948
rect 17064 -11372 17080 -10948
rect 16984 -11388 17080 -11372
<< properties >>
string FIXED_BBOX 16312 10920 16792 11400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 34 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
