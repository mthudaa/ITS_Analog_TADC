magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -194 -398 194 364
<< pmos >>
rect -100 -336 100 264
<< pdiff >>
rect -158 219 -100 264
rect -158 185 -146 219
rect -112 185 -100 219
rect -158 151 -100 185
rect -158 117 -146 151
rect -112 117 -100 151
rect -158 83 -100 117
rect -158 49 -146 83
rect -112 49 -100 83
rect -158 15 -100 49
rect -158 -19 -146 15
rect -112 -19 -100 15
rect -158 -53 -100 -19
rect -158 -87 -146 -53
rect -112 -87 -100 -53
rect -158 -121 -100 -87
rect -158 -155 -146 -121
rect -112 -155 -100 -121
rect -158 -189 -100 -155
rect -158 -223 -146 -189
rect -112 -223 -100 -189
rect -158 -257 -100 -223
rect -158 -291 -146 -257
rect -112 -291 -100 -257
rect -158 -336 -100 -291
rect 100 219 158 264
rect 100 185 112 219
rect 146 185 158 219
rect 100 151 158 185
rect 100 117 112 151
rect 146 117 158 151
rect 100 83 158 117
rect 100 49 112 83
rect 146 49 158 83
rect 100 15 158 49
rect 100 -19 112 15
rect 146 -19 158 15
rect 100 -53 158 -19
rect 100 -87 112 -53
rect 146 -87 158 -53
rect 100 -121 158 -87
rect 100 -155 112 -121
rect 146 -155 158 -121
rect 100 -189 158 -155
rect 100 -223 112 -189
rect 146 -223 158 -189
rect 100 -257 158 -223
rect 100 -291 112 -257
rect 146 -291 158 -257
rect 100 -336 158 -291
<< pdiffc >>
rect -146 185 -112 219
rect -146 117 -112 151
rect -146 49 -112 83
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect -146 -155 -112 -121
rect -146 -223 -112 -189
rect -146 -291 -112 -257
rect 112 185 146 219
rect 112 117 146 151
rect 112 49 146 83
rect 112 -19 146 15
rect 112 -87 146 -53
rect 112 -155 146 -121
rect 112 -223 146 -189
rect 112 -291 146 -257
<< poly >>
rect -58 345 58 361
rect -58 328 -17 345
rect -100 311 -17 328
rect 17 328 58 345
rect 17 311 100 328
rect -100 264 100 311
rect -100 -362 100 -336
<< polycont >>
rect -17 311 17 345
<< locali >>
rect -58 311 -17 345
rect 17 311 58 345
rect -146 233 -112 268
rect -146 161 -112 185
rect -146 89 -112 117
rect -146 17 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -89
rect -146 -189 -112 -161
rect -146 -257 -112 -233
rect -146 -340 -112 -305
rect 112 233 146 268
rect 112 161 146 185
rect 112 89 146 117
rect 112 17 146 49
rect 112 -53 146 -19
rect 112 -121 146 -89
rect 112 -189 146 -161
rect 112 -257 146 -233
rect 112 -340 146 -305
<< viali >>
rect -17 311 17 345
rect -146 219 -112 233
rect -146 199 -112 219
rect -146 151 -112 161
rect -146 127 -112 151
rect -146 83 -112 89
rect -146 55 -112 83
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect -146 -155 -112 -127
rect -146 -161 -112 -155
rect -146 -223 -112 -199
rect -146 -233 -112 -223
rect -146 -291 -112 -271
rect -146 -305 -112 -291
rect 112 219 146 233
rect 112 199 146 219
rect 112 151 146 161
rect 112 127 146 151
rect 112 83 146 89
rect 112 55 146 83
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
rect 112 -155 146 -127
rect 112 -161 146 -155
rect 112 -223 146 -199
rect 112 -233 146 -223
rect 112 -291 146 -271
rect 112 -305 146 -291
<< metal1 >>
rect -54 345 54 351
rect -54 311 -17 345
rect 17 311 54 345
rect -54 305 54 311
rect -152 233 -106 264
rect -152 199 -146 233
rect -112 199 -106 233
rect -152 161 -106 199
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -199 -106 -161
rect -152 -233 -146 -199
rect -112 -233 -106 -199
rect -152 -271 -106 -233
rect -152 -305 -146 -271
rect -112 -305 -106 -271
rect -152 -336 -106 -305
rect 106 233 152 264
rect 106 199 112 233
rect 146 199 152 233
rect 106 161 152 199
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -199 152 -161
rect 106 -233 112 -199
rect 146 -233 152 -199
rect 106 -271 152 -233
rect 106 -305 112 -271
rect 146 -305 152 -271
rect 106 -336 152 -305
<< end >>
