* PEX produced on Tue Sep 16 01:43:30 AM CST 2025 using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from tt_um_tsar_adc.ext - technology: sky130A

.subckt tt_um_tsar_adc clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_out[0]
+ uio_out[1] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] VDPWR VGND
X0 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_8403_19478# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_13164_28398# sar9b_0._06_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4 VGND sar9b_0.net5 a_7914_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 VDPWR a_10098_19171# a_9900_19047# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X8 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDPWR a_4749_27652# sar9b_0.net58 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X13 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X14 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X15 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 a_7926_23234# sar9b_0.net62 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X19 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=31.32 ps=341.28 w=0.5 l=0.5
X20 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X22 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X23 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X24 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X26 a_5896_22188# a_4755_22138# a_5739_22488# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X27 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X28 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X30 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X31 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X33 a_40321_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X34 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X35 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X37 VGND a_13011_24802# single_9b_cdac_0.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X38 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B a_16970_11404# VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X39 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X40 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X41 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X43 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X44 a_12047_26517# a_11842_26426# a_11382_26138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X45 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X46 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X48 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X49 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 a_8438_18958# a_8303_18859# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X53 a_3855_25792# a_4125_25958# a_4083_25852# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.05565 ps=0.685 w=0.42 l=0.15
X54 VGND a_12870_22267# a_12828_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X55 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X56 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X57 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X58 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X59 VGND sar9b_0.net52 a_12246_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X60 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VGND sar9b_0.clknet_1_1__leaf_CLK a_2835_24136# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X62 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X63 VGND a_13011_23238# single_9b_cdac_1.CF[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X64 a_5182_22567# sar9b_0.net64 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X65 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X66 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X67 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X68 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X69 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=282.12262 ps=2.58843k w=0.42 l=1
X70 a_12047_22521# a_11658_22138# a_11382_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X71 a_5196_19448# sar9b_0.net16 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X72 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X73 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X75 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X77 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X78 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X80 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X81 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X82 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X83 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X84 sar9b_0.net34 a_10284_25707# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X85 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X86 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X87 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VGND sar9b_0.net47 a_7062_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VGND a_11915_28371# uo_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X92 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X93 a_7890_26108# a_8345_26455# a_8294_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X94 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X96 VDPWR sar9b_0.net59 a_2847_26141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X97 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X98 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X99 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X100 a_12828_22145# a_11658_22138# a_12618_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X101 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X102 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X103 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 a_2918_20140# a_2739_20140# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X105 a_7343_27849# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X106 VDPWR a_11178_24802# a_11430_24931# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X107 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X108 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X109 VDPWR a_4771_18260# sar9b_0.net56 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X110 a_6634_18206# sar9b_0.net73 a_7155_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X111 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X112 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X113 a_10895_22855# a_10690_22806# a_10230_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X114 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X115 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10254_2858# dw_12589_1395# dw_12589_1395# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X116 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X117 a_26951_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X118 VGND a_6880_26815# sar9b_0.net21 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X119 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X120 single_9b_cdac_0.SW[7] a_10859_26330# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X121 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X122 a_2706_26108# a_3161_26455# a_3110_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X124 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X125 a_6534_27123# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X126 a_7978_22202# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X127 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X130 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 a_11842_19766# a_11658_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X132 VDPWR sar9b_0.net17 a_2931_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X133 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X135 a_11436_17742# sar9b_0.net2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X136 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X137 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 a_7155_18146# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X140 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X141 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X142 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 uo_out[0] a_11915_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X145 VGND a_4044_24776# sar9b_0.net72 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X146 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X147 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X148 sar9b_0.net40 a_6444_19448# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X149 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X153 VDPWR a_13216_23805# sar9b_0.net32 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X154 single_9b_cdac_1.SW[6] a_13011_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X155 VGND a_9588_27045# a_9593_26914# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X156 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X159 VGND sar9b_0.net52 a_10710_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X161 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X162 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=486.22675 ps=3.99183k w=1 l=1
X165 sar9b_0.net1 a_6867_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X166 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X167 a_5962_24151# a_5753_24250# a_5298_24499# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X168 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X169 VDPWR a_6834_20780# a_6636_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X170 a_10098_19171# a_10548_19053# a_10500_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X171 a_3561_22527# a_3027_22138# a_3454_22567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X172 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X176 a_12618_18142# a_11842_18434# a_12182_18427# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X177 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X178 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X179 a_8006_17229# a_7743_16817# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X180 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[1] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X182 a_9414_23127# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X183 a_6444_21738# sar9b_0._02_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X187 a_7404_17715# sar9b_0.net1 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24915 pd=2.37 as=0.15198 ps=1.17 w=0.55 l=0.15
X188 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VDPWR sar9b_0.net58 a_5046_27230# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X190 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X191 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X192 a_11568_24809# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X193 a_7831_22521# a_7402_22441# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X194 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X196 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X197 a_4072_19474# sar9b_0.net46 a_3994_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.20165 pd=1.285 as=0.0888 ps=0.98 w=0.74 l=0.15
X198 VGND a_8166_27595# a_8124_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X199 a_8842_16874# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X200 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X201 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 single_9b_cdac_0.SW[3] a_12491_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X204 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X205 sar9b_0.net18 a_2508_27440# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X206 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X207 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=93.96 ps=773.28003 w=1.5 l=0.5
X208 VDPWR sar9b_0._10_ a_4496_20468# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 th_dif_sw_0.CK a_10227_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X212 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X214 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X215 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X216 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X219 a_5459_22165# a_4934_22432# a_5289_22527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X220 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X222 VDPWR a_10932_25713# a_10937_25582# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X224 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X225 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X226 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X227 a_5506_17478# a_5322_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X228 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 a_8124_27473# a_6954_27466# a_7914_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X231 VDPWR a_7590_24931# a_7540_25221# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X232 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X233 a_10830_19068# a_10548_19053# a_11191_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X234 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDPWR a_5235_27466# uo_out[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X236 VGND a_4210_22378# a_4168_22188# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X237 a_6038_20140# a_5126_20140# a_5931_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X238 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X239 VDPWR sar9b_0.net22 a_8691_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X240 a_4011_22488# a_3206_22432# a_3713_22522# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X241 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X242 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X243 VDPWR sar9b_0.net35 a_3946_26198# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X244 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VDPWR sar9b_0.net54 a_7926_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X246 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X251 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X252 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X255 a_10926_17021# a_10649_17131# a_11256_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X256 a_11915_27039# sar9b_0.net30 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X257 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X258 sar9b_0.net36 a_9996_16784# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X259 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X260 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X261 a_2508_20780# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X262 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X266 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X267 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X268 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X270 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X271 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X272 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X273 a_5481_20185# a_5126_20140# a_5374_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X274 a_11382_18146# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X275 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X276 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X277 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X278 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X280 a_13216_19809# a_12618_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X281 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X282 a_7542_27530# a_7478_27751# a_7464_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X283 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VGND sar9b_0.net45 a_12647_27128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X285 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X286 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X287 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X288 VDPWR a_11030_22954# a_10985_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X289 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X290 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X291 a_11256_16874# a_10858_17113# a_11178_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X292 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X294 VGND sar9b_0.net68 a_3073_24815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X295 a_5289_22527# a_4934_22432# a_5182_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X296 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X297 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X298 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X299 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X301 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X302 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X303 VGND a_13011_24570# single_9b_cdac_1.CF[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X304 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 a_8303_23853# a_8098_23762# a_7638_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X306 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X307 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X308 a_12618_26134# a_11658_26134# a_12182_26419# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X309 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X310 VDPWR a_6579_18832# sar9b_0.net46 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X311 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X312 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A a_50962_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X313 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X316 a_11842_23762# a_11658_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X317 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 a_7464_27530# a_7138_27758# a_7343_27849# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X319 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X320 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X321 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X322 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X323 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X324 VGND sar9b_0.clknet_1_0__leaf_CLK a_4947_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X325 a_12870_19603# a_12618_19474# a_13008_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X326 VDPWR sar9b_0.net59 a_9279_27227# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 single_9b_cdac_0.SW[2] a_13067_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X329 VGND sar9b_0.net63 a_4811_23656# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2695 pd=2.08 as=0.13062 ps=1.025 w=0.55 l=0.15
X330 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X331 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A a_59529_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X332 a_11178_16874# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X333 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X334 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X335 a_3073_24815# sar9b_0._14_ sar9b_0._16_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X336 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X337 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X338 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X339 VGND a_7890_26108# a_7692_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X340 a_9935_24187# a_9730_24138# a_9270_24566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X341 VDPWR a_8595_17910# single_9b_cdac_1.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X342 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X343 VGND a_11776_27801# sar9b_0.net25 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X344 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X345 VDPWR a_10506_24506# a_10758_24459# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X346 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X347 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X348 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X349 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X351 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X352 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X353 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X354 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X355 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X356 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 a_21368_4076# th_dif_sw_0.th_sw_1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X358 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X359 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X360 a_9974_17626# a_9839_17527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X361 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X362 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X363 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X364 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X365 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X366 a_5151_28559# a_5010_28495# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X367 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X368 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X369 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X370 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X371 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X374 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X375 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X376 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDPWR tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X378 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 single_9b_cdac_1.SW[5] a_13011_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X380 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VGND a_7590_24931# a_7548_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X383 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X384 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X385 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X386 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X387 a_9634_17478# a_9450_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X388 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X391 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X392 VGND a_4811_23656# sar9b_0._13_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X393 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X394 a_12870_18271# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X396 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X397 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 a_9174_17906# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X400 VGND a_7347_24160# sar9b_0.net54 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X401 VDPWR a_12588_16784# sar9b_0.net2 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X402 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X403 a_16185_12837# tdc_0.phase_detector_0.pd_out_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X404 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X405 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X406 sar9b_0.net39 a_6540_22112# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X407 VGND a_12870_19603# a_12828_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X408 a_3454_22567# sar9b_0.net67 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X409 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X410 a_5832_27170# a_5506_26802# a_5711_26851# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X411 a_11466_23174# a_10690_22806# a_11030_22954# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X412 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X413 VGND a_8691_28566# uo_out[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X414 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X415 sar9b_0.clk_div_0.COUNT\[0\] a_5938_22378# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X416 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X419 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X420 VDPWR sar9b_0.net7 a_11658_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X421 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X424 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X425 a_11214_25728# a_10937_25582# a_11544_25838# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X426 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X429 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X430 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X433 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X434 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X435 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X436 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X437 a_9942_27470# sar9b_0.net43 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X438 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X440 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X441 a_11146_25483# a_10932_25713# a_10482_25831# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X442 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X445 a_12828_19481# a_11658_19474# a_12618_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X446 a_10926_17021# a_10644_16791# a_11287_17193# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X447 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X448 VGND sar9b_0.net59 a_8118_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X449 VDPWR a_10035_19474# sar9b_0.net48 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X451 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 a_10932_25713# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X453 a_6922_23534# sar9b_0.net10 a_7443_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X454 VGND sar9b_0.net43 a_11859_20574# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X455 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X456 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X457 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[2] a_55773_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X458 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X459 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X460 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VDPWR single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X462 a_11008_17491# a_10410_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X463 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X464 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X465 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X466 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X467 VGND a_5633_20244# a_5651_20547# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X468 a_64331_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X469 a_4330_27170# a_3545_26914# a_3822_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X470 VDPWR a_6880_26815# sar9b_0.net21 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X471 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X472 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X474 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X475 a_10690_22806# a_10506_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X476 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 sar9b_0.net44 a_6307_27584# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X478 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X479 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X480 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X481 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X482 VDPWR a_9974_17626# a_9929_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X483 VDPWR a_10742_27751# a_10697_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X484 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X485 VDPWR a_7890_26108# a_7692_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X486 VDPWR sar9b_0._07_ a_5628_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X487 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDPWR clk a_4332_23043# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X489 a_11382_22142# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X490 a_10607_21189# a_10402_21098# a_9942_20810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X491 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X492 a_13216_23805# a_12618_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X493 a_11287_17193# a_10858_17113# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X494 VDPWR sar9b_0.net44 a_6954_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X495 VDPWR a_5633_20244# a_5588_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X496 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 a_10098_19171# a_10553_18922# a_10502_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X498 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X499 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X500 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X502 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X503 VGND a_8595_17910# single_9b_cdac_1.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X504 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X505 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X507 a_4293_25852# a_4136_25584# a_3855_25792# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1181 ps=1.035 w=0.55 l=0.15
X508 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X509 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X510 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 a_9929_17527# a_9450_17846# a_9839_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X512 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] a_46159_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X515 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X516 VGND sar9b_0.net46 a_7830_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X517 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VDPWR sar9b_0.cyclic_flag_0.FINAL a_8883_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X519 a_10697_27849# a_10218_27466# a_10607_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X520 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X521 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X522 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X523 single_9b_cdac_1.SW[3] a_10803_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X524 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X525 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X526 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X527 a_7978_22202# a_7193_22459# a_7470_22349# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X528 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X531 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 a_9802_26815# a_9593_26914# a_9138_27163# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X533 a_7638_23474# sar9b_0.net11 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X534 a_9472_23805# a_8874_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X535 a_5588_20145# a_4947_20140# a_5481_20185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X536 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X537 a_11380_27885# a_10402_27758# a_11178_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X538 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X539 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X540 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X541 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X542 a_8842_16874# a_8057_17131# a_8334_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X543 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X544 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VGND sar9b_0.net21 a_7539_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X548 VGND a_10528_20155# sar9b_0.net38 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X549 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X550 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X551 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X552 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X553 single_9b_cdac_1.CF[7] a_12435_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X554 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X555 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X557 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X558 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X559 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 a_2940_25096# a_2893_24992# sar9b_0._16_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X561 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X562 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X563 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X564 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X565 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X567 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X568 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X571 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X573 VDPWR single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X574 VDPWR a_4811_23656# sar9b_0._13_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.3346 pd=1.76 as=0.3304 ps=2.83 w=1.12 l=0.15
X575 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X576 VGND a_5196_24776# sar9b_0.net68 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X577 VDPWR a_13011_16810# single_9b_cdac_1.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X578 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X579 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 single_9b_cdac_0.SW[8] a_9323_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X581 sar9b_0.net39 a_6540_22112# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X582 VDPWR sar9b_0.net47 a_6879_22145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X583 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X584 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X586 VDPWR a_10859_26330# single_9b_cdac_0.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X587 a_3180_19448# sar9b_0._09_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X588 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X589 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X590 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X591 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X592 a_8874_23470# a_7914_23470# a_8438_23755# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X593 a_3725_23194# a_3695_23038# a_3647_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X594 a_3273_20185# a_2739_20140# a_3166_20145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X595 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X598 VDPWR a_6534_27123# a_6484_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X599 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X600 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X601 VDPWR a_10182_20463# a_10132_20155# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X602 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X603 VGND a_3819_24136# a_4018_24235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X604 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X606 VDPWR a_8691_28566# uo_out[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X607 a_6738_22112# a_7193_22459# a_7142_22557# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X608 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X609 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A a_45123_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X610 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X611 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X612 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X614 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X615 VGND a_13011_24570# single_9b_cdac_1.CF[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X616 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X618 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X619 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 a_4236_21738# sar9b_0._05_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X621 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X622 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X623 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X624 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X626 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X627 a_11160_19178# a_10762_18823# a_11082_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X628 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X630 a_3539_24543# a_3014_24136# a_3369_24181# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X631 VDPWR sar9b_0.net10 a_11658_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X632 a_10218_21842# a_9258_21842# a_9782_21622# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X633 single_9b_cdac_1.CF[3] a_13011_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X634 a_8303_18859# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X635 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X637 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VDPWR a_12618_18142# a_12870_18271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X639 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X640 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X641 VDPWR a_12435_20806# single_9b_cdac_1.CF[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X642 VDPWR a_9126_23599# a_9076_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X643 single_9b_cdac_0.SW[1] a_13011_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X644 single_9b_cdac_1.SW[7] a_13011_19242# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X645 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X646 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X647 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X649 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X650 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 sar9b_0.net11 a_5484_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X652 sar9b_0._08_ a_4072_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.20905 ps=1.305 w=0.74 l=0.15
X653 a_6484_17491# a_5506_17478# a_6282_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X654 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X655 VGND a_13011_21906# single_9b_cdac_1.CF[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X656 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X657 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X658 a_11776_25137# a_11178_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X659 VDPWR a_9414_23127# a_9364_22819# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X660 sar9b_0.net35 a_7404_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X661 a_8013_23234# sar9b_0.net62 a_7926_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X662 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X663 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X664 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 a_11082_19178# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X666 a_10662_17799# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X667 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X668 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 a_9366_27227# a_9138_27163# a_9279_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X670 a_7284_20787# sar9b_0.net56 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X671 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X673 a_11842_22430# a_11658_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 VDPWR sar9b_0._07_ a_3795_19512# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2478 ps=2.27 w=0.84 l=0.15
X676 a_10194_16784# a_10649_17131# a_10598_17229# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X677 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X678 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X680 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X681 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X682 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X684 VDPWR a_3822_27060# a_3754_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X685 a_11722_25838# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X686 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X687 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X688 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X689 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X690 VGND sar9b_0.net20 a_8115_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X691 a_13008_23477# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X692 VGND a_10470_21795# a_10428_21899# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X693 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 uo_out[6] a_8115_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X695 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X696 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X697 single_9b_cdac_0.SW[0] a_13011_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X698 uo_out[7] a_5235_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X699 a_9138_27163# a_9588_27045# a_9540_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X700 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X701 VGND sar9b_0.clk_div_0.COUNT\[1\] a_3219_22860# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11312 pd=1.065 as=0.15675 ps=1.67 w=0.55 l=0.15
X702 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X703 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X704 VGND sar9b_0.net51 a_9363_20826# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X705 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X708 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X709 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X711 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X712 VGND sar9b_0.net66 sar9b_0._05_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X713 VDPWR sar9b_0.net8 a_8970_20510# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X714 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X716 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X717 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X718 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X719 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X721 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A a_41357_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X722 uio_out[1] a_2931_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X723 a_6744_23238# a_6484_22845# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X724 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X726 VDPWR single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X727 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X728 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VDPWR single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X730 a_10428_21899# a_9258_21842# a_10218_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X731 a_9323_27662# sar9b_0.net34 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X732 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X733 a_8512_27801# a_7914_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X734 VDPWR sar9b_0.net45 a_10218_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X735 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X736 VDPWR sar9b_0.net47 a_7374_19685# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X737 a_8006_18561# a_7743_18149# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X738 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X739 a_10070_24286# a_9935_24187# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X740 a_2892_23070# sar9b_0._18_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X741 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X743 a_5289_22527# a_4755_22138# a_5182_22567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X744 a_4496_20468# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X745 VDPWR a_3156_27447# a_3161_27787# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X746 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X747 a_2892_23070# sar9b_0._18_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X748 VGND a_5394_18116# a_5196_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X749 VDPWR sar9b_0.net49 a_10227_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X750 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X751 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X752 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X753 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X754 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X755 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X756 a_6538_24506# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X757 a_9494_20290# a_9359_20191# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X758 VGND sar9b_0.net48 a_8502_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X759 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X760 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 a_12243_25898# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X763 VDPWR a_3438_27677# a_3370_27769# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X764 sar9b_0.net45 a_8883_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X765 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X767 a_5046_17906# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X768 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X769 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 a_5506_26802# a_5322_27170# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X771 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X773 a_12182_18427# a_12047_18525# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X774 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X777 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X780 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X783 VGND sar9b_0.net37 a_8019_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X784 single_9b_cdac_1.SW[0] a_8595_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X785 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X786 VDPWR sar9b_0.net60 a_6678_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X787 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X788 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X789 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 VDPWR a_13011_20806# single_9b_cdac_1.CF[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X791 single_9b_cdac_1.SW[8] a_11859_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X792 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X793 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X794 a_15265_9613# th_dif_sw_0.VCP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X795 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X797 VDPWR a_12870_26263# a_12820_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X798 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X799 a_8502_19178# a_8438_18958# a_8424_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X800 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X801 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X802 tdc_0.phase_detector_0.INN a_16527_10454# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X803 VDPWR sar9b_0.net58 a_3438_27677# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X804 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X805 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X806 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X807 a_5414_28147# a_5151_28559# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X808 a_10816_21487# a_10218_21842# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X809 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X810 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X811 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X814 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X816 VDPWR a_3372_25734# sar9b_0.net69 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X817 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X819 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X820 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X822 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X823 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X824 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X826 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X827 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X828 a_7138_27758# a_6954_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X829 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X830 single_9b_cdac_0.SW[7] a_10859_26330# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X831 single_9b_cdac_0.SW[6] a_9323_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X832 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X833 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X834 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X835 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X836 a_8386_22806# a_8202_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X837 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X838 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X839 a_8424_19178# a_8098_18810# a_8303_18859# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X841 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X842 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X843 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X844 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X845 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X846 VGND a_11859_20574# single_9b_cdac_1.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X847 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X849 VDPWR tdc_0.OUTP tdc_0.OUTN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X850 uo_out[4] a_8691_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X851 VDPWR a_13011_24570# single_9b_cdac_1.CF[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X852 VDPWR sar9b_0.net47 a_6783_19481# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X853 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X854 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X855 sar9b_0._07_ a_3371_23106# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.4816 pd=3.1 as=0.203 ps=1.505 w=1.12 l=0.15
X856 single_9b_cdac_1.CF[5] a_13011_23238# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X857 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X858 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X859 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X860 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X861 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 a_5846_22572# a_4934_22432# a_5739_22488# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X863 a_12047_18525# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X864 tdc_0.OUTN tdc_0.phase_detector_0.pd_out_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X865 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X867 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X868 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X869 a_6052_19792# sar9b_0._07_ a_5581_19664# VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X870 a_21368_4076# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_18214_3039# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X871 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X872 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X874 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X875 a_8842_18206# sar9b_0.net5 a_9363_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X876 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X877 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X878 a_6642_19448# a_7097_19795# a_7046_19893# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X879 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X880 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X881 a_4330_27170# a_3540_27045# a_3822_27060# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X882 a_5002_23764# sar9b_0.net72 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.3346 ps=1.76 w=0.84 l=0.15
X883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X884 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X885 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X886 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 a_7343_27849# a_6954_27466# a_6678_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X888 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X889 a_5801_17527# a_5322_17846# a_5711_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X890 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X891 sar9b_0.net48 a_10035_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X892 VDPWR sar9b_0.net48 a_6126_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X893 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X896 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X897 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X898 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X899 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X900 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X901 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X902 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X903 VDPWR a_5394_18116# a_5196_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X904 a_21368_4076# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X905 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X906 VDPWR a_5580_24776# sar9b_0._03_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X907 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X908 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X909 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X910 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X912 a_5812_21028# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3685 pd=2.44 as=0.17462 ps=1.185 w=0.55 l=0.15
X913 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X914 a_3994_19474# sar9b_0._07_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.14457 ps=1.15 w=0.74 l=0.15
X915 a_11214_25728# a_10932_25713# a_11575_25519# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X916 a_9363_18146# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X918 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X919 uo_out[7] a_5235_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X920 VGND sar9b_0.net59 a_9366_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X921 a_9782_21622# a_9647_21523# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X922 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X924 sar9b_0._06_ a_12560_27128# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X925 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X926 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X927 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X928 VDPWR a_2603_17006# th_dif_sw_0.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X929 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X930 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X931 VGND sar9b_0.net52 a_8502_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X932 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X933 sar9b_0._15_ a_4467_24162# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X934 sar9b_0.net44 a_6307_27584# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X935 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X936 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X937 VDPWR tdc_0.phase_detector_0.pd_out_0.A a_16185_13034# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X938 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X939 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X940 VGND a_12491_27662# single_9b_cdac_0.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X941 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X942 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X943 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X944 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X945 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X946 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X947 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X948 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X949 a_11575_25519# a_11146_25483# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X950 a_12137_26517# a_11658_26134# a_12047_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X951 a_2508_23444# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X952 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X953 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 a_8502_23534# a_8438_23755# a_8424_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X955 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X956 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X957 a_9076_23889# a_8098_23762# a_8874_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X958 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X959 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X960 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X961 dw_17224_1400# a_18214_3039# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X962 VGND a_13011_21906# single_9b_cdac_1.CF[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X965 a_5711_26851# a_5322_27170# a_5046_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X966 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X967 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X968 a_12182_22423# a_12047_22521# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X969 a_6252_20780# sar9b_0._11_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X970 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X971 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 VGND sar9b_0.net12 a_12435_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X973 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X974 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X975 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X976 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X977 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X979 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X980 a_7590_24931# a_7338_24802# a_7728_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X981 a_6252_20780# sar9b_0._11_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X983 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X984 a_10598_17229# a_10335_16817# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X985 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X986 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X987 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X988 a_8424_23534# a_8098_23762# a_8303_23853# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X989 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X990 a_10623_25895# a_10482_25831# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 a_9552_23231# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X993 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X994 a_10985_22855# a_10506_23174# a_10895_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X995 a_6250_28502# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X996 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X997 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X999 VGND sar9b_0.net9 a_10506_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1000 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1001 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1002 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1003 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1004 VDPWR a_9930_20510# a_10182_20463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1005 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1006 VDPWR a_6282_27170# a_6534_27123# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1007 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1008 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1009 VDPWR sar9b_0.net61 a_7978_22202# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1010 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1011 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1012 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1013 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1014 a_5628_19768# a_5581_19664# sar9b_0._10_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X1015 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1016 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1017 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1018 sar9b_0._18_ sar9b_0._17_ a_5183_20819# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1019 a_9138_27163# a_9593_26914# a_9542_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X1020 VGND a_8622_26345# a_8554_26437# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1021 single_9b_cdac_1.SW[4] a_11859_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1022 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1023 a_9935_24187# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1024 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1025 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1026 a_11842_19766# a_11658_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1027 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1028 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1029 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1030 a_12047_22521# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1031 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1033 sar9b_0.net49 a_9363_20826# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X1034 sar9b_0.net6 a_7404_18116# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1035 th_dif_sw_0.VCN ua[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1036 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1037 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1039 a_11030_22954# a_10895_22855# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1040 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1041 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1043 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1044 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1045 a_7540_25221# a_6562_25094# a_7338_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1046 a_5183_20819# sar9b_0.net65 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X1047 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1048 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 a_10742_27751# a_10607_27849# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1050 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1051 a_5581_20992# a_5812_21028# a_5761_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1052 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1055 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1056 VDPWR a_12064_22819# sar9b_0.net30 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1057 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1058 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1060 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1061 a_7402_22441# a_7188_22119# a_6738_22112# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1062 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1063 VGND a_11915_27039# single_9b_cdac_0.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X1064 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1065 VDPWR a_9162_23174# a_9414_23127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1066 sar9b_0._12_ a_5523_21528# a_5765_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3182 pd=2.34 as=0.0888 ps=0.98 w=0.74 l=0.15
X1067 VGND a_12588_16784# sar9b_0.net2 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X1068 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1069 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1070 sar9b_0.net48 a_10035_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1071 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1072 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1074 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1075 a_6771_28562# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1076 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15182 ps=1.125 w=0.55 l=0.15
X1077 VDPWR sar9b_0.net12 a_12435_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1078 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1079 VDPWR sar9b_0.net61 a_8842_16874# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1080 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1081 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1082 VDPWR a_12491_27662# single_9b_cdac_0.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1083 a_3819_24136# a_3014_24136# a_3521_24240# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X1084 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1085 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1086 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1087 VGND a_9323_27662# single_9b_cdac_0.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X1088 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1089 VDPWR sar9b_0.clk_div_0.COUNT\[1\] sar9b_0._17_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3304 ps=2.83 w=1.12 l=0.15
X1090 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1091 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 VDPWR a_10227_18142# th_dif_sw_0.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1093 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1094 a_8622_26345# a_8340_26115# a_8983_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X1095 VDPWR a_4365_25770# a_4293_25852# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.2331 ps=1.395 w=0.84 l=0.15
X1096 VGND sar9b_0.net26 a_13011_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1097 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1098 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1099 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1100 a_3262_24141# sar9b_0.net70 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X1101 a_5765_21842# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.22412 ps=1.365 w=0.74 l=0.15
X1102 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1103 a_7566_21017# a_7284_20787# a_7927_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X1104 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1105 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1106 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1108 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1109 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1110 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1111 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1112 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1113 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1114 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1115 a_6102_24806# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1116 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1117 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1118 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1119 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1120 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1121 VGND sar9b_0.net10 a_13011_23238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1122 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1123 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1124 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1125 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1126 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1127 a_11338_19178# a_10553_18922# a_10830_19068# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1128 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1129 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1130 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1131 VDPWR a_10528_20155# sar9b_0.net38 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1132 a_5443_19074# sar9b_0.net4 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1133 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1134 uo_out[7] a_5235_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1135 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1136 VDPWR a_2706_27440# a_2508_27440# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1137 VGND a_11339_27039# single_9b_cdac_0.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1138 VDPWR a_10662_17799# a_10612_17491# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1139 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1140 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1141 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1142 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1143 a_8781_20570# sar9b_0.net61 a_8694_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1144 a_8266_17113# a_8052_16791# a_7602_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1145 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1146 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1147 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1148 VDPWR a_13216_18477# sar9b_0.net28 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1149 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1150 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1151 a_9846_21842# a_9782_21622# a_9768_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1152 a_7927_21189# a_7498_21109# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X1153 VDPWR a_11430_20935# a_11380_21225# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1154 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1155 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1156 VGND single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1157 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1158 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A a_65367_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1159 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1160 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1161 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1162 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1163 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1164 VDPWR single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1165 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1166 VDPWR sar9b_0.clknet_0_CLK a_2508_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1167 a_4934_22432# a_4755_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X1168 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1169 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1170 a_10859_26330# sar9b_0.net33 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X1171 VDPWR a_8438_23755# a_8393_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1172 a_4583_20468# sar9b_0.net60 a_4496_20468# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X1173 a_7046_19893# a_6783_19481# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1175 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1176 a_11008_17491# a_10410_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1177 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1178 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1179 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1180 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1181 a_5962_24151# a_5748_24381# a_5298_24499# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1182 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1183 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1184 VDPWR sar9b_0.net50 a_11382_18146# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1185 a_9768_21842# a_9442_21474# a_9647_21523# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1186 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1187 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1188 a_5581_20992# sar9b_0._08_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.19322 ps=1.32 w=0.55 l=0.15
X1189 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1190 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1191 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1192 VGND sar9b_0.net54 a_6966_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1194 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1195 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1196 VGND sar9b_0.net10 a_11658_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1197 single_9b_cdac_1.CF[0] a_13011_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1198 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1199 a_3946_26198# sar9b_0.net35 a_4467_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1200 a_8393_23853# a_7914_23470# a_8303_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1201 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1202 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1203 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1204 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1205 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1206 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 VGND sar9b_0.net68 a_2893_24992# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X1208 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1209 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1210 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1211 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1212 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1213 single_9b_cdac_1.CF[2] a_11859_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1214 VGND sar9b_0.net50 a_11469_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1215 a_10378_27170# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X1216 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1217 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1218 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1219 VDPWR sar9b_0.net26 a_13011_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1220 a_11842_23762# a_11658_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1221 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1222 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1223 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1224 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1225 VDPWR a_13067_27662# single_9b_cdac_0.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1226 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1227 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y a_54737_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1228 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1229 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1230 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1231 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1232 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1234 a_4293_25852# a_4125_25958# a_3855_25792# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.1428 ps=1.225 w=0.84 l=0.15
X1235 single_9b_cdac_1.SW[0] a_8595_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1236 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1237 a_4467_26138# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1238 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1239 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1240 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1241 a_9540_27227# a_9279_27227# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1242 a_12182_22423# a_12047_22521# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1243 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1244 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1245 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1246 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1247 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1248 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1249 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1250 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1251 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1252 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1253 VDPWR a_7566_21017# a_7498_21109# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1254 a_11469_19478# sar9b_0.net73 a_11382_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1255 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1256 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1257 VDPWR a_10926_17021# a_10858_17113# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1258 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1259 VGND a_3603_28156# sar9b_0.net59 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1260 VDPWR a_9323_27662# single_9b_cdac_0.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1261 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1262 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1263 VDPWR sar9b_0.net58 a_5151_28559# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1264 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1266 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1267 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1268 a_10470_21795# a_10218_21842# a_10608_21899# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1269 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1270 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1271 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1272 VGND a_11915_27039# single_9b_cdac_0.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1273 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1274 a_3166_20145# sar9b_0._00_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X1275 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1276 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1277 a_9647_21523# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1278 VGND a_7374_19685# a_7306_19777# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1280 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1281 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1282 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1283 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1284 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1285 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1286 a_5046_27230# sar9b_0.net39 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1287 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1288 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1289 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1290 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[1] a_60565_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1291 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1292 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1293 a_10528_20155# a_9930_20510# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1294 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1295 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1296 single_9b_cdac_1.SW[1] a_10803_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1297 VDPWR sar9b_0.net48 a_9174_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1298 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1299 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1300 VGND a_10098_19171# a_9900_19047# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1301 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1302 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1303 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1304 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1305 a_5238_28559# a_5010_28495# a_5151_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1306 VGND a_9323_27662# single_9b_cdac_0.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1307 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1308 a_9942_20810# sar9b_0.net7 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1309 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1310 a_50962_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1311 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1312 VGND a_13011_19242# single_9b_cdac_1.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1313 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1314 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1315 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1316 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1317 sar9b_0.net47 a_7443_21496# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X1318 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A a_36555_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1319 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1320 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1321 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1322 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1323 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1324 VDPWR single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1325 a_35519_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1326 a_11842_18434# a_11658_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1328 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1329 VDPWR single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1330 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1331 VDPWR a_5196_24776# sar9b_0.net68 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1332 VGND sar9b_0.clknet_0_CLK a_2508_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X1333 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1334 VDPWR a_6642_19448# a_6444_19448# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1335 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1336 a_7092_19455# sar9b_0.net10 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1337 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1338 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1339 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1340 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1341 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1342 VGND a_3438_27677# a_3370_27769# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1343 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1344 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1345 single_9b_cdac_0.SW[4] a_11915_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X1346 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1347 VDPWR sar9b_0.net72 sar9b_0._14_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1348 a_6534_17799# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1349 a_8074_20870# a_7289_21127# a_7566_21017# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1350 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VDPWR a_10482_3438# VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X1351 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1352 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1353 VDPWR a_13216_22473# sar9b_0.net31 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1354 VDPWR a_10742_21091# a_10697_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1355 a_11434_16874# a_10649_17131# a_10926_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1356 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1357 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1358 VGND sar9b_0.net44 a_6954_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1359 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1360 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1361 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1362 a_5481_20185# a_4947_20140# a_5374_20145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X1363 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1364 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1365 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1366 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1367 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1368 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1369 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1370 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1371 uio_out[0] a_4083_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1372 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1373 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1374 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1375 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1376 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1377 VDPWR a_11776_25137# sar9b_0.net13 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1378 a_8303_18859# a_7914_19178# a_7638_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1379 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1380 VGND sar9b_0._04_ a_3027_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1381 a_4811_23656# sar9b_0.net63 a_5002_23764# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1134 ps=1.11 w=0.84 l=0.15
X1382 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1383 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1384 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1385 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1387 a_3425_20244# a_3273_20185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X1388 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1389 VDPWR a_6307_27584# sar9b_0.net44 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1390 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1391 a_12820_23889# a_11842_23762# a_12618_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1392 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1393 a_6444_21738# sar9b_0._02_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1394 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1396 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1397 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1398 a_16555_12124# tdc_0.OUTN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1399 VGND sar9b_0.net17 a_2931_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1400 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1401 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1402 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1403 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1404 a_3156_27447# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1405 a_4332_23043# clk VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1406 VDPWR sar9b_0.net53 a_11382_22142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1407 a_10697_21189# a_10218_20806# a_10607_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1408 VGND a_10803_19474# single_9b_cdac_1.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1409 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1410 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1411 uio_out[1] a_2931_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1412 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1413 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1414 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1415 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1416 a_7138_27758# a_6954_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1418 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1419 sar9b_0.net56 a_4771_18260# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X1420 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1421 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1422 sar9b_0.net17 a_2508_26108# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1423 a_3822_27060# a_3545_26914# a_4152_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X1424 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1425 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1426 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1427 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1428 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1429 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1430 VDPWR th_dif_sw_0.th_sw_1.CKB a_18214_3039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X1431 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1432 a_9760_22819# a_9162_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1433 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1434 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1435 sar9b_0.net51 a_5811_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2051 ps=1.52 w=1.12 l=0.15
X1436 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1437 VGND sar9b_0.net46 a_7830_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1438 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1439 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1440 VGND single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1441 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1442 VGND sar9b_0.net53 a_11469_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1443 a_10132_20155# a_9154_20142# a_9930_20510# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1444 VGND a_6126_18353# a_6058_18445# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1445 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1446 VGND a_4011_22488# a_4210_22378# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X1447 a_4812_21738# sar9b_0.clk_div_0.COUNT\[3\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1448 th_dif_sw_0.VCN th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCN VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X1449 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1450 VDPWR sar9b_0.net52 a_7638_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1451 sar9b_0._05_ sar9b_0.net66 a_2828_22432# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X1452 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1453 VGND sar9b_0.net58 a_2934_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1454 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1455 a_7142_22557# a_6879_22145# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1456 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1457 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1458 a_9279_27227# a_9138_27163# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X1459 a_4152_27170# a_3754_26815# a_4074_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1460 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1461 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1462 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1463 a_3747_25724# a_3855_25792# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1229 ps=1.085 w=0.64 l=0.15
X1464 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 a_21368_4076# th_dif_sw_0.th_sw_1.CKB a_18214_3039# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X1466 VDPWR a_12435_24802# single_9b_cdac_1.CF[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1467 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1468 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1469 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] a_31753_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1470 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1471 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1472 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1474 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1475 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1476 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1477 single_9b_cdac_1.SW[6] a_13011_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1478 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1479 a_11469_23474# sar9b_0.net74 a_11382_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1480 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1481 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1483 VDPWR a_5010_28495# a_4812_28371# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1484 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1485 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1486 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11655 ps=1.055 w=0.74 l=0.15
X1487 a_5526_24563# a_5298_24499# a_5439_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1488 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1489 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1490 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1491 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1492 VDPWR a_9323_27662# single_9b_cdac_0.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1493 a_3443_20547# a_2918_20140# a_3273_20185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X1494 VDPWR a_8595_17910# single_9b_cdac_1.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1495 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1496 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1497 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1498 a_8074_20870# a_7284_20787# a_7566_21017# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1499 a_4074_27170# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X1500 a_10134_24506# a_10070_24286# a_10056_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1501 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1502 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1503 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1504 a_13216_18477# a_12618_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1505 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1506 sar9b_0._14_ sar9b_0.net72 a_2637_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1507 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1508 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1509 a_7478_27751# a_7343_27849# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1510 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1511 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1512 VDPWR a_5844_18123# a_5849_18463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1513 VGND sar9b_0.net22 a_8691_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1514 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1515 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1516 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1517 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1518 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1519 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1520 VDPWR a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
X1521 a_55773_15501# single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1522 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y a_49926_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1523 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1524 VDPWR clk a_15151_10456# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X1525 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1526 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1528 VGND a_9126_19131# a_9084_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1529 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1530 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1531 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1532 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1533 a_10056_24506# a_9730_24138# a_9935_24187# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1534 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1535 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1536 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1537 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1538 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1539 a_8303_23853# a_7914_23470# a_7638_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1540 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1541 a_11842_22430# a_11658_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1542 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1543 uo_out[5] a_7539_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1544 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1545 a_11338_19178# a_10548_19053# a_10830_19068# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1546 a_5506_17478# a_5322_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1547 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1549 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1550 VDPWR a_10803_19474# single_9b_cdac_1.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1551 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1552 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1553 VDPWR a_13011_19242# single_9b_cdac_1.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1554 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1555 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1556 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1557 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1558 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1559 single_9b_cdac_1.CF[8] a_13011_25902# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1560 VGND a_6744_23238# a_6861_22828# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11485 pd=1.085 as=0.2436 ps=2 w=0.42 l=0.18
X1561 VDPWR a_9472_18823# sar9b_0.net26 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1562 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1563 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1564 a_6346_23773# a_6132_23451# a_5682_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1565 VGND a_7470_22349# a_7402_22441# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1566 VDPWR a_11436_17742# sar9b_0.net61 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1567 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1568 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1570 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1571 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1572 a_3976_24520# a_2835_24136# a_3819_24136# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X1573 a_9084_19235# a_7914_19178# a_8874_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1574 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1575 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1576 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1577 a_5394_18116# a_5844_18123# a_5796_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X1578 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1579 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1580 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1581 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1582 VDPWR a_10410_17846# a_10662_17799# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1583 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1584 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1585 a_6250_28502# a_5460_28377# a_5742_28392# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1586 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1587 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1588 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1589 a_12618_26134# a_11842_26426# a_12182_26419# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1590 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1591 a_46159_15501# single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1592 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1593 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1594 a_9935_24187# a_9546_24506# a_9270_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1595 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1596 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1597 a_6767_25185# a_6562_25094# a_6102_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1598 VGND sar9b_0.net8 a_11658_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1599 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1600 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1601 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1602 uo_out[1] a_12531_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1603 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1604 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1605 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1606 a_13216_19809# a_12618_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1607 VGND sar9b_0.net35 a_8595_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1608 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1609 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1611 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1612 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1613 a_10420_21487# a_9442_21474# a_10218_21842# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1614 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1615 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1616 a_4211_19474# sar9b_0.net71 a_4072_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=1.55 as=0.20165 ps=1.285 w=0.74 l=0.15
X1617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1618 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1619 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1620 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1621 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1622 VDPWR a_8115_28566# uo_out[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1623 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1624 VDPWR a_13011_24802# single_9b_cdac_0.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1625 a_7188_22119# sar9b_0.net9 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1626 a_5796_18149# a_5535_18149# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1627 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1628 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1629 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.B a_16185_12837# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1630 a_6880_26815# a_6282_27170# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1631 VDPWR sar9b_0.net56 a_10218_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1632 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1633 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1634 a_11776_27801# a_11178_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1635 a_7882_19538# a_7092_19455# a_7374_19685# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1636 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1637 a_9154_20142# a_8970_20510# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1638 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1639 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1640 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1641 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1642 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1643 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1644 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1645 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1646 VGND a_8340_26115# a_8345_26455# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1647 sar9b_0.net57 a_5443_19074# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1648 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1649 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1650 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1651 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1652 a_12182_19759# a_12047_19857# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1653 VGND a_13011_19242# single_9b_cdac_1.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X1654 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1655 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1656 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1657 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1658 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1659 VDPWR clk a_4332_23043# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1660 VDPWR a_10830_19068# a_10762_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1661 VDPWR a_2931_28566# uio_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1662 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1663 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1664 a_4531_25875# a_4293_25852# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1648 ps=1.245 w=0.42 l=0.15
X1665 a_9839_17527# a_9634_17478# a_9174_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1666 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1667 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1668 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1669 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1670 VDPWR a_3540_27045# a_3545_26914# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1671 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1672 a_11178_24802# a_10218_24802# a_10742_25087# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1673 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1675 a_10402_27758# a_10218_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1676 a_11178_20806# a_10402_21098# a_10742_21091# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1677 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1678 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1679 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1680 a_10895_22855# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1681 VDPWR sar9b_0.net46 a_8334_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X1682 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1683 a_3156_27447# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1684 VDPWR a_7602_18116# a_7404_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1685 a_9126_23599# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1686 tdc_0.phase_detector_0.INP a_15151_10456# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X1687 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1688 VDPWR sar9b_0.net62 a_6538_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1689 a_7602_18116# a_8052_18123# a_8004_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X1690 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1691 a_3521_24240# a_3369_24181# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X1692 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1693 VDPWR a_8883_27466# sar9b_0.net45 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1694 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1695 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1696 single_9b_cdac_1.CF[4] a_13011_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1697 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1698 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1699 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1700 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1701 a_8554_26437# a_8345_26455# a_7890_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X1702 a_5580_24776# sar9b_0._15_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1703 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1704 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1705 VGND a_9939_28566# uo_out[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1706 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1707 VGND sar9b_0.clknet_0_CLK a_2508_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X1708 a_11434_16874# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X1709 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1710 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1711 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1712 a_5126_20140# a_4947_20140# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X1713 VGND a_5443_19074# sar9b_0.net57 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1714 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X1715 uo_out[6] a_8115_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1716 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1717 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1718 VDPWR a_3713_22522# a_3668_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X1719 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1720 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1721 a_11382_26138# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1722 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1723 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1724 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1725 a_6879_22145# a_6738_22112# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X1726 ua[3] th_dif_sw_0.th_sw_1.CK ua[3] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X1727 a_13008_18149# sar9b_0.net50 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1728 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1729 a_10402_21098# a_10218_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1730 VGND a_10803_19474# single_9b_cdac_1.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X1731 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1732 VGND sar9b_0.net11 a_13011_24570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1733 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1734 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1735 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1736 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1737 a_9634_17478# a_9450_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1738 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1739 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1740 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1741 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1742 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1743 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1744 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1745 a_8118_26141# a_7890_26108# a_8031_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1746 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1747 a_41357_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1748 VGND sar9b_0.net54 a_5526_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1749 VDPWR a_11430_27595# a_11380_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1750 VGND a_9472_23805# sar9b_0.net12 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1751 VDPWR a_10859_26330# single_9b_cdac_0.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1752 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1753 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1754 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1755 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1756 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1757 a_3668_22567# a_3027_22138# a_3561_22527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X1758 sar9b_0._04_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1759 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1760 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1761 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1762 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1763 VDPWR a_11859_17910# single_9b_cdac_1.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1764 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1765 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1766 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1767 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1768 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1769 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1770 a_9647_21523# a_9258_21842# a_8982_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1771 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1773 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1774 a_3713_22522# a_3561_22527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X1775 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1776 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1777 VDPWR a_8691_28566# uo_out[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1778 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1779 VDPWR sar9b_0.net47 a_6975_20813# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1780 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1781 uo_out[5] a_7539_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1782 VDPWR single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1783 VDPWR a_13011_23238# single_9b_cdac_1.CF[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1784 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1785 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1786 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1787 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1788 a_6252_19074# sar9b_0.net15 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1789 a_2828_22432# sar9b_0._12_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X1790 a_6634_18206# a_5844_18123# a_6126_18353# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1792 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1793 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1794 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1795 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1796 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1797 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1798 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1799 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1800 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1801 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1802 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1803 VDPWR a_13164_28398# sar9b_0.net14 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1804 single_9b_cdac_1.SW[2] a_8019_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1805 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1806 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1807 VGND sar9b_0.net53 a_11094_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1808 a_8842_16874# sar9b_0.net61 a_9363_16814# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1809 VDPWR single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1810 a_59529_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1812 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1813 VGND a_3372_25734# sar9b_0.net69 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X1814 VGND sar9b_0.net11 a_11658_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1815 VGND a_4083_28566# uio_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1816 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1817 VDPWR sar9b_0.clknet_1_1__leaf_CLK a_4755_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1819 a_3946_27530# sar9b_0.net36 a_4467_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1820 a_9323_27662# sar9b_0.net34 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X1821 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1822 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1823 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1824 a_13216_23805# a_12618_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1825 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1826 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1827 single_9b_cdac_0.SW[0] a_13011_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1828 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1829 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1830 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1831 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1832 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1833 a_13164_28398# sar9b_0._06_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1834 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1835 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1836 a_7936_25137# a_7338_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1837 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1838 a_12870_26263# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1839 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1840 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1841 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1842 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1843 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1844 a_11722_25838# a_10937_25582# a_11214_25728# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1845 a_11094_23174# a_11030_22954# a_11016_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1846 single_9b_cdac_1.CF[5] a_13011_23238# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1847 a_9363_16814# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1848 th_dif_sw_0.CKB a_2603_17006# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1849 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1850 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1851 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1852 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1853 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1854 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1856 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1857 a_4467_27470# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1858 a_8983_26517# a_8554_26437# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X1859 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1860 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1861 a_12182_23755# a_12047_23853# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1862 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1863 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1864 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1865 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1867 VDPWR sar9b_0.net12 a_11658_26134# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1868 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1869 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1870 a_10607_27849# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1871 VDPWR a_6534_17799# a_6484_17491# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1872 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1874 VDPWR a_5682_23444# a_5484_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1875 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1876 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1877 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1878 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1879 VDPWR sar9b_0.net59 a_9942_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1880 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1881 VDPWR a_3723_20140# a_3922_20239# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X1882 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1883 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1884 sar9b_0.net63 a_6861_22828# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.11485 ps=1.085 w=0.74 l=0.15
X1885 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1886 VDPWR sar9b_0.net36 a_10803_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1887 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1888 a_11030_22954# a_10895_22855# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1889 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1890 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1891 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1892 VGND sar9b_0.net58 a_3318_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1893 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1894 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1895 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1896 a_12064_22819# a_11466_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1897 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1898 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1899 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1900 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1901 a_9542_26815# a_9279_27227# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1902 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1903 a_5812_21028# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2898 ps=2.37 w=0.84 l=0.15
X1904 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1905 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1906 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1907 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[2] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1908 sar9b_0._11_ a_4496_20468# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X1909 VGND a_7092_19455# a_7097_19795# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1910 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1911 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1912 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1913 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1914 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1915 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1916 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1917 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1918 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1919 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1920 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1921 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1922 VGND a_11104_24151# sar9b_0.net42 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1923 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1924 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1925 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1926 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1927 sar9b_0.net34 a_10284_25707# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X1928 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1929 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1930 a_5910_23477# a_5682_23444# a_5823_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1931 a_13008_22145# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1932 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1933 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1935 VDPWR sar9b_0.net52 a_10623_25895# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1936 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1937 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1938 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1939 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1940 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1941 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1942 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1943 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1944 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1945 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1946 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1947 VDPWR sar9b_0.net18 a_4083_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1948 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1949 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1950 VDPWR sar9b_0.net61 a_11434_16874# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1952 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1953 VDPWR sar9b_0.net38 a_6250_28502# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1954 a_6966_24866# a_6902_25087# a_6888_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1955 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1956 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1957 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1958 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1959 VDPWR a_8340_26115# a_8345_26455# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1960 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1961 a_7236_20813# a_6975_20813# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1962 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1964 sar9b_0.net58 a_4749_27652# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1965 VDPWR a_11859_21906# single_9b_cdac_1.CF[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1966 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1967 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1968 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1969 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1970 VGND a_3156_27447# a_3161_27787# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1971 VGND tdc_0.RDY a_5331_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1972 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1973 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1974 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1975 VDPWR a_8622_26345# a_8554_26437# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1976 a_5711_26851# a_5506_26802# a_5046_27230# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1977 VDPWR a_11859_17910# single_9b_cdac_1.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1978 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1979 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1980 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1981 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1982 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1983 a_5133_27230# sar9b_0.net39 a_5046_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1984 a_10742_21091# a_10607_21189# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1985 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1986 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1987 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1988 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1989 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1990 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1991 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1992 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1993 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1994 VDPWR a_3156_26115# a_3161_26455# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1995 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1996 a_3723_20140# a_2918_20140# a_3425_20244# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X1997 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1998 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1999 a_6888_24866# a_6562_25094# a_6767_25185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2000 VDPWR a_9363_20826# sar9b_0.net49 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X2001 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2002 a_10482_25831# a_10932_25713# a_10884_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2003 single_9b_cdac_1.CF[7] a_12435_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2004 VGND sar9b_0.net50 a_12246_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2005 sar9b_0.net35 a_7404_16784# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2006 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2007 VDPWR a_3438_26345# a_3370_26437# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2008 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2009 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2010 VDPWR sar9b_0.net59 a_8622_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2011 a_4467_24162# sar9b_0._13_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X2012 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2013 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2014 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2015 a_5010_28495# a_5465_28246# a_5414_28147# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2016 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2017 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2018 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2019 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2020 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2021 sar9b_0.net53 a_10227_23490# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2022 a_3370_27769# a_3161_27787# a_2706_27440# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2023 VGND sar9b_0.net59 a_10806_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2024 a_5742_28392# a_5460_28377# a_6103_28183# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2025 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2026 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2027 a_9782_21622# a_9647_21523# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X2028 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2030 VGND a_12531_28566# uo_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2031 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2032 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2033 VDPWR sar9b_0.net59 a_3438_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2034 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2035 a_8591_22855# a_8386_22806# a_7926_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2036 single_9b_cdac_0.SW[3] a_12491_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2037 a_10884_25895# a_10623_25895# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2038 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2039 single_9b_cdac_0.SW[1] a_13011_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2040 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2041 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2042 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2043 VDPWR a_2706_26108# a_2508_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2044 a_5931_20140# a_4947_20140# a_5633_20244# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X2045 VDPWR sar9b_0.net41 a_13011_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2046 a_10422_16817# a_10194_16784# a_10335_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2047 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2048 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2049 VGND a_5739_22488# a_5938_22378# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X2050 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2051 a_9130_26198# a_8345_26455# a_8622_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X2052 VGND a_11859_21906# single_9b_cdac_1.CF[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2053 th_dif_sw_0.CK a_10227_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2055 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2056 th_dif_sw_0.CKB a_2603_17006# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2057 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2058 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2059 a_6103_28183# a_5674_28147# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2060 a_10806_27530# a_10742_27751# a_10728_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2061 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2062 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2063 VDPWR sar9b_0.net54 a_6102_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2064 VDPWR sar9b_0.net65 a_5083_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X2065 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2066 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2067 VDPWR sar9b_0.net47 a_6052_19792# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X2068 VDPWR a_12618_26134# a_12870_26263# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2069 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A a_54737_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2070 a_8304_27473# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2071 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2072 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2074 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2075 a_45123_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2076 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2077 VGND sar9b_0.net9 a_13011_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X2078 a_3180_19448# sar9b_0._09_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2079 VDPWR a_5196_19448# sar9b_0.net71 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2080 VGND a_10830_19068# a_10762_18823# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2081 VDPWR a_5235_27466# uo_out[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2082 a_7374_19685# a_7092_19455# a_7735_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2083 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2084 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2086 VGND a_10816_21487# sar9b_0.net9 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2087 a_9930_20510# a_9154_20142# a_9494_20290# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2088 a_5910_17846# a_5846_17626# a_5832_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2089 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2090 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2091 a_5374_20145# sar9b_0._01_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X2092 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2093 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2094 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2095 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2096 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2097 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2098 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2099 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[8] a_26951_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2100 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2101 a_10728_27530# a_10402_27758# a_10607_27849# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2102 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2103 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2104 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2105 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2106 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2107 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2108 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2109 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2110 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2111 a_7478_27751# a_7343_27849# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2112 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2113 a_5700_24563# a_5439_24563# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2114 a_6058_18445# a_5849_18463# a_5394_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2115 VGND th_dif_sw_0.th_sw_1.CK a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X2116 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2117 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2118 a_10830_19068# a_10553_18922# a_11160_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2119 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2120 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2121 a_2508_23444# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2122 VGND sar9b_0.net56 a_5322_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2123 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2124 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2125 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2126 a_10548_19053# sar9b_0.net7 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2127 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2128 a_15400_11316# tdc_0.phase_detector_0.INP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X2129 VGND a_4083_28566# uio_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2130 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2131 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2132 a_10816_21487# a_10218_21842# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2133 VGND clk a_4332_23043# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X2134 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2135 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2136 a_3438_27677# a_3156_27447# a_3799_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2137 VGND a_8883_27466# sar9b_0.net45 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2138 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2139 a_12246_26198# a_12182_26419# a_12168_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2140 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2141 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2142 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2143 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2144 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2145 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2146 a_5742_28392# a_5465_28246# a_6072_28502# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2147 a_9130_26198# a_8340_26115# a_8622_26345# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2148 a_6922_23534# a_6132_23451# a_6414_23681# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2149 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2150 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2151 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2152 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2153 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2154 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2155 a_35519_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2156 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2157 VDPWR sar9b_0.net25 a_12531_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2158 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2159 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2160 a_5846_17626# a_5711_17527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2161 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2162 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2163 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2164 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2165 VDPWR a_6744_23238# a_6861_22828# VDPWR sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.475 as=0.51 ps=3.02 w=1 l=0.25
X2166 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2167 VGND sar9b_0.net54 a_5910_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2168 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2169 a_10182_20463# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2170 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2171 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2172 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2173 a_10620_17903# a_9450_17846# a_10410_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2175 a_3799_27849# a_3370_27769# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2176 a_11339_27039# sar9b_0.net31 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X2177 VDPWR sar9b_0.net42 a_10378_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X2178 VDPWR a_11859_21906# single_9b_cdac_1.CF[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2180 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2182 a_2940_25096# sar9b_0.net68 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X2183 VGND a_7188_22119# a_7193_22459# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2185 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2186 a_12168_26198# a_11842_26426# a_12047_26517# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2187 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2188 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2189 a_6072_28502# a_5674_28147# a_5994_28502# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2190 single_9b_cdac_0.SW[2] a_13067_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2191 VDPWR a_7338_24802# a_7590_24931# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2192 a_5633_20244# a_5481_20185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X2193 a_5844_18123# sar9b_0.net6 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2194 VGND sar9b_0.net48 a_10038_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2195 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2196 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2197 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2198 a_7374_19685# a_7097_19795# a_7704_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2199 th_dif_sw_0.CKB a_2603_17006# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X2200 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2201 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2202 a_65367_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2203 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2204 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2205 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2206 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2207 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2208 sar9b_0.net43 a_5100_24375# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2210 VDPWR a_9870_27060# a_9802_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2211 a_12182_26419# a_12047_26517# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X2212 VGND sar9b_0.net53 a_12246_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2213 VDPWR a_4011_22488# a_4210_22378# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2214 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2215 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2216 VGND single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2217 VDPWR a_9939_28566# uo_out[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2218 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2219 single_9b_cdac_1.CF[7] a_12435_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2220 a_11430_20935# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2221 sar9b_0.net16 a_3922_20239# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X2222 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2223 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2224 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2225 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2226 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2227 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2228 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2229 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2230 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2231 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2232 a_2603_17006# sar9b_0.net16 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2235 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2236 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2237 uo_out[4] a_8691_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2238 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2239 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2240 a_5711_17527# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2241 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2242 VDPWR a_7092_19455# a_7097_19795# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2243 a_6126_18353# a_5844_18123# a_6487_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2244 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2245 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2246 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2247 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2248 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2249 a_7704_19538# a_7306_19777# a_7626_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2250 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2251 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2252 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2253 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2254 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2255 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2256 VDPWR a_7374_19685# a_7306_19777# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2257 VGND a_8334_18353# a_8266_18445# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2258 single_9b_cdac_1.SW[5] a_13011_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2259 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2260 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2261 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2262 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2263 VGND clk a_15197_10290# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X2264 VGND a_12064_22819# sar9b_0.net30 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2266 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2267 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2268 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2269 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2270 VDPWR sar9b_0.net9 a_13011_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2271 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2272 VGND a_2603_17006# th_dif_sw_0.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2273 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2274 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2275 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2276 sar9b_0.net23 a_7692_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X2277 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2278 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2279 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2280 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2281 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2282 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2283 a_6487_18525# a_6058_18445# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2284 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2286 VGND a_13011_17910# single_9b_cdac_1.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2287 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2288 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2289 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2290 VDPWR a_7443_21496# sar9b_0.net47 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X2291 a_7626_19538# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2292 VDPWR a_12182_19759# a_12137_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2293 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2294 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2295 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2296 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2297 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2298 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2299 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2300 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2301 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2302 a_7728_24809# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2303 a_2508_23444# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X2304 a_7483_23174# sar9b_0.clk_div_0.COUNT\[1\] sar9b_0._17_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X2305 VGND sar9b_0.net56 a_10218_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2306 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2307 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2308 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2309 a_10506_24506# a_9546_24506# a_10070_24286# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2310 a_8052_18123# sar9b_0.net56 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2311 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2312 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2313 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2314 a_11842_18434# a_11658_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2315 VDPWR sar9b_0.net39 a_11859_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2316 VGND sar9b_0.net48 a_10422_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2317 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2318 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2319 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2320 VGND sar9b_0.net56 a_9450_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2321 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2322 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2323 a_12047_26517# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2324 a_5651_20547# a_5126_20140# a_5481_20185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X2325 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2326 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y a_30717_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2327 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2328 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2329 a_6282_27170# a_5506_26802# a_5846_26950# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2330 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2331 VDPWR sar9b_0.clk_div_0.COUNT\[1\] a_3219_22860# VDPWR sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X2332 VDPWR a_6282_17846# a_6534_17799# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2333 a_9960_17846# a_9634_17478# a_9839_17527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2334 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2335 a_15197_10290# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_15151_10456# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X2336 a_13008_19481# sar9b_0.net50 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2337 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2338 a_7890_26108# a_8340_26115# a_8292_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2339 VDPWR a_5441_22522# a_5396_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X2340 VDPWR sar9b_0.net51 a_6579_18832# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X2341 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2342 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2344 VDPWR a_4083_28566# uio_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2345 a_7404_17715# sar9b_0.net1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2051 ps=1.52 w=0.84 l=0.15
X2346 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2347 a_8166_27595# a_7914_27466# a_8304_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X2348 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2349 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2350 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2352 a_6538_24506# sar9b_0.net62 a_7059_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2353 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2354 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2355 single_9b_cdac_1.CF[2] a_11859_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2356 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2357 a_6307_27584# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X2358 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2359 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2360 dw_12589_1395# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VDPWR dw_12589_1395# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X2361 a_6126_18353# a_5849_18463# a_6456_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2362 a_8694_20570# sar9b_0.net61 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2363 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2364 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2365 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2366 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2367 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2368 a_8292_26141# a_8031_26141# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2369 VGND a_10758_24459# a_10716_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2370 a_7830_18149# a_7602_18116# a_7743_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2371 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2373 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2374 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2375 VGND a_12531_28566# uo_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2376 a_5396_22567# a_4755_22138# a_5289_22527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X2377 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A a_49926_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2378 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2380 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2381 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2382 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2383 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2384 VGND th_dif_sw_0.th_sw_1.CK a_10482_3438# VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X2385 a_36555_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2387 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2388 VGND a_3713_22522# a_3731_22165# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X2389 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2390 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2391 a_9162_23174# a_8386_22806# a_8726_22954# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2392 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2393 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2394 a_7059_24566# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2395 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2396 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2397 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2398 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2399 a_3713_22522# a_3561_22527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2400 sar9b_0.net46 a_6579_18832# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2401 sar9b_0.net4 a_5331_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2402 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2403 a_6456_18206# a_6058_18445# a_6378_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2404 VDPWR a_5846_17626# a_5801_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2405 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2406 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2407 VDPWR a_6126_18353# a_6058_18445# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2408 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2410 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2411 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2412 a_10716_24563# a_9546_24506# a_10506_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2413 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2414 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2415 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2416 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2418 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2419 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2420 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2421 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2423 a_60565_15501# single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2424 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2425 single_9b_cdac_1.CF[7] a_12435_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2426 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2427 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2428 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2429 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2430 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2431 a_12491_27662# sar9b_0.net29 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2432 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2433 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2434 a_8004_18149# a_7743_18149# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2435 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2436 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2437 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2438 a_6378_18206# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2439 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2440 VDPWR a_13011_17910# single_9b_cdac_1.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2441 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2442 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2443 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2444 single_9b_cdac_1.CF[6] a_13011_24570# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2445 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2446 VDPWR a_2547_28132# sar9b_0.net60 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2447 a_7638_19238# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2448 VGND a_16159_13315# tdc_0.RDY VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X2449 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2450 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X2451 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2454 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2455 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2456 single_9b_cdac_0.SW[8] a_9323_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2457 a_6282_27170# a_5322_27170# a_5846_26950# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2458 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2459 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2460 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2461 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2462 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2463 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2464 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2465 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2467 a_4365_25770# a_4125_25958# a_4588_25473# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.0504 ps=0.66 w=0.42 l=0.15
X2468 VDPWR sar9b_0.net59 a_9870_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2469 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2470 VDPWR sar9b_0.net51 a_7443_21496# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X2471 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2472 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2473 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2474 VGND a_13216_22473# sar9b_0.net31 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2475 a_5844_18123# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2476 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2477 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2478 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2479 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2480 a_4771_18260# sar9b_0.net57 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2481 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2483 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2484 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2485 VGND sar9b_0.net1 a_10707_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2486 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2487 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2488 a_3880_20524# a_2739_20140# a_3723_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X2489 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2490 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2491 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2492 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2493 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2494 sar9b_0.net20 a_4812_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2495 a_3369_24181# a_2835_24136# a_3262_24141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X2496 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2497 sar9b_0._10_ a_5581_19664# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X2498 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2499 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2500 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2501 a_4588_25473# a_4293_25852# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.18985 ps=1.545 w=0.42 l=0.15
X2502 VDPWR a_12182_23755# a_12137_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2503 single_9b_cdac_1.SW[8] a_11859_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2504 VGND sar9b_0.net50 a_11469_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2505 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2506 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2507 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2508 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2509 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2510 a_6391_24187# a_5962_24151# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2511 VDPWR a_6902_25087# a_6857_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2512 a_6834_20780# a_7289_21127# a_7238_21225# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2513 VGND a_7404_17715# sar9b_0.net73 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X2514 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2515 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2516 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2517 a_7548_24809# a_6378_24802# a_7338_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2518 VGND a_8940_24402# sar9b_0.net62 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2519 VDPWR sar9b_0.net7 a_11859_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2520 single_9b_cdac_1.SW[1] a_10803_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2521 VGND tdc_0.OUTN a_6867_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2522 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2523 a_9162_23174# a_8202_23174# a_8726_22954# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2524 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2525 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2526 a_6307_27584# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2527 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2528 VGND a_10227_18142# th_dif_sw_0.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2529 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2530 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2531 sar9b_0._14_ sar9b_0.net63 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2532 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2533 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2534 sar9b_0.net52 a_9165_24988# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2535 VGND a_11776_25137# sar9b_0.net13 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2536 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2537 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2538 a_15052_11404# tdc_0.phase_detector_0.INN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X2539 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2540 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2541 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2542 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2543 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2544 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2545 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2546 sar9b_0.net16 a_3922_20239# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X2547 a_11469_18146# sar9b_0.net73 a_11382_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2550 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2551 VDPWR sar9b_0.net9 a_10506_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2552 a_11776_21141# a_11178_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2553 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2554 a_6857_25185# a_6378_24802# a_6767_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2555 VDPWR a_11104_24151# sar9b_0.net42 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2556 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2557 VDPWR a_12531_28566# uo_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2558 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2559 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2560 a_11544_25838# a_11146_25483# a_11466_25838# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2561 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2562 VDPWR clk a_16527_10454# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X2563 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2564 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2565 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2566 a_11178_27466# a_10402_27758# a_10742_27751# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2567 a_6767_25185# a_6378_24802# a_6102_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2568 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2569 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2570 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2571 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2572 VGND a_6252_19074# sar9b_0.net55 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2573 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2574 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2575 VGND tdc_0.phase_detector_0.pd_out_0.B a_16159_13315# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X2576 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2577 single_9b_cdac_0.SW[0] a_13011_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2578 sar9b_0.net47 a_7443_21496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2579 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2580 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2581 VGND sar9b_0.net47 a_5581_19664# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X2582 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2583 a_13067_27662# sar9b_0.net28 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2584 a_10402_21098# a_10218_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2585 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2586 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2587 a_9942_24806# sar9b_0.net12 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2588 a_7443_23474# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2589 sar9b_0.net74 a_10707_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2590 VGND sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X2591 single_9b_cdac_1.SW[3] a_10803_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2592 a_31753_15501# single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2593 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2594 a_3425_20244# a_3273_20185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2595 a_8842_18206# a_8052_18123# a_8334_18353# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2596 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2597 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2598 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2599 a_11016_23174# a_10690_22806# a_10895_22855# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2600 VDPWR a_5443_19074# sar9b_0.net57 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2601 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2602 a_6642_19448# a_7092_19455# a_7044_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2603 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2604 a_3747_25724# a_3855_25792# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1862 ps=1.475 w=0.84 l=0.15
X2605 VGND a_9165_24988# sar9b_0.net52 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X2606 a_8303_23853# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2607 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2608 a_11466_25838# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2609 a_3754_26815# a_3540_27045# a_3090_27163# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2610 VGND a_13011_17910# single_9b_cdac_1.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2611 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2612 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2613 a_16222_11316# tdc_0.phase_detector_0.INN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X2614 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2615 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2616 a_6250_28502# sar9b_0.net38 a_6771_28562# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2617 a_3540_27045# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2618 VDPWR single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2619 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2620 a_10608_21899# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2621 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2622 a_6880_17491# a_6282_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2623 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2624 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2625 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2626 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2627 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2628 VDPWR sar9b_0.net27 a_13011_27234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2629 a_3819_24136# a_2835_24136# a_3521_24240# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X2630 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2631 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2632 VDPWR a_9138_27163# a_8940_27039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2633 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2634 a_10402_27758# a_10218_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2635 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2636 VGND a_3438_26345# a_3370_26437# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2637 VDPWR a_13216_26469# sar9b_0.net33 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2638 sar9b_0.net51 a_5811_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15198 ps=1.17 w=0.74 l=0.15
X2639 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2640 a_5439_24563# a_5298_24499# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2641 VDPWR a_8874_23470# a_9126_23599# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2642 VGND a_12435_20806# single_9b_cdac_1.CF[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2643 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2644 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2645 a_6360_24506# a_5962_24151# a_6282_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2646 VGND sar9b_0.net49 a_10806_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2647 a_3690_27530# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2648 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2649 VDPWR a_12870_23599# a_12820_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2650 a_59529_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2651 VGND a_13067_27662# single_9b_cdac_0.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2652 a_7602_16784# a_8052_16791# a_8004_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2653 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2654 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2655 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2656 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2657 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2658 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2659 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2660 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2661 VDPWR a_13011_21906# single_9b_cdac_1.CF[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2662 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2663 a_2706_27440# a_3156_27447# a_3108_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2664 a_2508_20780# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X2665 VDPWR a_10548_19053# a_10553_18922# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2666 single_9b_cdac_1.SW[0] a_8595_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2667 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2668 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2670 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2671 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2672 VDPWR sar9b_0.net54 a_6030_24396# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2673 a_11434_16874# sar9b_0.net61 a_11955_16814# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2675 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2676 VDPWR sar9b_0.net3 a_2547_28132# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X2677 a_12820_22557# a_11842_22430# a_12618_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X2678 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2679 VDPWR sar9b_0.net52 a_11382_26138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2680 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2681 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2682 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2683 a_10482_25831# a_10937_25582# a_10886_25483# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2684 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2685 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2686 a_3156_26115# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2687 a_6282_24506# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2688 VGND a_10803_18142# single_9b_cdac_1.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2689 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2690 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2691 th_dif_sw_0.VCN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X2692 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2693 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2694 a_10806_20870# a_10742_21091# a_10728_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2695 a_7882_19538# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X2696 a_10607_27849# a_10218_27466# a_9942_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2697 VGND sar9b_0.net49 a_8781_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2698 VDPWR a_5931_20140# a_6130_20239# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2699 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2700 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2701 VDPWR a_4236_21738# sar9b_0.net67 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2702 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2703 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2704 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2705 a_12588_16784# tdc_0.OUTP VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2707 a_3108_27473# a_2847_27473# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2708 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2709 sar9b_0.net27 a_5196_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X2710 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2711 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2712 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2713 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2714 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2715 VGND a_6642_19448# a_6444_19448# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2716 a_9472_18823# a_8874_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2717 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2718 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2719 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X2720 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2721 VGND a_10548_19053# a_10553_18922# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2722 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2723 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2724 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2725 a_7498_21109# a_7284_20787# a_6834_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2726 VGND sar9b_0.net53 a_11469_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2727 a_10728_20870# a_10402_21098# a_10607_21189# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2728 a_10858_17113# a_10644_16791# a_10194_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2729 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2730 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2731 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2732 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2733 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2734 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2735 a_3371_23106# sar9b_0.clk_div_0.COUNT\[2\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X2736 VDPWR a_10816_21487# sar9b_0.net9 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2737 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2738 VGND sar9b_0.net59 a_2934_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2739 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2741 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2742 a_8622_26345# a_8345_26455# a_8952_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2743 a_3647_23194# a_3219_22860# a_3371_23106# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X2744 a_6414_23681# a_6137_23791# a_6744_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2746 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2747 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2748 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2749 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2750 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2751 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2752 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2753 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2754 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2755 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2756 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2757 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2758 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2759 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# a_16357_9613# VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X2760 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2761 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2762 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2763 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2764 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2765 sar9b_0.clk_div_0.COUNT\[3\] a_4210_22378# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X2766 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2767 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2768 a_11469_22142# sar9b_0.net73 a_11382_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2769 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2770 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2771 VGND a_2706_27440# a_2508_27440# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2772 VDPWR a_7478_27751# a_7433_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2773 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2774 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2775 VGND sar9b_0.net49 a_9069_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2776 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCP VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X2777 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2778 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2779 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2780 a_12047_26517# a_11658_26134# a_11382_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2781 a_4934_22432# a_4755_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2782 VGND a_5844_18123# a_5849_18463# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2783 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2784 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2785 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2786 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2787 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2788 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2789 VDPWR sar9b_0.net4 a_6378_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2790 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2791 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2792 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2793 a_7566_21017# a_7289_21127# a_7896_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2794 a_10607_21189# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2795 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2796 VGND a_13011_20806# single_9b_cdac_1.CF[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2797 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2798 VGND sar9b_0.net42 a_13011_19242# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X2799 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2800 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2801 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2802 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2803 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2804 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2805 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2806 a_2893_24992# sar9b_0._14_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X2807 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2808 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2809 a_7936_25137# a_7338_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2810 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2812 VDPWR sar9b_0.net49 a_9942_20810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2814 VGND a_13011_27234# single_9b_cdac_0.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2815 VDPWR a_2603_17006# th_dif_sw_0.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2816 a_9069_21902# sar9b_0.net8 a_8982_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2817 single_9b_cdac_1.CF[4] a_13011_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2818 a_5931_20140# a_5126_20140# a_5633_20244# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X2819 VDPWR sar9b_0.net12 a_9546_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2820 a_2918_20140# a_2739_20140# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2821 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2822 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2823 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2824 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2825 a_11430_27595# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2826 a_7338_24802# a_6562_25094# a_6902_25087# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2827 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2828 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2829 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2830 a_11842_26426# a_11658_26134# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2831 VGND a_12491_27662# single_9b_cdac_0.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X2832 a_7896_20870# a_7498_21109# a_7818_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2833 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2834 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2835 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2836 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2837 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2838 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2839 a_3014_24136# a_2835_24136# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X2840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2841 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2842 VDPWR a_5739_22488# a_5938_22378# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2843 VDPWR a_3795_19512# a_4292_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2557 pd=1.59 as=0.21 ps=1.42 w=1 l=0.15
X2844 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2845 VDPWR a_10803_18142# single_9b_cdac_1.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2846 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2847 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2848 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2849 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2850 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2851 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2852 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2853 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X2854 VGND a_10227_18142# th_dif_sw_0.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2856 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2857 VGND single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2858 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2859 VGND a_13216_19809# sar9b_0.net29 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2860 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2861 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2862 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2863 VDPWR a_10470_21795# a_10420_21487# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2864 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2865 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2866 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2867 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2868 a_7818_20870# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2869 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2870 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2871 VGND a_6534_17799# a_6492_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2872 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2873 VGND a_8052_18123# a_8057_18463# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2874 VGND sar9b_0.net7 a_11658_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2875 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2876 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2877 a_6562_25094# a_6378_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2878 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2879 sar9b_0.net54 a_7347_24160# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2880 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2882 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2883 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2884 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2885 a_9839_17527# a_9450_17846# a_9174_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2886 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2887 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2888 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2889 VDPWR single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2890 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2891 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2892 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2893 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2895 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2896 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2897 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2898 sar9b_0.net53 a_10227_23490# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X2899 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2900 a_8940_24402# sar9b_0.net2 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2901 VDPWR sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# VDPWR sky130_fd_pr__pfet_01v8 ad=0.27625 pd=1.625 as=0.1176 ps=1.4 w=0.42 l=0.15
X2902 VDPWR tdc_0.OUTN a_6867_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2903 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2904 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2905 a_5126_20140# a_4947_20140# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2906 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2907 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2908 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2909 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2910 a_6492_17903# a_5322_17846# a_6282_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2911 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2912 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2913 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2914 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2915 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2916 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2918 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2919 a_12182_18427# a_12047_18525# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2920 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2921 a_45123_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2922 a_8266_18445# a_8057_18463# a_7602_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2923 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2924 a_5801_26851# a_5322_27170# a_5711_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2925 a_9839_17527# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2926 single_9b_cdac_1.SW[4] a_11859_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2927 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2928 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2929 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2930 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2931 VDPWR sar9b_0.net58 a_5742_28392# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2932 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y a_25915_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2933 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2934 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2935 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2936 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2937 VGND sar9b_0.net63 sar9b_0._02_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2938 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2939 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2940 a_3156_26115# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2941 a_6975_20813# a_6834_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2942 VDPWR a_7602_16784# a_7404_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2943 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2944 a_5994_28502# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2945 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2946 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2947 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2948 VGND a_12435_20806# single_9b_cdac_1.CF[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2949 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2950 single_9b_cdac_0.SW[8] a_9323_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X2951 VGND a_9126_23599# a_9084_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2952 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2953 VGND a_3822_27060# a_3754_26815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2954 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2955 single_9b_cdac_1.CF[8] a_13011_25902# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2956 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2957 VDPWR sar9b_0._14_ a_4467_24162# VDPWR sky130_fd_pr__pfet_01v8 ad=0.36323 pd=1.84 as=0.126 ps=1.14 w=0.84 l=0.15
X2958 single_9b_cdac_1.CF[0] a_13011_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2959 VGND single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2960 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2961 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2962 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2963 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2964 VDPWR sar9b_0.net57 a_9258_21842# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2965 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2966 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X2967 a_6250_28502# a_5465_28246# a_5742_28392# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X2968 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X2969 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2970 a_13216_26469# a_12618_26134# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2971 VDPWR a_5523_21528# sar9b_0._12_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.196 ps=1.47 w=1.12 l=0.15
X2972 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2973 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2974 a_8681_22855# a_8202_23174# a_8591_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2975 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2976 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2977 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2978 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2979 VGND a_10803_18142# single_9b_cdac_1.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2980 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2981 VDPWR a_12491_27662# single_9b_cdac_0.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2982 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2983 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2984 a_10886_25483# a_10623_25895# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X2985 a_9084_23477# a_7914_23470# a_8874_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2986 a_5441_22522# a_5289_22527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2987 sar9b_0.net70 a_3027_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2988 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2989 VDPWR a_13011_27234# single_9b_cdac_0.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2990 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2992 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2993 a_3540_27045# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2994 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2995 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2996 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2997 VDPWR a_10227_18142# th_dif_sw_0.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2999 a_9154_20142# a_8970_20510# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3000 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3001 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3002 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3003 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3004 a_4811_23656# sar9b_0.net72 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.13062 pd=1.025 as=0.15198 ps=1.17 w=0.55 l=0.15
X3005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3006 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3007 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3008 a_12870_26263# a_12618_26134# a_13008_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3009 ua[4] th_dif_sw_0.th_sw_1.CK ua[4] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X3010 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3011 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3012 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3013 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3014 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3015 a_11380_25221# a_10402_25094# a_11178_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3016 a_7882_19538# a_7097_19795# a_7374_19685# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3017 a_8334_18353# a_8052_18123# a_8695_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3018 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3019 a_10742_21091# a_10607_21189# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3020 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3021 VGND a_11339_27039# single_9b_cdac_0.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X3022 a_12820_19893# a_11842_19766# a_12618_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3023 VGND a_4771_18260# sar9b_0.net56 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3024 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3025 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3026 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y a_40321_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3027 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3028 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3030 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3031 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3032 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3033 a_4698_25851# a_4136_25584# a_4365_25770# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X3034 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3035 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3036 VGND a_13216_23805# sar9b_0.net32 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3037 VDPWR a_6252_20780# sar9b_0._01_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3039 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3040 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3041 a_5702_24151# a_5439_24563# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3042 VGND a_5938_22378# a_5896_22188# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X3043 VGND sar9b_0.net54 a_6189_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3044 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3045 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3046 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3047 VDPWR sar9b_0.clknet_0_CLK a_2508_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3048 a_5739_22488# a_4934_22432# a_5441_22522# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X3049 VGND sar9b_0.net48 a_7725_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3050 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3051 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3052 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3054 a_8695_18525# a_8266_18445# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X3055 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3056 VGND a_6307_27584# sar9b_0.net44 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3057 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3058 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3059 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3060 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3061 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3062 a_4332_23043# clk VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X3063 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3064 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3065 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3066 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3067 a_3946_27530# a_3161_27787# a_3438_27677# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3068 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3069 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3070 VGND a_13011_20806# single_9b_cdac_1.CF[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3071 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3072 a_5182_22567# sar9b_0.net64 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X3073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3074 VGND a_5196_19448# sar9b_0.net71 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3075 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3076 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3077 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3078 VGND a_12870_26263# a_12828_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3079 a_6189_24806# sar9b_0.net13 a_6102_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3080 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3081 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3082 VGND a_13011_27234# single_9b_cdac_0.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3083 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3084 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3086 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3087 a_7725_19238# sar9b_0.net73 a_7638_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3088 th_dif_sw_0.CK a_10227_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3089 a_11104_24151# a_10506_24506# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3090 VDPWR clk a_14871_9671# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X3091 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3092 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3093 a_6902_25087# a_6767_25185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3094 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3095 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3096 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3097 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3098 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3099 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3100 a_4083_25852# a_3747_25724# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1197 ps=1.41 w=0.42 l=0.15
X3101 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3102 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3103 single_9b_cdac_1.CF[2] a_11859_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3104 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A a_30717_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3105 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3106 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3108 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3109 single_9b_cdac_0.SW[6] a_9323_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3110 VDPWR a_13067_27662# single_9b_cdac_0.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3111 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3112 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3113 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3114 a_8334_18353# a_8057_18463# a_8664_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X3115 VDPWR sar9b_0.net38 a_10803_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3116 a_10378_27170# sar9b_0.net42 a_10899_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3117 a_12828_26141# a_11658_26134# a_12618_26134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3118 a_10895_22855# a_10506_23174# a_10230_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3119 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3120 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3121 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3122 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3123 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3124 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3125 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3126 uo_out[3] a_9939_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3127 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3128 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3129 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3130 VDPWR a_11178_20806# a_11430_20935# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3131 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3132 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3133 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3134 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3135 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3136 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3137 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3138 single_9b_cdac_1.SW[2] a_8019_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3139 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3140 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3141 uo_out[2] a_10995_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3142 VDPWR sar9b_0._07_ a_5523_21528# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2786 pd=1.64 as=0.2478 ps=2.27 w=0.84 l=0.15
X3143 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3144 VGND a_11430_20935# a_11388_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3145 a_7092_19455# sar9b_0.net10 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3146 a_6634_18206# a_5849_18463# a_6126_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3147 VDPWR a_8052_18123# a_8057_18463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3148 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3149 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3150 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3151 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3152 VGND sar9b_0.net45 a_10218_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3153 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3154 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3155 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3156 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3157 a_8664_18206# a_8266_18445# a_8586_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3158 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3159 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3160 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3161 a_10899_27230# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3162 sar9b_0.net54 a_7347_24160# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X3163 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3164 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3165 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3166 VDPWR a_8334_18353# a_8266_18445# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3167 VDPWR a_5742_28392# a_5674_28147# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3168 VGND a_8334_17021# a_8266_17113# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3169 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3170 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3171 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3172 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3173 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3174 VGND a_10482_25831# a_10284_25707# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3175 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3176 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3177 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3178 a_26951_15501# single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3180 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3181 a_6767_25185# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3182 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3183 a_3318_27227# a_3090_27163# a_3231_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3184 VDPWR a_11214_25728# a_11146_25483# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3185 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3186 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3187 a_10254_2858# th_dif_sw_0.th_sw_1.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X3188 VGND a_5682_23444# a_5484_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3189 a_11388_20813# a_10218_20806# a_11178_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3190 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3191 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3192 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3193 VDPWR a_9494_20290# a_9449_20191# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3194 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3195 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3196 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3197 VDPWR a_11859_20574# single_9b_cdac_1.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3198 a_8586_18206# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3199 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3200 single_9b_cdac_0.SW[5] a_11339_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3201 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3202 VGND a_3156_26115# a_3161_26455# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3203 single_9b_cdac_0.SW[6] a_9323_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3204 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3205 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3206 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3207 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3208 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3209 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3210 a_8052_16791# sar9b_0.net5 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3211 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3212 VDPWR sar9b_0._03_ a_4698_25851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2972 pd=2.41 as=0.09835 ps=1.005 w=0.42 l=0.15
X3213 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3214 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3215 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3216 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3217 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3218 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3219 a_10254_2858# th_dif_sw_0.th_sw_1.CKB a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X3220 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3221 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3222 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3223 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3224 a_6870_19481# a_6642_19448# a_6783_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3225 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3226 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3227 VGND sar9b_0.net18 a_4083_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3228 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3229 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3230 VGND sar9b_0.net50 a_12246_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3231 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3232 uio_out[0] a_4083_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3233 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3235 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3236 VGND sar9b_0._14_ a_4673_24464# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.111 ps=1.045 w=0.64 l=0.15
X3237 a_10607_21189# a_10218_20806# a_9942_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3238 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3239 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3240 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3241 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3242 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3243 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3244 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3245 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3246 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3247 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3249 a_3370_26437# a_3161_26455# a_2706_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3250 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3251 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3252 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3253 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3254 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3255 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3256 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3257 VDPWR sar9b_0.net49 a_8694_20570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3258 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3259 uio_out[1] a_2931_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3260 sar9b_0.net24 a_8940_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3261 VGND a_9472_18823# sar9b_0.net26 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3262 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3263 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3264 a_9323_28371# sar9b_0.net32 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X3265 VGND a_11718_23127# a_11676_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3266 a_10029_20810# sar9b_0.net7 a_9942_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3267 a_7830_16817# a_7602_16784# a_7743_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3268 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3269 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3270 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3271 VGND a_8512_27801# sar9b_0.net22 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3272 single_9b_cdac_0.SW[5] a_11339_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X3273 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X3274 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3275 VDPWR a_11718_23127# a_11668_22819# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3276 a_2934_27473# a_2706_27440# a_2847_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3277 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3278 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3279 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3280 VGND a_3723_20140# a_3922_20239# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X3281 VDPWR sar9b_0.net63 a_6286_22804# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X3282 tdc_0.phase_detector_0.INP a_15151_10456# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3283 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3284 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3285 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3286 VGND a_11214_25728# a_11146_25483# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3287 VGND a_10194_16784# a_9996_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3288 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3289 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3290 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3291 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3292 sar9b_0.net15 a_6130_20239# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X3293 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3294 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3295 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3296 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3297 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3298 sar9b_0.net70 a_3027_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3299 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3300 a_8098_23762# a_7914_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3301 a_11676_23231# a_10506_23174# a_11466_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3302 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3303 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3304 VDPWR sar9b_0.net54 a_6414_23681# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X3305 sar9b_0.clk_div_0.COUNT\[0\] a_5938_22378# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X3306 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3307 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3308 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3309 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3310 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3312 a_7590_24931# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3313 a_21684_3438# VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X3314 VDPWR a_12435_24802# single_9b_cdac_1.CF[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3315 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3316 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3317 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[3] a_50962_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3318 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3319 a_5682_23444# a_6132_23451# a_6084_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3320 VGND a_6534_27123# a_6492_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3321 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3322 VGND th_dif_sw_0.VCN a_14897_9355# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3323 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3324 a_11718_23127# a_11466_23174# a_11856_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3325 VGND sar9b_0.net69 sar9b_0._04_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3326 VGND sar9b_0.net51 a_7443_21496# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X3327 a_8004_16817# a_7743_16817# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3328 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3329 uo_out[3] a_9939_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3330 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3331 VGND a_5812_21028# a_5581_20992# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17462 pd=1.185 as=0.077 ps=0.83 w=0.55 l=0.15
X3332 single_9b_cdac_1.SW[6] a_13011_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3333 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3334 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3335 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3336 a_10932_25713# sar9b_0.net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3337 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3338 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3339 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3340 VDPWR sar9b_0.net48 a_7638_19238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3341 VGND a_13011_20574# single_9b_cdac_1.CF[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3342 sar9b_0.net24 a_8940_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X3343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3344 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3345 a_11955_16814# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3346 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3347 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3348 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3349 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3350 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3352 VGND a_3521_24240# a_3539_24543# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X3353 VDPWR a_9126_19131# a_9076_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3354 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3355 a_3438_26345# a_3156_26115# a_3799_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3356 VGND a_6030_24396# a_5962_24151# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3357 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3358 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3359 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3360 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3361 a_6084_23477# a_5823_23477# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3362 sar9b_0.net1 a_6867_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X3363 a_6492_27227# a_5322_27170# a_6282_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3364 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3365 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3366 uo_out[4] a_8691_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3367 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3368 VGND single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3369 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3370 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3371 a_6744_23238# a_6484_22845# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.27625 ps=1.625 w=1 l=0.25
X3372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3373 VGND sar9b_0.net4 a_6378_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3374 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3375 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3376 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3377 VDPWR a_3521_24240# a_3476_24141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X3378 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3379 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3381 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3382 tdc_0.OUTN tdc_0.OUTP a_16555_12412# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3383 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3384 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3385 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3386 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3387 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3388 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3389 a_3799_26517# a_3370_26437# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X3390 VDPWR a_11859_20574# single_9b_cdac_1.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3391 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3392 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3393 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3394 VDPWR a_10803_19474# single_9b_cdac_1.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3395 a_15151_10456# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X3396 a_2508_20780# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X3397 a_12684_20379# sar9b_0.net51 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24915 pd=2.37 as=0.15198 ps=1.17 w=0.55 l=0.15
X3398 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3399 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3400 a_8952_26198# a_8554_26437# a_8874_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3401 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3402 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3403 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3404 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3405 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3406 a_3476_24141# a_2835_24136# a_3369_24181# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X3407 VGND sar9b_0.net53 a_12246_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3408 a_9264_19235# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3409 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3410 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3411 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3412 a_6902_25087# a_6767_25185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3413 VDPWR a_6444_21738# sar9b_0.net64 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3414 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3415 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3416 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3417 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3418 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3419 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3420 a_12047_19857# a_11842_19766# a_11382_19478# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3421 single_9b_cdac_1.SW[7] a_13011_19242# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3423 VGND sar9b_0.net25 a_12531_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3424 a_10690_22806# a_10506_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3425 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3426 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3427 uo_out[1] a_12531_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3428 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3429 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3430 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3431 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3432 a_10230_23234# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3433 a_8874_26198# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3434 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3435 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3436 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3437 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3438 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3439 VGND sar9b_0.net47 a_6870_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X3440 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3441 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3442 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3443 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3444 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y a_64331_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3445 VDPWR a_2892_23070# sar9b_0.net66 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3446 VDPWR a_13011_24802# single_9b_cdac_0.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3447 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3448 VDPWR sar9b_0.net13 a_13011_25902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3449 a_12491_27662# sar9b_0.net29 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X3450 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3453 VDPWR sar9b_0.net5 a_13011_20574# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3454 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3455 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3456 VDPWR a_7936_25137# sar9b_0.cyclic_flag_0.FINAL VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3457 VDPWR a_4812_21738# sar9b_0.net65 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3458 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3459 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3460 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3461 a_5443_19074# sar9b_0.net4 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X3462 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3463 a_3690_26198# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3464 a_12684_20379# sar9b_0.net51 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2051 ps=1.52 w=0.84 l=0.15
X3465 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X3467 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3468 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3469 a_3946_27530# a_3156_27447# a_3438_27677# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X3470 sar9b_0.net3 a_2451_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3471 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3472 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3473 sar9b_0._12_ sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2786 ps=1.64 w=1.12 l=0.15
X3474 VDPWR a_12182_18427# a_12137_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3475 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3476 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3477 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3478 sar9b_0.net10 a_6636_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3479 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3480 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3481 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3482 a_8074_20870# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3483 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3484 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3485 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3486 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3487 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3488 VGND sar9b_0.net60 a_6765_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3489 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3490 VGND sar9b_0.net36 a_10803_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3491 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3492 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3493 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3494 VGND a_3540_27045# a_3545_26914# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3495 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3496 a_9974_17626# a_9839_17527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3497 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3498 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3499 a_10607_25185# a_10402_25094# a_9942_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3500 VDPWR sar9b_0.net54 a_5439_24563# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X3501 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3502 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3503 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A a_55773_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3504 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3505 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3506 a_3166_20145# sar9b_0._00_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X3507 VGND sar9b_0.net8 a_8970_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3508 sar9b_0.net4 a_5331_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X3509 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3510 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3511 a_54737_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3512 a_6538_24506# a_5748_24381# a_6030_24396# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X3513 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3514 VGND th_dif_sw_0.VCP a_17125_9355# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3515 VGND a_9939_28566# uo_out[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3516 a_9480_20510# a_9154_20142# a_9359_20191# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3517 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3518 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3519 single_9b_cdac_1.CF[4] a_13011_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3520 a_10762_18823# a_10548_19053# a_10098_19171# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X3521 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[8] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3522 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3523 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3524 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3525 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3526 a_10548_19053# sar9b_0.net7 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3527 a_16357_9613# th_dif_sw_0.VCN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3528 a_7978_22202# sar9b_0.net61 a_8499_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3529 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3530 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3531 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3532 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3533 sar9b_0.net60 a_2547_28132# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3534 a_6765_27470# sar9b_0.net40 a_6678_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3535 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3536 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3537 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3538 VGND a_10995_28566# uo_out[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3539 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3540 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3541 VDPWR sar9b_0.net45 a_12560_27128# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X3542 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3543 VDPWR sar9b_0.net62 a_7882_19538# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X3544 VGND sar9b_0.net46 a_5910_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3545 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3546 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3547 VGND a_3180_19448# sar9b_0._00_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3550 a_3754_26815# a_3545_26914# a_3090_27163# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3551 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3552 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3553 tdc_0.RDY a_16159_13315# a_16185_13034# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X3554 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3555 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3556 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3557 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3558 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3559 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3560 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3561 single_9b_cdac_0.SW[5] a_11339_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3562 a_5298_24499# a_5748_24381# a_5700_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3563 a_8499_22142# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3564 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3565 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A a_46159_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3566 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3567 VGND sar9b_0._03_ a_4698_25851# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.23015 pd=2.1 as=0.15563 ps=1.215 w=0.42 l=0.15
X3568 a_4118_22572# a_3206_22432# a_4011_22488# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X3569 VGND a_7602_18116# a_7404_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3570 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3571 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3572 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3573 a_11668_22819# a_10690_22806# a_11466_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3574 VDPWR single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3575 VGND a_10227_23490# sar9b_0.net53 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3576 VDPWR single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3577 a_6286_22804# sar9b_0._12_ sar9b_0._02_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X3578 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3579 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3580 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3581 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3582 VDPWR sar9b_0.net65 a_3371_23106# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.26 as=0.126 ps=1.14 w=0.84 l=0.15
X3583 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3584 th_dif_sw_0.VCP ua[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3585 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3586 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3587 a_3370_27769# a_3156_27447# a_2706_27440# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X3588 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3589 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3590 a_2637_24802# sar9b_0.net63 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3591 sar9b_0._11_ a_4496_20468# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3592 a_13067_27662# sar9b_0.net28 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X3593 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3594 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3595 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3596 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3597 VGND a_5742_28392# a_5674_28147# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3598 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3599 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3600 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3601 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3602 a_12870_23599# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3603 VGND sar9b_0.net46 a_5133_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3604 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3606 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3607 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3608 a_12047_23853# a_11842_23762# a_11382_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3609 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3610 sar9b_0.net49 a_9363_20826# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X3611 VGND a_10662_17799# a_10620_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3612 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3613 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3614 VDPWR a_10482_25831# a_10284_25707# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3615 VDPWR sar9b_0.clknet_0_CLK a_2508_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3616 VGND a_11859_17910# single_9b_cdac_1.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3618 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3619 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3620 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3621 VGND a_13011_20574# single_9b_cdac_1.CF[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3622 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3623 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3624 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3625 single_9b_cdac_0.SW[0] a_13011_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3626 VDPWR sar9b_0.net57 a_7914_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3627 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3628 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X3629 VGND a_12684_20379# sar9b_0.net50 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X3630 a_11382_19478# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3631 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3632 a_6562_25094# a_6378_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3633 a_9126_19131# a_8874_19178# a_9264_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3634 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3635 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3636 VDPWR single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3637 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3638 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3639 a_5460_28377# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3640 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3641 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3642 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3643 VGND a_7539_28566# uo_out[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3644 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3645 VGND sar9b_0.net41 a_13011_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3646 a_9076_18823# a_8098_18810# a_8874_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3647 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3648 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3649 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3650 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3651 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3652 single_9b_cdac_1.CF[5] a_13011_23238# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3653 VDPWR a_4210_22378# a_4118_22572# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X3654 a_6282_17846# a_5322_17846# a_5846_17626# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3655 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3656 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3657 VDPWR sar9b_0.net24 a_10995_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3658 VGND a_13011_25902# single_9b_cdac_1.CF[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3659 VDPWR sar9b_0.net37 a_8019_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3660 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3661 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3662 a_9730_24138# a_9546_24506# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3663 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3664 VDPWR a_11178_27466# a_11430_27595# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3665 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3666 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3667 a_11776_21141# a_11178_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3668 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3670 VDPWR a_12182_22423# a_12137_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3671 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3672 a_9270_24566# sar9b_0.net62 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3673 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A a_25915_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3675 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3676 a_11842_26426# a_11658_26134# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3677 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3678 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3679 VDPWR sar9b_0.clknet_1_1__leaf_CLK a_2835_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3680 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3681 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3682 VDPWR sar9b_0.net51 a_9363_20826# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X3683 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3684 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3685 VDPWR sar9b_0.net43 a_11859_20574# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3686 single_9b_cdac_1.SW[3] a_10803_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3687 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3688 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3689 uo_out[0] a_11915_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3690 VDPWR a_5298_24499# a_5100_24375# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3691 a_12618_19474# a_11658_19474# a_12182_19759# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3692 VDPWR a_8512_27801# sar9b_0.net22 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3693 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3694 VGND sar9b_0.net49 a_10029_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3695 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3696 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] a_41357_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3697 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3698 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3699 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3700 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3701 a_3090_27163# a_3540_27045# a_3492_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3702 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3703 VDPWR a_10194_16784# a_9996_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3704 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3705 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3707 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3708 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3709 a_3110_27885# a_2847_27473# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3710 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3711 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3712 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3713 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3714 VGND a_10859_26330# single_9b_cdac_0.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3715 a_5739_22488# a_4755_22138# a_5441_22522# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X3716 a_11430_20935# a_11178_20806# a_11568_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3717 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3718 a_11776_25137# a_11178_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3719 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3720 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3721 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3722 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3723 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3724 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3725 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3726 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3727 a_7402_22441# a_7193_22459# a_6738_22112# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3728 sar9b_0.net48 a_10035_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3729 VGND a_8052_16791# a_8057_17131# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3730 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3731 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3732 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3733 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3734 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3735 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3736 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3737 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3738 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3739 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3741 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3742 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3743 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3744 a_9870_27060# a_9588_27045# a_10231_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3745 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3746 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3747 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3748 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3749 a_3492_27227# a_3231_27227# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3750 a_4922_20857# sar9b_0._17_ a_4886_21124# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3751 a_11338_19178# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3752 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3753 VDPWR a_10227_23490# sar9b_0.net53 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X3754 sar9b_0.net63 a_6861_22828# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.194 ps=1.475 w=1.12 l=0.15
X3755 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3756 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3757 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3758 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3759 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3760 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3761 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3762 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3763 a_5761_19487# sar9b_0._07_ sar9b_0._10_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X3764 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3765 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3766 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3767 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3768 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X3769 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3770 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3771 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3772 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3773 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3774 a_49926_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3775 VDPWR a_6252_19074# sar9b_0.net55 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3776 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3777 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3778 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3779 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3780 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3781 a_8266_17113# a_8057_17131# a_7602_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3783 VDPWR a_9323_28371# single_9b_cdac_0.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3784 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3785 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3787 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3788 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A a_40321_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3789 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3790 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3791 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3792 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3793 VGND sar9b_0.net52 a_10806_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3794 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3795 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3796 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3797 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3798 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3799 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3800 a_9130_26198# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3801 VDPWR a_12870_22267# a_12820_22557# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3802 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3803 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3804 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3805 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3806 VGND sar9b_0.net7 a_11859_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3807 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3808 VDPWR a_13011_25902# single_9b_cdac_1.CF[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3809 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3811 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3812 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3813 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3814 VDPWR a_13011_20574# single_9b_cdac_1.CF[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3815 a_9261_17906# sar9b_0.net6 a_9174_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3816 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3817 a_10470_21795# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3818 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3819 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3820 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3821 a_2706_26108# a_3156_26115# a_3108_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3822 a_9442_21474# a_9258_21842# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3823 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3824 VGND a_6880_17491# sar9b_0.net5 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3826 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3827 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3828 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3829 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3830 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3831 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3832 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3833 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3834 a_10806_24866# a_10742_25087# a_10728_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3835 a_8982_21902# sar9b_0.net8 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3836 a_5628_19768# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X3837 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3838 VDPWR single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3839 VGND a_10995_28566# uo_out[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3840 a_5506_26802# a_5322_27170# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3841 a_11382_23474# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3842 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3843 a_8512_27801# a_7914_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3844 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3845 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3846 a_10742_27751# a_10607_27849# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3847 VGND a_6414_23681# a_6346_23773# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3848 VDPWR a_12618_23470# a_12870_23599# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3849 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3850 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3851 single_9b_cdac_0.SW[1] a_13011_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3852 a_5441_22522# a_5289_22527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X3853 single_9b_cdac_1.SW[5] a_13011_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3854 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3856 sar9b_0.net23 a_7692_26108# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3857 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3858 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3859 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3860 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3861 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3862 VDPWR sar9b_0.net23 a_9939_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3863 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3864 VGND a_4922_20857# sar9b_0._18_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X3865 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3866 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3867 a_3108_26141# a_2847_26141# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3868 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3869 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3870 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3871 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3872 VGND a_4236_21738# sar9b_0.net67 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3873 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3874 a_7343_27849# a_7138_27758# a_6678_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3875 a_8098_23762# a_7914_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3876 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3877 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3878 VGND sar9b_0.net52 a_11469_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3879 a_10728_24866# a_10402_25094# a_10607_25185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3880 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3881 VGND a_8019_17910# single_9b_cdac_1.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3882 VGND sar9b_0.net49 a_10227_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3884 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3885 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3886 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3887 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.th_sw_main_0.VGS ua[4] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X3888 uio_out[0] a_4083_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3889 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3890 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3891 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3892 a_3855_25792# a_4136_25584# a_4091_25468# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.09975 ps=0.895 w=0.42 l=0.15
X3893 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3894 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3895 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3896 a_9165_24988# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.2102 ps=1.505 w=1 l=0.15
X3897 VGND a_4018_24235# a_3976_24520# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X3898 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3899 a_6132_23451# sar9b_0.net57 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3900 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3901 a_8842_18206# a_8057_18463# a_8334_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3902 single_9b_cdac_1.SW[4] a_11859_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3903 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3904 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3905 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3906 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3907 VGND a_9138_27163# a_8940_27039# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3908 a_12618_23470# a_11658_23470# a_12182_23755# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3909 VGND a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.2109 ps=2.05 w=0.74 l=0.15
X3910 a_8874_23470# a_8098_23762# a_8438_23755# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3911 a_8386_22806# a_8202_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3912 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3913 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3914 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3915 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3916 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3917 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3918 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3919 single_9b_cdac_1.CF[1] a_12435_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3920 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3921 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3922 VGND sar9b_0._07_ a_5523_21528# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.22412 pd=1.365 as=0.15675 ps=1.67 w=0.55 l=0.15
X3923 VDPWR a_9782_21622# a_9737_21523# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3924 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3925 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3926 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3928 a_11469_26138# sar9b_0.net74 a_11382_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3929 a_11146_25483# a_10937_25582# a_10482_25831# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3930 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3931 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3932 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3933 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3935 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3936 VGND a_2706_26108# a_2508_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3937 VGND a_6252_20780# sar9b_0._01_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3938 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3939 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3940 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3941 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3942 a_6030_24396# a_5748_24381# a_6391_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3943 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3944 a_3231_27227# a_3090_27163# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X3945 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3946 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3947 sar9b_0._17_ sar9b_0.net63 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2352 ps=1.54 w=1.12 l=0.15
X3948 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3949 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3950 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3952 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3953 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3954 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3955 a_9930_20510# a_8970_20510# a_9494_20290# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3956 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3957 tdc_0.RDY tdc_0.phase_detector_0.pd_out_0.B a_16542_13134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X3958 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3959 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3960 VDPWR sar9b_0.net54 a_10227_23490# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X3961 sar9b_0.net10 a_6636_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X3962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3964 VDPWR a_8166_27595# a_8116_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3965 VDPWR sar9b_0.net52 a_9942_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3966 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3967 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3968 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3969 VGND a_10926_17021# a_10858_17113# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3970 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3971 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3972 a_2847_27473# a_2706_27440# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X3973 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3974 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3975 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3976 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3977 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3978 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_4947_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3979 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3980 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X3981 VGND a_13011_25902# single_9b_cdac_1.CF[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3983 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3984 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3985 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3986 VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# dw_17224_1400# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X3987 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3988 a_8438_23755# a_8303_23853# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3989 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3990 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3991 VDPWR a_5581_20992# sar9b_0._09_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.3304 ps=2.83 w=1.12 l=0.15
X3992 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3993 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3994 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3995 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3996 a_10800_17903# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3997 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3999 VGND a_11430_27595# a_11388_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4000 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4001 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4002 VGND sar9b_0.net6 a_12435_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4003 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4004 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4005 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4006 VGND sar9b_0.net53 a_9357_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4007 sar9b_0.net74 a_10707_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4008 a_7306_19777# a_7097_19795# a_6642_19448# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4009 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4010 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4011 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4012 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4013 VDPWR a_9323_28371# single_9b_cdac_0.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4014 VDPWR sar9b_0.net58 a_4467_24162# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X4015 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4016 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4017 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4018 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4019 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4020 sar9b_0.net59 a_3603_28156# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X4021 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4022 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4023 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4024 VDPWR a_9939_28566# uo_out[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4025 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4026 VGND a_13216_18477# sar9b_0.net28 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4027 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4028 sar9b_0.net43 a_5100_24375# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4029 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4030 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4031 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4032 a_3438_27677# a_3161_27787# a_3768_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4033 sar9b_0._07_ a_3371_23106# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.11312 ps=1.065 w=0.74 l=0.15
X4034 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4035 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4036 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4037 a_11388_27473# a_10218_27466# a_11178_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4038 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4039 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4040 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4041 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INN a_15400_11316# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4042 VGND sar9b_0.net58 a_5238_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4043 VDPWR a_10995_28566# uo_out[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4044 a_9357_24566# sar9b_0.net62 a_9270_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4045 VDPWR a_8019_17910# single_9b_cdac_1.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4046 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4047 a_8052_18123# sar9b_0.net56 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4048 a_10859_26330# sar9b_0.net33 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X4049 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4050 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4051 VDPWR a_7347_24160# sar9b_0.net54 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X4052 VGND sar9b_0.net53 a_10317_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4053 a_6088_20524# a_4947_20140# a_5931_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X4054 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4055 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4056 VDPWR sar9b_0.net10 a_6922_23534# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4057 sar9b_0._04_ sar9b_0.net69 a_2540_22432# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X4058 a_5535_18149# a_5394_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4059 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4060 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4061 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4062 a_9802_26815# a_9588_27045# a_9138_27163# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4063 a_6030_24396# a_5753_24250# a_6360_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4064 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4065 single_9b_cdac_1.CF[3] a_13011_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4066 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4067 a_3768_27530# a_3370_27769# a_3690_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4068 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4069 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4070 a_9359_20191# a_8970_20510# a_8694_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4071 a_12246_19538# a_12182_19759# a_12168_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4072 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4073 a_11915_28371# sar9b_0.net14 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X4074 a_5748_24381# sar9b_0.net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4075 VGND a_2603_17006# th_dif_sw_0.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4076 a_4886_21124# sar9b_0.net65 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4077 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4078 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4079 a_3991_19768# sar9b_0._07_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.4075 pd=1.815 as=0.1853 ps=1.385 w=1 l=0.15
X4080 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4081 VDPWR a_3180_19448# sar9b_0._00_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4082 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4083 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4084 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4086 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4087 a_10506_24506# a_9730_24138# a_10070_24286# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4088 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4089 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4090 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4091 VDPWR a_11339_27039# single_9b_cdac_0.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4092 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4093 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4094 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4095 a_12560_27128# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X4096 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X4097 a_10317_23234# sar9b_0.net74 a_10230_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4098 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4099 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4100 VDPWR single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4101 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4102 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4103 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4104 a_10194_16784# a_10644_16791# a_10596_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X4105 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4106 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4107 VDPWR a_5460_28377# a_5465_28246# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4108 a_12168_19538# a_11842_19766# a_12047_19857# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4109 VGND sar9b_0.net23 a_9939_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4110 uo_out[1] a_12531_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4111 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4112 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4113 a_10029_27470# sar9b_0.net43 a_9942_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4114 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4115 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4116 a_10326_19235# a_10098_19171# a_10239_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X4117 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4118 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4119 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4120 uo_out[2] a_10995_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4121 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4122 single_9b_cdac_1.CF[6] a_13011_24570# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4123 a_16970_11404# tdc_0.phase_detector_0.INP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X4124 VDPWR a_4083_28566# uio_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4125 VDPWR sar9b_0.net55 a_5811_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X4126 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4127 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4128 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4129 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4130 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4131 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4132 VGND sar9b_0.net8 a_13011_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4133 a_10596_16817# a_10335_16817# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4134 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4135 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4136 a_3731_22165# a_3206_22432# a_3561_22527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X4137 single_9b_cdac_1.CF[2] a_11859_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4138 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4139 a_10200_27170# a_9802_26815# a_10122_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4140 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4141 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4142 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4143 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4144 a_7735_19857# a_7306_19777# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4145 VDPWR a_7539_28566# uo_out[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4146 a_8438_18958# a_8303_18859# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4147 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4148 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4149 VGND sar9b_0.net27 a_13011_27234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4150 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4151 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4152 a_5832_17846# a_5506_17478# a_5711_17527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4153 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4154 a_7914_27466# a_6954_27466# a_7478_27751# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4155 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] a_65367_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4156 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4157 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4158 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4159 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4160 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4161 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4162 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4163 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4164 VGND sar9b_0.net52 a_7725_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4165 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4166 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4167 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4168 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4169 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4170 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4171 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4172 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4173 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4174 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4175 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4176 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4177 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4178 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4179 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4180 VDPWR a_11430_24931# a_11380_25221# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4181 single_9b_cdac_1.SW[1] a_10803_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4182 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4183 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4184 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4185 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4186 VDPWR a_12870_19603# a_12820_19893# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4187 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4188 a_10122_27170# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4189 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4190 VGND sar9b_0._10_ a_4583_20468# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X4191 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4192 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4194 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4195 a_5711_26851# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4196 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4197 VGND a_5460_28377# a_5465_28246# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4198 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4199 a_10896_24563# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4200 a_7725_23474# sar9b_0.net11 a_7638_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4201 VGND a_11859_21906# single_9b_cdac_1.CF[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4202 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4203 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4204 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4205 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4206 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4207 a_5298_24499# a_5753_24250# a_5702_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X4208 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4210 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4211 a_12820_18561# a_11842_18434# a_12618_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4212 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4213 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4214 VDPWR a_3922_20239# a_3830_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4215 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4216 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4217 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4218 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4219 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4220 a_6634_18206# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4221 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4222 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4223 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4224 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4225 VGND sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X4226 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4227 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4228 a_10762_18823# a_10553_18922# a_10098_19171# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4229 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4230 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4231 a_3561_22527# a_3206_22432# a_3454_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X4232 a_10662_17799# a_10410_17846# a_10800_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4235 a_4749_27652# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.2102 ps=1.505 w=1 l=0.15
X4236 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4237 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4238 a_9494_20290# a_9359_20191# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4239 VDPWR a_13011_17910# single_9b_cdac_1.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4240 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4241 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4242 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4243 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4244 VGND sar9b_0.net60 a_7542_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4245 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4246 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4247 VGND sar9b_0.net12 a_11658_26134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4248 single_9b_cdac_1.CF[6] a_13011_24570# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4249 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4250 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4251 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4252 sar9b_0.net60 a_2547_28132# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4253 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4254 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4255 a_10218_21842# a_9442_21474# a_9782_21622# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4256 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4257 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4258 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A a_64331_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4259 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4260 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4261 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4262 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4263 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4264 a_10038_17846# a_9974_17626# a_9960_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4266 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4267 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4268 a_5674_28147# a_5465_28246# a_5010_28495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4269 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4270 a_7743_16817# a_7602_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4271 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4272 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4273 a_3946_26198# a_3161_26455# a_3438_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4274 a_8591_22855# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4275 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4276 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4277 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4278 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4279 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4280 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1295 ps=1.09 w=0.74 l=0.15
X4281 a_16881_10256# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16527_10454# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4282 a_12246_23534# a_12182_23755# a_12168_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4283 sar9b_0.net27 a_5196_18116# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4284 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4285 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4286 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4287 VDPWR a_7188_22119# a_7193_22459# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4288 a_13216_18477# a_12618_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4290 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4291 a_21684_3438# th_dif_sw_0.th_sw_1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X4292 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4293 a_3380_20145# a_2739_20140# a_3273_20185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X4294 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4295 a_8116_27885# a_7138_27758# a_7914_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4296 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4297 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4298 a_7800_22202# a_7402_22441# a_7722_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4299 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4300 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4301 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4302 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4303 a_12182_26419# a_12047_26517# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4304 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4305 a_11718_23127# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4306 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4307 VGND clk a_16881_10256# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X4308 VDPWR a_7470_22349# a_7402_22441# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4309 a_5374_20145# sar9b_0._01_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X4310 VDPWR sar9b_0.net49 a_10035_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4312 sar9b_0.net20 a_4812_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4313 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4314 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4315 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4316 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4317 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4318 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4319 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4320 single_9b_cdac_1.SW[8] a_11859_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4321 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4322 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4323 VGND a_2547_28132# sar9b_0.net60 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4324 VDPWR a_6130_20239# a_6038_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4325 a_12168_23534# a_11842_23762# a_12047_23853# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4326 VDPWR a_7404_17715# sar9b_0.net73 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4328 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4329 sar9b_0.net17 a_2508_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4330 a_54737_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4331 VGND a_5235_27466# uo_out[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4332 a_10231_26851# a_9802_26815# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4333 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] a_36555_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4334 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4335 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4336 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4337 VDPWR sar9b_0.net47 a_7470_22349# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4338 a_7722_22202# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4339 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4340 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4341 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4342 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4343 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4344 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4345 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4346 VGND a_13011_16810# single_9b_cdac_1.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4347 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4348 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4349 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4350 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4351 a_6738_22112# a_7188_22119# a_7140_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X4352 sar9b_0._18_ a_4922_20857# a_5083_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X4353 a_9359_20191# a_9154_20142# a_8694_20570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4354 VDPWR sar9b_0.net46 a_8334_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4355 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4356 VDPWR a_9588_27045# a_9593_26914# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4357 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4358 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4359 a_4091_25468# a_3747_25724# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1239 ps=1.43 w=0.42 l=0.15
X4360 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4361 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4362 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4363 a_12137_19857# a_11658_19474# a_12047_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4364 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4365 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4366 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4367 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4368 VGND a_11430_24931# a_11388_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4369 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4370 VDPWR a_10644_16791# a_10649_17131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4371 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4372 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4373 single_9b_cdac_1.SW[6] a_13011_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4374 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4375 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4376 VDPWR a_12531_28566# uo_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4377 VDPWR a_5846_26950# a_5801_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4378 VDPWR a_8052_16791# a_8057_17131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4379 a_3946_26198# a_3156_26115# a_3438_26345# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4381 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4382 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4383 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4384 VDPWR sar9b_0.net53 a_10230_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4385 VGND sar9b_0.net48 a_10326_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4386 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4387 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4388 sar9b_0.clk_div_0.COUNT\[2\] a_4018_24235# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X4389 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4390 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4391 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4392 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A a_60565_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4393 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4394 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4396 a_5910_27170# a_5846_26950# a_5832_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4397 VGND sar9b_0.clknet_0_CLK a_2508_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4398 a_9126_19131# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4399 VDPWR tdc_0.RDY a_5331_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4400 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4401 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4402 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4403 a_50962_15501# single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4404 a_3494_26815# a_3231_27227# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4405 VDPWR a_9472_23805# sar9b_0.net12 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4406 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4407 VDPWR a_10742_25087# a_10697_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4408 a_11388_24809# a_10218_24802# a_11178_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4409 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4410 a_16527_10454# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X4411 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4412 a_4072_19474# sar9b_0.net71 a_3991_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.4075 ps=1.815 w=1 l=0.15
X4413 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4414 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4415 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4416 VGND a_2892_23070# sar9b_0.net66 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4417 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4418 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4419 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4420 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4421 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4422 VGND sar9b_0.net44 a_5322_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4423 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4424 a_4330_27170# sar9b_0.net37 a_4851_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4425 VGND a_3795_19512# a_4211_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.20905 pd=1.305 as=0.2997 ps=1.55 w=0.74 l=0.15
X4426 VGND a_9870_27060# a_9802_26815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X4427 VDPWR sar9b_0.net9 a_8074_20870# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4428 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4429 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4430 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4431 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4432 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4433 VDPWR sar9b_0.net40 a_13011_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4434 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4435 VDPWR a_8726_22954# a_8681_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4436 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4437 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4438 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4439 a_10697_25185# a_10218_24802# a_10607_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4440 a_8303_18859# a_8098_18810# a_7638_19238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4441 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4442 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4443 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A a_15052_11404# VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X4444 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4445 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4446 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4447 a_12588_16784# tdc_0.OUTP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4448 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4449 a_6880_26815# a_6282_27170# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4450 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4451 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4454 VGND a_13067_27662# single_9b_cdac_0.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4455 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4456 a_8790_23174# a_8726_22954# a_8712_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4457 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4458 a_10607_25185# a_10218_24802# a_9942_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4459 VDPWR a_10758_24459# a_10708_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4460 VGND a_6738_22112# a_6540_22112# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4461 VDPWR a_13011_21906# single_9b_cdac_1.CF[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4462 VDPWR tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4463 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4464 a_5846_26950# a_5711_26851# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4465 a_3364_25120# sar9b_0._14_ a_2893_24992# VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4466 a_10758_24459# a_10506_24506# a_10896_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4467 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4468 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4469 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4470 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4471 tdc_0.OUTP tdc_0.OUTN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4472 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4473 VGND a_6132_23451# a_6137_23791# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4474 VGND clk a_4332_23043# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4475 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4476 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4477 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4478 VGND sar9b_0.net11 a_8202_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4479 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4480 a_10029_24806# sar9b_0.net12 a_9942_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4481 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4482 VGND a_13164_28398# sar9b_0.net14 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4483 a_8712_23174# a_8386_22806# a_8591_22855# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4484 VDPWR sar9b_0.net6 a_12435_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4485 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4486 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4487 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4488 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4489 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4490 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4491 a_13216_22473# a_12618_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4492 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4493 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4494 sar9b_0.net15 a_6130_20239# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X4495 a_3946_27530# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4496 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4497 a_2934_26141# a_2706_26108# a_2847_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X4498 a_8031_26141# a_7890_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4499 VDPWR a_9165_24988# sar9b_0.net52 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X4500 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4501 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4502 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4503 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4504 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4505 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4506 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP a_16222_11316# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4507 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4508 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4509 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4510 a_9760_22819# a_9162_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4511 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4512 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4513 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4514 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4515 VGND a_7602_16784# a_7404_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4516 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4517 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4518 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4519 VGND a_10035_19474# sar9b_0.net48 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4520 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4521 a_6346_23773# a_6137_23791# a_5682_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4522 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4523 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4524 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4525 a_55773_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4526 VDPWR sar9b_0.net55 a_7347_24160# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X4527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4528 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4529 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4530 VGND sar9b_0.net57 a_7914_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4531 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4532 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4533 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4534 VGND a_10182_20463# a_10140_20567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4535 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A a_31753_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4536 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4537 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4538 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4539 VDPWR a_5748_24381# a_5753_24250# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4540 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4541 a_30717_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4542 a_4332_23043# clk VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4543 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4544 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4545 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4546 sar9b_0.net45 a_8883_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4547 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4548 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4549 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4550 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4551 a_12137_23853# a_11658_23470# a_12047_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4552 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4553 VGND sar9b_0.net47 a_6966_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4554 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4555 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4556 a_11776_27801# a_11178_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4557 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4558 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4559 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4560 VGND a_10932_25713# a_10937_25582# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4561 a_2508_20780# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4562 sar9b_0.net40 a_6444_19448# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4563 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4564 single_9b_cdac_0.SW[3] a_12491_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X4565 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4567 VDPWR sar9b_0.net1 a_10707_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4568 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4570 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4571 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4572 a_8438_23755# a_8303_23853# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4573 VDPWR sar9b_0.net50 a_11382_19478# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4574 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4575 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4576 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4577 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4578 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4579 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4580 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4581 VGND sar9b_0.net59 a_10029_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4582 a_46159_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4583 VGND a_7936_25137# sar9b_0.cyclic_flag_0.FINAL VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4584 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4585 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4586 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4587 VGND sar9b_0.net54 a_10227_23490# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X4588 a_49926_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4589 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4590 single_9b_cdac_1.CF[4] a_13011_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4591 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4592 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4593 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4594 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4595 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4596 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4597 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4598 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4599 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4600 a_11430_27595# a_11178_27466# a_11568_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4601 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4602 uo_out[0] a_11915_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4603 a_4330_27170# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4604 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4605 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4606 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4607 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4609 VDPWR sar9b_0.net53 a_9270_24566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4610 a_5196_19448# sar9b_0.net16 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4611 VGND a_11436_17742# sar9b_0.net61 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4612 a_12618_22138# a_11842_22430# a_12182_22423# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4613 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4614 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4615 a_3014_24136# a_2835_24136# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4616 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4617 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4618 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4619 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4620 VDPWR sar9b_0.net8 a_13011_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4621 VDPWR a_10803_18142# single_9b_cdac_1.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4622 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4623 a_6414_23681# a_6132_23451# a_6775_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X4624 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4625 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4626 VDPWR a_11915_28371# uo_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4627 VGND a_5748_24381# a_5753_24250# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4628 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4629 single_9b_cdac_0.SW[4] a_11915_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4630 VGND a_5235_27466# uo_out[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4631 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4632 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4633 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4634 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4635 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4637 a_9165_24988# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X4638 VDPWR sar9b_0.net57 a_10218_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4639 a_7044_19481# a_6783_19481# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4640 VGND a_13011_16810# single_9b_cdac_1.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4641 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4642 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4643 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4644 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4645 VGND a_7443_21496# sar9b_0.net47 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4646 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4647 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4648 VGND a_7566_21017# a_7498_21109# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X4649 VGND sar9b_0.net51 a_6579_18832# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X4650 a_12047_18525# a_11842_18434# a_11382_18146# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4651 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4652 VGND a_5580_24776# sar9b_0._03_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4653 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4654 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4655 VGND a_6444_21738# sar9b_0.net64 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4656 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4657 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4658 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4659 a_3830_20140# a_2918_20140# a_3723_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X4660 VDPWR a_10035_19474# sar9b_0.net48 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4661 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4662 a_12047_19857# a_11658_19474# a_11382_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4663 VGND a_11008_17491# sar9b_0.net7 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4664 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4665 a_6775_23853# a_6346_23773# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4666 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4667 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4668 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4670 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4671 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4672 a_10378_27170# a_9593_26914# a_9870_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4673 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4676 a_11178_24802# a_10402_25094# a_10742_25087# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4677 a_3369_24181# a_3014_24136# a_3262_24141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X4678 a_5823_23477# a_5682_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4679 sar9b_0._08_ a_4072_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2557 ps=1.59 w=1.12 l=0.15
X4680 VDPWR sar9b_0.net11 a_13011_24570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4681 a_11178_20806# a_10218_20806# a_10742_21091# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4682 VDPWR sar9b_0.net61 a_11338_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4683 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4684 VDPWR a_6030_24396# a_5962_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4685 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4686 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4687 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4688 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4689 uo_out[0] a_11915_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X4690 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4691 a_6672_17903# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4692 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4693 VDPWR a_3695_23038# a_3371_23106# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.147 ps=1.19 w=0.84 l=0.15
X4694 a_7284_20787# sar9b_0.net56 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4695 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4696 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4697 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4698 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4699 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4700 a_10644_16791# sar9b_0.net6 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4701 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4702 single_9b_cdac_0.SW[2] a_13067_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X4703 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4704 VGND a_4812_21738# sar9b_0.net65 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4705 a_5711_17527# a_5322_17846# a_5046_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4706 a_11722_25838# sar9b_0.net74 a_12243_25898# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4707 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4708 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4709 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4710 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4711 VGND a_11859_20574# single_9b_cdac_1.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4712 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4713 a_4561_24464# sar9b_0.net58 a_4467_24162# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1312 pd=1.05 as=0.1824 ps=1.85 w=0.64 l=0.15
X4714 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4715 VGND sar9b_0.clknet_0_CLK a_2508_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4716 a_10500_19235# a_10239_19235# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4717 VGND sar9b_0.net38 a_10803_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4718 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4719 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4720 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4721 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4722 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4723 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4724 a_5581_19664# sar9b_0._07_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X4725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4726 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4727 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4728 a_10402_25094# a_10218_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4729 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4730 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4731 tdc_0.phase_detector_0.INN a_16527_10454# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X4732 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4733 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4734 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4735 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4736 VDPWR sar9b_0.net41 a_9130_26198# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4737 VGND a_5298_24499# a_5100_24375# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4738 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4739 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4740 single_9b_cdac_1.CF[8] a_13011_25902# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4741 VGND sar9b_0.net5 a_13011_20574# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4742 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4743 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4744 single_9b_cdac_1.CF[0] a_13011_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4746 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4747 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4748 VDPWR a_10218_21842# a_10470_21795# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X4749 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4750 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4751 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4752 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4753 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4754 VDPWR a_11776_21141# sar9b_0.net8 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4755 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4756 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4757 a_10708_24151# a_9730_24138# a_10506_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4758 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4759 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4760 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4761 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4762 VDPWR a_6132_23451# a_6137_23791# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4763 a_2603_17006# sar9b_0.net16 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X4764 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4765 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4766 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4767 a_3521_24240# a_3369_24181# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X4768 a_16542_13134# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X4769 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4770 VDPWR sar9b_0.net53 a_11382_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4771 VDPWR sar9b_0.net49 a_8982_21902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4772 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4773 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4774 a_6744_23534# a_6346_23773# a_6666_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4775 a_12870_23599# a_12618_23470# a_13008_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4776 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4777 VDPWR a_6414_23681# a_6346_23773# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4778 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4779 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4780 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4781 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4782 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4783 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4784 VDPWR a_13011_27234# single_9b_cdac_0.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4785 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4786 a_9264_23477# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4787 a_4168_22188# a_3027_22138# a_4011_22488# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X4788 VDPWR a_13011_16810# single_9b_cdac_1.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4789 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4790 a_41357_15501# single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4792 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4793 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4794 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4795 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4796 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4797 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4798 a_11191_18859# a_10762_18823# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4799 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4800 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4801 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4802 a_8554_26437# a_8340_26115# a_7890_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4803 VDPWR sar9b_0.net5 a_7914_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4804 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4805 VGND sar9b_0.net3 a_2547_28132# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4806 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4807 a_7433_27849# a_6954_27466# a_7343_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4808 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4809 a_8098_18810# a_7914_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4810 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4812 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4813 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4814 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4815 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4816 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4817 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4818 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4819 a_6666_23534# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4820 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4821 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4822 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4823 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4824 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4825 VGND a_10035_19474# sar9b_0.net48 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4826 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4827 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4828 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4829 a_3370_26437# a_3156_26115# a_2706_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4830 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4831 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4832 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4833 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4834 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4835 VGND a_4365_25770# a_4293_25852# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.10905 ps=1.025 w=0.55 l=0.15
X4836 a_3372_25734# sar9b_0._16_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4837 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4838 single_9b_cdac_1.CF[3] a_13011_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4839 VDPWR a_11915_28371# uo_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4840 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4841 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4842 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4843 VGND a_9760_22819# sar9b_0.net41 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4844 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4845 a_7238_21225# a_6975_20813# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4846 a_5633_20244# a_5481_20185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X4847 a_7743_18149# a_7602_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4848 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4849 a_12647_27128# sar9b_0.net52 a_12560_27128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4850 VDPWR a_12435_20806# single_9b_cdac_1.CF[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4851 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4852 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4853 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4854 a_12870_22267# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4856 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4857 single_9b_cdac_0.SW[1] a_13011_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4858 single_9b_cdac_1.SW[7] a_13011_19242# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4859 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4860 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4861 VGND a_5010_28495# a_4812_28371# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4862 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4863 a_12047_22521# a_11842_22430# a_11382_22142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4864 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4865 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4867 VGND a_12870_23599# a_12828_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4868 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4869 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4870 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4871 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4872 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4874 a_6538_24506# a_5753_24250# a_6030_24396# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4875 a_12047_23853# a_11658_23470# a_11382_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4876 VDPWR a_6738_22112# a_6540_22112# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X4877 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4878 single_9b_cdac_0.SW[3] a_12491_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X4879 VDPWR sar9b_0.net58 a_3231_27227# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4880 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4881 a_8940_24402# sar9b_0.net2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4882 a_12064_22819# a_11466_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4884 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4885 a_3372_25734# sar9b_0._16_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4886 VDPWR sar9b_0.clk_div_0.COUNT\[2\] sar9b_0._17_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.42 pd=2.99 as=0.168 ps=1.42 w=1.12 l=0.15
X4887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4888 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4889 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4890 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4891 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4892 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4893 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4895 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4896 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X4897 VGND a_10859_26330# single_9b_cdac_0.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4898 VGND a_3090_27163# a_2892_27039# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4899 a_10320_20567# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4900 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4901 a_5083_21100# sar9b_0._17_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X4902 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4903 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4904 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4905 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4906 sar9b_0.net18 a_2508_27440# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4907 VDPWR sar9b_0.net58 a_2847_27473# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4908 sar9b_0.net3 a_2451_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4909 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4910 VDPWR a_4044_24776# sar9b_0.net72 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4911 a_12828_23477# a_11658_23470# a_12618_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4912 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4913 th_dif_sw_0.CK a_10227_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4914 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4915 uo_out[6] a_8115_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4916 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4917 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4918 VDPWR a_12182_26419# a_12137_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4919 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4920 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4921 a_3438_26345# a_3161_26455# a_3768_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4922 a_2540_22432# sar9b_0._12_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X4923 a_7140_22145# a_6879_22145# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4924 a_10239_19235# a_10098_19171# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4925 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4926 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4927 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4928 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4929 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4930 a_8294_26553# a_8031_26141# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4931 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4932 a_2706_27440# a_3161_27787# a_3110_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X4933 a_5580_24776# sar9b_0._15_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4934 a_8842_16874# a_8052_16791# a_8334_17021# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4935 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4936 single_9b_cdac_0.SW[6] a_9323_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4937 VGND sar9b_0.net52 a_10029_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4938 a_12618_18142# a_11658_18142# a_12182_18427# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4939 a_6534_17799# a_6282_17846# a_6672_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4940 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4941 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4942 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4943 uio_out[1] a_2931_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4944 a_4749_27652# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X4945 a_13008_26141# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4946 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4947 VDPWR a_3603_28156# sar9b_0.net59 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X4948 VDPWR a_5938_22378# a_5846_22572# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4949 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4950 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4951 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4952 VDPWR sar9b_0.net48 a_10830_19068# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4953 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4954 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4955 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4956 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4957 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4958 a_11430_24931# a_11178_24802# a_11568_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4959 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4960 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4961 a_3110_26553# a_2847_26141# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4962 a_3768_26198# a_3370_26437# a_3690_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4963 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4964 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4965 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4966 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4967 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4968 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4969 VGND sar9b_0.net24 a_10995_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4970 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4971 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4972 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4973 a_3262_24141# sar9b_0.net70 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X4974 VGND sar9b_0.net49 a_9558_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4975 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4976 uo_out[2] a_10995_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4977 single_9b_cdac_1.SW[2] a_8019_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4978 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4979 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4980 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4981 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4982 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4983 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4984 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4985 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4986 a_4851_27230# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4987 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4988 VGND a_5441_22522# a_5459_22165# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X4989 sar9b_0.net36 a_9996_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4990 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4992 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4993 VDPWR sar9b_0.net48 a_5535_18149# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4994 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4995 a_10742_25087# a_10607_25185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4996 a_12618_19474# a_11842_19766# a_12182_19759# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4997 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4998 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4999 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5000 single_9b_cdac_1.SW[8] a_11859_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5001 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5002 VDPWR a_13011_20806# single_9b_cdac_1.CF[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5003 a_8166_27595# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5004 a_6966_22145# a_6738_22112# a_6879_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5005 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5006 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5007 a_11915_27039# sar9b_0.net30 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X5008 a_9558_20510# a_9494_20290# a_9480_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5009 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5010 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5011 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5012 a_4771_18260# sar9b_0.net57 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X5013 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5014 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5015 a_11568_20813# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5016 a_8842_18206# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5017 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5018 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5019 a_9730_24138# a_9546_24506# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5020 single_9b_cdac_1.CF[1] a_12435_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5021 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5022 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.11655 ps=1.055 w=0.74 l=0.15
X5023 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5024 single_9b_cdac_0.SW[2] a_13067_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5025 single_9b_cdac_0.SW[5] a_11339_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5026 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5027 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5028 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5030 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5031 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5032 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5033 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5034 a_10410_17846# a_9450_17846# a_9974_17626# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5035 a_9126_23599# a_8874_23470# a_9264_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5036 a_8591_22855# a_8202_23174# a_7926_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5037 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5039 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5040 a_5674_28147# a_5460_28377# a_5010_28495# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5041 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5042 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5043 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5044 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5045 a_5460_28377# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5046 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5047 a_8098_18810# a_7914_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5048 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5049 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5050 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5051 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5052 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5054 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5055 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5056 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5057 VGND single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5058 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5059 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5060 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5061 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5062 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5063 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5064 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5065 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5066 VDPWR a_13011_24570# single_9b_cdac_1.CF[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5067 single_9b_cdac_1.CF[5] a_13011_23238# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5068 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5069 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5070 a_5846_17626# a_5711_17527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5071 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5072 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5074 VGND sar9b_0.clk_div_0.COUNT\[2\] a_7597_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5075 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5076 a_7306_19777# a_7092_19455# a_6642_19448# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5077 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5078 sar9b_0.net11 a_5484_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5079 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5080 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5081 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5082 a_9359_20191# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5083 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5084 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5086 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5087 VDPWR a_3090_27163# a_2892_27039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X5088 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5089 VGND a_9323_28371# single_9b_cdac_0.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X5090 a_11915_28371# sar9b_0.net14 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X5091 uo_out[5] a_7539_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5092 a_10378_27170# a_9588_27045# a_9870_27060# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5093 a_11466_23174# a_10506_23174# a_11030_22954# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5094 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5095 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5096 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5097 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5098 VGND sar9b_0.net13 a_13011_25902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5099 VDPWR a_12618_22138# a_12870_22267# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5100 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5101 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5102 a_8074_20870# sar9b_0.net9 a_8595_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5103 a_10335_16817# a_10194_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5104 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5105 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5106 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5108 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5109 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5110 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5111 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5112 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5113 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5114 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5115 a_7597_23174# sar9b_0.net63 a_7483_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X5116 a_9647_21523# a_9442_21474# a_8982_21902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5117 a_10140_20567# a_8970_20510# a_9930_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5118 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5119 a_10070_24286# a_9935_24187# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5120 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5121 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5122 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5123 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5124 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5125 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5126 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5127 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5128 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5129 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5130 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5131 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5132 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5133 VDPWR sar9b_0.net60 a_3603_28156# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X5134 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5135 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5136 VGND sar9b_0.net55 a_7347_24160# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X5137 VGND sar9b_0.net49 a_9846_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5138 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5139 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5140 sar9b_0.net58 a_4749_27652# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.756 ps=3.59 w=1.12 l=0.15
X5141 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5142 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y a_35519_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5143 a_4673_24464# sar9b_0._13_ a_4561_24464# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.045 as=0.1312 ps=1.05 w=0.64 l=0.15
X5144 a_11856_23231# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5145 a_10182_20463# a_9930_20510# a_10320_20567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5146 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5147 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5148 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5149 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5150 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5151 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5152 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5153 a_8595_20810# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5154 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5155 a_12618_22138# a_11658_22138# a_12182_22423# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5156 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A a_26951_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5157 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5158 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5159 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5160 VDPWR sar9b_0.net73 a_6634_18206# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5161 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5162 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5163 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5164 a_25915_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5165 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5166 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X5167 single_9b_cdac_0.SW[7] a_10859_26330# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X5168 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5169 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5170 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5171 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5172 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5173 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5175 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5176 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5177 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5178 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5180 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5181 VDPWR sar9b_0.net48 a_10926_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5182 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5183 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5185 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5186 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5187 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5188 a_9442_21474# a_9258_21842# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5189 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5190 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5191 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5192 VGND a_9414_23127# a_9372_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5193 sar9b_0._05_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5194 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5195 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5196 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5197 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5198 VDPWR sar9b_0.net46 a_7743_16817# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5199 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5200 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5201 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B a_16555_12124# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5202 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5203 a_12618_23470# a_11842_23762# a_12182_23755# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5204 a_6672_27227# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5205 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5206 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5207 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5208 a_6922_23534# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5209 a_8726_22954# a_8591_22855# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5210 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5211 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5212 a_9130_26198# sar9b_0.net41 a_9651_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5213 sar9b_0._15_ a_4467_24162# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.36323 ps=1.84 w=1.12 l=0.15
X5214 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5215 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5216 a_7188_22119# sar9b_0.net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5217 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5218 a_2847_26141# a_2706_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5219 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5220 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5221 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5222 a_6058_18445# a_5844_18123# a_5394_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5224 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5225 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5226 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5227 VDPWR a_11466_23174# a_11718_23127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5228 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5229 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5230 VDPWR a_9760_22819# sar9b_0.net41 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5231 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5232 a_11430_24931# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5233 a_7978_22202# a_7188_22119# a_7470_22349# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5234 sar9b_0.net56 a_4771_18260# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5235 a_7602_16784# a_8057_17131# a_8006_17229# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5236 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5237 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5238 a_9372_23231# a_8202_23174# a_9162_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5239 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5240 single_9b_cdac_1.CF[1] a_12435_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5241 a_12870_19603# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5242 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5243 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5244 sar9b_0.net59 a_3603_28156# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X5245 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5246 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5247 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5249 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5250 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5251 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5252 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5253 a_65367_15501# single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5254 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5255 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5256 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5257 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5258 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5259 a_3371_23106# a_3219_22860# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X5260 a_9414_23127# a_9162_23174# a_9552_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5261 VDPWR sar9b_0.net8 a_11658_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5262 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5263 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5264 a_11178_27466# a_10218_27466# a_10742_27751# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5265 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5266 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5267 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5268 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X5269 VGND a_7284_20787# a_7289_21127# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X5270 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5271 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5272 a_3723_20140# a_2739_20140# a_3425_20244# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X5273 VGND a_10644_16791# a_10649_17131# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X5274 VGND sar9b_0.net47 a_5761_19487# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X5275 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5276 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5277 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5278 a_5846_26950# a_5711_26851# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5279 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5280 a_10025_24187# a_9546_24506# a_9935_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5281 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5282 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5283 a_9588_27045# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5284 a_40321_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5285 a_9449_20191# a_8970_20510# a_9359_20191# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5286 single_9b_cdac_0.SW[8] a_9323_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5287 a_9472_23805# a_8874_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5288 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5290 single_9b_cdac_1.SW[7] a_13011_19242# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5291 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5292 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5293 a_10644_16791# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5294 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5295 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5296 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5297 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5298 VGND sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X5299 VDPWR a_11008_17491# sar9b_0.net7 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5300 VDPWR a_4125_25958# a_4136_25584# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5301 a_8052_16791# sar9b_0.net5 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5302 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5303 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5304 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5305 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5306 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5307 VGND sar9b_0.net57 a_10218_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5308 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5309 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5310 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5311 uo_out[5] a_7539_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5312 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5313 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5314 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5315 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5316 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5317 VGND a_9323_28371# single_9b_cdac_0.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5318 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5319 VDPWR a_8874_19178# a_9126_19131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5320 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5321 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5322 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5323 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5324 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5325 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5326 a_12246_18206# a_12182_18427# a_12168_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5327 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5328 VGND a_5581_20992# sar9b_0._09_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.19322 pd=1.32 as=0.2109 ps=2.05 w=0.74 l=0.15
X5329 a_7498_21109# a_7289_21127# a_6834_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X5330 VDPWR a_8438_18958# a_8393_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5331 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5332 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5333 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5334 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5335 sar9b_0._02_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5336 VDPWR sar9b_0._04_ a_3027_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5337 VGND sar9b_0.net48 a_9261_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5338 a_10858_17113# a_10649_17131# a_10194_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X5339 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5340 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5341 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5342 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5344 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5345 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5346 a_8726_22954# a_8591_22855# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5347 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5348 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5349 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5350 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5352 VGND a_8115_28566# uo_out[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5353 VDPWR a_11776_27801# sar9b_0.net25 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5354 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5355 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5356 a_10410_17846# a_9634_17478# a_9974_17626# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5357 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5358 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5359 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5360 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5361 a_12168_18206# a_11842_18434# a_12047_18525# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5362 a_30717_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5363 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5364 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5365 single_9b_cdac_1.SW[1] a_10803_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5366 a_10502_18823# a_10239_19235# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5367 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5368 a_8393_18859# a_7914_19178# a_8303_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5369 VDPWR sar9b_0.net56 a_5322_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5370 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5371 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5372 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5373 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5374 a_4698_25851# a_4125_25958# a_4365_25770# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.07875 ps=0.865 w=0.42 l=0.15
X5375 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5376 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5377 VGND a_2931_28566# uio_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5378 uo_out[7] a_5235_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5380 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5381 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5382 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5383 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5384 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5385 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5386 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5387 a_3946_26198# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5388 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5389 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5390 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5391 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5392 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5393 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5394 a_60565_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5395 VDPWR sar9b_0._14_ a_2940_25096# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X5396 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5397 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5398 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5399 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5400 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5401 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5402 VGND ui_in[0] a_2451_27234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X5403 a_11339_27039# sar9b_0.net31 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X5404 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5405 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5406 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5407 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5408 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5409 a_36555_15501# single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5410 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5411 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5412 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5413 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5414 VDPWR a_4018_24235# a_3926_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X5415 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5416 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5417 VDPWR sar9b_0.net42 a_13011_19242# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5418 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5419 VDPWR sar9b_0.net36 a_3946_27530# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5420 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5421 VDPWR sar9b_0.net59 a_8031_26141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5422 single_9b_cdac_1.SW[3] a_10803_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5423 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5424 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5425 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5426 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5427 VDPWR a_12870_18271# a_12820_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X5428 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5429 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5430 VGND sar9b_0.net39 a_11859_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5431 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5432 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5433 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5434 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.B VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X5435 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5436 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5437 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5438 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5439 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5440 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5441 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5442 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5443 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5444 a_6534_27123# a_6282_27170# a_6672_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5445 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5446 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5447 single_9b_cdac_1.CF[0] a_13011_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5448 a_8874_19178# a_8098_18810# a_8438_18958# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5449 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5451 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5454 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5455 a_4236_21738# sar9b_0._05_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5456 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5457 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5458 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5459 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5460 a_7914_27466# a_7138_27758# a_7478_27751# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5461 a_6484_26815# a_5506_26802# a_6282_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5462 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5463 sar9b_0.net46 a_6579_18832# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X5464 a_3206_22432# a_3027_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5465 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5466 VDPWR sar9b_0.net11 a_11658_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5467 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5468 VGND a_13216_26469# sar9b_0.net33 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5469 a_5748_24381# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5470 VGND a_3922_20239# a_3880_20524# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X5471 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5472 VDPWR sar9b_0.net20 a_8115_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5473 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5474 VDPWR a_12618_19474# a_12870_19603# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5475 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5476 VGND sar9b_0.net53 a_10134_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5477 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5478 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5479 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5480 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5481 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5482 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5483 a_10758_24459# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5484 single_9b_cdac_1.SW[0] a_8595_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5485 VGND a_8691_28566# uo_out[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5486 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5487 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5488 a_8334_17021# a_8057_17131# a_8664_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5489 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5490 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5491 VDPWR sar9b_0.clknet_0_CLK a_2508_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5492 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5493 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5494 a_3839_23194# sar9b_0.clk_div_0.COUNT\[2\] a_3725_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.1344 ps=1.06 w=0.64 l=0.15
X5495 sar9b_0.net6 a_7404_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5496 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5497 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5498 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5499 VGND single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5500 VGND a_7539_28566# uo_out[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5501 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5502 VDPWR a_12684_20379# sar9b_0.net50 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5503 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5504 a_3454_22567# sar9b_0.net67 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X5505 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5506 VDPWR ui_in[0] a_2451_27234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5507 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5508 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5509 a_12246_22202# a_12182_22423# a_12168_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5510 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5511 a_9364_22819# a_8386_22806# a_9162_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5512 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5513 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5514 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5515 a_8664_16874# a_8266_17113# a_8586_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5516 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5517 VDPWR sar9b_0.net56 a_9450_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5518 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5519 VDPWR sar9b_0.net37 a_4330_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5520 VDPWR a_3819_24136# a_4018_24235# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X5521 VGND a_11776_21141# sar9b_0.net8 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5522 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5523 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5524 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5525 single_9b_cdac_0.SW[4] a_11915_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5526 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5527 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5528 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5529 a_31753_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5531 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5532 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5533 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5534 a_12168_22202# a_11842_22430# a_12047_22521# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5535 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5536 a_6922_23534# a_6137_23791# a_6414_23681# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X5537 a_3273_20185# a_2918_20140# a_3166_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X5538 a_5622_18149# a_5394_18116# a_5535_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5539 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5540 VDPWR a_8940_24402# sar9b_0.net62 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5541 VGND a_6130_20239# a_6088_20524# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X5542 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5543 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5544 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5545 VDPWR a_11915_27039# single_9b_cdac_0.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5546 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5547 a_8586_16874# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X5548 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5549 sar9b_0._06_ a_12560_27128# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X5550 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5551 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5552 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5553 VGND a_8595_17910# single_9b_cdac_1.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5554 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5555 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5556 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5557 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5558 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5559 a_10402_25094# a_10218_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5560 VGND sar9b_0.net12 a_9546_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5561 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5562 VGND a_5931_20140# a_6130_20239# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X5563 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5564 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5565 VGND sar9b_0.net55 a_5811_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.24915 ps=2.37 w=0.55 l=0.15
X5566 sar9b_0.clk_div_0.COUNT\[2\] a_4018_24235# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X5567 a_12137_18525# a_11658_18142# a_12047_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5568 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y a_59529_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5569 VGND a_4749_27652# sar9b_0.net58 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X5570 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5571 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5572 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5573 sar9b_0.net48 a_10035_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5574 a_3090_27163# a_3545_26914# a_3494_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5575 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5576 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5577 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5578 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5579 a_12182_19759# a_12047_19857# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5580 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5581 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5582 a_3822_27060# a_3540_27045# a_4183_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5583 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X5584 a_14897_9355# clk a_14871_9671# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5585 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5586 VDPWR sar9b_0.net54 a_5823_23477# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5587 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5588 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5589 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5590 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5591 VDPWR sar9b_0.net74 a_11722_25838# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5592 a_11436_17742# sar9b_0.net2 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5593 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5594 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5595 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5596 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5597 VDPWR sar9b_0.net10 a_13011_23238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5598 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5599 VGND a_12435_24802# single_9b_cdac_1.CF[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5600 a_6252_19074# sar9b_0.net15 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5601 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5602 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5603 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5604 a_4332_23043# clk VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X5605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5606 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5607 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5608 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5609 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5610 a_4011_22488# a_3027_22138# a_3713_22522# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X5611 a_11338_19178# sar9b_0.net61 a_11859_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5612 sar9b_0.net52 a_9165_24988# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.756 ps=3.59 w=1.12 l=0.15
X5613 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5614 a_5682_23444# a_6137_23791# a_6086_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5615 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5616 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5617 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5618 VDPWR sar9b_0.net52 a_11214_25728# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5619 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5620 uo_out[3] a_9939_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5621 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5622 a_9870_27060# a_9593_26914# a_10200_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5623 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5624 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5625 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5626 VGND a_8115_28566# uo_out[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5627 a_4183_26851# a_3754_26815# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X5628 sar9b_0.net57 a_5443_19074# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5629 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5630 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5631 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5632 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5633 a_9588_27045# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5634 a_12820_26553# a_11842_26426# a_12618_26134# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5635 a_16555_12412# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5636 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5637 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5638 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5639 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5640 VDPWR sar9b_0.net68 a_3364_25120# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5641 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5642 a_10607_27849# a_10402_27758# a_9942_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5643 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5644 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5645 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5646 VGND sar9b_0._07_ a_3795_19512# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14457 pd=1.15 as=0.15675 ps=1.67 w=0.55 l=0.15
X5647 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5648 a_7470_22349# a_7188_22119# a_7831_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5649 a_11859_19238# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5650 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5651 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5652 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5653 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5654 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5655 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5656 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5657 VGND a_2931_28566# uio_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5658 VDPWR a_13011_25902# single_9b_cdac_1.CF[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5659 a_8334_17021# a_8052_16791# a_8695_17193# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5660 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5661 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5662 VDPWR a_13011_20574# single_9b_cdac_1.CF[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5663 a_12047_19857# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5664 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5665 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5666 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5667 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5668 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5669 VDPWR sar9b_0.net46 a_5046_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X5670 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5671 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5672 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5673 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5674 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5675 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5676 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5677 a_6132_23451# sar9b_0.net57 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5678 a_6880_17491# a_6282_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5679 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5680 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5681 VDPWR single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5682 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5683 a_5394_18116# a_5849_18463# a_5798_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5684 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5685 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5686 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5687 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5688 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5689 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5690 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5691 a_13216_26469# a_12618_26134# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5692 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5693 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5694 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5695 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5696 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5697 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5698 a_8695_17193# a_8266_17113# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X5699 single_9b_cdac_1.SW[5] a_13011_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5700 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5701 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5702 single_9b_cdac_0.SW[7] a_10859_26330# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5703 a_64331_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5704 a_5133_17906# sar9b_0.net46 a_5046_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5705 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5706 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5707 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5708 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5709 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5710 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5711 VDPWR a_10070_24286# a_10025_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5712 VGND a_8019_17910# single_9b_cdac_1.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5713 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5714 VGND sar9b_0.net57 a_9258_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5716 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5717 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5718 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5719 uo_out[4] a_8691_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5720 VGND a_3425_20244# a_3443_20547# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X5721 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5722 VGND sar9b_0.net19 a_5235_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5723 a_4812_21738# sar9b_0.clk_div_0.COUNT\[3\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5724 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5726 uio_out[0] a_4083_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5727 sar9b_0.net19 a_2892_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5728 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5729 VGND a_9363_20826# sar9b_0.net49 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5730 VGND sar9b_0.net40 a_13011_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5731 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5732 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5733 single_9b_cdac_1.SW[4] a_11859_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5734 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5735 sar9b_0._16_ a_2893_24992# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X5736 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5737 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5738 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5739 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1764 ps=1.26 w=0.84 l=0.15
X5740 a_11434_16874# a_10644_16791# a_10926_17021# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5741 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5742 a_10607_25185# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5743 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5744 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5746 VGND a_13011_24802# single_9b_cdac_0.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5747 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5748 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5749 VDPWR sar9b_0.net46 a_7743_18149# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5750 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5751 VDPWR a_11915_27039# single_9b_cdac_0.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5752 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5753 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5754 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5755 single_9b_cdac_1.CF[1] a_12435_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5756 VDPWR a_3425_20244# a_3380_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X5757 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5758 VGND single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5759 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5760 a_9651_26138# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5761 a_7470_22349# a_7193_22459# a_7800_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5762 sar9b_0.net37 a_9900_19047# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5763 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5764 a_9323_28371# sar9b_0.net32 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X5765 VDPWR a_13011_19242# single_9b_cdac_1.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5766 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5767 a_10254_2858# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X5768 single_9b_cdac_1.CF[8] a_13011_25902# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5769 a_12137_22521# a_11658_22138# a_12047_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5770 VGND sar9b_0.cyclic_flag_0.FINAL a_8883_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5771 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5772 VGND a_13011_23238# single_9b_cdac_1.CF[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5773 VDPWR sar9b_0.net58 a_3822_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5774 VGND sar9b_0.net48 a_5622_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X5775 a_7602_18116# a_8057_18463# a_8006_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5776 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5777 a_7338_24802# a_6378_24802# a_6902_25087# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5778 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5779 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5780 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5781 a_12182_23755# a_12047_23853# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5782 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5783 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5784 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5785 VDPWR a_7284_20787# a_7289_21127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5786 a_12870_18271# a_12618_18142# a_13008_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5787 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5788 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5789 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5790 ua[4] th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X5791 a_17125_9355# clk a_16331_9671# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5792 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5793 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5794 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5795 VGND a_11859_17910# single_9b_cdac_1.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5796 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5797 VGND sar9b_0._17_ a_4922_20857# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X5798 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5799 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5800 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5801 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5802 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5803 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5804 VDPWR clk a_16331_9671# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X5805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5806 VDPWR a_8334_17021# a_8266_17113# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X5807 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5808 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5809 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5811 VDPWR a_8115_28566# uo_out[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5812 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5814 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5815 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5816 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5817 sar9b_0.net19 a_2892_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5818 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5819 VDPWR sar9b_0.net48 a_10239_19235# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5820 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5821 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5822 VDPWR sar9b_0.net21 a_7539_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5823 VGND sar9b_0.net65 a_3839_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15182 pd=1.125 as=0.1152 ps=1 w=0.64 l=0.15
X5824 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5825 uo_out[3] a_9939_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5826 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5827 VDPWR sar9b_0.net47 a_7566_21017# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5828 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5829 a_8874_19178# a_7914_19178# a_8438_18958# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5830 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5831 VGND sar9b_0.net58 a_5910_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5832 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y a_45123_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5833 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5834 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5835 VDPWR a_2931_28566# uio_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5836 sar9b_0.net37 a_9900_19047# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5837 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5838 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5839 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5840 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5841 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5842 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5843 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X5844 VGND sar9b_0.clknet_1_1__leaf_CLK a_4755_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X5845 th_dif_sw_0.CKB a_2603_17006# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X5846 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5847 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5848 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5849 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5850 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5851 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5852 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5853 a_7062_20813# a_6834_20780# a_6975_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5854 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5856 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5857 a_11568_27473# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5858 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1739 ps=1.21 w=0.74 l=0.15
X5859 a_12047_23853# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5860 sar9b_0.clk_div_0.COUNT\[3\] a_4210_22378# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X5861 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5862 VGND a_12870_18271# a_12828_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5863 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5864 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5865 a_5010_28495# a_5460_28377# a_5412_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X5866 VDPWR a_10995_28566# uo_out[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5867 a_4365_25770# a_4136_25584# a_4531_25875# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.0441 ps=0.63 w=0.42 l=0.15
X5868 VDPWR a_8019_17910# single_9b_cdac_1.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5869 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5870 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5871 a_9472_18823# a_8874_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5872 a_12047_18525# a_11658_18142# a_11382_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5873 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5874 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5875 VDPWR sar9b_0.net44 a_5322_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5876 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5877 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5878 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5879 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X5880 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5882 a_6834_20780# a_7284_20787# a_7236_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X5883 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5884 uo_out[6] a_8115_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5885 VDPWR sar9b_0.net19 a_5235_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5886 a_6678_27470# sar9b_0.net40 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5888 VGND a_11915_28371# uo_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X5889 single_9b_cdac_1.CF[3] a_13011_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5890 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5891 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5892 VDPWR a_7914_27466# a_8166_27595# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5893 VGND sar9b_0.net54 a_8790_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5894 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5895 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5896 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5897 single_9b_cdac_0.SW[4] a_11915_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5898 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5899 VGND a_12435_24802# single_9b_cdac_1.CF[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5900 VGND sar9b_0.net49 a_10035_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5901 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5902 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5903 a_5412_28559# a_5151_28559# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X5904 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5905 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5906 a_12828_18149# a_11658_18142# a_12618_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5907 VGND sar9b_0.net58 a_5133_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5908 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5909 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5910 VDPWR sar9b_0.net5 a_8842_18206# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5911 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5912 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5913 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5914 a_11722_25838# a_10932_25713# a_11214_25728# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5915 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5916 a_5761_21100# sar9b_0._08_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2382 ps=1.555 w=1 l=0.15
X5917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A a_35519_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5918 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5919 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5920 VDPWR a_11339_27039# single_9b_cdac_0.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5921 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5922 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5923 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5924 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5925 a_6086_23889# a_5823_23477# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5926 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5928 a_10710_25895# a_10482_25831# a_10623_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5929 a_4922_20857# sar9b_0.net65 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X5930 a_10528_20155# a_9930_20510# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5931 a_25915_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5932 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5933 VDPWR sar9b_0.net11 a_8202_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5935 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5936 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5937 uo_out[1] a_12531_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5938 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5939 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5940 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5941 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5942 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5943 a_13216_22473# a_12618_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5944 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5945 a_2508_23444# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5946 a_3206_22432# a_3027_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X5947 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5948 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5949 uo_out[2] a_10995_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5950 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5951 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5952 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5953 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5954 single_9b_cdac_1.CF[6] a_13011_24570# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5955 a_6783_19481# a_6642_19448# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5956 VDPWR a_6880_17491# sar9b_0.net5 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5957 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5958 VDPWR tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X5959 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5960 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5961 VDPWR a_13011_23238# single_9b_cdac_1.CF[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5963 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5964 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5965 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5966 VGND a_6579_18832# sar9b_0.net46 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5967 a_8266_18445# a_8052_18123# a_7602_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5968 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5969 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5970 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5971 VDPWR single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5972 VDPWR a_13216_19809# sar9b_0.net29 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5973 VGND sar9b_0.net54 a_8013_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5974 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5975 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5976 a_3926_24136# a_3014_24136# a_3819_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X5977 a_4292_19768# sar9b_0.net46 a_4072_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.195 ps=1.39 w=1 l=0.15
X5978 a_7882_19538# sar9b_0.net62 a_8403_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5979 single_9b_cdac_1.SW[2] a_8019_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5980 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5981 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5982 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5983 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5984 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5985 VDPWR a_7539_28566# uo_out[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5986 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5987 a_11104_24151# a_10506_24506# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5988 a_12870_22267# a_12618_22138# a_13008_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5989 a_10612_17491# a_9634_17478# a_10410_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5990 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5991 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5992 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# a_15265_9613# VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X5993 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5994 VGND sar9b_0.net60 a_3603_28156# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X5995 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5996 VGND a_6834_20780# a_6636_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5997 a_5711_17527# a_5506_17478# a_5046_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5999 a_10742_25087# a_10607_25185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6000 a_5798_18561# a_5535_18149# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X6001 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6002 a_11380_21225# a_10402_21098# a_11178_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X6003 VDPWR sar9b_0.net48 a_10335_16817# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X6004 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6006 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6007 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6008 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6009 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6010 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6011 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6012 a_9737_21523# a_9258_21842# a_9647_21523# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X6013 VDPWR sar9b_0.net35 a_8595_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X6014 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6015 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6016 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6017 VGND a_4125_25958# a_4136_25584# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2553 ps=2.17 w=0.74 l=0.15
X6018 a_6282_17846# a_5506_17478# a_5846_17626# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X6019 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6020 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6021 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 a_10227_23490# sar9b_0.net38 0.02331f
C1 a_8098_23762# a_8874_23470# 0.3578f
C2 sar9b_0.net58 a_5046_27230# 0.26485f
C3 VDPWR sar9b_0.net44 0.51556f
C4 sar9b_0.net13 a_10402_25094# 0.01895f
C5 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[5] 7.94111f
C6 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[4] 0.02008f
C7 a_10218_27466# a_10742_27751# 0.05022f
C8 a_7478_27751# sar9b_0.net36 0.06675f
C9 a_7882_19538# sar9b_0.net47 0.23112f
C10 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[1] 16.8012f
C11 a_10859_26330# sar9b_0.net42 0.04314f
C12 a_5322_17846# a_5046_17906# 0.1263f
C13 a_4812_28371# sar9b_0.net58 0.02979f
C14 a_8019_17910# sar9b_0.net37 0.20475f
C15 sar9b_0.net18 sar9b_0.net58 0.33351f
C16 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.05472f
C17 sar9b_0.net63 sar9b_0.net69 0.04307f
C18 sar9b_0.net8 sar9b_0.net40 0.02953f
C19 a_11338_19178# sar9b_0.net73 0.01335f
C20 sar9b_0.net8 a_11842_19766# 0.02187f
C21 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.05105f
C22 sar9b_0.net18 a_2706_27440# 0.06755f
C23 sar9b_0.net9 single_9b_cdac_1.CF[2] 0.25447f
C24 sar9b_0.net8 sar9b_0.net51 0.28615f
C25 a_12435_24802# single_9b_cdac_1.CF[7] 0.35432f
C26 sar9b_0.clk_div_0.COUNT\[0\] clk 0.21954f
C27 sar9b_0.net42 sar9b_0.net5 0.01903f
C28 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.7611f
C29 a_6414_23681# a_6922_23534# 0.19065f
C30 VDPWR a_7936_25137# 0.20887f
C31 a_8842_18206# sar9b_0.net37 0.01698f
C32 single_9b_cdac_1.SW[1] a_57946_16877# 0.28324f
C33 sar9b_0.net60 sar9b_0.net4 0.69419f
C34 sar9b_0.net49 a_9930_20510# 0.25469f
C35 a_38738_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.23864f
C36 a_3561_22527# a_3454_22567# 0.14439f
C37 sar9b_0.net60 sar9b_0._15_ 0.04165f
C38 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.3196f
C39 a_5046_27230# sar9b_0.net37 0.04431f
C40 VDPWR a_8438_23755# 0.20949f
C41 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.76578f
C42 sar9b_0.net27 a_5196_18116# 0.2837f
C43 a_11382_23474# sar9b_0.net53 0.25588f
C44 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.45521f
C45 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C46 VDPWR a_11776_21141# 0.20631f
C47 a_4755_22138# a_5739_22488# 0.08669f
C48 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] 1.15121f
C49 a_13011_21906# sar9b_0.net9 0.22439f
C50 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 ua[0] 0.13178f
C51 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.31534f
C52 a_7097_19795# a_7374_19685# 0.09983f
C53 sar9b_0.net23 a_7692_26108# 0.27877f
C54 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[2\] 0.03174f
C55 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.01003f
C56 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 1.71649f
C57 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.6919f
C58 a_57946_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.23864f
C59 sar9b_0.net4 a_5753_24250# 0.02172f
C60 sar9b_0.net65 a_3027_22138# 0.01967f
C61 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.S[0] 0.01492f
C62 a_44418_17740# single_9b_cdac_1.SW[4] 0.18991f
C63 VDPWR single_9b_cdac_0.SW[8] 2.48304f
C64 sar9b_0._15_ a_5753_24250# 0.05531f
C65 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[4] 10.6485f
C66 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.19325f
C67 a_11338_19178# sar9b_0.net48 0.20192f
C68 sar9b_0.net69 sar9b_0.clknet_1_1__leaf_CLK 0.08399f
C69 sar9b_0.net26 sar9b_0.net53 0.06847f
C70 sar9b_0.net8 a_10742_21091# 0.03386f
C71 sar9b_0.net25 uo_out[0] 0.27942f
C72 single_9b_cdac_1.CF[7] a_13011_24570# 0.03372f
C73 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.19125f
C74 VDPWR sar9b_0._00_ 0.73774f
C75 sar9b_0.net12 a_11842_26426# 0.02738f
C76 a_21368_4076# ua[0] 0.17332f
C77 sar9b_0.net35 tdc_0.OUTN 0.05242f
C78 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.VCP 0.31462f
C79 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[4] 0.01997f
C80 a_10218_24802# sar9b_0.net12 0.06895f
C81 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.10626f
C82 sar9b_0.net57 a_5535_18149# 0.01663f
C83 sar9b_0.net40 sar9b_0._02_ 0.48012f
C84 a_8057_18463# a_8334_18353# 0.09983f
C85 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.36013f
C86 a_5289_22527# sar9b_0.net39 0.0302f
C87 sar9b_0.net49 sar9b_0.net5 0.51189f
C88 sar9b_0._09_ sar9b_0._07_ 0.58193f
C89 a_6058_18445# a_6126_18353# 0.35559f
C90 a_5849_18463# a_6634_18206# 0.26257f
C91 m2_23774_17236# VDPWR 0.19016f
C92 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.17533f
C93 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[6] 0.0313f
C94 sar9b_0.net56 sar9b_0.net73 0.05473f
C95 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.03484f
C96 VDPWR a_2893_24992# 0.23635f
C97 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C98 single_9b_cdac_0.SW[6] th_dif_sw_0.VCN 0.09468f
C99 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[7] 14.2348f
C100 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.6205f
C101 a_2893_24992# sar9b_0._14_ 0.34774f
C102 sar9b_0.net72 sar9b_0.net68 0.02728f
C103 VDPWR a_4749_27652# 0.4017f
C104 a_11008_17491# sar9b_0.net61 0.03855f
C105 sar9b_0._18_ sar9b_0.clknet_1_1__leaf_CLK 0.02875f
C106 a_7926_23234# sar9b_0.net62 0.21091f
C107 a_5823_23477# sar9b_0.net11 0.05916f
C108 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02552f
C109 sar9b_0._09_ sar9b_0._08_ 0.0865f
C110 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36555_29911# 0.01076f
C111 VDPWR a_10227_23490# 0.4365f
C112 a_5581_20992# a_5812_21028# 0.10754f
C113 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.12431f
C114 sar9b_0.net13 a_6767_25185# 0.07236f
C115 a_5196_24776# sar9b_0._03_ 0.10899f
C116 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[0] 0.03109f
C117 th_dif_sw_0.th_sw_1.CK ua[3] 0.42268f
C118 sar9b_0.net58 a_5674_28147# 0.12675f
C119 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[0] 18.6433f
C120 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] 3.1021f
C121 sar9b_0.net66 sar9b_0.clknet_1_0__leaf_CLK 0.08897f
C122 sar9b_0.net59 sar9b_0.net45 0.55332f
C123 single_9b_cdac_0.SW[7] a_29134_26999# 0.28324f
C124 a_10707_23470# sar9b_0.net36 0.02924f
C125 a_11338_19178# sar9b_0.net50 0.01132f
C126 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0._12_ 0.30315f
C127 a_10816_21487# sar9b_0.net36 0.02497f
C128 a_11339_27039# sar9b_0.net52 0.07246f
C129 a_8266_17113# sar9b_0.net27 0.02296f
C130 sar9b_0.net63 sar9b_0.net60 0.09293f
C131 a_10227_23490# sar9b_0.net1 0.13989f
C132 sar9b_0.net2 a_10758_24459# 0.07084f
C133 single_9b_cdac_0.SW[7] sar9b_0.net38 0.18897f
C134 a_2931_28566# sar9b_0.net60 0.09891f
C135 a_10803_18142# sar9b_0.net73 0.13298f
C136 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[2] 0.01637f
C137 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[0] 18.6879f
C138 a_8031_26141# sar9b_0.cyclic_flag_0.FINAL 0.03467f
C139 a_6783_19481# sar9b_0.net40 0.05886f
C140 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR 0.84061f
C141 sar9b_0.net24 a_8940_27039# 0.28492f
C142 a_8303_18859# sar9b_0.net48 0.22623f
C143 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C144 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 3.10626f
C145 sar9b_0.net45 a_8883_27466# 0.30828f
C146 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.84426f
C147 sar9b_0.net48 single_9b_cdac_1.SW[0] 0.1553f
C148 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36555_15501# 0.01076f
C149 a_10218_27466# a_10607_27849# 0.06034f
C150 ui_in[2] ui_in[1] 0.03102f
C151 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C152 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[2] 0.01297f
C153 sar9b_0.net56 sar9b_0.net48 0.26514f
C154 sar9b_0.net47 a_6879_22145# 0.17478f
C155 sar9b_0.net41 sar9b_0.net37 0.12296f
C156 a_2835_24136# a_2508_23444# 0.01422f
C157 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 a_63626_26990# 0.14695f
C158 a_7638_19238# a_8098_18810# 0.26257f
C159 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.10429f
C160 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[7] 0.02364f
C161 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[4] 0.02019f
C162 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.0313f
C163 th_dif_sw_0.CK sar9b_0.net38 0.21539f
C164 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.95338f
C165 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62553f
C166 sar9b_0.net7 a_11008_17491# 0.27173f
C167 a_10858_17113# a_10644_16791# 0.04522f
C168 a_4755_22138# sar9b_0._18_ 0.01306f
C169 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.07517f
C170 single_9b_cdac_1.SW[3] clk 0.10355f
C171 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS ua[4] 0.93546f
C172 sar9b_0.net59 a_9870_27060# 0.26796f
C173 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[0] 0.01464f
C174 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 a_49221_17740# 0.14695f
C175 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP a_62748_26999# 0.04592f
C176 sar9b_0.net32 a_12182_23755# 0.01954f
C177 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.01003f
C178 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.84425f
C179 sar9b_0.net17 sar9b_0.net19 0.01908f
C180 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62573f
C181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.7611f
C182 a_7566_21017# a_8074_20870# 0.19065f
C183 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 2.71729f
C184 a_10762_18823# sar9b_0.net36 0.01606f
C185 a_10506_24506# a_11104_24151# 0.06623f
C186 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INP 0.06558f
C187 a_7638_23474# a_6922_23534# 0.03811f
C188 a_10218_24802# a_9942_24806# 0.1263f
C189 VDPWR a_5739_22488# 0.09539f
C190 a_10690_22806# sar9b_0.net53 0.11211f
C191 sar9b_0.net41 a_9730_24138# 0.02215f
C192 a_12870_26263# a_12618_26134# 0.27388f
C193 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.93403f
C194 single_9b_cdac_0.SW[6] uo_out[0] 0.04513f
C195 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 0.19266f
C196 sar9b_0.net27 single_9b_cdac_0.SW[0] 0.01491f
C197 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[0] 0.0223f
C198 a_8595_17910# sar9b_0.net5 0.02485f
C199 a_7097_19795# sar9b_0.net10 0.06701f
C200 sar9b_0.net56 sar9b_0.net46 2.24988f
C201 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.02513f
C202 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[8] 0.03927f
C203 a_4922_20857# sar9b_0.net65 0.08585f
C204 a_8166_27595# a_8512_27801# 0.07649f
C205 a_3206_22432# a_3713_22522# 0.21226f
C206 a_8057_18463# sar9b_0.net61 0.01568f
C207 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.105f
C208 a_9162_23174# sar9b_0.net54 0.27476f
C209 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[3] 0.04427f
C210 single_9b_cdac_0.SW[2] sar9b_0.net28 0.04952f
C211 VDPWR sar9b_0._13_ 0.47588f
C212 a_11842_18434# sar9b_0.net27 0.01125f
C213 a_7404_16784# sar9b_0.net6 0.01335f
C214 sar9b_0.net19 a_3822_27060# 0.0307f
C215 sar9b_0._13_ sar9b_0._14_ 0.15271f
C216 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.62443f
C217 sar9b_0.net42 sar9b_0.net74 0.61827f
C218 sar9b_0.net9 single_9b_cdac_1.CF[4] 0.01701f
C219 a_6678_27470# sar9b_0.net44 0.04249f
C220 sar9b_0.net56 a_9154_20142# 0.01042f
C221 a_10607_25185# sar9b_0.net12 0.06942f
C222 a_2892_27039# sar9b_0.net19 0.29845f
C223 VDPWR a_9126_19131# 0.28669f
C224 a_11658_18142# a_11842_18434# 0.44532f
C225 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C226 sar9b_0.clknet_1_0__leaf_CLK a_2918_20140# 0.12018f
C227 sar9b_0.net43 sar9b_0.net59 0.30303f
C228 th_dif_sw_0.CK sar9b_0.net6 0.02947f
C229 VDPWR a_5711_17527# 0.25721f
C230 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.22879f
C231 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.03729f
C232 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.07579f
C233 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.95338f
C234 VDPWR sar9b_0._10_ 0.48054f
C235 a_10803_18142# single_9b_cdac_1.SW[3] 0.3509f
C236 VDPWR a_13011_23238# 0.48316f
C237 sar9b_0.net42 sar9b_0.net31 0.08505f
C238 dw_12589_1395# a_10482_3438# 0.05479f
C239 a_11842_26426# a_12047_26517# 0.09983f
C240 sar9b_0.net49 a_10035_19474# 0.26854f
C241 VDPWR single_9b_cdac_0.SW[7] 2.68913f
C242 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[5] 0.0313f
C243 a_4755_22138# sar9b_0.net60 0.01468f
C244 VDPWR a_9546_24506# 0.86145f
C245 a_2835_24136# sar9b_0.net70 0.06896f
C246 single_9b_cdac_1.CF[3] single_9b_cdac_1.CF[0] 0.04014f
C247 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.22597f
C248 sar9b_0.net23 uo_out[3] 0.10721f
C249 sar9b_0.net28 single_9b_cdac_1.CF[0] 0.0432f
C250 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.3196f
C251 a_7289_21127# a_7284_20787# 0.44098f
C252 a_10528_20155# sar9b_0.net51 0.04328f
C253 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[8] 2.12011f
C254 sar9b_0.net16 a_2603_17006# 0.22549f
C255 a_11859_17910# sar9b_0.net39 0.20696f
C256 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.27713f
C257 VDPWR a_7404_16784# 0.19127f
C258 a_11859_20574# single_9b_cdac_1.SW[8] 0.35377f
C259 VDPWR sar9b_0.net69 1.21061f
C260 sar9b_0._09_ a_3991_19768# 0.01296f
C261 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.10499f
C262 VDPWR a_11382_22142# 0.28804f
C263 VDPWR th_dif_sw_0.CK 1.56597f
C264 single_9b_cdac_0.SW[8] single_9b_cdac_0.SW[3] 0.026f
C265 a_6954_27466# sar9b_0.net45 0.02051f
C266 sar9b_0.net52 sar9b_0.net37 0.74767f
C267 sar9b_0._14_ sar9b_0.net69 0.03025f
C268 sar9b_0.net48 a_5394_18116# 0.26617f
C269 sar9b_0.net17 a_2706_26108# 0.01317f
C270 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0313f
C271 sar9b_0.net58 a_3231_27227# 0.17354f
C272 a_5235_27466# a_5460_28377# 0.01146f
C273 single_9b_cdac_1.SW[1] sar9b_0.net6 0.04631f
C274 single_9b_cdac_1.cdac_sw_9b_0.S[4] a_43540_16877# 0.59531f
C275 sar9b_0.net22 uo_out[4] 0.11108f
C276 single_9b_cdac_1.CF[3] single_9b_cdac_1.SW[2] 0.01297f
C277 a_11382_18146# sar9b_0.net61 0.02131f
C278 sar9b_0.net59 a_3540_27045# 0.0106f
C279 a_2739_20140# a_3166_20145# 0.04602f
C280 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.51772f
C281 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.10984p
C282 a_10218_24802# a_11430_24931# 0.07766f
C283 sar9b_0.net49 a_9942_20810# 0.28171f
C284 a_7404_17715# sar9b_0.net73 0.12657f
C285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C286 sar9b_0.net41 sar9b_0.net57 0.02983f
C287 sar9b_0.net8 sar9b_0.net42 0.01991f
C288 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C289 VDPWR sar9b_0._18_ 1.75124f
C290 th_dif_sw_0.th_sw_1.CKB a_10166_3438# 0.06536f
C291 a_11382_23474# a_12047_23853# 0.19065f
C292 a_8340_26115# sar9b_0.net59 0.17782f
C293 sar9b_0.net26 a_12047_22521# 0.01371f
C294 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 ua[0] 0.12076f
C295 VDPWR sar9b_0._01_ 0.28816f
C296 a_10649_17131# single_9b_cdac_1.SW[2] 0.0163f
C297 sar9b_0.net30 sar9b_0.net26 0.11005f
C298 sar9b_0.net43 sar9b_0.net12 0.38567f
C299 single_9b_cdac_1.SW[5] a_38738_16877# 0.28324f
C300 a_8345_26455# a_9130_26198# 0.26257f
C301 VDPWR a_5046_17906# 0.28567f
C302 a_3454_22567# a_3027_22138# 0.04602f
C303 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.69086f
C304 sar9b_0.net67 sar9b_0._05_ 0.21501f
C305 uo_out[3] ui_in[0] 0.06786f
C306 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.42014f
C307 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C308 VDPWR single_9b_cdac_1.SW[1] 2.46863f
C309 a_3540_27045# a_4330_27170# 0.1263f
C310 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.22655f
C311 single_9b_cdac_1.SW[4] ua[0] 0.13619f
C312 sar9b_0.net13 sar9b_0.net12 0.39165f
C313 a_10607_25185# a_9942_24806# 0.19065f
C314 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.42784f
C315 sar9b_0.net28 single_9b_cdac_1.SW[8] 0.04546f
C316 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[4] 0.03482f
C317 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.28575f
C318 sar9b_0._07_ a_5126_20140# 0.02529f
C319 a_7092_19455# sar9b_0.net47 0.18759f
C320 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[6] 8.40786f
C321 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.81428f
C322 a_7470_22349# a_7978_22202# 0.19065f
C323 sar9b_0.net10 a_7402_22441# 0.01467f
C324 a_5628_19768# sar9b_0._07_ 0.03465f
C325 sar9b_0.net7 a_11382_18146# 0.05241f
C326 a_5460_28377# a_5742_28392# 0.06034f
C327 a_13011_23238# sar9b_0.net29 0.02021f
C328 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.03729f
C329 single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.26707f
C330 sar9b_0.net35 sar9b_0.net39 0.0534f
C331 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.81428f
C332 a_10402_25094# sar9b_0.net38 0.0296f
C333 sar9b_0.net3 sar9b_0.net17 0.49213f
C334 a_10548_19053# a_10553_18922# 0.44532f
C335 sar9b_0.net8 sar9b_0.net49 0.4261f
C336 a_4755_22138# a_4934_22432# 0.54361f
C337 sar9b_0.net2 sar9b_0.net39 0.23235f
C338 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.83441f
C339 a_9126_19131# a_9472_18823# 0.07649f
C340 sar9b_0.net24 sar9b_0.net36 0.37491f
C341 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C342 tdc_0.OUTP th_dif_sw_0.CKB 0.30524f
C343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[3] 0.01887f
C344 VDPWR a_6126_18353# 0.26525f
C345 single_9b_cdac_0.cdac_sw_9b_0.S[5] a_39616_26990# 0.22512f
C346 a_5711_26851# a_5322_27170# 0.05462f
C347 a_9839_17527# a_9974_17626# 0.35559f
C348 single_9b_cdac_0.SW[1] clk 0.13072f
C349 a_9363_20826# a_9258_21842# 0.02481f
C350 a_8202_23174# a_9414_23127# 0.07766f
C351 a_8386_22806# a_8726_22954# 0.24088f
C352 a_6132_23451# a_5823_23477# 0.07766f
C353 a_5711_17527# a_5846_17626# 0.35559f
C354 a_8052_18123# sar9b_0.net37 0.01856f
C355 VDPWR a_3795_19512# 0.60141f
C356 VDPWR a_3180_19448# 0.26779f
C357 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.19266f
C358 a_6880_17491# sar9b_0.net56 0.0197f
C359 sar9b_0.net44 a_5711_26851# 0.06353f
C360 a_10553_18922# sar9b_0.net38 0.02338f
C361 VDPWR sar9b_0.net60 2.99913f
C362 a_10816_21487# sar9b_0.net9 0.31769f
C363 sar9b_0._07_ sar9b_0.net4 0.13017f
C364 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.71729f
C365 sar9b_0.net40 sar9b_0.net73 0.05965f
C366 sar9b_0.net11 sar9b_0.net54 0.36694f
C367 a_7092_19455# a_6642_19448# 0.03471f
C368 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[5] 0.02008f
C369 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[4] 0.20642f
C370 sar9b_0.net36 a_10623_25895# 0.01701f
C371 a_7404_17715# sar9b_0.net46 0.03295f
C372 sar9b_0.net51 sar9b_0.net73 0.03243f
C373 a_9546_24506# a_9270_24566# 0.1263f
C374 a_12618_23470# clk 0.0119f
C375 a_10649_17131# sar9b_0.net61 0.01074f
C376 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.6919f
C377 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.01402f
C378 a_2892_23070# a_3219_22860# 0.09161f
C379 a_10895_22855# sar9b_0.net2 0.01734f
C380 a_6484_22845# sar9b_0.clk_div_0.COUNT\[2\] 0.0424f
C381 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[2\] 0.04613f
C382 a_7284_20787# sar9b_0.net47 0.17237f
C383 VDPWR a_5753_24250# 0.21444f
C384 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.05472f
C385 th_dif_sw_0.th_sw_1.CKB a_10254_2858# 0.42927f
C386 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.01664f
C387 a_6252_20780# sar9b_0._17_ 0.05545f
C388 a_10218_27466# a_10995_28566# 0.01498f
C389 sar9b_0.net48 a_9174_17906# 0.2009f
C390 VDPWR a_12618_26134# 0.35483f
C391 sar9b_0.net43 a_9942_24806# 0.01787f
C392 a_8052_18123# a_7602_18116# 0.03471f
C393 sar9b_0.net53 a_12047_22521# 0.22562f
C394 single_9b_cdac_0.SW[1] a_57946_26999# 0.28324f
C395 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[0] 0.02907f
C396 sar9b_0.net52 sar9b_0.net57 0.87251f
C397 sar9b_0.net27 clk 0.04404f
C398 a_6975_20813# sar9b_0.net40 0.01008f
C399 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.0187f
C400 single_9b_cdac_0.SW[5] clk 0.153f
C401 sar9b_0.net30 sar9b_0.net53 0.04133f
C402 sar9b_0.net35 a_6902_25087# 0.0142f
C403 sar9b_0.net13 a_9942_24806# 0.08367f
C404 sar9b_0.net23 single_9b_cdac_0.SW[8] 0.02815f
C405 sar9b_0.net33 sar9b_0.net52 0.30065f
C406 a_3561_22527# sar9b_0._12_ 0.03484f
C407 sar9b_0.clknet_0_CLK sar9b_0._12_ 0.02864f
C408 sar9b_0.net40 sar9b_0.net48 0.10648f
C409 sar9b_0.net53 a_12047_23853# 0.22582f
C410 sar9b_0.net41 a_10410_17846# 0.06272f
C411 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.26707f
C412 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.43767f
C413 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.11216f
C414 a_11382_22142# a_11658_22138# 0.1263f
C415 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[3] 0.026f
C416 a_10623_25895# a_10937_25582# 0.07826f
C417 a_4083_28566# sar9b_0.net60 0.05402f
C418 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.02149f
C419 sar9b_0.net27 single_9b_cdac_1.SW[0] 0.02138f
C420 a_10506_23174# sar9b_0.net11 0.06113f
C421 a_7338_24802# sar9b_0.net54 0.26564f
C422 a_3369_24181# a_3521_24240# 0.22338f
C423 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[2] 0.01297f
C424 a_2931_28566# a_3156_27447# 0.01146f
C425 VDPWR uio_out[0] 0.76516f
C426 sar9b_0.net74 sar9b_0.net11 0.42192f
C427 a_40321_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.01076f
C428 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.A 0.10129f
C429 VDPWR a_10402_25094# 0.21159f
C430 sar9b_0.net56 sar9b_0.net27 0.19838f
C431 a_8098_23762# sar9b_0.net54 0.02919f
C432 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.22609f
C433 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C434 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[3] 0.12359f
C435 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.01175f
C436 VDPWR a_5506_26802# 0.2219f
C437 sar9b_0.net63 a_6484_22845# 0.05368f
C438 sar9b_0.net31 sar9b_0.net11 0.38707f
C439 a_7188_22119# a_7470_22349# 0.05462f
C440 sar9b_0.net2 sar9b_0.net36 1.60268f
C441 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 3.27788f
C442 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.1717f
C443 sar9b_0.net19 a_5046_27230# 0.02764f
C444 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[7] 5.94919f
C445 sar9b_0.net27 a_13011_20806# 0.04065f
C446 a_10218_27466# a_9588_27045# 0.01007f
C447 tdc_0.OUTP single_9b_cdac_1.SW[0] 0.86423f
C448 sar9b_0.net40 sar9b_0.net50 0.30217f
C449 a_5484_23444# sar9b_0.net57 0.04904f
C450 VDPWR a_10553_18922# 0.21937f
C451 th_dif_sw_0.th_sw_1.CKB ua[3] 0.08416f
C452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46159_29911# 0.01076f
C453 VDPWR a_4934_22432# 0.89137f
C454 sar9b_0.net40 single_9b_cdac_1.SW[3] 0.03187f
C455 a_12870_18271# sar9b_0.net50 0.17284f
C456 a_11842_19766# sar9b_0.net50 0.10082f
C457 th_dif_sw_0.th_sw_1.CKB clk 0.0198f
C458 sar9b_0.net46 sar9b_0.net51 0.64278f
C459 VDPWR a_48343_26999# 1.81495f
C460 VDPWR a_9974_17626# 0.19746f
C461 sar9b_0.net40 a_12618_18142# 0.01397f
C462 sar9b_0.net65 sar9b_0._17_ 0.17308f
C463 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.31534f
C464 sar9b_0.net50 sar9b_0.net51 0.03079f
C465 a_12870_18271# a_12618_18142# 0.27388f
C466 a_11842_18434# a_12047_18525# 0.09983f
C467 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] 1.55949f
C468 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.17533f
C469 a_7890_26108# a_8340_26115# 0.03529f
C470 a_8031_26141# a_7692_26108# 0.07649f
C471 uo_out[4] uo_out[3] 2.93276f
C472 sar9b_0.net63 a_5823_23477# 0.05368f
C473 sar9b_0.net60 a_5682_23444# 0.04812f
C474 sar9b_0._10_ sar9b_0.net71 0.01246f
C475 sar9b_0.net32 uo_out[1] 0.22658f
C476 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.01152f
C477 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C478 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.42014f
C479 a_9154_20142# sar9b_0.net51 0.06402f
C480 a_8874_19178# sar9b_0.net5 0.01167f
C481 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.08672f
C482 a_4083_28566# uio_out[0] 0.37232f
C483 sar9b_0.net36 a_10758_24459# 0.02391f
C484 a_11338_19178# sar9b_0.net26 0.05306f
C485 sar9b_0.net52 a_11178_24802# 0.24274f
C486 sar9b_0._07_ sar9b_0.clknet_1_1__leaf_CLK 0.02605f
C487 clk single_9b_cdac_1.SW[7] 0.08277f
C488 a_9126_23599# a_8874_23470# 0.27388f
C489 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 ua[0] 0.12378f
C490 sar9b_0.net13 a_11430_24931# 0.03609f
C491 a_10218_27466# a_11178_27466# 0.03432f
C492 single_9b_cdac_1.cdac_sw_9b_0.S[1] ua[0] 1.19426f
C493 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._05_ 0.03201f
C494 a_7914_27466# sar9b_0.net36 0.06473f
C495 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] 3.10218f
C496 a_7926_23234# sar9b_0.net11 0.05391f
C497 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.07579f
C498 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[4] 1.90184f
C499 sar9b_0.net20 sar9b_0.net58 0.46059f
C500 sar9b_0.net32 a_9939_28566# 0.04595f
C501 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C502 VDPWR a_14897_9355# 0.01057f
C503 a_21684_3438# th_dif_sw_0.th_sw_1.CK 0.12114f
C504 a_5100_24375# a_4467_24162# 0.01351f
C505 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.26709f
C506 VDPWR sar9b_0.net67 0.30253f
C507 sar9b_0.net31 sar9b_0.net45 0.06702f
C508 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP a_29134_26999# 0.04592f
C509 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.01515f
C510 single_9b_cdac_0.cdac_sw_9b_0.S[5] th_dif_sw_0.VCN 6.58553f
C511 sar9b_0.net18 a_3161_27787# 0.01348f
C512 sar9b_0.net55 a_6484_22845# 0.01609f
C513 sar9b_0._07_ sar9b_0.net55 0.01037f
C514 a_21368_4076# dw_17224_1400# 26.7601f
C515 single_9b_cdac_1.SW[0] single_9b_cdac_1.SW[7] 0.02168f
C516 a_14871_9671# th_dif_sw_0.VCP 0.07081f
C517 sar9b_0.net26 clk 0.04511f
C518 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] 3.10214f
C519 a_6880_17491# a_7404_17715# 0.01194f
C520 sar9b_0.net43 sar9b_0.net54 0.53075f
C521 VDPWR a_6767_25185# 0.26598f
C522 sar9b_0.clknet_1_0__leaf_CLK sar9b_0.clknet_1_1__leaf_CLK 0.01438f
C523 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.07517f
C524 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.02638f
C525 a_10858_17113# single_9b_cdac_1.SW[1] 0.01467f
C526 sar9b_0.net48 a_7914_19178# 0.17382f
C527 VDPWR a_8874_23470# 0.39649f
C528 sar9b_0.net58 a_6250_28502# 0.20323f
C529 a_4011_22488# sar9b_0.clknet_0_CLK 0.01809f
C530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.SW[2] 0.17199f
C531 single_9b_cdac_1.CF[8] a_13011_24802# 0.02059f
C532 sar9b_0.net13 sar9b_0.net54 1.09911f
C533 sar9b_0.net59 sar9b_0.net38 0.05434f
C534 sar9b_0.net58 a_5322_27170# 0.17211f
C535 a_4755_22138# sar9b_0._07_ 0.01014f
C536 a_7374_19685# sar9b_0.net35 0.01051f
C537 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.06503f
C538 a_7097_19795# a_7882_19538# 0.26257f
C539 single_9b_cdac_1.SW[6] ua[0] 0.13161f
C540 a_13011_16810# single_9b_cdac_1.SW[5] 0.35162f
C541 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.22875f
C542 a_4755_22138# a_5441_22522# 0.27693f
C543 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.05472f
C544 a_6678_27470# sar9b_0.net60 0.21743f
C545 sar9b_0.net72 sar9b_0._16_ 0.06363f
C546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[5] 0.02149f
C547 a_8970_20510# a_8694_20570# 0.1263f
C548 sar9b_0.net58 sar9b_0.net44 1.08603f
C549 a_3946_27530# sar9b_0.net36 0.17818f
C550 a_9802_26815# a_9138_27163# 0.16939f
C551 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.10499f
C552 VDPWR sar9b_0.net25 0.46378f
C553 single_9b_cdac_0.SW[6] sar9b_0.net38 0.16268f
C554 sar9b_0.net8 a_11178_20806# 0.05383f
C555 a_5289_22527# a_5182_22567# 0.14439f
C556 VDPWR a_8694_20570# 0.32519f
C557 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.03729f
C558 single_9b_cdac_1.CF[8] a_13011_25902# 0.35919f
C559 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 ua[0] 0.12378f
C560 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.3545f
C561 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0313f
C562 a_8057_18463# a_8842_18206# 0.26257f
C563 a_6540_22112# sar9b_0.net39 0.30426f
C564 sar9b_0.net36 a_7343_27849# 0.04959f
C565 a_10239_19235# a_10098_19171# 0.27388f
C566 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.06503f
C567 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.12898f
C568 ui_in[7] ui_in[6] 0.03102f
C569 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.02632f
C570 sar9b_0.net46 a_7914_19178# 0.07106f
C571 a_4922_20857# sar9b_0._17_ 0.32016f
C572 single_9b_cdac_0.SW[2] sar9b_0._06_ 0.01711f
C573 a_5298_24499# sar9b_0.net54 0.25564f
C574 sar9b_0.net41 a_11008_17491# 0.03875f
C575 sar9b_0.net37 a_5322_27170# 0.05304f
C576 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[4] 0.36316f
C577 sar9b_0.net68 a_2940_25096# 0.01396f
C578 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.26709f
C579 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.31809f
C580 sar9b_0.net43 sar9b_0.net74 0.18429f
C581 a_3795_19512# a_4072_19474# 0.26693f
C582 a_16159_13315# tdc_0.RDY 0.14369f
C583 sar9b_0.net35 single_9b_cdac_1.SW[2] 0.05528f
C584 a_6132_23451# sar9b_0.net54 0.17758f
C585 a_5581_20992# sar9b_0._11_ 0.06877f
C586 sar9b_0.net71 a_3795_19512# 0.03166f
C587 sar9b_0.net44 sar9b_0.net37 0.76756f
C588 sar9b_0.net13 sar9b_0.net74 0.34392f
C589 th_dif_sw_0.CKB th_dif_sw_0.VCP 0.21902f
C590 sar9b_0.net40 a_6414_23681# 0.0209f
C591 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01152f
C592 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.84082f
C593 sar9b_0.net42 sar9b_0.net73 1.30182f
C594 sar9b_0.net18 sar9b_0.net3 0.04914f
C595 sar9b_0.net13 sar9b_0.net31 0.02786f
C596 a_10470_21795# sar9b_0.net49 0.17598f
C597 sar9b_0.net12 sar9b_0.net38 0.02887f
C598 sar9b_0.net24 a_9279_27227# 0.03138f
C599 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR 3.27795f
C600 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C601 sar9b_0.net45 sar9b_0.net34 0.19873f
C602 sar9b_0.net53 clk 0.10487f
C603 sar9b_0.net30 a_12047_23853# 0.03166f
C604 sar9b_0.net33 a_12182_26419# 0.06698f
C605 a_10690_22806# clk 0.02916f
C606 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.17533f
C607 sar9b_0.net70 a_2508_23444# 0.08416f
C608 a_16222_11316# tdc_0.phase_detector_0.INP 0.02778f
C609 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C610 sar9b_0.net60 a_6030_24396# 0.02375f
C611 single_9b_cdac_0.SW[4] a_13011_27234# 0.05684f
C612 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.38397f
C613 a_9323_27662# single_9b_cdac_0.SW[8] 0.35813f
C614 single_9b_cdac_0.SW[8] uo_out[4] 0.18749f
C615 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.69086f
C616 VDPWR sar9b_0.net59 4.515f
C617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02813f
C618 single_9b_cdac_0.SW[3] a_48343_26999# 0.28324f
C619 sar9b_0.net64 sar9b_0._18_ 0.2077f
C620 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.SW[5] 0.17355f
C621 VDPWR a_3156_27447# 0.84513f
C622 sar9b_0.net54 sar9b_0.net4 0.17203f
C623 sar9b_0.net32 a_12618_23470# 0.0684f
C624 sar9b_0.net58 a_4749_27652# 0.34567f
C625 a_3027_22138# sar9b_0._12_ 0.16198f
C626 sar9b_0._15_ sar9b_0.net54 0.08938f
C627 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[6] 0.02024f
C628 a_5753_24250# a_6030_24396# 0.09983f
C629 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.04988f
C630 sar9b_0.net65 sar9b_0._12_ 0.02841f
C631 a_5938_22378# sar9b_0._12_ 0.07878f
C632 VDPWR a_8883_27466# 0.46906f
C633 sar9b_0.net43 sar9b_0.net8 0.04888f
C634 a_10830_19068# single_9b_cdac_1.SW[1] 0.01619f
C635 sar9b_0.net42 sar9b_0.net48 0.07688f
C636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP a_33936_16877# 0.04592f
C637 VDPWR a_6738_22112# 0.36714f
C638 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 a_30012_26990# 0.14695f
C639 a_11030_22954# sar9b_0.net53 0.14085f
C640 a_3819_24136# a_3014_24136# 0.29221f
C641 sar9b_0.net49 sar9b_0.net73 0.10388f
C642 sar9b_0.net34 a_9870_27060# 0.01531f
C643 sar9b_0.net60 sar9b_0._03_ 0.02848f
C644 single_9b_cdac_0.SW[6] VDPWR 2.34024f
C645 a_4018_24235# a_2835_24136# 0.0649f
C646 VDPWR a_6484_22845# 0.26318f
C647 VDPWR sar9b_0._07_ 0.94013f
C648 a_10506_23174# a_11718_23127# 0.07766f
C649 a_10690_22806# a_11030_22954# 0.24088f
C650 a_12618_26134# a_13216_26469# 0.06623f
C651 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C652 a_4332_23043# sar9b_0.net39 0.05206f
C653 sar9b_0.net9 sar9b_0.net2 0.0459f
C654 sar9b_0.net12 a_9165_24988# 0.01031f
C655 VDPWR a_5441_22522# 0.10419f
C656 sar9b_0.net35 sar9b_0.net61 0.03955f
C657 sar9b_0.net32 sar9b_0.net27 0.2123f
C658 sar9b_0.net35 sar9b_0.net10 1.66696f
C659 sar9b_0.net32 single_9b_cdac_0.SW[5] 0.11624f
C660 sar9b_0.net40 sar9b_0.net21 0.06941f
C661 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] 1.15121f
C662 a_12064_22819# sar9b_0.net10 0.06469f
C663 VDPWR a_4330_27170# 0.29064f
C664 a_7284_20787# a_6834_20780# 0.03471f
C665 a_6636_20780# a_6975_20813# 0.07649f
C666 sar9b_0.net2 sar9b_0.net61 0.18227f
C667 sar9b_0.net2 sar9b_0.net10 0.02528f
C668 VDPWR sar9b_0._08_ 0.41847f
C669 a_3206_22432# a_4210_22378# 0.06302f
C670 a_11718_23127# sar9b_0.net31 0.01022f
C671 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[0] 0.02666f
C672 sar9b_0.net40 sar9b_0.net27 0.81488f
C673 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.14962f
C674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.7611f
C675 single_9b_cdac_1.cdac_sw_9b_0.S[0] th_dif_sw_0.VCP 0.21807p
C676 a_11915_28371# a_12531_28566# 0.03551f
C677 a_7602_16784# sar9b_0.net6 0.04668f
C678 a_12870_18271# sar9b_0.net27 0.02288f
C679 sar9b_0.net36 sar9b_0.net39 0.02403f
C680 a_7284_20787# a_7443_21496# 0.02666f
C681 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[2] 0.01887f
C682 clk th_dif_sw_0.VCP 1.62194f
C683 sar9b_0.net61 tdc_0.OUTN 0.01037f
C684 a_5633_20244# a_5931_20140# 0.02614f
C685 a_3231_27227# sar9b_0.net19 0.04509f
C686 a_18214_3039# w_17430_1606# 0.14276f
C687 VDPWR a_9900_19047# 0.20374f
C688 a_11658_18142# a_12870_18271# 0.07766f
C689 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.19147f
C690 a_13011_24802# a_13011_24570# 0.02551f
C691 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[8] 16.1938f
C692 VDPWR a_5823_23477# 0.26508f
C693 sar9b_0.net38 a_9930_20510# 0.02335f
C694 a_8591_22855# clk 0.02075f
C695 a_8940_24402# sar9b_0.net62 0.23108f
C696 a_3922_20239# a_2739_20140# 0.0649f
C697 a_4812_28371# a_5151_28559# 0.07649f
C698 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP a_62748_16877# 0.04592f
C699 a_4083_28566# sar9b_0.net59 0.10812f
C700 sar9b_0.net52 a_10284_25707# 0.02758f
C701 sar9b_0.net42 sar9b_0.net50 0.03413f
C702 a_5580_24776# a_6102_24806# 0.01519f
C703 VDPWR sar9b_0.clknet_1_0__leaf_CLK 2.99385f
C704 a_9942_24806# sar9b_0.net38 0.01422f
C705 sar9b_0.net49 sar9b_0.net48 0.59286f
C706 sar9b_0.net64 sar9b_0.net60 0.08504f
C707 a_10995_28566# single_9b_cdac_0.SW[5] 0.01783f
C708 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.CF[4] 0.12358f
C709 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[2] 0.01297f
C710 sar9b_0.net43 sar9b_0.net34 0.26137f
C711 tdc_0.OUTP sar9b_0.net40 0.02274f
C712 VDPWR sar9b_0.net12 1.09949f
C713 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 ua[0] 0.11907f
C714 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR 0.84061f
C715 a_10644_16791# a_10194_16784# 0.03493f
C716 a_9996_16784# a_10335_16817# 0.07649f
C717 VDPWR a_7602_16784# 0.3319f
C718 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C719 a_10895_22855# sar9b_0.net36 0.01323f
C720 a_6562_25094# a_7590_24931# 0.07826f
C721 sar9b_0.net7 sar9b_0.net2 0.26633f
C722 sar9b_0.net40 a_6444_19448# 0.30912f
C723 sar9b_0.net1 sar9b_0.net12 0.03139f
C724 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] 0.12898f
C725 sar9b_0._09_ a_5196_19448# 0.04256f
C726 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.03488f
C727 a_7138_27758# sar9b_0.net45 0.01918f
C728 sar9b_0.net48 a_5849_18463# 0.10592f
C729 a_6102_24806# a_6378_24802# 0.1263f
C730 sar9b_0.net38 sar9b_0.net5 0.08475f
C731 a_9760_22819# sar9b_0.net74 0.01641f
C732 sar9b_0._13_ sar9b_0.net58 0.09533f
C733 a_2739_20140# a_3273_20185# 0.35097f
C734 a_2918_20140# a_3425_20244# 0.21226f
C735 sar9b_0._00_ a_3166_20145# 0.13532f
C736 sar9b_0.net27 a_13011_20574# 0.04061f
C737 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.24199f
C738 sar9b_0.net38 a_9323_28371# 0.03711f
C739 a_10402_25094# a_10742_25087# 0.24088f
C740 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[7] 4.16011f
C741 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.17533f
C742 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.28523f
C743 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.3545f
C744 a_8438_23755# sar9b_0.net57 0.02145f
C745 a_13011_17910# sar9b_0.net27 0.03831f
C746 a_10644_16791# a_10410_17846# 0.01861f
C747 a_10926_17021# sar9b_0.net6 0.05497f
C748 a_5506_26802# a_5711_26851# 0.09983f
C749 sar9b_0.net43 a_9935_24187# 0.09338f
C750 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[5] 0.01482f
C751 VDPWR a_6954_27466# 0.83781f
C752 sar9b_0.net49 a_9154_20142# 0.09704f
C753 a_4011_22488# a_3027_22138# 0.08669f
C754 sar9b_0.net6 a_6634_18206# 0.09307f
C755 a_10227_18142# sar9b_0.net73 0.11717f
C756 sar9b_0.net40 single_9b_cdac_1.SW[7] 0.05122f
C757 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C758 single_9b_cdac_1.cdac_sw_9b_0.S[8] ua[0] 16.2977f
C759 a_3540_27045# a_3156_26115# 0.15019f
C760 a_4011_22488# sar9b_0.net65 0.01096f
C761 a_9930_20510# a_8970_20510# 0.03529f
C762 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[7] 0.02052f
C763 a_4922_20857# a_4886_21124# 0.01114f
C764 a_9126_19131# sar9b_0.net37 0.058f
C765 a_10218_20806# a_10402_21098# 0.44532f
C766 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.22879f
C767 sar9b_0.net32 sar9b_0.net26 0.27199f
C768 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C769 a_3521_24240# sar9b_0.clk_div_0.COUNT\[1\] 0.01149f
C770 VDPWR a_9930_20510# 0.34995f
C771 sar9b_0.net55 sar9b_0.net54 0.51028f
C772 sar9b_0.net6 sar9b_0.net5 0.134f
C773 sar9b_0.net42 a_10482_25831# 0.02488f
C774 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.15242f
C775 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[4] 0.06019f
C776 VDPWR a_10926_17021# 0.26037f
C777 a_10166_3438# a_10254_2858# 0.99857f
C778 uio_out[0] ui_in[0] 0.06786f
C779 VDPWR a_9942_24806# 0.28868f
C780 a_10553_18922# a_10830_19068# 0.09983f
C781 single_9b_cdac_0.cdac_sw_9b_0.S[5] a_38738_26999# 0.59531f
C782 single_9b_cdac_0.cdac_sw_9b_0.S[6] th_dif_sw_0.VCN 3.33405f
C783 a_4934_22432# sar9b_0.net64 0.25605f
C784 a_7638_23474# sar9b_0.net62 0.01517f
C785 a_9472_18823# a_9900_19047# 0.01872f
C786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.07579f
C787 sar9b_0.net40 sar9b_0.net26 0.02504f
C788 VDPWR a_6634_18206# 0.28909f
C789 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.26625f
C790 VDPWR a_10859_26330# 0.42645f
C791 a_9634_17478# a_10410_17846# 0.3578f
C792 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.SW[8] 0.17661f
C793 sar9b_0.net26 a_11842_19766# 0.02027f
C794 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.10429f
C795 a_48343_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.23864f
C796 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[0] 0.02356f
C797 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.28813f
C798 sar9b_0.net40 a_6534_27123# 0.03801f
C799 sar9b_0.net26 sar9b_0.net51 0.02947f
C800 a_5682_23444# a_5823_23477# 0.27388f
C801 a_5506_17478# a_6282_17846# 0.3578f
C802 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.38397f
C803 VDPWR a_7890_26108# 0.33944f
C804 a_10227_18142# sar9b_0.net48 0.02398f
C805 tdc_0.phase_detector_0.INN a_15400_11316# 0.02778f
C806 a_11178_27466# single_9b_cdac_0.SW[5] 0.03553f
C807 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[1] 4.15038f
C808 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C809 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.3196f
C810 sar9b_0._11_ sar9b_0.net10 0.01541f
C811 sar9b_0.net30 clk 0.0304f
C812 sar9b_0._02_ sar9b_0.net4 0.02372f
C813 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.03729f
C814 a_7092_19455# a_7097_19795# 0.44098f
C815 single_9b_cdac_0.SW[2] a_54032_26990# 0.18991f
C816 a_21684_3438# th_dif_sw_0.th_sw_1.CKB 0.03405f
C817 VDPWR sar9b_0.net5 1.99906f
C818 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] 3.10218f
C819 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.95338f
C820 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[3] 0.026f
C821 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C822 sar9b_0.net36 a_10937_25582# 0.02011f
C823 a_8115_28566# uo_out[5] 0.03775f
C824 a_9546_24506# a_9730_24138# 0.43747f
C825 sar9b_0.net7 a_10218_20806# 0.06569f
C826 a_13011_27234# sar9b_0._06_ 0.21168f
C827 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.02666f
C828 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.42784f
C829 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[2] 0.01297f
C830 a_9270_24566# sar9b_0.net12 0.04846f
C831 sar9b_0._02_ sar9b_0.clk_div_0.COUNT\[2\] 0.09854f
C832 sar9b_0.net14 uo_out[1] 0.127f
C833 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.S[1] 16.8012f
C834 single_9b_cdac_1.SW[6] sar9b_0.net28 0.14409f
C835 VDPWR a_9323_28371# 0.43901f
C836 single_9b_cdac_0.SW[0] clk 0.23595f
C837 sar9b_0.net1 sar9b_0.net5 0.83129f
C838 a_11382_26138# sar9b_0.net12 0.03109f
C839 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C840 VDPWR a_12047_26517# 0.26706f
C841 a_5748_24381# a_6538_24506# 0.1263f
C842 a_11859_17910# single_9b_cdac_1.SW[4] 0.35232f
C843 a_8052_18123# a_8057_18463# 0.44098f
C844 a_5196_18116# a_5394_18116# 0.06623f
C845 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.38037f
C846 a_8052_16791# a_7602_16784# 0.03471f
C847 a_7404_16784# a_7743_16817# 0.07649f
C848 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 a_44418_17740# 0.14695f
C849 a_8940_27039# a_9279_27227# 0.07649f
C850 a_3454_22567# sar9b_0._12_ 0.02006f
C851 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.0303f
C852 sar9b_0.net24 sar9b_0.cyclic_flag_0.FINAL 0.01327f
C853 a_10218_27466# sar9b_0.net45 0.24807f
C854 clk a_14871_9671# 0.36908f
C855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C856 a_11382_22142# a_11842_22430# 0.26257f
C857 a_11178_20806# sar9b_0.net73 0.01344f
C858 sar9b_0.net58 sar9b_0.net60 0.88421f
C859 a_10932_25713# a_11214_25728# 0.06034f
C860 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.17461f
C861 sar9b_0.net32 sar9b_0.net53 0.15479f
C862 a_11722_25838# a_10937_25582# 0.26257f
C863 a_8982_21902# a_9442_21474# 0.26257f
C864 a_9258_21842# a_9647_21523# 0.05462f
C865 a_6282_17846# a_5322_17846# 0.03529f
C866 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A 2.29405f
C867 VDPWR a_11430_24931# 0.26219f
C868 a_9126_23599# sar9b_0.net54 0.05162f
C869 a_10506_23174# sar9b_0.net38 0.02378f
C870 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCN 1.01731f
C871 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] 0.12898f
C872 sar9b_0._07_ a_4072_19474# 0.1462f
C873 sar9b_0.net74 sar9b_0.net38 0.03312f
C874 sar9b_0.net32 uo_out[2] 0.09101f
C875 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.3196f
C876 VDPWR a_5846_26950# 0.20642f
C877 sar9b_0._07_ sar9b_0.net71 0.05408f
C878 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0303f
C879 sar9b_0.net9 sar9b_0.net39 0.52789f
C880 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[7] 0.24198f
C881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.26942f
C882 sar9b_0.net63 sar9b_0._02_ 0.07961f
C883 a_7188_22119# a_7978_22202# 0.1263f
C884 a_6738_22112# a_7193_22459# 0.3578f
C885 sar9b_0.net38 a_9942_20810# 0.01655f
C886 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.62443f
C887 a_5374_20145# a_5481_20185# 0.14439f
C888 sar9b_0.net42 a_10506_24506# 0.01765f
C889 sar9b_0._08_ a_4072_19474# 0.09389f
C890 sar9b_0.net10 sar9b_0.net39 0.16291f
C891 sar9b_0.net61 sar9b_0.net39 0.42188f
C892 sar9b_0._09_ sar9b_0.net46 0.01177f
C893 sar9b_0._08_ sar9b_0.net71 0.35019f
C894 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.27713f
C895 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.22352f
C896 sar9b_0.net60 sar9b_0.net37 0.02643f
C897 a_12870_19603# sar9b_0.net50 0.17286f
C898 sar9b_0.net56 a_9363_20826# 0.12663f
C899 sar9b_0.net42 sar9b_0.net27 0.03289f
C900 a_8691_28566# a_8883_27466# 0.01221f
C901 sar9b_0._10_ sar9b_0.net57 0.02676f
C902 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.06503f
C903 a_10644_16791# a_11008_17491# 0.0165f
C904 sar9b_0.net42 single_9b_cdac_0.SW[5] 0.01977f
C905 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C906 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 1.71649f
C907 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.17533f
C908 single_9b_cdac_1.SW[3] th_dif_sw_0.VCN 0.09454f
C909 a_8345_26455# a_8340_26115# 0.43491f
C910 VDPWR sar9b_0.net54 3.92712f
C911 sar9b_0._17_ clk 0.03014f
C912 sar9b_0.net40 a_6562_25094# 0.02042f
C913 a_8074_20870# sar9b_0.net9 0.16977f
C914 sar9b_0.net33 single_9b_cdac_0.SW[7] 0.01742f
C915 single_9b_cdac_1.SW[4] sar9b_0.net2 0.03719f
C916 a_10995_28566# uo_out[2] 0.42572f
C917 a_8098_18810# sar9b_0.net61 0.02618f
C918 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C919 a_4211_19474# a_4072_19474# 0.02538f
C920 sar9b_0.net60 a_6137_23791# 0.02305f
C921 sar9b_0.net8 a_11382_19478# 0.03762f
C922 sar9b_0.net36 single_9b_cdac_1.SW[2] 0.1913f
C923 a_10859_26330# a_11382_26138# 0.04056f
C924 single_9b_cdac_1.SW[5] th_dif_sw_0.CK 0.23096f
C925 a_9494_20290# sar9b_0.net51 0.05999f
C926 a_9472_18823# sar9b_0.net5 0.02035f
C927 sar9b_0.net23 sar9b_0.net59 1.32079f
C928 a_8074_20870# sar9b_0.net61 0.0249f
C929 sar9b_0.net1 sar9b_0.net54 0.49885f
C930 sar9b_0.net19 a_5322_27170# 0.02142f
C931 a_8874_23470# a_9472_23805# 0.06623f
C932 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[0] 0.01887f
C933 a_6678_27470# a_6954_27466# 0.1263f
C934 sar9b_0.net58 a_5506_26802# 0.08623f
C935 a_10218_24802# a_10482_25831# 0.02278f
C936 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.SW[7] 0.05167f
C937 sar9b_0.net13 a_11776_25137# 0.29958f
C938 a_10402_27758# a_11430_27595# 0.07826f
C939 th_dif_sw_0.CKB clk 0.11297f
C940 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C941 VDPWR a_10035_19474# 0.46118f
C942 sar9b_0.net35 sar9b_0.cyclic_flag_0.FINAL 0.0808f
C943 sar9b_0.net8 sar9b_0.net38 0.02476f
C944 sar9b_0.net7 sar9b_0.net39 0.0839f
C945 sar9b_0.net35 sar9b_0.net15 0.01154f
C946 a_18214_3039# dw_17224_1400# 1.98311f
C947 a_6307_27584# sar9b_0.net36 0.04789f
C948 a_10218_20806# a_10607_21189# 0.06034f
C949 sar9b_0.net44 sar9b_0.net19 0.14271f
C950 uo_out[5] uo_out[6] 2.98352f
C951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.CF[5] 0.03484f
C952 VDPWR a_9132_7271# 1.60705f
C953 sar9b_0._13_ a_4467_24162# 0.11876f
C954 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.24223f
C955 sar9b_0.net53 sar9b_0.net62 0.14142f
C956 clk a_15151_10456# 0.19995f
C957 sar9b_0.net43 sar9b_0.net73 0.14358f
C958 sar9b_0.net21 uo_out[6] 0.34168f
C959 a_8052_16791# sar9b_0.net5 0.21543f
C960 single_9b_cdac_1.cdac_sw_9b_0.S[4] th_dif_sw_0.VCP 13.5521f
C961 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C962 sar9b_0.net18 a_3370_27769# 0.02082f
C963 sar9b_0.net55 sar9b_0._02_ 0.49529f
C964 sar9b_0._18_ sar9b_0.net57 0.25105f
C965 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS th_dif_sw_0.VCP 0.14643f
C966 VDPWR a_62748_16877# 1.81495f
C967 a_15265_9613# th_dif_sw_0.VCP 0.10972f
C968 uio_in[4] uio_in[3] 0.03102f
C969 a_11382_26138# a_12047_26517# 0.19065f
C970 th_dif_sw_0.CKB single_9b_cdac_1.SW[0] 0.0171f
C971 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42784f
C972 single_9b_cdac_0.SW[5] a_39616_26990# 0.18991f
C973 sar9b_0._01_ sar9b_0.net57 0.02763f
C974 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.12898f
C975 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[1] 0.2176f
C976 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[0] 0.02149f
C977 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.17533f
C978 VDPWR a_10506_23174# 0.8367f
C979 single_9b_cdac_0.SW[8] ua[0] 0.20384f
C980 a_3206_22432# sar9b_0.net70 0.04299f
C981 VDPWR sar9b_0.net74 1.07986f
C982 a_8019_17910# sar9b_0.net35 0.16492f
C983 a_5506_26802# sar9b_0.net37 0.11789f
C984 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.clknet_0_CLK 0.08397f
C985 sar9b_0.net64 sar9b_0._07_ 0.04413f
C986 sar9b_0.net9 sar9b_0.net36 0.33969f
C987 sar9b_0.net14 a_13164_28398# 0.14522f
C988 VDPWR a_9942_20810# 0.29503f
C989 single_9b_cdac_0.cdac_sw_9b_0.S[7] th_dif_sw_0.VCN 1.61586f
C990 VDPWR sar9b_0.net31 1.59832f
C991 sar9b_0._10_ a_4496_20468# 0.16691f
C992 a_2940_25096# sar9b_0._16_ 0.11593f
C993 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95338f
C994 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C995 a_12588_16784# a_13011_16810# 0.05125f
C996 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36044f
C997 sar9b_0.net10 sar9b_0.net36 0.03634f
C998 sar9b_0.net36 sar9b_0.net61 0.03284f
C999 sar9b_0.net42 single_9b_cdac_1.SW[7] 0.01299f
C1000 sar9b_0.net36 a_10402_21098# 0.0105f
C1001 sar9b_0.net38 sar9b_0.net34 0.38358f
C1002 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.3601f
C1003 a_9802_26815# a_9588_27045# 0.05022f
C1004 a_10858_17113# a_10926_17021# 0.35559f
C1005 sar9b_0.net44 a_3161_27787# 0.02151f
C1006 sar9b_0.net8 sar9b_0.net6 0.09366f
C1007 sar9b_0.net42 a_11382_23474# 0.02429f
C1008 a_10742_25087# sar9b_0.net12 0.06525f
C1009 single_9b_cdac_0.SW[5] sar9b_0.net14 0.06325f
C1010 a_10553_18922# a_10098_19171# 0.3578f
C1011 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C1012 sar9b_0._05_ a_3027_21906# 0.07466f
C1013 sar9b_0.net41 a_11859_17910# 0.05709f
C1014 a_5460_28377# uo_out[6] 0.03666f
C1015 a_2508_20780# a_2739_20140# 0.01678f
C1016 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02784f
C1017 sar9b_0.net68 a_5196_24776# 0.14653f
C1018 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[6] 0.01482f
C1019 sar9b_0.net42 sar9b_0.net26 0.59576f
C1020 sar9b_0.net60 sar9b_0.net57 0.11607f
C1021 sar9b_0.net8 a_8970_20510# 0.23591f
C1022 uo_out[0] uo_out[1] 3.57901f
C1023 sar9b_0.net30 a_11658_26134# 0.01536f
C1024 a_6414_23681# sar9b_0.net11 0.02893f
C1025 a_4072_19474# a_3991_19768# 0.03072f
C1026 a_3795_19512# a_4292_19768# 0.02251f
C1027 tdc_0.phase_detector_0.pd_out_0.B tdc_0.RDY 0.0496f
C1028 a_5682_23444# sar9b_0.net54 0.24995f
C1029 VDPWR a_11859_21906# 0.45768f
C1030 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[5] 4.15421f
C1031 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C1032 a_10662_17799# sar9b_0.net48 0.1748f
C1033 sar9b_0.net52 single_9b_cdac_0.SW[4] 0.35739f
C1034 VDPWR sar9b_0.net8 1.26787f
C1035 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.SW[0] 0.22983f
C1036 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.net4 0.27294f
C1037 sar9b_0.net69 sar9b_0.clk_div_0.COUNT\[1\] 0.04869f
C1038 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.45521f
C1039 VDPWR a_7926_23234# 0.30357f
C1040 sar9b_0.net7 sar9b_0.net36 0.02886f
C1041 sar9b_0.net40 a_6922_23534# 0.01201f
C1042 a_9996_16784# sar9b_0.net27 0.02177f
C1043 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.27803f
C1044 clk single_9b_cdac_1.SW[0] 0.21166f
C1045 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[2] 0.34042f
C1046 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.CF[3] 0.01346f
C1047 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24495f
C1048 a_8554_26437# sar9b_0.cyclic_flag_0.FINAL 0.06206f
C1049 a_7306_19777# sar9b_0.net40 0.02675f
C1050 sar9b_0.net8 sar9b_0.net1 0.02481f
C1051 a_8874_19178# sar9b_0.net48 0.29136f
C1052 sar9b_0.net24 a_9593_26914# 0.11222f
C1053 sar9b_0.net49 a_9258_21842# 0.19249f
C1054 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.71729f
C1055 sar9b_0.clk_div_0.COUNT\[3\] a_4812_21738# 0.29499f
C1056 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.clk_div_0.COUNT\[2\] 0.31022f
C1057 a_11030_22954# clk 0.01673f
C1058 sar9b_0.net33 a_12618_26134# 0.07184f
C1059 a_11842_26426# sar9b_0.net27 0.01173f
C1060 a_10742_27751# a_10607_27849# 0.35559f
C1061 sar9b_0.net27 a_13216_19809# 0.01127f
C1062 a_12684_20379# sar9b_0.net5 0.051f
C1063 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 ua[0] 0.12076f
C1064 a_8098_18810# a_8438_18958# 0.24088f
C1065 sar9b_0.net32 sar9b_0.net30 1.27934f
C1066 sar9b_0._18_ sar9b_0.clk_div_0.COUNT\[1\] 0.17343f
C1067 a_8874_23470# sar9b_0.net37 0.02487f
C1068 sar9b_0.net49 sar9b_0.net26 0.02489f
C1069 single_9b_cdac_1.SW[2] a_9450_17846# 0.01334f
C1070 sar9b_0.net31 sar9b_0.net29 0.0246f
C1071 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C1072 VDPWR a_2847_27473# 0.29759f
C1073 sar9b_0.net56 single_9b_cdac_1.SW[0] 0.04752f
C1074 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1075 single_9b_cdac_0.SW[1] th_dif_sw_0.VCN 0.09453f
C1076 sar9b_0._04_ sar9b_0._12_ 0.12021f
C1077 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 1.56111f
C1078 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C1079 single_9b_cdac_1.SW[8] single_9b_cdac_1.CF[0] 3.87975f
C1080 a_8691_28566# a_9323_28371# 0.0245f
C1081 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.45521f
C1082 VDPWR sar9b_0.net34 0.38274f
C1083 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.69086f
C1084 a_10402_25094# sar9b_0.net57 0.01621f
C1085 single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.10499f
C1086 VDPWR sar9b_0._02_ 0.67644f
C1087 sar9b_0._18_ a_3371_23106# 0.05658f
C1088 a_5506_17478# sar9b_0.net46 0.1904f
C1089 a_8694_20570# sar9b_0.net37 0.01919f
C1090 a_8334_17021# sar9b_0.net61 0.06633f
C1091 sar9b_0.net27 sar9b_0.net11 0.03459f
C1092 sar9b_0._12_ clk 0.1358f
C1093 a_6579_18832# a_5844_18123# 0.01182f
C1094 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.71649f
C1095 sar9b_0.cyclic_flag_0.FINAL a_8940_27039# 0.01546f
C1096 sar9b_0.net23 a_7890_26108# 0.05346f
C1097 a_7374_19685# sar9b_0.net10 0.04605f
C1098 sar9b_0.net41 sar9b_0.net2 0.36918f
C1099 sar9b_0.net74 a_11382_26138# 0.17525f
C1100 sar9b_0.net48 sar9b_0.net4 0.02286f
C1101 a_9472_23805# sar9b_0.net12 0.27258f
C1102 sar9b_0.net60 a_4496_20468# 0.09564f
C1103 VDPWR a_3156_26115# 0.78981f
C1104 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[0\] 0.2165f
C1105 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.28523f
C1106 a_8334_18353# sar9b_0.net61 0.02726f
C1107 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[2] 0.21903f
C1108 single_9b_cdac_0.SW[7] ua[0] 0.25507f
C1109 sar9b_0.net42 sar9b_0.net53 0.62196f
C1110 a_12870_19603# sar9b_0.net27 0.0267f
C1111 sar9b_0.net31 a_11382_26138# 0.01042f
C1112 a_10690_22806# sar9b_0.net42 0.01178f
C1113 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] 0.93526f
C1114 sar9b_0.net40 a_11658_19474# 0.07402f
C1115 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C1116 a_11842_18434# a_12870_18271# 0.07826f
C1117 a_11658_19474# a_11842_19766# 0.44532f
C1118 sar9b_0.net38 a_10528_20155# 0.31876f
C1119 VDPWR a_6282_17846# 0.34765f
C1120 sar9b_0.net59 sar9b_0.net58 0.82667f
C1121 single_9b_cdac_0.SW[5] th_dif_sw_0.VCN 0.09454f
C1122 sar9b_0.net20 a_5151_28559# 0.06913f
C1123 a_5010_28495# a_5460_28377# 0.03432f
C1124 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[1\] 0.02478f
C1125 a_10803_19474# single_9b_cdac_1.SW[1] 0.35106f
C1126 sar9b_0.net58 a_3156_27447# 0.17605f
C1127 sar9b_0.net52 a_10623_25895# 0.21039f
C1128 sar9b_0.net31 a_11658_22138# 0.02838f
C1129 sar9b_0.net18 a_3946_27530# 0.02978f
C1130 VDPWR a_3438_26345# 0.27271f
C1131 VDPWR a_6783_19481# 0.27053f
C1132 VDPWR a_9935_24187# 0.26083f
C1133 a_3156_27447# a_2706_27440# 0.03471f
C1134 a_2508_27440# a_2847_27473# 0.07649f
C1135 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.11216f
C1136 a_13011_24802# single_9b_cdac_1.CF[7] 0.05123f
C1137 a_10166_3438# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.16499f
C1138 a_14871_9671# a_15265_9613# 0.12812f
C1139 sar9b_0.net61 a_9450_17846# 0.04773f
C1140 sar9b_0.net46 sar9b_0.net4 0.06536f
C1141 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.42784f
C1142 a_7566_21017# a_7284_20787# 0.05462f
C1143 tdc_0.OUTN tdc_0.phase_detector_0.pd_out_0.A 0.11925f
C1144 sar9b_0.net61 single_9b_cdac_1.SW[2] 0.04325f
C1145 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR 3.27795f
C1146 a_7638_23474# sar9b_0.net11 0.23589f
C1147 a_10644_16791# a_10649_17131# 0.43869f
C1148 single_9b_cdac_1.SW[4] sar9b_0.net39 0.01225f
C1149 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[7] 0.01482f
C1150 VDPWR a_7743_18149# 0.25964f
C1151 VDPWR ua[4] 1.80222f
C1152 a_9363_20826# sar9b_0.net51 0.24159f
C1153 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[3] 0.31534f
C1154 VDPWR a_8057_17131# 0.24259f
C1155 sar9b_0.net21 sar9b_0.net45 0.04091f
C1156 VDPWR a_12182_22423# 0.19338f
C1157 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.24399f
C1158 a_8166_27595# sar9b_0.net45 0.03834f
C1159 sar9b_0.net58 a_4330_27170# 0.28291f
C1160 sar9b_0.net48 a_6058_18445# 0.14602f
C1161 single_9b_cdac_1.cdac_sw_9b_0.S[0] a_63626_17740# 0.22513f
C1162 a_8883_27466# a_9323_27662# 0.03138f
C1163 sar9b_0.net59 sar9b_0.net37 0.15299f
C1164 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.84426f
C1165 sar9b_0.net45 single_9b_cdac_0.SW[5] 0.0907f
C1166 a_5322_17846# sar9b_0.net46 0.23175f
C1167 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.10626f
C1168 sar9b_0.net36 a_10607_21189# 0.02616f
C1169 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.95338f
C1170 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.SW[2] 0.01427f
C1171 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.02632f
C1172 single_9b_cdac_0.SW[6] uo_out[4] 0.02556f
C1173 a_6738_22112# sar9b_0.net47 0.26419f
C1174 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.10626f
C1175 sar9b_0.net47 sar9b_0._07_ 0.17483f
C1176 sar9b_0.net54 a_6030_24396# 0.22581f
C1177 a_2739_20140# a_3723_20140# 0.08669f
C1178 sar9b_0._00_ a_3273_20185# 0.04988f
C1179 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.12898f
C1180 VDPWR a_12182_23755# 0.19519f
C1181 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.26942f
C1182 a_10378_27170# sar9b_0.net36 0.05314f
C1183 a_10402_25094# a_11178_24802# 0.3578f
C1184 a_13164_28398# uo_out[0] 0.0371f
C1185 single_9b_cdac_1.SW[1] ua[0] 0.15672f
C1186 VDPWR a_3425_20244# 0.10699f
C1187 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.42509f
C1188 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[0\] 0.01636f
C1189 a_26951_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C1190 single_9b_cdac_0.SW[4] a_43540_26999# 0.28324f
C1191 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.VCN 0.21849f
C1192 sar9b_0.net40 sar9b_0._17_ 0.02904f
C1193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 a_54032_17740# 0.14695f
C1194 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[8] 1.89002f
C1195 a_5711_26851# a_5846_26950# 0.35559f
C1196 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[5] 0.01887f
C1197 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.1236f
C1198 a_11434_16874# sar9b_0.net6 0.07229f
C1199 a_3370_26437# sar9b_0.net59 0.14542f
C1200 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C1201 a_11382_23474# sar9b_0.net11 0.04486f
C1202 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[2] 0.22161f
C1203 VDPWR a_7138_27758# 0.2246f
C1204 single_9b_cdac_1.SW[0] a_63626_17740# 0.18991f
C1205 sar9b_0.net49 a_9494_20290# 0.1204f
C1206 sar9b_0.net43 a_8940_24402# 0.06556f
C1207 a_8622_26345# a_9130_26198# 0.19065f
C1208 a_4330_27170# sar9b_0.net37 0.17592f
C1209 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C1210 sar9b_0.net52 sar9b_0.net2 0.02335f
C1211 a_8303_23853# sar9b_0.net11 0.02489f
C1212 a_3219_22860# sar9b_0.clknet_1_1__leaf_CLK 0.01128f
C1213 sar9b_0.net9 sar9b_0.net10 0.65359f
C1214 sar9b_0.net9 sar9b_0.net61 0.58982f
C1215 single_9b_cdac_0.SW[5] uo_out[0] 0.08425f
C1216 a_10470_21795# sar9b_0.net38 0.02191f
C1217 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.net65 0.16477f
C1218 a_7638_23474# a_8098_23762# 0.26257f
C1219 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C1220 VDPWR a_3027_21906# 0.29917f
C1221 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.01751f
C1222 single_9b_cdac_0.SW[2] a_13011_27234# 0.04188f
C1223 sar9b_0.net10 sar9b_0.net61 0.02017f
C1224 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.04988f
C1225 th_dif_sw_0.VCN single_9b_cdac_1.SW[7] 0.09453f
C1226 a_9900_19047# sar9b_0.net37 0.27085f
C1227 sar9b_0.net26 sar9b_0.net11 0.03443f
C1228 a_10218_20806# a_11430_20935# 0.07766f
C1229 a_5465_28246# a_5674_28147# 0.24088f
C1230 a_5460_28377# sar9b_0.net45 0.20577f
C1231 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 2.82171f
C1232 VDPWR a_10528_20155# 0.20299f
C1233 a_11915_27039# sar9b_0.net52 0.03127f
C1234 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.02149f
C1235 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C1236 a_11382_19478# sar9b_0.net73 0.17436f
C1237 VDPWR a_11434_16874# 0.27783f
C1238 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10254_2858# 1.3306f
C1239 a_10548_19053# sar9b_0.net73 0.01967f
C1240 a_9900_19047# a_10098_19171# 0.06623f
C1241 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 ua[0] 0.12088f
C1242 a_7978_22202# sar9b_0.net62 0.01108f
C1243 a_6282_27170# a_5322_27170# 0.03529f
C1244 a_9974_17626# a_10410_17846# 0.16939f
C1245 sar9b_0.net60 a_6378_24802# 0.01004f
C1246 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.19266f
C1247 a_8386_22806# a_9414_23127# 0.07826f
C1248 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[4] 0.42014f
C1249 sar9b_0.net43 a_10506_24506# 0.07702f
C1250 a_6132_23451# a_6414_23681# 0.05462f
C1251 a_5823_23477# a_6137_23791# 0.07826f
C1252 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[6] 2.01497f
C1253 a_5846_17626# a_6282_17846# 0.16939f
C1254 a_10218_27466# sar9b_0.net38 0.01643f
C1255 VDPWR a_5196_19448# 0.22579f
C1256 sar9b_0.net51 a_6252_19074# 0.05727f
C1257 a_5046_27230# sar9b_0.net39 0.19915f
C1258 VDPWR a_8345_26455# 0.25217f
C1259 VDPWR a_43540_16877# 1.81495f
C1260 single_9b_cdac_0.cdac_sw_9b_0.S[4] a_43540_26999# 0.59531f
C1261 a_7404_17715# sar9b_0.net56 0.02799f
C1262 sar9b_0.net38 sar9b_0.net73 0.26685f
C1263 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.42509f
C1264 a_5235_27466# uo_out[7] 0.39295f
C1265 sar9b_0.net44 a_6282_27170# 0.02958f
C1266 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.42016f
C1267 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.3196f
C1268 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[8] 0.31534f
C1269 sar9b_0.net7 sar9b_0.net9 0.36253f
C1270 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.28813f
C1271 a_13011_19242# sar9b_0.net27 0.02433f
C1272 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.0303f
C1273 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP a_43540_16877# 0.04592f
C1274 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26955f
C1275 sar9b_0.net13 sar9b_0.net27 0.04207f
C1276 sar9b_0.net7 sar9b_0.net61 0.28001f
C1277 a_8303_23853# a_8098_23762# 0.09983f
C1278 a_9270_24566# a_9935_24187# 0.19065f
C1279 a_9546_24506# a_10070_24286# 0.04522f
C1280 sar9b_0.net7 a_10402_21098# 0.08721f
C1281 a_11466_23174# a_12064_22819# 0.06623f
C1282 a_10335_16817# sar9b_0.net6 0.04672f
C1283 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C1284 a_9730_24138# sar9b_0.net12 0.06386f
C1285 a_10548_19053# sar9b_0.net48 0.16225f
C1286 sar9b_0.net48 a_9839_17527# 0.2029f
C1287 VDPWR a_13067_27662# 0.51166f
C1288 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02666f
C1289 sar9b_0.net36 sar9b_0.cyclic_flag_0.FINAL 0.23039f
C1290 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.22875f
C1291 sar9b_0.net27 a_12560_27128# 0.02362f
C1292 a_5844_18123# a_5535_18149# 0.07766f
C1293 single_9b_cdac_1.cdac_sw_9b_0.S[5] a_38738_16877# 0.59531f
C1294 a_8052_16791# a_8057_17131# 0.44098f
C1295 a_7602_16784# a_7743_16817# 0.27388f
C1296 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1297 sar9b_0.net40 clk 0.03834f
C1298 single_9b_cdac_1.SW[0] a_9174_17906# 0.04125f
C1299 a_2893_24992# sar9b_0.net68 0.07409f
C1300 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.43767f
C1301 sar9b_0.net48 sar9b_0.net38 0.55083f
C1302 a_16222_11316# tdc_0.phase_detector_0.pd_out_0.A 0.48692f
C1303 a_9138_27163# a_9588_27045# 0.03432f
C1304 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.02666f
C1305 a_4011_22488# sar9b_0._12_ 0.04991f
C1306 sar9b_0.net56 a_9174_17906# 0.04252f
C1307 tdc_0.RDY tdc_0.OUTN 0.07358f
C1308 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.12898f
C1309 VDPWR a_10470_21795# 0.2699f
C1310 a_8031_26141# sar9b_0.net59 0.20849f
C1311 clk a_15265_9613# 0.01191f
C1312 VDPWR a_10335_16817# 0.2584f
C1313 sar9b_0.clknet_1_0__leaf_CLK a_3166_20145# 0.02652f
C1314 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[6] 4.16175f
C1315 sar9b_0.net52 a_7914_23470# 0.15191f
C1316 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C1317 a_11658_22138# a_12182_22423# 0.05022f
C1318 sar9b_0.net6 sar9b_0.net73 0.44042f
C1319 sar9b_0._07_ sar9b_0.net57 1.15961f
C1320 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] 1.15133f
C1321 sar9b_0.net53 sar9b_0.net11 0.33023f
C1322 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[2\] 1.2616f
C1323 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.03729f
C1324 a_10690_22806# sar9b_0.net11 0.12946f
C1325 a_11382_19478# sar9b_0.net50 0.23074f
C1326 a_10470_21795# a_10218_21842# 0.27388f
C1327 a_10548_19053# sar9b_0.net50 0.02815f
C1328 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.SW[3] 0.01382f
C1329 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.07517f
C1330 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.7611f
C1331 single_9b_cdac_1.cdac_sw_9b_0.S[6] th_dif_sw_0.VCP 3.33405f
C1332 VDPWR a_11776_25137# 0.19971f
C1333 a_3014_24136# a_3262_24141# 0.05308f
C1334 a_2835_24136# a_3521_24240# 0.27693f
C1335 a_9472_23805# sar9b_0.net54 0.08291f
C1336 VDPWR sar9b_0.clk_div_0.COUNT\[0\] 0.52537f
C1337 sar9b_0.net15 a_5844_18123# 0.0119f
C1338 sar9b_0.net24 uo_out[3] 0.06521f
C1339 a_5331_16810# sar9b_0.net4 0.1431f
C1340 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.12431f
C1341 sar9b_0.net56 sar9b_0.net40 0.02195f
C1342 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.CF[2] 0.10503f
C1343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.12358f
C1344 sar9b_0.net43 a_5962_24151# 0.02064f
C1345 sar9b_0._08_ sar9b_0.net57 0.62749f
C1346 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24779f
C1347 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.05472f
C1348 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.28523f
C1349 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.01003f
C1350 VDPWR a_16185_13034# 0.19332f
C1351 sar9b_0.net41 sar9b_0.net39 0.25189f
C1352 sar9b_0.net56 sar9b_0.net51 0.81695f
C1353 sar9b_0.net17 uio_out[1] 0.1629f
C1354 a_10218_27466# VDPWR 0.8229f
C1355 sar9b_0.net42 a_11104_24151# 0.30428f
C1356 a_6867_16810# sar9b_0.net27 0.04386f
C1357 a_33936_16877# single_9b_cdac_1.SW[6] 0.28324f
C1358 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[7] 0.21593f
C1359 a_6540_22112# a_6879_22145# 0.07649f
C1360 a_11430_20935# sar9b_0.net39 0.02333f
C1361 VDPWR sar9b_0.net73 1.85779f
C1362 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.81428f
C1363 a_5823_23477# sar9b_0.net57 0.0298f
C1364 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.62443f
C1365 a_13011_19242# single_9b_cdac_1.SW[7] 0.36033f
C1366 a_6879_22145# sar9b_0.net39 0.04509f
C1367 sar9b_0.net43 a_5439_24563# 0.02732f
C1368 a_9323_28371# a_9323_27662# 0.0246f
C1369 a_7188_22119# sar9b_0.net62 0.04051f
C1370 sar9b_0.net48 sar9b_0.net6 1.12384f
C1371 a_24332_26999# single_9b_cdac_0.SW[8] 0.28324f
C1372 a_6130_20239# sar9b_0.net15 0.12036f
C1373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C1374 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02513f
C1375 sar9b_0.net5 sar9b_0.net37 0.14722f
C1376 th_dif_sw_0.CK a_11382_18146# 0.05375f
C1377 sar9b_0.net1 sar9b_0.net73 0.94195f
C1378 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.45521f
C1379 dw_12589_1395# th_dif_sw_0.CK 0.01665f
C1380 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[1] 0.22097f
C1381 clk sar9b_0.net62 0.06683f
C1382 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.69086f
C1383 sar9b_0.net12 sar9b_0.net57 0.27108f
C1384 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[1] 1.81416f
C1385 sar9b_0.net27 sar9b_0.net4 0.23295f
C1386 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.19147f
C1387 sar9b_0._10_ a_5581_19664# 0.13526f
C1388 a_8438_18958# sar9b_0.net61 0.0222f
C1389 sar9b_0.net29 a_13067_27662# 0.10621f
C1390 sar9b_0.net63 a_6414_23681# 0.04702f
C1391 a_6052_19792# a_5581_19664# 0.01114f
C1392 VDPWR a_3219_22860# 0.26196f
C1393 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C1394 sar9b_0.net33 sar9b_0.net12 0.05295f
C1395 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[7] 0.01471f
C1396 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38317f
C1397 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[0] 0.45278f
C1398 VDPWR a_6975_20813# 0.25935f
C1399 a_5298_24499# a_5962_24151# 0.16939f
C1400 sar9b_0.net60 a_3922_20239# 0.01343f
C1401 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.95338f
C1402 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.26707f
C1403 a_10218_24802# a_10932_25713# 0.04762f
C1404 sar9b_0.net58 a_5846_26950# 0.13488f
C1405 a_6678_27470# a_7138_27758# 0.26257f
C1406 sar9b_0._05_ sar9b_0.clknet_0_CLK 0.03678f
C1407 a_10742_27751# a_11178_27466# 0.16939f
C1408 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0313f
C1409 a_8591_22855# sar9b_0.net11 0.05189f
C1410 sar9b_0.net27 a_5322_17846# 0.0316f
C1411 VDPWR sar9b_0.net48 5.69977f
C1412 a_8202_23174# sar9b_0.net54 0.18332f
C1413 sar9b_0.net23 sar9b_0.net34 0.07163f
C1414 sar9b_0.net46 sar9b_0.net6 0.09629f
C1415 a_4136_25584# a_4293_25852# 0.21226f
C1416 a_10402_21098# a_10607_21189# 0.09983f
C1417 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 2.82181f
C1418 sar9b_0.net56 sar9b_0.net62 0.01262f
C1419 sar9b_0.net50 sar9b_0.net6 0.16111f
C1420 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.02149f
C1421 VDPWR th_dif_sw_0.th_sw_1.CK 2.01535f
C1422 a_9942_27470# sar9b_0.net59 0.22307f
C1423 a_7602_18116# sar9b_0.net5 0.04179f
C1424 a_5298_24499# a_5439_24563# 0.27388f
C1425 single_9b_cdac_1.SW[3] sar9b_0.net6 0.2526f
C1426 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[2] 0.22184f
C1427 a_12618_18142# sar9b_0.net6 0.01945f
C1428 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.0303f
C1429 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38397f
C1430 a_7338_24802# a_6562_25094# 0.3578f
C1431 a_6767_25185# a_6378_24802# 0.06034f
C1432 a_9939_28566# sar9b_0.net38 0.04052f
C1433 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.6919f
C1434 sar9b_0.net1 sar9b_0.net48 0.20331f
C1435 a_13011_20806# a_13011_20574# 0.02551f
C1436 single_9b_cdac_0.SW[4] single_9b_cdac_0.SW[8] 0.03894f
C1437 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[1] 0.2162f
C1438 single_9b_cdac_0.SW[5] a_38738_26999# 0.28324f
C1439 single_9b_cdac_0.cdac_sw_9b_0.S[7] a_29134_26999# 0.59531f
C1440 a_11339_27039# sar9b_0.net31 0.19953f
C1441 th_dif_sw_0.VCN th_dif_sw_0.VCP 0.69759f
C1442 sar9b_0.net3 sar9b_0.net60 0.11243f
C1443 sar9b_0._11_ a_4947_20140# 0.14426f
C1444 VDPWR a_7498_21109# 0.19831f
C1445 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# 0.18915f
C1446 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.95338f
C1447 a_3561_22527# sar9b_0.clknet_1_1__leaf_CLK 0.04276f
C1448 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.84381f
C1449 sar9b_0.clknet_0_CLK sar9b_0.clknet_1_1__leaf_CLK 0.04779f
C1450 a_6484_22845# sar9b_0.clk_div_0.COUNT\[1\] 0.04883f
C1451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 3.10626f
C1452 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[1\] 1.08101f
C1453 a_5846_26950# sar9b_0.net37 0.0568f
C1454 single_9b_cdac_0.SW[6] a_33936_26999# 0.28324f
C1455 a_9363_20826# sar9b_0.net49 0.32854f
C1456 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.0303f
C1457 a_8334_17021# a_8842_16874# 0.19065f
C1458 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.6205f
C1459 VDPWR sar9b_0.net46 2.39016f
C1460 th_dif_sw_0.CK sar9b_0.net28 0.15795f
C1461 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 1.56012f
C1462 sar9b_0.net38 a_10482_25831# 0.01616f
C1463 VDPWR sar9b_0.net50 2.24819f
C1464 uo_out[2] uo_out[0] 0.01052f
C1465 a_7374_19685# a_7882_19538# 0.19065f
C1466 a_9930_20510# a_10182_20463# 0.27388f
C1467 sar9b_0.net41 sar9b_0.net36 0.03019f
C1468 VDPWR single_9b_cdac_1.SW[3] 2.54341f
C1469 a_8303_18859# a_7914_19178# 0.05462f
C1470 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[6] 0.01887f
C1471 a_4947_20140# a_5374_20145# 0.04602f
C1472 a_4496_20468# sar9b_0.clknet_1_0__leaf_CLK 0.10004f
C1473 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C1474 VDPWR a_12618_18142# 0.35481f
C1475 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C1476 a_7478_27751# sar9b_0.net60 0.13192f
C1477 sar9b_0.net55 a_6414_23681# 0.0176f
C1478 a_8970_20510# a_9154_20142# 0.43491f
C1479 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.6919f
C1480 sar9b_0.net7 a_10607_21189# 0.06928f
C1481 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[8] 0.05215f
C1482 sar9b_0.net1 sar9b_0.net46 0.42025f
C1483 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C1484 a_9802_26815# a_9870_27060# 0.35559f
C1485 VDPWR a_15400_11316# 0.52162f
C1486 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38702f
C1487 a_3371_23106# sar9b_0._07_ 0.18693f
C1488 a_9942_24806# sar9b_0.net57 0.04118f
C1489 sar9b_0.net17 a_2892_27039# 0.01295f
C1490 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1491 VDPWR a_9154_20142# 0.24213f
C1492 a_13067_27662# single_9b_cdac_0.SW[3] 0.02544f
C1493 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C1494 a_11178_24802# sar9b_0.net12 0.08132f
C1495 a_6252_20780# sar9b_0.net4 0.02886f
C1496 sar9b_0.net54 sar9b_0.net37 0.24974f
C1497 a_8334_18353# a_8842_18206# 0.19065f
C1498 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 2.82223f
C1499 sar9b_0._05_ a_4812_21738# 0.01191f
C1500 a_5439_24563# sar9b_0._15_ 0.06796f
C1501 a_10859_26330# sar9b_0.net33 0.22653f
C1502 sar9b_0.net1 a_9154_20142# 0.01157f
C1503 sar9b_0.net27 a_12870_26263# 0.0306f
C1504 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1505 a_8019_17910# single_9b_cdac_1.SW[2] 0.35523f
C1506 VDPWR uo_out[1] 0.933f
C1507 sar9b_0.net43 sar9b_0.net53 0.57297f
C1508 a_10182_20463# sar9b_0.net5 0.04725f
C1509 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[3] 0.22098f
C1510 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.38397f
C1511 a_5812_21028# sar9b_0._01_ 0.14953f
C1512 sar9b_0.net30 a_11842_26426# 0.01579f
C1513 a_6922_23534# sar9b_0.net11 0.05827f
C1514 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.38037f
C1515 a_6137_23791# sar9b_0.net54 0.06976f
C1516 a_7890_26108# a_8031_26141# 0.27388f
C1517 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] 1.15122f
C1518 sar9b_0.net44 a_3161_26455# 0.01837f
C1519 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.SW[6] 0.17155f
C1520 sar9b_0.net71 a_5196_19448# 0.14653f
C1521 sar9b_0.net13 sar9b_0.net53 0.0108f
C1522 a_5100_24375# sar9b_0.net39 0.0223f
C1523 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP 0.04344f
C1524 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.84061f
C1525 sar9b_0.net36 a_9593_26914# 0.11605f
C1526 a_21684_3438# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.63339f
C1527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[2] 0.31534f
C1528 a_3090_27163# a_3545_26914# 0.3578f
C1529 sar9b_0.net4 a_5443_19074# 0.31469f
C1530 sar9b_0.net43 a_9802_26815# 0.01853f
C1531 sar9b_0.net60 a_5151_28559# 0.02736f
C1532 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.02638f
C1533 a_9939_28566# VDPWR 0.44769f
C1534 a_11338_19178# sar9b_0.net42 0.02024f
C1535 a_10649_17131# single_9b_cdac_1.SW[1] 0.0197f
C1536 a_9472_18823# sar9b_0.net48 0.04471f
C1537 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR 0.38397f
C1538 sar9b_0.net33 a_12047_26517# 0.04976f
C1539 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07579f
C1540 sar9b_0.net35 sar9b_0.net44 0.01492f
C1541 a_16527_10454# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.09051f
C1542 single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR 4.1608f
C1543 VDPWR a_11436_17742# 0.21601f
C1544 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.11216f
C1545 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.42784f
C1546 sar9b_0.net13 a_6562_25094# 0.12325f
C1547 sar9b_0.net30 sar9b_0.net11 0.14416f
C1548 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.12898f
C1549 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.363f
C1550 a_8202_23174# a_7926_23234# 0.1263f
C1551 single_9b_cdac_0.SW[6] ua[0] 0.22043f
C1552 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[5] 0.244f
C1553 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.12358f
C1554 VDPWR a_10482_25831# 0.34041f
C1555 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.5604f
C1556 sar9b_0.net42 clk 0.03904f
C1557 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24399f
C1558 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.93403f
C1559 a_5812_21028# sar9b_0.net60 0.24213f
C1560 sar9b_0.net59 sar9b_0.net19 0.15362f
C1561 single_9b_cdac_1.SW[8] a_12618_19474# 0.02801f
C1562 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] 0.12898f
C1563 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C1564 sar9b_0.net52 sar9b_0.net36 0.10328f
C1565 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.69086f
C1566 sar9b_0.net38 uo_out[5] 0.25815f
C1567 a_8019_17910# sar9b_0.net61 0.01405f
C1568 a_11718_23127# sar9b_0.net53 0.17359f
C1569 sar9b_0._18_ a_3695_23038# 0.02716f
C1570 sar9b_0.net38 a_10506_24506# 0.02782f
C1571 a_10690_22806# a_11718_23127# 0.07826f
C1572 a_5846_17626# sar9b_0.net46 0.19277f
C1573 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.0303f
C1574 sar9b_0.net38 sar9b_0.net21 0.04603f
C1575 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.02149f
C1576 a_8842_16874# sar9b_0.net61 0.2111f
C1577 a_13011_23238# single_9b_cdac_1.CF[5] 0.35518f
C1578 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[2\] 0.26122f
C1579 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.71729f
C1580 a_7882_19538# sar9b_0.net61 0.01172f
C1581 a_7882_19538# sar9b_0.net10 0.05509f
C1582 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[4] 0.03897f
C1583 sar9b_0.net55 a_6444_19448# 0.01836f
C1584 VDPWR a_2847_26141# 0.31739f
C1585 a_5196_24776# sar9b_0.net39 0.03191f
C1586 sar9b_0.net36 sar9b_0.net22 0.02611f
C1587 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 1.71649f
C1588 single_9b_cdac_0.SW[0] th_dif_sw_0.VCN 0.09453f
C1589 sar9b_0.net19 a_4330_27170# 0.04522f
C1590 a_11030_22954# sar9b_0.net42 0.0141f
C1591 a_8052_16791# sar9b_0.net46 0.1629f
C1592 sar9b_0.net60 a_6282_27170# 0.04032f
C1593 sar9b_0.net40 a_12870_18271# 0.02062f
C1594 sar9b_0.net40 a_11842_19766# 0.1379f
C1595 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C1596 a_11658_19474# a_12870_19603# 0.07766f
C1597 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1598 sar9b_0.net40 sar9b_0.net51 0.02551f
C1599 sar9b_0.net32 a_10995_28566# 0.04889f
C1600 VDPWR a_6414_23681# 0.26663f
C1601 VDPWR a_6880_17491# 0.19624f
C1602 a_9162_23174# clk 0.02449f
C1603 sar9b_0.net8 sar9b_0.net37 0.15963f
C1604 sar9b_0.net16 sar9b_0._00_ 0.01551f
C1605 sar9b_0.net20 a_5465_28246# 0.10985f
C1606 sar9b_0.net15 a_6579_18832# 0.01202f
C1607 sar9b_0.net57 sar9b_0.net54 1.01482f
C1608 VDPWR a_3561_22527# 0.14464f
C1609 sar9b_0.net30 sar9b_0.net45 0.11616f
C1610 sar9b_0.net58 a_2847_27473# 0.17334f
C1611 sar9b_0.net52 a_10937_25582# 0.11747f
C1612 sar9b_0.net31 a_11842_22430# 0.01313f
C1613 VDPWR a_29134_16877# 1.81495f
C1614 VDPWR sar9b_0.clknet_0_CLK 2.46803f
C1615 VDPWR a_3946_26198# 0.30347f
C1616 sar9b_0.net41 single_9b_cdac_1.SW[2] 0.0369f
C1617 a_11722_25838# sar9b_0.net52 0.22698f
C1618 th_dif_sw_0.CK a_13216_18477# 0.04814f
C1619 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A a_54737_15495# 0.01076f
C1620 a_2835_24136# sar9b_0.net69 0.01995f
C1621 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C1622 a_2706_27440# a_2847_27473# 0.27388f
C1623 sar9b_0.net13 a_10932_25713# 0.23395f
C1624 a_3156_27447# a_3161_27787# 0.44098f
C1625 a_11146_25483# a_10937_25582# 0.24088f
C1626 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.03729f
C1627 a_12182_19759# single_9b_cdac_1.SW[8] 0.01333f
C1628 a_16331_9671# a_16357_9613# 0.12812f
C1629 a_14871_9671# th_dif_sw_0.VCN 0.11478f
C1630 a_6880_17491# sar9b_0.net1 0.01138f
C1631 a_8074_20870# a_7284_20787# 0.1263f
C1632 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[0] 0.74373f
C1633 single_9b_cdac_0.SW[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.24198f
C1634 VDPWR a_8940_24402# 0.29362f
C1635 sar9b_0.net67 a_4236_21738# 0.14162f
C1636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C1637 single_9b_cdac_0.SW[1] VDPWR 2.63243f
C1638 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.CF[3] 0.18985f
C1639 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96835f
C1640 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.42784f
C1641 a_10858_17113# sar9b_0.net48 0.12168f
C1642 sar9b_0.net18 uio_out[1] 0.0124f
C1643 VDPWR a_5331_16810# 0.25165f
C1644 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.6919f
C1645 single_9b_cdac_1.cdac_sw_9b_0.S[7] ua[0] 1.97892f
C1646 sar9b_0.net56 sar9b_0.net49 0.45655f
C1647 VDPWR a_12618_22138# 0.32654f
C1648 a_6250_28502# a_5465_28246# 0.26257f
C1649 sar9b_0.net25 a_12531_28566# 0.21118f
C1650 sar9b_0.net58 a_3156_26115# 0.01128f
C1651 a_3027_22138# sar9b_0._05_ 0.07932f
C1652 a_8512_27801# sar9b_0.net45 0.03235f
C1653 sar9b_0.net27 sar9b_0.net6 1.39158f
C1654 sar9b_0.net4 a_6562_25094# 0.01993f
C1655 a_9323_27662# sar9b_0.net34 0.21484f
C1656 sar9b_0.net59 a_2706_26108# 0.26567f
C1657 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[1] 0.22097f
C1658 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C1659 sar9b_0.net65 sar9b_0._05_ 0.31289f
C1660 sar9b_0.net24 single_9b_cdac_0.SW[7] 0.05134f
C1661 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[2] 0.21948f
C1662 single_9b_cdac_1.cdac_sw_9b_0.S[3] a_49221_17740# 0.22497f
C1663 a_3946_27530# sar9b_0.net44 0.05385f
C1664 VDPWR a_13164_28398# 0.25851f
C1665 VDPWR a_12618_23470# 0.32668f
C1666 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.26707f
C1667 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.01003f
C1668 a_11430_24931# a_11178_24802# 0.27388f
C1669 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01402f
C1670 clk tdc_0.phase_detector_0.INN 0.04168f
C1671 sar9b_0.net55 a_5443_19074# 0.03144f
C1672 VDPWR uo_out[5] 0.89589f
C1673 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.36006f
C1674 a_13011_20574# sar9b_0.net51 0.0305f
C1675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 3.10626f
C1676 sar9b_0.net40 sar9b_0.net62 0.08027f
C1677 VDPWR a_10506_24506# 0.34709f
C1678 VDPWR sar9b_0.net21 0.42201f
C1679 sar9b_0._09_ sar9b_0._17_ 0.04079f
C1680 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.08121f
C1681 tdc_0.OUTP sar9b_0.net6 0.49725f
C1682 a_5506_26802# a_6282_27170# 0.3578f
C1683 sar9b_0.net51 sar9b_0.net62 0.49495f
C1684 sar9b_0.net33 sar9b_0.net74 0.12313f
C1685 sar9b_0.net41 sar9b_0.net9 0.02887f
C1686 a_3027_22138# sar9b_0.clknet_1_1__leaf_CLK 0.03197f
C1687 sar9b_0.net40 a_13011_17910# 0.02505f
C1688 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[2] 0.3633f
C1689 VDPWR a_8166_27595# 0.26961f
C1690 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02632f
C1691 VDPWR sar9b_0.net27 3.63493f
C1692 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.03488f
C1693 VDPWR single_9b_cdac_0.SW[5] 2.59365f
C1694 sar9b_0.net65 sar9b_0.clknet_1_1__leaf_CLK 0.19718f
C1695 a_10548_19053# sar9b_0.net26 0.06094f
C1696 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.69086f
C1697 VDPWR a_11658_18142# 0.82655f
C1698 sar9b_0.net41 sar9b_0.net10 0.02787f
C1699 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.12431f
C1700 sar9b_0.net41 sar9b_0.net61 0.74807f
C1701 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C1702 sar9b_0.net46 a_4072_19474# 0.32046f
C1703 a_7914_23470# a_8438_23755# 0.05022f
C1704 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.30106f
C1705 sar9b_0.net33 sar9b_0.net31 0.02107f
C1706 VDPWR a_4812_21738# 0.27108f
C1707 sar9b_0.net71 sar9b_0.net46 0.29319f
C1708 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.04988f
C1709 sar9b_0.net1 sar9b_0.net27 0.07267f
C1710 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[8] 0.03384f
C1711 a_6783_19481# sar9b_0.net47 0.24046f
C1712 a_4947_20140# a_6130_20239# 0.0649f
C1713 a_5126_20140# a_5931_20140# 0.29221f
C1714 a_10402_21098# a_11430_20935# 0.07826f
C1715 th_dif_sw_0.CKB th_dif_sw_0.VCN 0.12032f
C1716 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 1.55942f
C1717 sar9b_0.net26 sar9b_0.net38 0.02477f
C1718 sar9b_0.net18 sar9b_0.net17 0.03659f
C1719 a_3370_26437# a_3156_26115# 0.04522f
C1720 single_9b_cdac_0.cdac_sw_9b_0.S[1] ua[0] 1.18579f
C1721 VDPWR tdc_0.OUTP 0.58425f
C1722 sar9b_0.net13 sar9b_0.net30 0.0911f
C1723 sar9b_0.net50 a_12684_20379# 0.11466f
C1724 a_10553_18922# a_10762_18823# 0.24088f
C1725 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C1726 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.0303f
C1727 single_9b_cdac_0.SW[1] sar9b_0.net29 0.30909f
C1728 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.04988f
C1729 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C1730 sar9b_0.net43 a_11104_24151# 0.02813f
C1731 a_8595_17910# single_9b_cdac_1.SW[0] 0.35058f
C1732 a_6132_23451# a_6922_23534# 0.1263f
C1733 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.01515f
C1734 VDPWR a_6444_19448# 0.20267f
C1735 sar9b_0.net51 a_7914_19178# 0.05227f
C1736 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.51772f
C1737 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.12898f
C1738 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 3.10626f
C1739 a_8595_17910# sar9b_0.net56 0.09371f
C1740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.05472f
C1741 VDPWR a_7638_23474# 0.28218f
C1742 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.CF[8] 0.19143f
C1743 VDPWR a_7470_22349# 0.26136f
C1744 sar9b_0.net8 sar9b_0.net57 0.16844f
C1745 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1746 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C1747 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.12431f
C1748 VDPWR a_5460_28377# 0.81693f
C1749 a_4934_22432# a_5289_22527# 0.18757f
C1750 a_4755_22138# a_5938_22378# 0.0649f
C1751 sar9b_0.net41 sar9b_0.net7 0.05595f
C1752 a_3370_26437# a_3438_26345# 0.35559f
C1753 sar9b_0.net41 a_9442_21474# 0.01846f
C1754 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.28523f
C1755 a_7926_23234# sar9b_0.net57 0.01631f
C1756 a_6642_19448# a_6783_19481# 0.27388f
C1757 a_7092_19455# a_7374_19685# 0.05462f
C1758 sar9b_0.net16 sar9b_0._10_ 0.06203f
C1759 sar9b_0.net66 sar9b_0._04_ 0.02178f
C1760 a_2893_24992# sar9b_0._16_ 0.18199f
C1761 VDPWR th_dif_sw_0.th_sw_1.CKB 3.04581f
C1762 a_3922_20239# sar9b_0.clknet_1_0__leaf_CLK 0.09413f
C1763 a_5931_20140# sar9b_0.net4 0.01405f
C1764 a_3855_25792# a_4136_25584# 0.29207f
C1765 a_9730_24138# a_9935_24187# 0.09983f
C1766 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.24207f
C1767 a_8940_24402# a_9270_24566# 0.04271f
C1768 sar9b_0.net2 a_9546_24506# 0.05795f
C1769 VDPWR a_5962_24151# 0.19439f
C1770 a_10830_19068# sar9b_0.net48 0.22344f
C1771 sar9b_0.net35 a_7404_16784# 0.26643f
C1772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C1773 sar9b_0.net11 clk 0.17325f
C1774 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42509f
C1775 a_3014_24136# sar9b_0.clknet_1_1__leaf_CLK 0.09139f
C1776 a_11178_24802# sar9b_0.net74 0.03041f
C1777 a_13011_23238# a_13216_22473# 0.01043f
C1778 sar9b_0.net26 sar9b_0.net6 0.75213f
C1779 a_8052_18123# a_8334_18353# 0.05462f
C1780 a_7602_18116# a_7743_18149# 0.27388f
C1781 sar9b_0.net27 sar9b_0.net29 0.42418f
C1782 sar9b_0.net39 a_5322_27170# 0.02945f
C1783 a_5394_18116# a_5849_18463# 0.3578f
C1784 VDPWR a_6252_20780# 0.26608f
C1785 VDPWR single_9b_cdac_1.SW[7] 2.36972f
C1786 a_13011_25902# a_13011_24802# 0.0246f
C1787 a_7743_16817# a_8057_17131# 0.07826f
C1788 sar9b_0.net31 a_11178_24802# 0.01626f
C1789 sar9b_0.net2 th_dif_sw_0.CK 0.02407f
C1790 VDPWR a_5439_24563# 0.25892f
C1791 a_9279_27227# a_9593_26914# 0.07826f
C1792 tdc_0.OUTN a_7404_16784# 0.05215f
C1793 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0._12_ 0.05952f
C1794 VDPWR a_11382_23474# 0.29464f
C1795 a_13011_23238# a_13216_23805# 0.01179f
C1796 sar9b_0.net44 sar9b_0.net39 0.24822f
C1797 ua[3] th_dif_sw_0.VCN 3.30291f
C1798 a_10742_27751# sar9b_0.net45 0.02244f
C1799 a_18214_3039# a_21368_4076# 0.99857f
C1800 VDPWR a_9258_21842# 0.86858f
C1801 clk th_dif_sw_0.VCN 2.08719f
C1802 VDPWR a_8303_23853# 0.26302f
C1803 sar9b_0.clknet_1_0__leaf_CLK a_3273_20185# 0.06919f
C1804 th_dif_sw_0.CK tdc_0.OUTN 0.07179f
C1805 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.42014f
C1806 a_11658_22138# a_12618_22138# 0.03432f
C1807 a_11842_22430# a_12182_22423# 0.24088f
C1808 a_11030_22954# sar9b_0.net11 0.0681f
C1809 a_9546_24506# a_10758_24459# 0.07766f
C1810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_55773_15501# 0.01076f
C1811 a_9442_21474# a_9782_21622# 0.24088f
C1812 a_9258_21842# a_10218_21842# 0.03471f
C1813 a_9258_21842# sar9b_0.net1 0.01455f
C1814 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02519f
C1815 sar9b_0.net53 sar9b_0.net38 0.33144f
C1816 VDPWR sar9b_0.net26 0.97073f
C1817 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C1818 VDPWR a_5443_19074# 0.34039f
C1819 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[3] 0.02468f
C1820 sar9b_0._07_ a_5581_19664# 0.33323f
C1821 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.10626f
C1822 a_7289_21127# a_6975_20813# 0.07826f
C1823 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR 0.62443f
C1824 VDPWR a_6534_27123# 0.27103f
C1825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.19266f
C1826 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[2] 0.0313f
C1827 th_dif_sw_0.VCN single_9b_cdac_1.SW[0] 0.15316f
C1828 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] 27.3302f
C1829 a_6738_22112# a_7402_22441# 0.16939f
C1830 sar9b_0.net26 sar9b_0.net1 0.04547f
C1831 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C1832 sar9b_0.net2 single_9b_cdac_1.SW[1] 0.77878f
C1833 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.6919f
C1834 a_8052_16791# sar9b_0.net27 0.01294f
C1835 a_8098_23762# clk 0.01832f
C1836 a_8345_26455# sar9b_0.net37 0.02763f
C1837 VDPWR a_48343_16877# 1.81495f
C1838 a_11776_21141# sar9b_0.net39 0.01141f
C1839 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.62443f
C1840 a_11842_23762# a_12182_23755# 0.24088f
C1841 sar9b_0.net43 a_9138_27163# 0.01333f
C1842 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.26684f
C1843 sar9b_0.net54 a_6378_24802# 0.1648f
C1844 sar9b_0.net23 a_9939_28566# 0.20828f
C1845 a_62748_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.23864f
C1846 sar9b_0.net40 sar9b_0.net42 0.0514f
C1847 sar9b_0.net66 sar9b_0._12_ 0.16928f
C1848 VDPWR a_3027_22138# 0.44684f
C1849 a_8622_26345# a_8340_26115# 0.05462f
C1850 a_7289_21127# a_7498_21109# 0.24088f
C1851 sar9b_0.net42 sar9b_0.net51 0.01622f
C1852 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.01751f
C1853 VDPWR sar9b_0.net65 0.94256f
C1854 a_9165_24988# sar9b_0.net53 0.20816f
C1855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C1856 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02778f
C1857 VDPWR a_5938_22378# 0.38557f
C1858 sar9b_0.net16 a_3795_19512# 0.0476f
C1859 a_10506_23174# a_10230_23234# 0.1263f
C1860 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[3] 0.06162f
C1861 a_7743_18149# a_7404_18116# 0.07649f
C1862 a_10230_23234# sar9b_0.net74 0.2089f
C1863 a_6678_27470# sar9b_0.net21 0.01436f
C1864 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR 2.81428f
C1865 sar9b_0.net35 sar9b_0.net60 0.02971f
C1866 a_7092_19455# sar9b_0.net10 0.25701f
C1867 a_11466_23174# sar9b_0.net10 0.05039f
C1868 sar9b_0.net60 sar9b_0.net16 0.01459f
C1869 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C1870 single_9b_cdac_0.cdac_sw_9b_0.S[0] a_62748_26999# 0.59531f
C1871 uo_out[1] ui_in[0] 0.06797f
C1872 uo_out[0] clk 0.48415f
C1873 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.01879f
C1874 a_6954_27466# a_7478_27751# 0.05022f
C1875 a_11430_27595# a_11776_27801# 0.07649f
C1876 a_6636_20780# sar9b_0.net40 0.02169f
C1877 sar9b_0._08_ a_5812_21028# 0.05999f
C1878 a_24332_16877# single_9b_cdac_1.SW[8] 0.28324f
C1879 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.19266f
C1880 a_8057_18463# sar9b_0.net5 0.10125f
C1881 a_12047_18525# sar9b_0.net6 0.01853f
C1882 sar9b_0.net44 sar9b_0.net36 0.21739f
C1883 sar9b_0.net49 sar9b_0.net40 0.16393f
C1884 a_7338_24802# a_7590_24931# 0.27388f
C1885 sar9b_0._16_ sar9b_0.net69 0.04762f
C1886 a_4365_25770# a_4698_25851# 0.14439f
C1887 sar9b_0.net49 sar9b_0.net51 0.50265f
C1888 a_8340_26115# a_9138_27163# 0.01342f
C1889 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS th_dif_sw_0.VCN 0.14643f
C1890 sar9b_0._11_ sar9b_0._10_ 0.03596f
C1891 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16357_9613# 0.16728f
C1892 a_9942_27470# sar9b_0.net34 0.03758f
C1893 VDPWR sar9b_0.net53 3.3527f
C1894 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 a_34814_17740# 0.14695f
C1895 a_10858_17113# sar9b_0.net27 0.025f
C1896 VDPWR a_10690_22806# 0.22042f
C1897 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.3196f
C1898 single_9b_cdac_0.SW[1] a_13216_26469# 0.02143f
C1899 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[4] 0.02149f
C1900 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.SW[5] 0.02506f
C1901 sar9b_0._02_ sar9b_0.clk_div_0.COUNT\[1\] 0.01796f
C1902 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07517f
C1903 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.01003f
C1904 sar9b_0.net45 a_10607_27849# 0.05607f
C1905 VDPWR uo_out[2] 0.90561f
C1906 ui_in[6] ui_in[5] 0.03102f
C1907 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.02149f
C1908 sar9b_0.net1 sar9b_0.net53 0.19803f
C1909 a_9472_18823# sar9b_0.net26 0.27337f
C1910 a_10182_20463# a_10528_20155# 0.07649f
C1911 sar9b_0.net43 clk 0.04165f
C1912 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.12431f
C1913 a_5126_20140# a_5633_20244# 0.21226f
C1914 a_4947_20140# a_5481_20185# 0.35097f
C1915 a_7284_20787# sar9b_0.net61 0.01281f
C1916 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.7611f
C1917 VDPWR a_12047_18525# 0.26725f
C1918 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.SW[8] 0.22497f
C1919 a_7914_27466# sar9b_0.net60 0.24386f
C1920 sar9b_0._17_ sar9b_0.net4 0.77945f
C1921 a_8970_20510# a_9494_20290# 0.04522f
C1922 a_8694_20570# a_9359_20191# 0.19065f
C1923 sar9b_0.net73 sar9b_0.net37 0.02388f
C1924 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.83441f
C1925 VDPWR a_3014_24136# 0.9015f
C1926 VDPWR a_9802_26815# 0.20303f
C1927 sar9b_0.net32 sar9b_0.net14 0.14467f
C1928 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[1] 0.22097f
C1929 a_10378_27170# a_9593_26914# 0.26257f
C1930 a_10858_17113# tdc_0.OUTP 0.06033f
C1931 sar9b_0.net27 a_12684_20379# 0.01643f
C1932 VDPWR a_6562_25094# 0.22221f
C1933 a_3695_23038# sar9b_0._07_ 0.02799f
C1934 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.28523f
C1935 VDPWR a_9494_20290# 0.20426f
C1936 a_5289_22527# sar9b_0._07_ 0.01435f
C1937 sar9b_0.net49 a_10742_21091# 0.13511f
C1938 sar9b_0.net60 a_5523_21528# 0.24769f
C1939 a_12435_24802# sar9b_0.net12 0.22022f
C1940 sar9b_0._17_ sar9b_0.clk_div_0.COUNT\[2\] 0.57711f
C1941 a_6975_20813# sar9b_0.net47 0.17348f
C1942 single_9b_cdac_0.cdac_sw_9b_0.S[5] ua[0] 1.56372f
C1943 a_11658_26134# a_11842_26426# 0.44532f
C1944 a_5441_22522# a_5289_22527# 0.22517f
C1945 a_5739_22488# sar9b_0.net39 0.01448f
C1946 sar9b_0.net36 single_9b_cdac_0.SW[8] 0.07497f
C1947 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.01751f
C1948 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.05472f
C1949 single_9b_cdac_0.SW[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.363f
C1950 sar9b_0.net57 a_5196_19448# 0.01615f
C1951 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.28523f
C1952 a_10402_27758# single_9b_cdac_0.SW[7] 0.01715f
C1953 sar9b_0.net41 single_9b_cdac_1.SW[4] 0.24901f
C1954 sar9b_0.net1 a_9494_20290# 0.02028f
C1955 sar9b_0._11_ sar9b_0._18_ 0.03308f
C1956 sar9b_0.net27 a_13216_26469# 0.01058f
C1957 sar9b_0.net64 sar9b_0.clknet_0_CLK 0.01151f
C1958 a_11859_21906# single_9b_cdac_1.CF[2] 0.35504f
C1959 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] 1.15122f
C1960 sar9b_0.net43 a_11030_22954# 0.01262f
C1961 a_11859_20574# sar9b_0.net5 0.03891f
C1962 sar9b_0._11_ sar9b_0._01_ 0.04965f
C1963 a_6346_23773# sar9b_0.net54 0.1286f
C1964 VDPWR a_4922_20857# 0.22486f
C1965 sar9b_0.net72 a_2893_24992# 0.03569f
C1966 a_8031_26141# a_8345_26455# 0.07826f
C1967 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C1968 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.38397f
C1969 a_3545_26914# a_3754_26815# 0.24088f
C1970 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C1971 a_7602_18116# sar9b_0.net73 0.08061f
C1972 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.SW[4] 0.1498f
C1973 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP a_29134_16877# 0.04592f
C1974 VDPWR th_dif_sw_0.VCP 6.87158f
C1975 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.75853f
C1976 sar9b_0.net48 sar9b_0.net37 0.18456f
C1977 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.CF[2] 0.19321f
C1978 a_3540_27045# a_3545_26914# 0.44532f
C1979 sar9b_0.net4 a_6252_19074# 0.05708f
C1980 sar9b_0.net36 a_4749_27652# 0.07973f
C1981 VDPWR a_8591_22855# 0.29655f
C1982 a_2892_27039# a_3231_27227# 0.07649f
C1983 a_7498_21109# sar9b_0.net47 0.15768f
C1984 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.6919f
C1985 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C1986 a_6132_23451# clk 0.01117f
C1987 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.02784f
C1988 a_7347_24160# sar9b_0.net54 0.37926f
C1989 a_7193_22459# a_7470_22349# 0.09983f
C1990 sar9b_0.net60 a_5465_28246# 0.02116f
C1991 sar9b_0._01_ a_5374_20145# 0.13551f
C1992 sar9b_0.net32 a_11842_26426# 0.01684f
C1993 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[6] 1.94202f
C1994 a_10098_19171# sar9b_0.net48 0.29653f
C1995 sar9b_0.net49 a_9647_21523# 0.22799f
C1996 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[6] 0.09845f
C1997 single_9b_cdac_0.SW[7] single_9b_cdac_1.CF[7] 1.81115f
C1998 a_11718_23127# clk 0.01747f
C1999 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96985f
C2000 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[4] 0.03895f
C2001 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 2.82215f
C2002 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C2003 a_2508_23444# sar9b_0.net69 0.06549f
C2004 sar9b_0.net60 a_7343_27849# 0.20041f
C2005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.03729f
C2006 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[0] 0.06503f
C2007 sar9b_0.net63 sar9b_0._17_ 0.1985f
C2008 sar9b_0.net13 a_7590_24931# 0.04157f
C2009 a_8098_18810# a_9126_19131# 0.07826f
C2010 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C2011 VDPWR a_5196_18116# 0.20215f
C2012 a_9450_17846# a_9634_17478# 0.43869f
C2013 a_12182_19759# a_12618_19474# 0.16939f
C2014 single_9b_cdac_1.SW[2] a_9634_17478# 0.01591f
C2015 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C2016 a_10926_17021# a_10649_17131# 0.09983f
C2017 sar9b_0.net46 sar9b_0.net37 0.07123f
C2018 sar9b_0.net56 a_8874_19178# 0.01259f
C2019 VDPWR a_10932_25713# 0.81346f
C2020 VDPWR a_3438_27677# 0.25451f
C2021 a_7602_18116# sar9b_0.net48 0.06506f
C2022 a_11382_22142# sar9b_0.net39 0.03507f
C2023 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.84425f
C2024 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.12898f
C2025 a_5506_17478# sar9b_0.net56 0.03523f
C2026 th_dif_sw_0.CK sar9b_0.net39 0.03714f
C2027 tdc_0.phase_detector_0.pd_out_0.A a_16970_11404# 0.18949f
C2028 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.08121f
C2029 sar9b_0._11_ sar9b_0.net60 0.60917f
C2030 single_9b_cdac_1.SW[8] a_12047_19857# 0.03035f
C2031 a_6030_24396# a_5962_24151# 0.35559f
C2032 sar9b_0.net32 sar9b_0.net11 0.02514f
C2033 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.17185f
C2034 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[0\] 0.01565f
C2035 a_11382_19478# a_11658_19474# 0.1263f
C2036 a_9270_24566# sar9b_0.net53 0.22967f
C2037 a_2892_23070# sar9b_0.net66 0.14576f
C2038 sar9b_0.net4 clk 0.04636f
C2039 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 1.55982f
C2040 a_9154_20142# sar9b_0.net37 0.02634f
C2041 a_10644_16791# sar9b_0.net61 0.02207f
C2042 uo_out[5] ui_in[0] 0.06786f
C2043 a_8266_17113# sar9b_0.net6 0.01365f
C2044 VDPWR a_5931_20140# 0.09106f
C2045 uo_out[6] uo_out[7] 2.95271f
C2046 a_7188_22119# sar9b_0.clk_div_0.COUNT\[2\] 0.01175f
C2047 sar9b_0.net40 sar9b_0.net11 0.02451f
C2048 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C2049 sar9b_0._18_ sar9b_0.net39 0.295f
C2050 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[8] 0.01791f
C2051 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C2052 sar9b_0.net24 sar9b_0.net59 0.29571f
C2053 a_5748_24381# a_5753_24250# 0.44532f
C2054 sar9b_0.clk_div_0.COUNT\[2\] clk 0.11336f
C2055 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[5] 0.31534f
C2056 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] 0.17948f
C2057 sar9b_0.net53 a_11658_22138# 0.16567f
C2058 a_7602_18116# sar9b_0.net46 0.27602f
C2059 a_7743_16817# sar9b_0.net46 0.17057f
C2060 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.75853f
C2061 sar9b_0.net73 a_7404_18116# 0.09233f
C2062 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07517f
C2063 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C2064 sar9b_0.net26 a_12684_20379# 0.01826f
C2065 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[7] 0.01887f
C2066 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C2067 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[1] 0.22097f
C2068 sar9b_0.net40 a_12870_19603# 0.07154f
C2069 a_3819_24136# sar9b_0.clk_div_0.COUNT\[2\] 0.01683f
C2070 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] 1.15121f
C2071 a_13011_20574# a_13216_19809# 0.01043f
C2072 sar9b_0._13_ sar9b_0.net72 0.1941f
C2073 a_11842_19766# a_12870_19603# 0.07826f
C2074 a_6307_27584# sar9b_0.net44 0.23235f
C2075 VDPWR a_6922_23534# 0.2895f
C2076 sar9b_0.net56 sar9b_0.net4 0.03241f
C2077 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.17717f
C2078 a_9760_22819# clk 0.01624f
C2079 VDPWR a_3454_22567# 0.01572f
C2080 a_8115_28566# uo_out[6] 0.42188f
C2081 VDPWR a_8266_17113# 0.19893f
C2082 sar9b_0.net31 a_12870_22267# 0.03044f
C2083 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.07579f
C2084 sar9b_0.net55 sar9b_0._17_ 0.77591f
C2085 VDPWR a_7306_19777# 0.20423f
C2086 sar9b_0.net70 sar9b_0.net69 0.12146f
C2087 a_3156_27447# a_3370_27769# 0.04522f
C2088 a_2847_27473# a_3161_27787# 0.07826f
C2089 a_2547_28132# a_2931_28566# 0.09678f
C2090 sar9b_0.net61 a_9634_17478# 0.16934f
C2091 a_10194_16784# a_10335_16817# 0.27388f
C2092 VDPWR a_8266_18445# 0.19813f
C2093 a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK 1.89917f
C2094 sar9b_0.net56 a_5322_17846# 0.23955f
C2095 sar9b_0.net34 a_10284_25707# 0.27185f
C2096 sar9b_0.net32 sar9b_0.net45 0.02882f
C2097 single_9b_cdac_0.SW[7] sar9b_0.net36 0.33484f
C2098 VDPWR a_12047_22521# 0.24932f
C2099 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.84061f
C2100 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C2101 sar9b_0._04_ sar9b_0._05_ 0.2432f
C2102 sar9b_0.net48 a_7404_18116# 0.02507f
C2103 a_8266_18445# sar9b_0.net1 0.0136f
C2104 sar9b_0.net59 a_3161_26455# 0.10291f
C2105 sar9b_0.net70 sar9b_0._18_ 0.03792f
C2106 VDPWR sar9b_0.net30 0.61341f
C2107 sar9b_0.net63 clk 0.08413f
C2108 sar9b_0.net40 sar9b_0.net45 0.05943f
C2109 sar9b_0.net60 sar9b_0.net39 0.1395f
C2110 sar9b_0.net72 sar9b_0.net69 0.04519f
C2111 sar9b_0.net11 sar9b_0.net62 0.20455f
C2112 a_11842_18434# sar9b_0.net6 0.02355f
C2113 sar9b_0._12_ sar9b_0.net4 0.24818f
C2114 a_11339_27039# single_9b_cdac_0.SW[5] 0.36476f
C2115 sar9b_0.net22 sar9b_0.cyclic_flag_0.FINAL 0.02996f
C2116 th_dif_sw_0.CK sar9b_0.net36 0.03321f
C2117 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.02632f
C2118 VDPWR a_12047_23853# 0.26429f
C2119 a_11178_24802# a_11776_25137# 0.06623f
C2120 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.42784f
C2121 sar9b_0._18_ a_4332_23043# 0.03742f
C2122 sar9b_0.net55 a_6252_19074# 0.17527f
C2123 VDPWR single_9b_cdac_0.SW[0] 3.07511f
C2124 VDPWR a_11104_24151# 0.19368f
C2125 sar9b_0._12_ sar9b_0.clk_div_0.COUNT\[2\] 0.06165f
C2126 sar9b_0.net49 sar9b_0.net42 0.02948f
C2127 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.SW[7] 0.17154f
C2128 a_33936_26999# single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.59531f
C2129 a_5846_26950# a_6282_27170# 0.16939f
C2130 sar9b_0.net32 uo_out[0] 0.0917f
C2131 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.10429f
C2132 sar9b_0.net8 single_9b_cdac_1.CF[1] 0.12551f
C2133 sar9b_0.net35 sar9b_0.net59 0.93479f
C2134 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[3] 0.08999f
C2135 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.3196f
C2136 sar9b_0.net57 sar9b_0.net46 0.19212f
C2137 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.62443f
C2138 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] 3.10207f
C2139 VDPWR a_8512_27801# 0.19986f
C2140 a_3156_26115# a_2706_26108# 0.03471f
C2141 a_2508_26108# a_2847_26141# 0.07649f
C2142 a_4044_24776# sar9b_0.clk_div_0.COUNT\[2\] 0.01228f
C2143 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.clk_div_0.COUNT\[1\] 0.46155f
C2144 a_7638_19238# sar9b_0.net5 0.03793f
C2145 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.10499f
C2146 a_16159_13315# a_16185_13034# 0.19021f
C2147 VDPWR a_5235_27466# 0.38926f
C2148 a_10830_19068# sar9b_0.net26 0.04966f
C2149 VDPWR a_11842_18434# 0.23262f
C2150 VDPWR a_11658_19474# 0.84186f
C2151 a_5581_20992# sar9b_0._01_ 0.01832f
C2152 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.42014f
C2153 a_7914_23470# a_8874_23470# 0.03432f
C2154 a_10182_20463# a_9154_20142# 0.07826f
C2155 a_5010_28495# uo_out[7] 0.02505f
C2156 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.45521f
C2157 a_9942_27470# a_10218_27466# 0.1263f
C2158 a_6738_22112# sar9b_0.net35 0.02157f
C2159 VDPWR a_10166_3438# 0.07956f
C2160 VDPWR a_14871_9671# 0.67026f
C2161 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62538f
C2162 a_10742_21091# a_11178_20806# 0.16939f
C2163 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C2164 sar9b_0._07_ sar9b_0.net16 0.16722f
C2165 sar9b_0.net36 single_9b_cdac_1.SW[1] 0.03305f
C2166 m2_23774_17236# single_9b_cdac_1.SW[8] 0.02037f
C2167 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.45521f
C2168 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C2169 a_33936_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.23864f
C2170 VDPWR a_9363_20826# 0.44006f
C2171 a_3819_24136# sar9b_0.clknet_1_1__leaf_CLK 0.01525f
C2172 sar9b_0.net4 a_5394_18116# 0.02958f
C2173 a_10548_19053# a_11338_19178# 0.1263f
C2174 uio_in[3] uio_in[2] 0.03102f
C2175 a_10194_16784# sar9b_0.net48 0.24027f
C2176 a_8098_23762# sar9b_0.net62 0.02357f
C2177 sar9b_0._08_ sar9b_0.net16 0.13446f
C2178 a_12491_27662# sar9b_0.net32 0.02118f
C2179 sar9b_0.net41 single_9b_cdac_1.SW[6] 0.01701f
C2180 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.45521f
C2181 a_8940_24402# sar9b_0.net37 0.01757f
C2182 sar9b_0.net55 clk 0.03649f
C2183 a_9363_20826# sar9b_0.net1 0.02566f
C2184 a_6137_23791# a_6414_23681# 0.09983f
C2185 a_6282_17846# a_6534_17799# 0.27388f
C2186 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 3.04383f
C2187 VDPWR a_8622_26345# 0.28256f
C2188 sar9b_0.net8 a_11859_20574# 0.0265f
C2189 sar9b_0.net20 a_7539_28566# 0.08083f
C2190 a_3219_22860# sar9b_0.clk_div_0.COUNT\[1\] 0.21033f
C2191 sar9b_0.net63 sar9b_0._12_ 0.07563f
C2192 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.26942f
C2193 sar9b_0.net60 a_4332_23043# 0.05573f
C2194 sar9b_0.net5 a_9359_20191# 0.0567f
C2195 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[2] 0.01791f
C2196 sar9b_0.net31 single_9b_cdac_1.CF[3] 0.01828f
C2197 sar9b_0.net32 sar9b_0.net13 0.02694f
C2198 VDPWR a_7978_22202# 0.29273f
C2199 VDPWR a_5742_28392# 0.25649f
C2200 a_10707_23470# sar9b_0.net74 0.16592f
C2201 sar9b_0.net41 a_9782_21622# 0.02219f
C2202 sar9b_0.net43 sar9b_0.net40 0.02302f
C2203 sar9b_0.net45 a_9588_27045# 0.25117f
C2204 sar9b_0.net63 a_4044_24776# 0.04322f
C2205 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[8] 0.2453f
C2206 a_7092_19455# a_7882_19538# 0.1263f
C2207 a_6783_19481# a_7097_19795# 0.07826f
C2208 sar9b_0._05_ sar9b_0._12_ 0.12977f
C2209 a_13011_19242# sar9b_0.net40 0.03f
C2210 sar9b_0.net16 sar9b_0.clknet_1_0__leaf_CLK 0.0448f
C2211 uo_out[5] uo_out[4] 2.90315f
C2212 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 1.71649f
C2213 a_4934_22432# sar9b_0.net39 0.0126f
C2214 a_3855_25792# a_4293_25852# 0.02614f
C2215 a_4125_25958# a_4365_25770# 0.35097f
C2216 sar9b_0.net43 sar9b_0.net51 0.39434f
C2217 a_9935_24187# a_10070_24286# 0.35559f
C2218 a_5581_20992# sar9b_0.net60 0.06229f
C2219 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C2220 sar9b_0.net13 sar9b_0.net40 0.24488f
C2221 sar9b_0.net60 sar9b_0.net36 0.25636f
C2222 a_13011_16810# single_9b_cdac_1.SW[4] 0.01587f
C2223 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.28523f
C2224 a_10803_19474# sar9b_0.net73 0.03401f
C2225 a_8266_17113# a_8052_16791# 0.04522f
C2226 VDPWR sar9b_0._17_ 1.32705f
C2227 sar9b_0.net29 single_9b_cdac_0.SW[0] 0.03951f
C2228 a_3371_23106# a_3219_22860# 0.24998f
C2229 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.05472f
C2230 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.SW[7] 0.14951f
C2231 sar9b_0.net48 a_10410_17846# 0.27687f
C2232 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.3186f
C2233 sar9b_0.net2 sar9b_0.net12 0.20768f
C2234 sar9b_0.net32 a_12560_27128# 0.01666f
C2235 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.84426f
C2236 sar9b_0.net21 sar9b_0.net37 0.06888f
C2237 sar9b_0.net38 clk 0.04449f
C2238 single_9b_cdac_0.cdac_sw_9b_0.S[6] ua[0] 1.66285f
C2239 single_9b_cdac_0.cdac_sw_9b_0.S[8] th_dif_sw_0.VCN 0.85562f
C2240 a_7743_18149# a_8057_18463# 0.07826f
C2241 a_8052_18123# a_8842_18206# 0.1263f
C2242 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.07579f
C2243 a_6834_20780# a_6975_20813# 0.27388f
C2244 a_5394_18116# a_6058_18445# 0.16939f
C2245 a_5844_18123# a_6126_18353# 0.05462f
C2246 single_9b_cdac_1.SW[0] a_9839_17527# 0.03009f
C2247 sar9b_0._07_ a_5523_21528# 0.18199f
C2248 VDPWR a_9138_27163# 0.37075f
C2249 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.71729f
C2250 sar9b_0._12_ sar9b_0.clknet_1_1__leaf_CLK 0.30353f
C2251 VDPWR th_dif_sw_0.CKB 1.43024f
C2252 a_9588_27045# a_9870_27060# 0.06034f
C2253 tdc_0.OUTN a_7602_16784# 0.07198f
C2254 sar9b_0.net45 uo_out[7] 0.02028f
C2255 sar9b_0.net8 single_9b_cdac_1.CF[3] 0.02324f
C2256 sar9b_0.net41 sar9b_0.net52 0.09293f
C2257 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.10499f
C2258 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36044f
C2259 VDPWR a_10254_2858# 0.51112f
C2260 a_8554_26437# sar9b_0.net59 0.1439f
C2261 sar9b_0.clknet_1_0__leaf_CLK a_3723_20140# 0.07189f
C2262 sar9b_0.net44 a_3822_27060# 0.01345f
C2263 a_11658_22138# a_12047_22521# 0.06034f
C2264 a_11842_22430# a_12618_22138# 0.3578f
C2265 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.10429f
C2266 VDPWR a_15151_10456# 0.3789f
C2267 sar9b_0.net58 a_5460_28377# 0.15559f
C2268 VDPWR a_5633_20244# 0.10568f
C2269 a_9730_24138# a_10506_24506# 0.3578f
C2270 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.26625f
C2271 a_10803_19474# sar9b_0.net48 0.02063f
C2272 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.62443f
C2273 a_3946_27530# a_3156_27447# 0.1263f
C2274 sar9b_0.net40 a_6132_23451# 0.01344f
C2275 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C2276 VDPWR a_6252_19074# 0.21971f
C2277 sar9b_0.net47 a_6444_19448# 0.06747f
C2278 a_10548_19053# a_10803_18142# 0.04032f
C2279 a_7498_21109# a_6834_20780# 0.16939f
C2280 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.42509f
C2281 sar9b_0.net43 sar9b_0.net62 0.65145f
C2282 single_9b_cdac_0.SW[6] single_9b_cdac_1.CF[6] 1.79589f
C2283 th_dif_sw_0.CK single_9b_cdac_1.SW[2] 0.04691f
C2284 sar9b_0.net47 a_7470_22349# 0.22357f
C2285 a_10402_25094# sar9b_0.net36 0.0133f
C2286 a_10742_27751# VDPWR 0.20368f
C2287 sar9b_0.net42 sar9b_0.net11 0.02571f
C2288 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.0313f
C2289 a_7743_16817# sar9b_0.net27 0.02921f
C2290 uo_out[2] ui_in[0] 0.0679f
C2291 a_4934_22432# a_4332_23043# 0.01428f
C2292 a_4755_22138# sar9b_0._12_ 0.15278f
C2293 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[0] 0.30922f
C2294 a_11842_23762# a_12618_23470# 0.3578f
C2295 a_10803_18142# sar9b_0.net38 0.20613f
C2296 sar9b_0.net49 a_10227_18142# 0.20483f
C2297 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.81428f
C2298 a_6414_23681# sar9b_0.net57 0.05577f
C2299 VDPWR a_11338_19178# 0.29105f
C2300 sar9b_0.net27 a_11842_22430# 0.01034f
C2301 dw_12589_1395# ua[4] 1.41177f
C2302 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 2.824f
C2303 VDPWR a_2547_28132# 0.36522f
C2304 sar9b_0.clknet_0_CLK sar9b_0.net57 0.03539f
C2305 a_6484_22845# a_6744_23238# 0.17405f
C2306 a_3425_20244# a_3273_20185# 0.22338f
C2307 th_dif_sw_0.CK a_12182_18427# 0.06686f
C2308 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.71729f
C2309 single_9b_cdac_0.SW[3] single_9b_cdac_0.SW[0] 0.01042f
C2310 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.58106f
C2311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C2312 VDPWR sar9b_0._04_ 0.59309f
C2313 a_9130_26198# a_8340_26115# 0.1263f
C2314 a_10553_18922# sar9b_0.net36 0.01892f
C2315 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP a_38738_26999# 0.04592f
C2316 sar9b_0.net27 a_11842_23762# 0.01034f
C2317 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.42784f
C2318 a_6642_19448# a_6444_19448# 0.06623f
C2319 sar9b_0.net6 single_9b_cdac_1.SW[0] 0.10368f
C2320 sar9b_0.net40 sar9b_0.net4 0.05476f
C2321 VDPWR a_7188_22119# 0.85695f
C2322 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.02149f
C2323 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[0] 4.15031f
C2324 sar9b_0._11_ sar9b_0._07_ 0.03254f
C2325 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] 3.10215f
C2326 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[2] 17.4687f
C2327 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[0] 0.31534f
C2328 a_9472_23805# sar9b_0.net53 0.01787f
C2329 VDPWR ua[3] 1.80857f
C2330 a_13011_23238# sar9b_0.net10 0.22279f
C2331 sar9b_0.net56 sar9b_0.net6 0.14505f
C2332 sar9b_0.net51 sar9b_0.net4 0.21881f
C2333 sar9b_0.net67 sar9b_0.net70 0.05082f
C2334 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[4] 0.03478f
C2335 single_9b_cdac_0.SW[1] sar9b_0.net33 0.06514f
C2336 VDPWR clk 4.0924f
C2337 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP a_38738_16877# 0.04592f
C2338 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C2339 a_6954_27466# a_7914_27466# 0.03432f
C2340 sar9b_0.net58 a_6534_27123# 0.17315f
C2341 sar9b_0.net40 sar9b_0.clk_div_0.COUNT\[2\] 0.02492f
C2342 a_7138_27758# a_7478_27751# 0.24088f
C2343 sar9b_0.net35 sar9b_0.net5 0.0951f
C2344 VDPWR a_3545_26914# 0.22169f
C2345 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.03543f
C2346 sar9b_0._08_ sar9b_0._11_ 0.26992f
C2347 a_9162_23174# sar9b_0.net11 0.06676f
C2348 a_8386_22806# sar9b_0.net54 0.10034f
C2349 VDPWR a_2451_27234# 0.27934f
C2350 VDPWR a_3819_24136# 0.09178f
C2351 sar9b_0.net1 clk 0.04871f
C2352 a_64331_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.01076f
C2353 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.01134f
C2354 sar9b_0.net2 sar9b_0.net5 0.0239f
C2355 a_10402_27758# sar9b_0.net59 0.08863f
C2356 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.75853f
C2357 a_9258_21842# sar9b_0.net37 0.02924f
C2358 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.84061f
C2359 VDPWR a_8303_18859# 0.2747f
C2360 sar9b_0.net10 a_11382_22142# 0.06561f
C2361 a_6767_25185# a_6902_25087# 0.35559f
C2362 th_dif_sw_0.CK sar9b_0.net61 0.02316f
C2363 a_4365_25770# sar9b_0.clknet_1_1__leaf_CLK 0.06633f
C2364 VDPWR single_9b_cdac_1.SW[0] 3.84179f
C2365 sar9b_0.net42 sar9b_0.net45 0.14568f
C2366 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[7] 0.02552f
C2367 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[3] 4.15101f
C2368 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.12898f
C2369 single_9b_cdac_1.SW[3] ua[0] 0.14032f
C2370 a_11146_25483# sar9b_0.net52 0.17111f
C2371 VDPWR sar9b_0.net56 1.95434f
C2372 a_3369_24181# a_3014_24136# 0.18752f
C2373 sar9b_0._11_ sar9b_0.clknet_1_0__leaf_CLK 0.08207f
C2374 a_11658_26134# a_12870_26263# 0.07766f
C2375 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[8] 0.21771f
C2376 sar9b_0.net26 sar9b_0.net37 0.22151f
C2377 a_4011_22488# sar9b_0.clknet_1_1__leaf_CLK 0.06293f
C2378 VDPWR a_11030_22954# 0.20335f
C2379 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C2380 a_17125_9355# th_dif_sw_0.VCP 0.05474f
C2381 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.10499f
C2382 sar9b_0.net57 sar9b_0.net27 0.10308f
C2383 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR 0.62443f
C2384 a_6534_27123# sar9b_0.net37 0.0697f
C2385 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C2386 VDPWR a_57946_26999# 1.81495f
C2387 sar9b_0.net33 sar9b_0.net27 0.03715f
C2388 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22352f
C2389 sar9b_0.net56 sar9b_0.net1 0.26215f
C2390 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.SW[0] 0.17156f
C2391 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.S[3] 16.7662f
C2392 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[2] 0.24301f
C2393 VDPWR a_13011_20806# 0.49978f
C2394 a_10098_19171# sar9b_0.net26 0.06434f
C2395 a_8874_19178# a_7914_19178# 0.03471f
C2396 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] 3.10048f
C2397 sar9b_0.net59 sar9b_0.net39 0.21806f
C2398 VDPWR a_10803_18142# 0.46102f
C2399 sar9b_0.net63 sar9b_0.net40 0.26974f
C2400 a_6307_27584# sar9b_0.net60 0.03874f
C2401 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP a_48343_16877# 0.04592f
C2402 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02545f
C2403 sar9b_0.net61 single_9b_cdac_1.SW[1] 0.13622f
C2404 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.SW[2] 0.17157f
C2405 a_6540_22112# a_6738_22112# 0.06623f
C2406 VDPWR a_7590_24931# 0.27042f
C2407 sar9b_0.net49 a_11178_20806# 0.26056f
C2408 sar9b_0.net7 th_dif_sw_0.CK 0.17128f
C2409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.12431f
C2410 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22526f
C2411 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net62 0.03763f
C2412 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.01173f
C2413 a_6954_27466# a_7343_27849# 0.06034f
C2414 a_6738_22112# sar9b_0.net39 0.05411f
C2415 VDPWR sar9b_0._12_ 1.04527f
C2416 single_9b_cdac_0.SW[6] single_9b_cdac_1.CF[7] 0.12064f
C2417 sar9b_0._07_ sar9b_0.net39 0.04027f
C2418 VDPWR a_10607_27849# 0.26664f
C2419 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP a_48343_26999# 0.04592f
C2420 single_9b_cdac_1.cdac_sw_9b_0.S[2] th_dif_sw_0.VCP 54.8348f
C2421 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[1\] 0.17923f
C2422 a_5441_22522# sar9b_0.net39 0.01163f
C2423 a_10218_20806# a_9930_20510# 0.01059f
C2424 sar9b_0.net29 clk 0.03602f
C2425 sar9b_0.net45 uo_out[6] 0.06932f
C2426 a_11382_23474# a_11842_23762# 0.26257f
C2427 sar9b_0.net26 a_11842_22430# 0.02923f
C2428 a_7638_23474# sar9b_0.net57 0.06419f
C2429 VDPWR a_4044_24776# 0.26952f
C2430 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.17209f
C2431 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.84426f
C2432 sar9b_0._14_ a_4044_24776# 0.04883f
C2433 a_2893_24992# a_2940_25096# 0.19021f
C2434 a_7890_26108# a_8554_26437# 0.16939f
C2435 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.19266f
C2436 a_8057_18463# sar9b_0.net73 0.07314f
C2437 a_43540_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.23864f
C2438 sar9b_0.net35 sar9b_0.net54 0.19733f
C2439 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.S[7] 1.06635f
C2440 VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.17946f
C2441 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.22352f
C2442 single_9b_cdac_0.cdac_sw_9b_0.S[7] ua[0] 1.97045f
C2443 a_3090_27163# a_3754_26815# 0.16939f
C2444 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[3] 0.12359f
C2445 sar9b_0.net26 a_11842_23762# 0.0241f
C2446 a_4812_28371# sar9b_0.net20 0.3101f
C2447 a_3090_27163# a_3540_27045# 0.03432f
C2448 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 1.71649f
C2449 a_10194_16784# sar9b_0.net27 0.05895f
C2450 a_5682_23444# clk 0.01117f
C2451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.07517f
C2452 sar9b_0.net7 single_9b_cdac_1.SW[1] 0.70147f
C2453 sar9b_0.net43 sar9b_0.net42 0.4289f
C2454 a_7193_22459# a_7978_22202# 0.26257f
C2455 sar9b_0._01_ a_5481_20185# 0.0279f
C2456 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.22939f
C2457 a_13011_19242# sar9b_0.net42 0.22277f
C2458 a_7936_25137# sar9b_0.cyclic_flag_0.FINAL 0.26867f
C2459 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[7] 0.06961f
C2460 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[4] 18.8692f
C2461 sar9b_0.net13 sar9b_0.net42 0.02401f
C2462 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.1588f
C2463 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.02638f
C2464 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A a_25915_15495# 0.01076f
C2465 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.07579f
C2466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.03729f
C2467 VDPWR a_5394_18116# 0.35368f
C2468 sar9b_0.net40 sar9b_0.net55 1.09485f
C2469 sar9b_0.net29 a_13011_20806# 0.01682f
C2470 a_5046_27230# a_5322_27170# 0.1263f
C2471 a_9174_17906# a_9839_17527# 0.19065f
C2472 a_9450_17846# a_9974_17626# 0.04522f
C2473 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A a_59529_15495# 0.01076f
C2474 a_12182_19759# a_12047_19857# 0.35559f
C2475 a_12870_19603# a_13216_19809# 0.07649f
C2476 sar9b_0.net60 uio_out[1] 0.27455f
C2477 a_7926_23234# a_8386_22806# 0.26257f
C2478 a_8202_23174# a_8591_22855# 0.05462f
C2479 single_9b_cdac_1.SW[2] a_9974_17626# 0.02309f
C2480 sar9b_0.net70 sar9b_0._07_ 0.01892f
C2481 a_11434_16874# a_10649_17131# 0.26257f
C2482 tdc_0.OUTP a_10194_16784# 0.02444f
C2483 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.22879f
C2484 a_9258_21842# sar9b_0.net57 0.22486f
C2485 sar9b_0.net55 sar9b_0.net51 0.50241f
C2486 a_8303_23853# sar9b_0.net57 0.04177f
C2487 VDPWR a_11214_25728# 0.25894f
C2488 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 ua[0] 0.12069f
C2489 a_8057_18463# sar9b_0.net48 0.01239f
C2490 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.42509f
C2491 a_5846_17626# sar9b_0.net56 0.02562f
C2492 sar9b_0.net44 a_5046_27230# 0.06448f
C2493 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.11216f
C2494 a_5753_24250# a_6538_24506# 0.26257f
C2495 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.42784f
C2496 sar9b_0.net59 sar9b_0.net36 0.44441f
C2497 sar9b_0.net40 a_11382_19478# 0.06135f
C2498 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.02149f
C2499 sar9b_0._07_ a_4332_23043# 0.07997f
C2500 a_11382_18146# sar9b_0.net73 0.16947f
C2501 sar9b_0.net57 a_5443_19074# 0.25423f
C2502 a_11382_19478# a_11842_19766# 0.26257f
C2503 a_7404_17715# sar9b_0.net6 0.01668f
C2504 sar9b_0.net43 sar9b_0.net49 0.0215f
C2505 a_9730_24138# sar9b_0.net53 0.08408f
C2506 a_6534_17799# sar9b_0.net46 0.2223f
C2507 a_5182_22567# sar9b_0._18_ 0.01534f
C2508 sar9b_0.net32 sar9b_0.net38 0.02088f
C2509 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 3.26837f
C2510 sar9b_0.net14 uo_out[0] 0.26202f
C2511 a_13067_27662# sar9b_0.net28 0.22031f
C2512 sar9b_0.net23 a_8622_26345# 0.03011f
C2513 single_9b_cdac_0.SW[3] clk 0.13418f
C2514 tdc_0.OUTP a_16159_13315# 0.05276f
C2515 sar9b_0.net2 sar9b_0.net74 0.26355f
C2516 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.12358f
C2517 sar9b_0.net36 a_8883_27466# 0.05427f
C2518 a_11008_17491# a_11436_17742# 0.01819f
C2519 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.19143f
C2520 a_5581_20992# sar9b_0._07_ 0.02281f
C2521 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.SW[4] 0.17303f
C2522 sar9b_0.net40 sar9b_0.net38 0.028f
C2523 sar9b_0.net70 sar9b_0.clknet_1_0__leaf_CLK 0.28843f
C2524 sar9b_0.net53 a_11842_22430# 0.09838f
C2525 a_8057_18463# sar9b_0.net46 0.10239f
C2526 a_10378_27170# single_9b_cdac_0.SW[7] 0.01306f
C2527 VDPWR a_4365_25770# 0.1412f
C2528 sar9b_0.net38 sar9b_0.net51 0.1037f
C2529 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0303f
C2530 sar9b_0.net24 sar9b_0.net34 0.14505f
C2531 a_5581_20992# sar9b_0._08_ 0.16775f
C2532 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.19266f
C2533 a_10607_25185# a_10218_24802# 0.06034f
C2534 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.22939f
C2535 VDPWR a_7404_17715# 0.22602f
C2536 single_9b_cdac_0.SW[1] ua[0] 0.14864f
C2537 sar9b_0.net20 a_5674_28147# 0.06614f
C2538 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C2539 VDPWR a_4011_22488# 0.08627f
C2540 sar9b_0.net58 a_3438_27677# 0.2256f
C2541 sar9b_0.net53 a_11842_23762# 0.09947f
C2542 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[4] 0.24199f
C2543 uio_out[1] uio_out[0] 2.82713f
C2544 sar9b_0.net41 a_9634_17478# 0.06387f
C2545 sar9b_0.net31 a_13216_22473# 0.28434f
C2546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A a_45123_15495# 0.01076f
C2547 a_3747_25724# a_4125_25958# 0.0649f
C2548 sar9b_0.net55 sar9b_0.net62 0.19573f
C2549 a_8591_22855# sar9b_0.net37 0.01032f
C2550 a_10284_25707# a_10482_25831# 0.06623f
C2551 sar9b_0.net31 a_11915_27039# 0.03331f
C2552 sar9b_0.net17 sar9b_0.net60 0.14205f
C2553 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[4] 0.0149f
C2554 sar9b_0.net61 a_9974_17626# 0.04925f
C2555 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C2556 a_10470_21795# a_10816_21487# 0.07649f
C2557 a_7404_17715# sar9b_0.net1 0.27002f
C2558 sar9b_0.net6 a_9174_17906# 0.18423f
C2559 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[2] 0.03797f
C2560 VDPWR a_11658_26134# 0.83989f
C2561 a_10335_16817# a_10649_17131# 0.07826f
C2562 a_8098_23762# sar9b_0.net11 0.05862f
C2563 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR 0.75853f
C2564 a_7914_23470# sar9b_0.net54 0.03451f
C2565 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.0303f
C2566 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.3196f
C2567 sar9b_0.net64 sar9b_0._17_ 0.0131f
C2568 sar9b_0.net36 sar9b_0.net12 0.02707f
C2569 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.27795f
C2570 a_7188_22119# a_7193_22459# 0.43491f
C2571 sar9b_0.net52 a_12182_26419# 0.14359f
C2572 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C2573 VDPWR a_3603_28156# 0.4289f
C2574 sar9b_0.net8 sar9b_0.net2 0.02074f
C2575 sar9b_0.net40 sar9b_0.net6 0.05038f
C2576 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.03488f
C2577 ua[4] w_12795_1601# 0.89427f
C2578 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 1.71649f
C2579 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.55985f
C2580 a_11842_19766# sar9b_0.net6 0.01376f
C2581 sar9b_0.net6 sar9b_0.net51 0.0241f
C2582 a_11382_18146# sar9b_0.net50 0.23307f
C2583 sar9b_0.net5 sar9b_0.net39 0.02145f
C2584 VDPWR a_9174_17906# 0.28468f
C2585 single_9b_cdac_1.SW[3] a_11382_18146# 0.03693f
C2586 single_9b_cdac_0.SW[5] ua[0] 0.1911f
C2587 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.17533f
C2588 sar9b_0.net53 sar9b_0.net57 0.08138f
C2589 a_12531_28566# uo_out[1] 0.38317f
C2590 a_10553_18922# sar9b_0.net7 0.06335f
C2591 sar9b_0.net32 VDPWR 1.40875f
C2592 sar9b_0.net27 single_9b_cdac_1.CF[2] 0.07174f
C2593 sar9b_0.net50 a_11859_20574# 0.05205f
C2594 VDPWR a_2892_23070# 0.30728f
C2595 sar9b_0.net63 a_4811_23656# 0.08526f
C2596 a_5748_24381# sar9b_0.net54 0.18387f
C2597 a_21177_7457# th_dif_sw_0.th_sw_1.CKB 2.27999f
C2598 sar9b_0.net38 a_9588_27045# 0.02021f
C2599 a_3156_26115# a_3161_26455# 0.44098f
C2600 a_2706_26108# a_2847_26141# 0.27388f
C2601 a_12588_16784# single_9b_cdac_1.SW[3] 0.02701f
C2602 a_8098_18810# sar9b_0.net5 0.01301f
C2603 single_9b_cdac_0.cdac_sw_9b_0.S[0] a_63626_26990# 0.22513f
C2604 sar9b_0.net43 a_10218_24802# 0.01463f
C2605 VDPWR sar9b_0.net40 1.99954f
C2606 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.B 0.0174f
C2607 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[2] 0.01791f
C2608 a_3206_22432# sar9b_0.net67 0.25532f
C2609 VDPWR a_12870_18271# 0.27198f
C2610 a_13011_19242# a_13216_19809# 0.01179f
C2611 a_25210_17740# single_9b_cdac_1.SW[8] 0.18991f
C2612 sar9b_0.net12 a_10937_25582# 0.02312f
C2613 VDPWR a_11842_19766# 0.23652f
C2614 single_9b_cdac_1.SW[4] th_dif_sw_0.CK 0.04291f
C2615 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[4] 4.15153f
C2616 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C2617 VDPWR sar9b_0.net51 1.04918f
C2618 a_11722_25838# sar9b_0.net12 0.01432f
C2619 sar9b_0.net13 a_10218_24802# 0.02005f
C2620 a_13011_21906# sar9b_0.net27 0.03613f
C2621 a_6954_27466# sar9b_0.net36 0.07226f
C2622 a_7306_19777# sar9b_0.net47 0.19638f
C2623 VDPWR th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.17946f
C2624 VDPWR a_15265_9613# 0.18873f
C2625 a_11430_20935# a_11776_21141# 0.07649f
C2626 sar9b_0.net40 sar9b_0.net1 0.0276f
C2627 uo_out[0] th_dif_sw_0.VCN 0.08774f
C2628 single_9b_cdac_1.cdac_sw_9b_0.S[8] a_24332_16877# 0.59531f
C2629 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 1.55982f
C2630 a_9942_20810# a_10218_20806# 0.1263f
C2631 sar9b_0.net1 sar9b_0.net51 0.16069f
C2632 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 a_58824_26990# 0.14695f
C2633 a_3603_28156# a_4083_28566# 0.03385f
C2634 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] 0.14551f
C2635 a_3438_26345# a_3161_26455# 0.09983f
C2636 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.11216f
C2637 a_10995_28566# VDPWR 0.45062f
C2638 sar9b_0.net4 a_5849_18463# 0.01533f
C2639 a_10830_19068# a_11338_19178# 0.19065f
C2640 a_10649_17131# sar9b_0.net48 0.06775f
C2641 VDPWR a_53154_26999# 1.81495f
C2642 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[5] 0.01887f
C2643 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.04988f
C2644 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_26951_15501# 0.01076f
C2645 a_9162_23174# a_9760_22819# 0.06623f
C2646 sar9b_0.net43 sar9b_0.net11 0.02461f
C2647 sar9b_0.net61 a_8694_20570# 0.18235f
C2648 a_6346_23773# a_6414_23681# 0.35559f
C2649 a_6137_23791# a_6922_23534# 0.26257f
C2650 a_6534_17799# a_6880_17491# 0.07649f
C2651 single_9b_cdac_0.SW[4] a_13067_27662# 0.0479f
C2652 VDPWR a_9130_26198# 0.30205f
C2653 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_60565_15501# 0.01076f
C2654 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[1\] 0.02971f
C2655 a_11008_17491# sar9b_0.net27 0.01194f
C2656 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.01003f
C2657 a_3713_22522# a_3561_22527# 0.22517f
C2658 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[3] 1.84733f
C2659 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 2.82231f
C2660 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[1] 0.21792f
C2661 VDPWR a_10742_21091# 0.20336f
C2662 a_10859_26330# sar9b_0.net36 0.01882f
C2663 a_4934_22432# a_5182_22567# 0.05308f
C2664 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.7611f
C2665 a_53154_26999# single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.59531f
C2666 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.71729f
C2667 a_8591_22855# sar9b_0.net57 0.01229f
C2668 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_1.CF[8] 0.01879f
C2669 a_6642_19448# a_7306_19777# 0.16939f
C2670 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C2671 VDPWR a_13011_20574# 0.42461f
C2672 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07579f
C2673 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.01664f
C2674 ua[0] single_9b_cdac_1.SW[7] 0.13071f
C2675 a_2739_20140# sar9b_0._00_ 0.0764f
C2676 sar9b_0.net31 a_11658_23470# 0.02378f
C2677 sar9b_0.net2 a_9935_24187# 0.06094f
C2678 a_10762_18823# sar9b_0.net48 0.14f
C2679 VDPWR sar9b_0.net62 2.17291f
C2680 a_3747_25724# sar9b_0.clknet_1_1__leaf_CLK 0.10609f
C2681 a_4125_25958# a_4698_25851# 0.04602f
C2682 a_3219_22860# a_3695_23038# 0.08279f
C2683 a_3371_23106# sar9b_0.net65 0.03052f
C2684 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C2685 sar9b_0.net32 sar9b_0.net29 0.02003f
C2686 sar9b_0.net38 a_8115_28566# 0.08106f
C2687 sar9b_0.net8 a_10218_20806# 0.04227f
C2688 sar9b_0.net36 sar9b_0.net5 0.02542f
C2689 VDPWR a_3372_25734# 0.23391f
C2690 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.07517f
C2691 a_11382_26138# a_11658_26134# 0.1263f
C2692 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.01003f
C2693 VDPWR a_13011_17910# 0.46728f
C2694 sar9b_0.net57 a_5196_18116# 0.09147f
C2695 a_7638_19238# sar9b_0.net73 0.17598f
C2696 a_7602_18116# a_8266_18445# 0.16939f
C2697 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.17533f
C2698 a_5849_18463# a_6058_18445# 0.24088f
C2699 a_5844_18123# a_6634_18206# 0.1263f
C2700 a_21684_3438# VDPWR 0.07087f
C2701 ui_in[0] clk 0.23226f
C2702 VDPWR a_9588_27045# 0.85382f
C2703 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.36041f
C2704 tdc_0.OUTN a_8057_17131# 0.03327f
C2705 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C2706 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.04988f
C2707 a_10859_26330# a_10937_25582# 0.01019f
C2708 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C2709 a_6132_23451# sar9b_0.net11 0.06939f
C2710 VDPWR a_9647_21523# 0.27298f
C2711 a_2451_27234# ui_in[0] 0.24933f
C2712 VDPWR a_53154_16877# 1.81495f
C2713 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.7611f
C2714 sar9b_0.net13 a_7338_24802# 0.07649f
C2715 sar9b_0.net52 a_8438_23755# 0.13752f
C2716 sar9b_0.net43 a_11178_20806# 0.01951f
C2717 a_11842_22430# a_12047_22521# 0.09983f
C2718 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[4] 0.02005f
C2719 a_12870_22267# a_12618_22138# 0.27388f
C2720 sar9b_0.net43 sar9b_0.net45 0.12328f
C2721 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[1] 2.07974f
C2722 sar9b_0.net58 a_5742_28392# 0.19468f
C2723 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46159_15501# 0.01076f
C2724 sar9b_0.net26 single_9b_cdac_1.CF[2] 0.03846f
C2725 a_17125_9355# clk 0.02939f
C2726 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C2727 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.05472f
C2728 a_11718_23127# sar9b_0.net11 0.03005f
C2729 a_10070_24286# a_10506_24506# 0.16939f
C2730 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 2.82223f
C2731 tdc_0.phase_detector_0.pd_out_0.B a_15400_11316# 0.48689f
C2732 a_9647_21523# sar9b_0.net1 0.02115f
C2733 a_3014_24136# sar9b_0.clk_div_0.COUNT\[1\] 0.0121f
C2734 VDPWR a_7914_19178# 0.75628f
C2735 a_9363_20826# sar9b_0.net37 0.01328f
C2736 sar9b_0.net42 a_11382_19478# 0.02021f
C2737 a_10548_19053# sar9b_0.net42 0.05396f
C2738 sar9b_0.net8 a_8982_21902# 0.17036f
C2739 sar9b_0._09_ a_5126_20140# 0.01059f
C2740 a_7638_19238# sar9b_0.net48 0.22589f
C2741 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 2.71729f
C2742 sar9b_0.net13 a_10607_25185# 0.06161f
C2743 sar9b_0.net47 a_7978_22202# 0.20624f
C2744 sar9b_0.net30 a_11842_23762# 0.02126f
C2745 sar9b_0.clknet_0_CLK a_4236_21738# 0.03044f
C2746 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.94202f
C2747 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.17533f
C2748 VDPWR uo_out[7] 1.05965f
C2749 a_11178_27466# VDPWR 0.35818f
C2750 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22352f
C2751 a_8622_26345# sar9b_0.net37 0.01006f
C2752 a_12531_28566# a_13164_28398# 0.02384f
C2753 sar9b_0.net64 sar9b_0._12_ 0.3293f
C2754 sar9b_0.net45 a_12560_27128# 0.20749f
C2755 a_12870_23599# a_12618_23470# 0.27388f
C2756 a_11842_23762# a_12047_23853# 0.09983f
C2757 a_6922_23534# sar9b_0.net57 0.06619f
C2758 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[1] 17.5055f
C2759 sar9b_0.net27 a_12870_22267# 0.02852f
C2760 sar9b_0.net43 a_9870_27060# 0.01268f
C2761 sar9b_0.net54 a_6902_25087# 0.12912f
C2762 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07579f
C2763 sar9b_0.net22 single_9b_cdac_0.SW[8] 0.02541f
C2764 sar9b_0.net29 a_13011_20574# 0.02075f
C2765 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.70254f
C2766 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.42784f
C2767 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 ua[0] 0.13461f
C2768 sar9b_0.net11 sar9b_0.net4 0.02493f
C2769 sar9b_0.net59 a_9279_27227# 0.1788f
C2770 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[8] 0.058f
C2771 a_6861_22828# sar9b_0._17_ 0.01915f
C2772 a_3425_20244# a_3723_20140# 0.02614f
C2773 single_9b_cdac_1.CF[1] sar9b_0.net27 0.07881f
C2774 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[8] 4.16613f
C2775 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.0303f
C2776 sar9b_0.net32 single_9b_cdac_0.SW[3] 0.04904f
C2777 a_7498_21109# a_7566_21017# 0.35559f
C2778 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C2779 a_7289_21127# sar9b_0.net56 0.01572f
C2780 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.SW[7] 0.15499f
C2781 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.42015f
C2782 sar9b_0.net27 a_12870_23599# 0.02852f
C2783 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net11 0.01289f
C2784 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 a_39616_26990# 0.14695f
C2785 a_7638_19238# sar9b_0.net46 0.03287f
C2786 single_9b_cdac_0.SW[5] a_12531_28566# 0.03035f
C2787 a_10230_23234# sar9b_0.net53 0.22171f
C2788 VDPWR a_8115_28566# 0.46684f
C2789 sar9b_0.net16 a_5196_19448# 0.27599f
C2790 a_10230_23234# a_10690_22806# 0.26257f
C2791 a_10506_23174# a_10895_22855# 0.05462f
C2792 sar9b_0.net41 a_9546_24506# 0.01299f
C2793 a_10218_27466# sar9b_0.net24 0.03703f
C2794 a_10895_22855# sar9b_0.net74 0.02448f
C2795 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C2796 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22655f
C2797 a_5083_21100# sar9b_0._18_ 0.10881f
C2798 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0._05_ 0.02778f
C2799 a_8334_17021# sar9b_0.net5 0.01036f
C2800 a_11178_24802# a_10932_25713# 0.02278f
C2801 a_7138_27758# a_7914_27466# 0.3578f
C2802 a_9760_22819# sar9b_0.net11 0.04919f
C2803 a_9138_27163# sar9b_0.net37 0.04632f
C2804 a_8726_22954# sar9b_0.net54 0.14f
C2805 sar9b_0.net40 a_6678_27470# 0.17609f
C2806 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C2807 VDPWR a_3090_27163# 0.37894f
C2808 a_3206_22432# sar9b_0.clknet_1_0__leaf_CLK 0.05926f
C2809 sar9b_0.net33 sar9b_0.net30 0.02513f
C2810 sar9b_0.net49 sar9b_0.net38 0.54905f
C2811 a_11859_21906# sar9b_0.net39 0.01794f
C2812 sar9b_0._07_ a_5481_20185# 0.02028f
C2813 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C2814 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[5] 0.0149f
C2815 a_11430_27595# sar9b_0.net59 0.17391f
C2816 a_8334_18353# sar9b_0.net5 0.06948f
C2817 a_10926_17021# single_9b_cdac_1.SW[2] 0.01526f
C2818 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.38397f
C2819 single_9b_cdac_1.CF[8] sar9b_0.net27 0.09104f
C2820 a_9270_24566# sar9b_0.net62 0.16799f
C2821 sar9b_0.net8 sar9b_0.net39 0.1827f
C2822 sar9b_0.net5 single_9b_cdac_1.CF[0] 0.02589f
C2823 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.75853f
C2824 a_11382_18146# a_11658_18142# 0.1263f
C2825 single_9b_cdac_1.cdac_sw_9b_0.S[3] a_48343_16877# 0.59531f
C2826 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[5] 0.01513f
C2827 sar9b_0.net36 a_10035_19474# 0.01195f
C2828 sar9b_0.net42 sar9b_0.net6 0.02813f
C2829 VDPWR a_4811_23656# 0.24092f
C2830 a_4812_28371# sar9b_0.net60 0.02169f
C2831 sar9b_0.net38 uo_out[6] 0.72968f
C2832 a_8202_23174# clk 0.02077f
C2833 sar9b_0.net43 sar9b_0.net13 0.02924f
C2834 sar9b_0.net18 sar9b_0.net60 0.03658f
C2835 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.12898f
C2836 a_12618_18142# a_13216_18477# 0.06623f
C2837 a_4698_25851# sar9b_0.clknet_1_1__leaf_CLK 0.02594f
C2838 a_10402_27758# sar9b_0.net34 0.01319f
C2839 a_11842_26426# a_12870_26263# 0.07826f
C2840 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.clknet_1_1__leaf_CLK 0.04637f
C2841 a_21177_7457# th_dif_sw_0.VCP 0.0867f
C2842 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[3] 0.01995f
C2843 single_9b_cdac_0.SW[1] sar9b_0.net28 0.04119f
C2844 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.7611f
C2845 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[3] 0.06019f
C2846 sar9b_0.net63 sar9b_0.net11 0.60944f
C2847 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22497f
C2848 sar9b_0.net5 single_9b_cdac_1.SW[2] 0.0302f
C2849 single_9b_cdac_1.SW[6] th_dif_sw_0.CK 0.11297f
C2850 a_6378_24802# a_6562_25094# 0.44532f
C2851 sar9b_0.net36 sar9b_0.net74 0.21507f
C2852 sar9b_0.net41 single_9b_cdac_1.SW[1] 0.01957f
C2853 VDPWR a_3747_25724# 0.37697f
C2854 a_9154_20142# a_9359_20191# 0.09983f
C2855 sar9b_0.net58 a_3545_26914# 0.10032f
C2856 VDPWR sar9b_0.net42 1.57366f
C2857 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.01751f
C2858 sar9b_0.net66 sar9b_0._05_ 0.18138f
C2859 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.02666f
C2860 sar9b_0._06_ a_13067_27662# 0.01122f
C2861 a_12588_16784# tdc_0.OUTP 0.28954f
C2862 sar9b_0.net43 a_5298_24499# 0.06128f
C2863 a_7188_22119# sar9b_0.net47 0.17293f
C2864 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.3601f
C2865 a_6540_22112# sar9b_0._02_ 0.02465f
C2866 sar9b_0.net8 a_12435_20806# 0.08962f
C2867 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.0303f
C2868 a_7138_27758# a_7343_27849# 0.09983f
C2869 m2_23774_17236# a_24332_16877# 0.01541f
C2870 a_3262_24141# sar9b_0.clknet_1_1__leaf_CLK 0.01978f
C2871 th_dif_sw_0.VCP ua[0] 1.04697f
C2872 a_6861_22828# clk 0.01643f
C2873 sar9b_0._02_ sar9b_0.net39 0.04135f
C2874 dw_12589_1395# th_dif_sw_0.th_sw_1.CKB 0.24188f
C2875 a_12684_20379# sar9b_0.net51 0.25465f
C2876 a_11658_23470# a_12182_23755# 0.05022f
C2877 sar9b_0.clk_div_0.COUNT\[3\] a_4755_22138# 0.02068f
C2878 sar9b_0.net27 single_9b_cdac_1.CF[3] 0.12277f
C2879 sar9b_0.net27 sar9b_0.net28 0.01665f
C2880 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.12431f
C2881 sar9b_0.net35 sar9b_0.net73 0.26229f
C2882 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_50962_29911# 0.01076f
C2883 a_5046_27230# a_5506_26802# 0.26257f
C2884 single_9b_cdac_1.SW[8] sar9b_0.net5 0.04994f
C2885 VDPWR a_6636_20780# 0.20851f
C2886 a_7978_22202# sar9b_0.net57 0.01265f
C2887 sar9b_0.net18 uio_out[0] 0.11108f
C2888 clk sar9b_0.net37 0.04254f
C2889 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C2890 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[1] 0.21746f
C2891 sar9b_0.net49 a_8970_20510# 0.17751f
C2892 a_8345_26455# a_8554_26437# 0.24088f
C2893 sar9b_0.net2 sar9b_0.net73 0.03106f
C2894 sar9b_0.net6 a_5849_18463# 0.01813f
C2895 a_3713_22522# a_3027_22138# 0.27693f
C2896 a_3822_27060# a_4330_27170# 0.19065f
C2897 single_9b_cdac_1.CF[1] sar9b_0.net26 0.05711f
C2898 a_11859_17910# single_9b_cdac_1.SW[3] 0.01458f
C2899 sar9b_0.net46 a_4771_18260# 0.03699f
C2900 sar9b_0.net74 a_10937_25582# 0.05953f
C2901 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] 3.10229f
C2902 a_3540_27045# a_3754_26815# 0.05022f
C2903 a_3713_22522# sar9b_0.net65 0.02109f
C2904 a_11722_25838# sar9b_0.net74 0.21463f
C2905 VDPWR sar9b_0.net49 2.96485f
C2906 a_3695_23038# sar9b_0.clknet_0_CLK 0.01593f
C2907 VDPWR a_9162_23174# 0.37599f
C2908 sar9b_0.net56 sar9b_0.net47 0.18012f
C2909 a_10649_17131# sar9b_0.net27 0.01161f
C2910 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42509f
C2911 sar9b_0.net57 sar9b_0._17_ 0.02056f
C2912 sar9b_0.net32 sar9b_0.net23 0.04971f
C2913 a_6137_23791# clk 0.01311f
C2914 a_7402_22441# a_7470_22349# 0.35559f
C2915 sar9b_0.net60 a_5674_28147# 0.02547f
C2916 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C2917 a_5151_28559# a_5460_28377# 0.07766f
C2918 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.12367f
C2919 sar9b_0.net55 sar9b_0.net11 0.02067f
C2920 single_9b_cdac_1.SW[0] sar9b_0.net37 0.06363f
C2921 a_10378_27170# sar9b_0.net59 0.22839f
C2922 VDPWR uo_out[6] 0.80816f
C2923 sar9b_0.net8 sar9b_0.net36 0.02461f
C2924 sar9b_0.net49 a_10218_21842# 0.2811f
C2925 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.0313f
C2926 a_11722_25838# sar9b_0.net31 0.01201f
C2927 sar9b_0.net49 sar9b_0.net1 0.10608f
C2928 sar9b_0.net61 sar9b_0.net5 0.55611f
C2929 a_10227_18142# sar9b_0.net38 0.06078f
C2930 a_10218_24802# sar9b_0.net38 0.02016f
C2931 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C2932 sar9b_0.net1 a_9162_23174# 0.01832f
C2933 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.S[8] 0.58106f
C2934 sar9b_0.net56 sar9b_0.net37 1.42615f
C2935 a_12435_24802# sar9b_0.net27 0.01432f
C2936 sar9b_0.net43 sar9b_0.net4 0.0207f
C2937 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C2938 sar9b_0.net35 sar9b_0.net48 0.03579f
C2939 sar9b_0.net43 sar9b_0._15_ 0.16183f
C2940 a_12684_20379# a_13011_20574# 0.08132f
C2941 VDPWR a_5849_18463# 0.21922f
C2942 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.12431f
C2943 a_7193_22459# sar9b_0.net62 0.02169f
C2944 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.02778f
C2945 sar9b_0.net13 sar9b_0.net4 0.20455f
C2946 sar9b_0.net20 a_6250_28502# 0.0646f
C2947 tdc_0.OUTP a_10649_17131# 0.06549f
C2948 sar9b_0.net13 sar9b_0._15_ 0.03815f
C2949 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.7611f
C2950 sar9b_0.net2 sar9b_0.net48 0.03105f
C2951 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.07579f
C2952 a_4947_20140# sar9b_0._10_ 0.0624f
C2953 a_9939_28566# sar9b_0.net24 0.05176f
C2954 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.03729f
C2955 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.64863f
C2956 a_8595_17910# sar9b_0.net6 0.03608f
C2957 VDPWR tdc_0.phase_detector_0.INN 0.51155f
C2958 a_10070_24286# sar9b_0.net53 0.1338f
C2959 VDPWR sar9b_0.net14 0.26926f
C2960 sar9b_0.net38 sar9b_0.net11 0.02613f
C2961 single_9b_cdac_1.cdac_sw_9b_0.S[3] th_dif_sw_0.VCP 27.3302f
C2962 a_11842_23762# clk 0.01052f
C2963 single_9b_cdac_0.SW[8] uo_out[3] 0.28955f
C2964 a_9996_16784# sar9b_0.net6 0.05001f
C2965 a_35519_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.01076f
C2966 sar9b_0.net23 a_9130_26198# 0.03663f
C2967 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.22879f
C2968 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B 0.36961f
C2969 sar9b_0.net27 a_13011_24570# 0.04167f
C2970 sar9b_0.net35 sar9b_0.net46 0.32715f
C2971 sar9b_0.net7 sar9b_0.net5 0.0215f
C2972 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C2973 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.7611f
C2974 sar9b_0.net36 sar9b_0.net34 0.04627f
C2975 sar9b_0.net16 sar9b_0.net46 0.16498f
C2976 a_6954_27466# a_7539_28566# 0.03399f
C2977 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.71649f
C2978 a_11436_17742# a_11859_17910# 0.05125f
C2979 sar9b_0.net28 single_9b_cdac_1.SW[7] 0.0883f
C2980 a_5298_24499# sar9b_0._15_ 0.079f
C2981 sar9b_0.net53 a_12870_22267# 0.17311f
C2982 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[5] 0.02021f
C2983 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[4] 0.05054f
C2984 sar9b_0.net2 single_9b_cdac_1.SW[3] 0.19941f
C2985 sar9b_0.net65 a_4236_21738# 0.08898f
C2986 a_5506_17478# sar9b_0.net4 0.03413f
C2987 a_29134_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.23864f
C2988 sar9b_0.net44 a_5322_27170# 0.25565f
C2989 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.33229f
C2990 tdc_0.OUTN sar9b_0.net46 0.09655f
C2991 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[8] 0.26707f
C2992 VDPWR a_4698_25851# 0.01249f
C2993 VDPWR a_8595_17910# 0.49252f
C2994 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[6] 4.16106f
C2995 VDPWR sar9b_0.clk_div_0.COUNT\[3\] 0.34467f
C2996 sar9b_0.net53 a_12870_23599# 0.17313f
C2997 sar9b_0.net41 a_9974_17626# 0.06988f
C2998 th_dif_sw_0.CK tdc_0.RDY 0.05459f
C2999 VDPWR a_9996_16784# 0.1892f
C3000 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.26707f
C3001 sar9b_0.net43 sar9b_0.net63 0.0282f
C3002 a_10482_25831# a_10623_25895# 0.27388f
C3003 a_7188_22119# sar9b_0.net57 0.01211f
C3004 a_3161_27787# a_3438_27677# 0.09983f
C3005 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.71729f
C3006 single_9b_cdac_1.SW[5] clk 0.08628f
C3007 single_9b_cdac_0.SW[4] a_13164_28398# 0.01356f
C3008 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C3009 sar9b_0._01_ a_4947_20140# 0.16646f
C3010 a_5506_17478# a_5322_17846# 0.43491f
C3011 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 3.04383f
C3012 sar9b_0.net57 clk 0.05645f
C3013 VDPWR a_11842_26426# 0.23378f
C3014 VDPWR a_10227_18142# 0.43915f
C3015 a_2508_20780# sar9b_0.clknet_0_CLK 0.47881f
C3016 VDPWR a_10218_24802# 0.81345f
C3017 VDPWR a_13216_19809# 0.21451f
C3018 sar9b_0._17_ sar9b_0.clk_div_0.COUNT\[1\] 0.15221f
C3019 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.12431f
C3020 sar9b_0.net10 sar9b_0.net54 0.15482f
C3021 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.22879f
C3022 sar9b_0.net59 sar9b_0.cyclic_flag_0.FINAL 0.74539f
C3023 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.28523f
C3024 uo_out[0] uio_in[7] 0.03102f
C3025 sar9b_0.net38 sar9b_0.net45 0.14791f
C3026 a_7289_21127# sar9b_0.net51 0.06342f
C3027 single_9b_cdac_1.CF[5] sar9b_0.net27 0.03004f
C3028 single_9b_cdac_0.SW[4] sar9b_0.net27 0.05602f
C3029 sar9b_0.net52 a_12618_26134# 0.26209f
C3030 single_9b_cdac_0.SW[0] ua[0] 0.15351f
C3031 VDPWR a_5010_28495# 0.34506f
C3032 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[5] 1.8421f
C3033 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[0] 0.02181f
C3034 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[4] 10.4962f
C3035 sar9b_0.cyclic_flag_0.FINAL a_8883_27466# 0.28976f
C3036 VDPWR a_3262_24141# 0.01376f
C3037 sar9b_0.net54 a_6538_24506# 0.22653f
C3038 sar9b_0.net58 a_4365_25770# 0.01101f
C3039 a_10607_25185# sar9b_0.net38 0.01125f
C3040 a_12435_24802# sar9b_0.net26 0.09225f
C3041 single_9b_cdac_1.CF[2] single_9b_cdac_0.SW[0] 0.35203f
C3042 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.42509f
C3043 sar9b_0.net56 sar9b_0.net57 0.1667f
C3044 a_11382_18146# a_12047_18525# 0.19065f
C3045 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net4 0.02026f
C3046 sar9b_0._06_ uo_out[1] 0.0432f
C3047 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.05472f
C3048 VDPWR sar9b_0.net11 1.08113f
C3049 a_30717_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.01076f
C3050 VDPWR sar9b_0.net66 0.70022f
C3051 sar9b_0.net70 a_3027_21906# 0.15443f
C3052 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.28033f
C3053 th_dif_sw_0.th_sw_1.CKB dw_17224_1400# 0.24436f
C3054 a_11436_17742# sar9b_0.net2 0.28173f
C3055 a_6282_27170# a_6534_27123# 0.27388f
C3056 a_5322_17846# sar9b_0.net4 0.02133f
C3057 sar9b_0.net60 a_5484_23444# 0.01027f
C3058 sar9b_0.net9 a_10506_23174# 0.21399f
C3059 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.38397f
C3060 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.01751f
C3061 sar9b_0.net9 sar9b_0.net74 0.10219f
C3062 a_2847_26141# a_3161_26455# 0.07826f
C3063 a_13011_16810# th_dif_sw_0.CK 0.0156f
C3064 sar9b_0.net60 a_4947_20140# 0.08548f
C3065 sar9b_0.net1 sar9b_0.net11 0.03134f
C3066 a_10762_18823# sar9b_0.net26 0.06684f
C3067 sar9b_0.net52 a_10402_25094# 0.0792f
C3068 sar9b_0.net43 sar9b_0.net55 0.27955f
C3069 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.84061f
C3070 VDPWR sar9b_0._09_ 0.86773f
C3071 VDPWR a_12870_19603# 0.27172f
C3072 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C3073 a_8098_23762# a_9126_23599# 0.07826f
C3074 a_11915_28371# sar9b_0.net25 0.11385f
C3075 a_10218_27466# a_10402_27758# 0.44532f
C3076 a_7138_27758# sar9b_0.net36 0.13653f
C3077 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.3601f
C3078 a_5235_27466# sar9b_0.net19 0.19875f
C3079 sar9b_0.net59 a_5046_27230# 0.01797f
C3080 VDPWR th_dif_sw_0.VCN 1.99513f
C3081 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[6] 0.0149f
C3082 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.81428f
C3083 a_7289_21127# sar9b_0.net62 0.02399f
C3084 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.0174f
C3085 sar9b_0.net59 a_4812_28371# 0.01553f
C3086 a_9942_20810# a_10402_21098# 0.26257f
C3087 sar9b_0.net31 sar9b_0.net10 0.16278f
C3088 sar9b_0.net57 sar9b_0._12_ 0.01983f
C3089 sar9b_0.net18 sar9b_0.net59 0.09486f
C3090 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.19266f
C3091 a_3946_26198# a_3161_26455# 0.26257f
C3092 sar9b_0.net18 a_3156_27447# 0.02909f
C3093 a_21177_7457# th_dif_sw_0.CKB 0.6816f
C3094 sar9b_0.net29 a_13216_19809# 0.27892f
C3095 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] 54.8348f
C3096 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C3097 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.net39 0.07149f
C3098 sar9b_0.net36 a_10528_20155# 0.0105f
C3099 single_9b_cdac_0.SW[7] uo_out[3] 0.06777f
C3100 VDPWR a_7338_24802# 0.35888f
C3101 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C3102 sar9b_0.net63 sar9b_0.net4 0.04374f
C3103 sar9b_0.net8 single_9b_cdac_1.SW[8] 0.05906f
C3104 sar9b_0.net60 a_6102_24806# 0.02205f
C3105 a_11859_17910# sar9b_0.net27 0.05667f
C3106 a_10194_16784# single_9b_cdac_1.SW[0] 0.02286f
C3107 sar9b_0.net63 sar9b_0._15_ 0.04597f
C3108 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.71729f
C3109 sar9b_0.net43 sar9b_0.net38 0.17602f
C3110 ui_in[5] ui_in[4] 0.03102f
C3111 uo_out[7] ui_in[0] 0.06786f
C3112 a_5046_27230# a_4330_27170# 0.03811f
C3113 VDPWR a_8098_23762# 0.25671f
C3114 a_4210_22378# sar9b_0.clknet_0_CLK 0.03169f
C3115 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.62443f
C3116 a_10707_23470# sar9b_0.net53 0.05847f
C3117 sar9b_0.net27 a_4771_18260# 0.02095f
C3118 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.71729f
C3119 VDPWR a_11178_20806# 0.35985f
C3120 a_29134_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.23864f
C3121 VDPWR sar9b_0.net45 1.95717f
C3122 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02652f
C3123 a_3946_26198# sar9b_0.net35 0.17078f
C3124 clk sar9b_0.clk_div_0.COUNT\[1\] 0.08722f
C3125 a_11859_21906# sar9b_0.net9 0.06677f
C3126 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[2\] 1.06971f
C3127 sar9b_0.net13 sar9b_0.net38 0.02597f
C3128 a_7097_19795# a_7306_19777# 0.24088f
C3129 sar9b_0.net40 sar9b_0.net58 0.01707f
C3130 sar9b_0.net73 sar9b_0.net39 0.09841f
C3131 sar9b_0.net9 sar9b_0.net8 0.25322f
C3132 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.81428f
C3133 a_3014_24136# sar9b_0.net68 0.11549f
C3134 a_8595_17910# a_8052_16791# 0.03549f
C3135 VDPWR a_10607_25185# 0.25735f
C3136 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C3137 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0303f
C3138 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 ua[0] 0.12088f
C3139 a_8334_17021# a_8057_17131# 0.09983f
C3140 sar9b_0.net7 a_9942_20810# 0.21228f
C3141 a_9174_17906# sar9b_0.net37 0.03941f
C3142 th_dif_sw_0.CKB ua[0] 0.02532f
C3143 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK 0.31513f
C3144 a_3695_23038# sar9b_0.net65 0.11374f
C3145 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.03729f
C3146 sar9b_0.net8 sar9b_0.net61 0.19337f
C3147 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 3.10626f
C3148 sar9b_0.net8 a_10402_21098# 0.16495f
C3149 a_8940_24402# sar9b_0.net2 0.24809f
C3150 a_11382_26138# a_11842_26426# 0.26257f
C3151 VDPWR a_2918_20140# 0.90101f
C3152 sar9b_0.net57 a_5394_18116# 0.02101f
C3153 sar9b_0.net47 sar9b_0.net40 0.3867f
C3154 sar9b_0.net40 a_6861_22828# 0.01547f
C3155 a_8057_18463# a_8266_18445# 0.24088f
C3156 single_9b_cdac_1.cdac_sw_9b_0.S[2] a_53154_16877# 0.59531f
C3157 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[2] 0.42016f
C3158 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.23864f
C3159 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C3160 m2_23774_26966# VDPWR 0.19016f
C3161 sar9b_0.net47 sar9b_0.net51 0.49323f
C3162 sar9b_0._02_ a_6444_21738# 0.25486f
C3163 single_9b_cdac_1.SW[0] a_10410_17846# 0.04572f
C3164 VDPWR a_9870_27060# 0.26408f
C3165 VDPWR uo_out[0] 0.86559f
C3166 sar9b_0.net40 sar9b_0.net37 0.05789f
C3167 sar9b_0.net42 a_10742_25087# 0.02075f
C3168 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.45521f
C3169 a_8202_23174# sar9b_0.net62 0.02827f
C3170 a_5682_23444# sar9b_0.net11 0.04944f
C3171 sar9b_0.net41 sar9b_0.net59 0.1373f
C3172 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.84423f
C3173 sar9b_0.net48 sar9b_0.net39 0.0236f
C3174 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.clknet_1_1__leaf_CLK 0.19127f
C3175 sar9b_0.net51 sar9b_0.net37 0.03332f
C3176 sar9b_0.net13 a_9165_24988# 0.11202f
C3177 sar9b_0.net52 a_8874_23470# 0.26484f
C3178 a_12618_22138# a_13216_22473# 0.06623f
C3179 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36322f
C3180 a_8691_28566# uo_out[6] 0.03562f
C3181 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.17533f
C3182 sar9b_0.net55 sar9b_0.net4 0.82102f
C3183 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.36044f
C3184 sar9b_0.net7 a_11859_21906# 0.21737f
C3185 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.05279f
C3186 sar9b_0.clk_div_0.COUNT\[0\] a_4332_23043# 0.84737f
C3187 sar9b_0.net40 a_6137_23791# 0.01879f
C3188 sar9b_0.net2 a_10506_24506# 0.076f
C3189 a_10335_16817# sar9b_0.net36 0.02026f
C3190 sar9b_0.net35 sar9b_0.net27 0.08696f
C3191 a_11776_27801# sar9b_0.net25 0.26874f
C3192 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.03436f
C3193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C3194 sar9b_0.net7 sar9b_0.net8 0.39284f
C3195 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] 3.11836f
C3196 sar9b_0.net16 sar9b_0.net27 0.02393f
C3197 single_9b_cdac_0.SW[1] a_58824_26990# 0.18991f
C3198 a_7890_26108# sar9b_0.cyclic_flag_0.FINAL 0.083f
C3199 a_6642_19448# sar9b_0.net40 0.06124f
C3200 a_8098_18810# sar9b_0.net48 0.09937f
C3201 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[2\] 0.02107f
C3202 sar9b_0.net2 sar9b_0.net27 0.34591f
C3203 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[7] 0.02149f
C3204 a_10230_23234# clk 0.01685f
C3205 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.12077f
C3206 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C3207 a_9942_27470# a_10607_27849# 0.19065f
C3208 a_12491_27662# VDPWR 0.49074f
C3209 a_9130_26198# sar9b_0.net37 0.01529f
C3210 a_6738_22112# a_6879_22145# 0.27388f
C3211 a_13164_28398# sar9b_0._06_ 0.28405f
C3212 sar9b_0.net43 VDPWR 3.08648f
C3213 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[0] 0.47599f
C3214 tdc_0.OUTN sar9b_0.net27 0.2611f
C3215 a_12618_23470# a_13216_23805# 0.06623f
C3216 single_9b_cdac_1.CF[1] single_9b_cdac_0.SW[0] 0.32684f
C3217 sar9b_0.net70 a_3219_22860# 0.03435f
C3218 VDPWR a_13011_19242# 0.48316f
C3219 sar9b_0.net27 a_13216_22473# 0.01241f
C3220 sar9b_0.net50 sar9b_0.net39 0.78191f
C3221 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] 0.26612f
C3222 single_9b_cdac_1.cdac_sw_9b_0.S[0] ua[0] 1.20078f
C3223 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[7] 0.0149f
C3224 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A a_40321_15495# 0.01076f
C3225 single_9b_cdac_1.SW[3] sar9b_0.net39 0.0537f
C3226 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.36674f
C3227 sar9b_0.net47 sar9b_0.net62 0.38866f
C3228 sar9b_0.net59 a_9593_26914# 0.11113f
C3229 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.6919f
C3230 VDPWR sar9b_0.net13 2.18619f
C3231 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.12431f
C3232 sar9b_0.net41 a_9900_19047# 0.01957f
C3233 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.28523f
C3234 sar9b_0.net36 sar9b_0.net73 0.03096f
C3235 tdc_0.OUTP sar9b_0.net2 0.24126f
C3236 a_10506_24506# a_10758_24459# 0.27388f
C3237 sar9b_0.net27 sar9b_0._06_ 0.01706f
C3238 sar9b_0.net27 a_13216_23805# 0.01206f
C3239 sar9b_0.net63 sar9b_0.clknet_1_1__leaf_CLK 0.02378f
C3240 a_8098_18810# sar9b_0.net46 0.03666f
C3241 single_9b_cdac_0.SW[5] sar9b_0._06_ 0.01662f
C3242 sar9b_0.net62 sar9b_0.net37 0.04598f
C3243 single_9b_cdac_1.CF[2] clk 0.09194f
C3244 a_12182_26419# a_12618_26134# 0.16939f
C3245 sar9b_0.net33 a_11658_26134# 0.07465f
C3246 tdc_0.OUTP tdc_0.OUTN 1.54073f
C3247 a_8019_17910# sar9b_0.net5 0.03181f
C3248 sar9b_0.net41 sar9b_0.net12 0.51525f
C3249 VDPWR a_10662_17799# 0.26449f
C3250 VDPWR a_12560_27128# 0.33605f
C3251 single_9b_cdac_1.SW[0] ua[0] 1.99402f
C3252 a_8842_16874# sar9b_0.net5 0.04569f
C3253 single_9b_cdac_0.cdac_sw_9b_0.S[3] ua[0] 1.59042f
C3254 a_8166_27595# a_7914_27466# 0.27388f
C3255 VDPWR a_3754_26815# 0.20695f
C3256 single_9b_cdac_0.SW[3] th_dif_sw_0.VCN 0.09453f
C3257 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[0] 3.80682f
C3258 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[6] 0.02056f
C3259 VDPWR a_3540_27045# 0.77744f
C3260 sar9b_0.net63 sar9b_0.net55 0.27808f
C3261 sar9b_0.net58 uo_out[7] 0.13384f
C3262 VDPWR a_5298_24499# 0.32802f
C3263 single_9b_cdac_0.SW[2] a_13067_27662# 0.3597f
C3264 sar9b_0.net61 a_8057_17131# 0.03749f
C3265 sar9b_0.net19 a_3545_26914# 0.17405f
C3266 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[8] 4.67496f
C3267 single_9b_cdac_1.CF[2] single_9b_cdac_1.SW[0] 0.22502f
C3268 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0313f
C3269 a_8842_18206# sar9b_0.net5 0.21948f
C3270 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[7] 0.31534f
C3271 a_9942_20810# a_10607_21189# 0.19065f
C3272 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.3196f
C3273 VDPWR a_8874_19178# 0.41712f
C3274 sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# 0.35818f
C3275 a_11382_18146# a_11842_18434# 0.26257f
C3276 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.30106f
C3277 sar9b_0.net36 sar9b_0.net48 0.17317f
C3278 VDPWR a_5506_17478# 0.21624f
C3279 VDPWR a_6132_23451# 0.78916f
C3280 sar9b_0.net20 sar9b_0.net60 0.0552f
C3281 VDPWR a_8340_26115# 0.87266f
C3282 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.25152f
C3283 a_6767_25185# a_6102_24806# 0.19065f
C3284 VDPWR a_5126_20140# 0.84448f
C3285 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[7] 0.363f
C3286 sar9b_0.net17 a_2847_27473# 0.02024f
C3287 sar9b_0.net42 a_11339_27039# 0.01795f
C3288 VDPWR a_5628_19768# 0.19326f
C3289 dw_12589_1395# a_10166_3438# 26.7601f
C3290 uo_out[6] ui_in[0] 0.06786f
C3291 single_9b_cdac_1.SW[5] sar9b_0.net40 0.09333f
C3292 sar9b_0.net32 sar9b_0.net33 0.02518f
C3293 sar9b_0._03_ a_4698_25851# 0.11739f
C3294 VDPWR a_11718_23127# 0.26767f
C3295 a_11658_19474# a_11859_20574# 0.03761f
C3296 a_2835_24136# a_3014_24136# 0.54426f
C3297 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.22513f
C3298 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.42784f
C3299 single_9b_cdac_1.CF[2] a_13011_20806# 0.01099f
C3300 a_10182_20463# sar9b_0.net51 0.04388f
C3301 sar9b_0.net40 sar9b_0.net57 0.02758f
C3302 a_12491_27662# sar9b_0.net29 0.22249f
C3303 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C3304 a_11436_17742# sar9b_0.net39 0.01601f
C3305 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.95338f
C3306 VDPWR a_6867_16810# 0.26271f
C3307 a_9546_24506# a_10227_23490# 0.02456f
C3308 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.95338f
C3309 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.47485f
C3310 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C3311 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.75853f
C3312 a_6378_24802# a_7590_24931# 0.07766f
C3313 sar9b_0.net60 a_6250_28502# 0.06687f
C3314 single_9b_cdac_1.CF[6] sar9b_0.net27 0.05684f
C3315 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 2.81718f
C3316 VDPWR a_4125_25958# 0.4305f
C3317 sar9b_0._09_ a_4072_19474# 0.06295f
C3318 a_9359_20191# a_9494_20290# 0.35559f
C3319 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[5] 0.09395f
C3320 a_6678_27470# sar9b_0.net45 0.08442f
C3321 sar9b_0._09_ sar9b_0.net71 0.06932f
C3322 sar9b_0.net48 a_5844_18123# 0.18591f
C3323 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.28523f
C3324 sar9b_0.cyclic_flag_0.FINAL sar9b_0.net54 0.09984f
C3325 sar9b_0.net1 a_6867_16810# 0.1431f
C3326 a_13011_21906# a_13011_20806# 0.0246f
C3327 sar9b_0.net58 a_3090_27163# 0.26444f
C3328 sar9b_0.net22 a_8883_27466# 0.02815f
C3329 single_9b_cdac_1.SW[3] sar9b_0.net36 0.01142f
C3330 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.12431f
C3331 sar9b_0.net8 a_10607_21189# 0.01911f
C3332 sar9b_0.net60 sar9b_0.net44 0.64939f
C3333 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.28523f
C3334 sar9b_0.net26 sar9b_0.net2 0.02343f
C3335 single_9b_cdac_1.CF[3] single_9b_cdac_0.SW[0] 0.40374f
C3336 VDPWR sar9b_0.net4 1.04258f
C3337 sar9b_0.net41 a_9930_20510# 0.02662f
C3338 sar9b_0.net28 single_9b_cdac_0.SW[0] 0.1354f
C3339 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 1.71649f
C3340 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 2.81428f
C3341 a_10218_24802# a_10742_25087# 0.05022f
C3342 VDPWR sar9b_0._15_ 0.37538f
C3343 a_4755_22138# sar9b_0.clknet_1_1__leaf_CLK 0.22079f
C3344 sar9b_0.net24 uo_out[2] 0.09027f
C3345 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 3.27833f
C3346 sar9b_0._14_ sar9b_0._15_ 0.01749f
C3347 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.7611f
C3348 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.69086f
C3349 a_11658_23470# a_12618_23470# 0.03432f
C3350 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.net64 0.02988f
C3351 a_7692_26108# sar9b_0.net59 0.04276f
C3352 VDPWR sar9b_0.clk_div_0.COUNT\[2\] 1.36928f
C3353 sar9b_0.net20 uio_out[0] 0.01201f
C3354 sar9b_0.net1 sar9b_0.net4 0.01778f
C3355 a_11434_16874# sar9b_0.net61 0.25057f
C3356 sar9b_0.net43 a_9270_24566# 0.05226f
C3357 VDPWR a_5761_21100# 0.01372f
C3358 single_9b_cdac_1.SW[5] a_39616_17740# 0.18991f
C3359 sar9b_0._14_ sar9b_0.clk_div_0.COUNT\[2\] 0.02642f
C3360 sar9b_0.net24 a_9802_26815# 0.01411f
C3361 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0313f
C3362 tdc_0.phase_detector_0.INP a_15400_11316# 0.02415f
C3363 a_4210_22378# a_3027_22138# 0.0649f
C3364 VDPWR a_5322_17846# 0.85398f
C3365 sar9b_0.net52 sar9b_0.net12 0.59278f
C3366 a_8334_18353# sar9b_0.net73 0.02504f
C3367 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C3368 sar9b_0.clknet_0_CLK a_2508_23444# 0.46608f
C3369 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C3370 w_17430_1606# ua[3] 0.88896f
C3371 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 2.71729f
C3372 a_11008_17491# a_10803_18142# 0.01179f
C3373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.19266f
C3374 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.26427f
C3375 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.42509f
C3376 a_7638_23474# a_7914_23470# 0.1263f
C3377 VDPWR a_9760_22819# 0.20965f
C3378 single_9b_cdac_1.cdac_sw_9b_0.S[8] a_25210_17740# 0.22352f
C3379 sar9b_0._07_ a_4947_20140# 0.02502f
C3380 sar9b_0.net57 sar9b_0.net62 0.5484f
C3381 single_9b_cdac_1.SW[5] a_13011_17910# 0.02888f
C3382 sar9b_0.net41 sar9b_0.net5 0.02649f
C3383 VDPWR a_38738_26999# 1.81495f
C3384 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.75815f
C3385 a_5460_28377# a_5465_28246# 0.44532f
C3386 sar9b_0.clknet_0_CLK sar9b_0.net39 0.08885f
C3387 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.81428f
C3388 dw_12589_1395# a_10254_2858# 1.98316f
C3389 VDPWR a_57946_16877# 1.81495f
C3390 uio_in[2] uio_in[1] 0.03102f
C3391 sar9b_0.net21 a_6880_26815# 0.2711f
C3392 sar9b_0.net1 a_9760_22819# 0.0139f
C3393 sar9b_0.net3 a_2547_28132# 0.27678f
C3394 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.95338f
C3395 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.84061f
C3396 a_12491_27662# single_9b_cdac_0.SW[3] 0.38351f
C3397 a_10239_19235# a_10553_18922# 0.07826f
C3398 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.69086f
C3399 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[0] 0.01887f
C3400 a_8874_19178# a_9472_18823# 0.06623f
C3401 VDPWR a_6058_18445# 0.20217f
C3402 a_3180_19448# sar9b_0._00_ 0.1679f
C3403 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.62443f
C3404 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.42509f
C3405 a_5506_26802# a_5322_27170# 0.43491f
C3406 a_9634_17478# a_9974_17626# 0.24088f
C3407 a_10378_27170# sar9b_0.net34 0.01673f
C3408 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[7] 0.02109f
C3409 a_8386_22806# a_8591_22855# 0.09983f
C3410 a_8202_23174# a_9162_23174# 0.03529f
C3411 a_5484_23444# a_5823_23477# 0.07649f
C3412 a_6132_23451# a_5682_23444# 0.03529f
C3413 a_5506_17478# a_5846_17626# 0.24088f
C3414 a_2892_23070# sar9b_0.clk_div_0.COUNT\[1\] 0.01011f
C3415 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C3416 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] 1.20704f
C3417 a_8334_18353# sar9b_0.net48 0.04696f
C3418 a_6534_17799# sar9b_0.net56 0.02731f
C3419 a_10402_27758# single_9b_cdac_0.SW[5] 0.013f
C3420 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_41357_15501# 0.01076f
C3421 sar9b_0.net44 a_5506_26802# 0.08971f
C3422 VDPWR sar9b_0.net63 1.51034f
C3423 a_10548_19053# sar9b_0.net38 0.01246f
C3424 VDPWR a_2931_28566# 0.47184f
C3425 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.01492f
C3426 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.06503f
C3427 a_10470_21795# sar9b_0.net9 0.03298f
C3428 sar9b_0.net40 sar9b_0.clk_div_0.COUNT\[1\] 0.0227f
C3429 a_4947_20140# sar9b_0.clknet_1_0__leaf_CLK 0.21937f
C3430 sar9b_0.net63 sar9b_0._14_ 0.30459f
C3431 single_9b_cdac_1.CF[4] clk 0.14003f
C3432 single_9b_cdac_1.CF[1] clk 0.08196f
C3433 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C3434 sar9b_0.net36 a_10482_25831# 0.02816f
C3435 VDPWR sar9b_0._05_ 0.50167f
C3436 a_8303_23853# a_7914_23470# 0.06034f
C3437 sar9b_0.net3 a_2451_27234# 0.15641f
C3438 sar9b_0.net56 a_8057_18463# 0.01557f
C3439 sar9b_0.net2 sar9b_0.net53 0.39622f
C3440 a_8334_17021# sar9b_0.net46 0.19846f
C3441 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.12358f
C3442 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.69086f
C3443 a_5812_21028# sar9b_0._17_ 0.04354f
C3444 sar9b_0.net48 a_9450_17846# 0.17495f
C3445 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.84427f
C3446 VDPWR a_12870_26263# 0.2717f
C3447 sar9b_0.net58 uo_out[6] 0.11715f
C3448 a_5748_24381# a_5962_24151# 0.05022f
C3449 sar9b_0.net23 sar9b_0.net45 0.02681f
C3450 sar9b_0.net48 single_9b_cdac_1.SW[2] 0.7306f
C3451 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.24779f
C3452 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[0] 0.22459f
C3453 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.01514f
C3454 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 3.10626f
C3455 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[0] 0.23282f
C3456 a_8334_18353# sar9b_0.net46 0.22365f
C3457 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 2.81139f
C3458 single_9b_cdac_1.CF[7] sar9b_0.net27 0.14896f
C3459 sar9b_0.net52 a_9942_24806# 0.20968f
C3460 a_6834_20780# sar9b_0.net40 0.01162f
C3461 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] 0.17948f
C3462 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[5] 0.02016f
C3463 a_6252_20780# sar9b_0._11_ 0.27844f
C3464 sar9b_0.net35 a_6562_25094# 0.02907f
C3465 a_11658_18142# sar9b_0.net39 0.02313f
C3466 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[0] 0.37948f
C3467 single_9b_cdac_0.SW[6] a_34814_26990# 0.18991f
C3468 sar9b_0.net9 sar9b_0.net73 0.02088f
C3469 a_3713_22522# sar9b_0._12_ 0.04441f
C3470 VDPWR sar9b_0.clknet_1_1__leaf_CLK 3.19348f
C3471 a_10607_25185# a_10742_25087# 0.35559f
C3472 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[4] 0.0313f
C3473 a_5439_24563# a_5748_24381# 0.07766f
C3474 sar9b_0.clknet_0_CLK a_4332_23043# 1.32864f
C3475 sar9b_0.net30 single_9b_cdac_0.SW[4] 0.11168f
C3476 ui_in[0] th_dif_sw_0.VCN 0.22659f
C3477 single_9b_cdac_1.CF[8] clk 0.12991f
C3478 sar9b_0.net40 a_10803_19474# 0.07638f
C3479 sar9b_0._14_ sar9b_0.clknet_1_1__leaf_CLK 0.02074f
C3480 sar9b_0.net49 sar9b_0.net37 0.07403f
C3481 single_9b_cdac_1.SW[1] a_58824_17740# 0.18991f
C3482 a_9162_23174# sar9b_0.net37 0.02849f
C3483 a_11382_23474# a_11658_23470# 0.1263f
C3484 sar9b_0.net10 sar9b_0.net73 0.07697f
C3485 sar9b_0.net61 sar9b_0.net73 0.22051f
C3486 sar9b_0.net51 a_7443_21496# 0.28357f
C3487 a_10402_21098# sar9b_0.net73 0.01426f
C3488 a_10482_25831# a_10937_25582# 0.3578f
C3489 a_10623_25895# a_10932_25713# 0.07766f
C3490 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] 1.15122f
C3491 single_9b_cdac_1.CF[1] a_13011_20806# 0.06696f
C3492 a_3370_27769# a_3438_27677# 0.35559f
C3493 sar9b_0.net53 a_10758_24459# 0.16837f
C3494 sar9b_0._01_ sar9b_0._10_ 0.03463f
C3495 a_10470_21795# a_9442_21474# 0.07826f
C3496 a_3369_24181# a_3262_24141# 0.14439f
C3497 sar9b_0.net41 sar9b_0.net54 0.04048f
C3498 a_5711_17527# a_5046_17906# 0.19065f
C3499 a_5846_17626# a_5322_17846# 0.04522f
C3500 sar9b_0.clknet_0_CLK sar9b_0.net72 0.06286f
C3501 a_9258_21842# a_8982_21902# 0.1263f
C3502 w_17430_1606# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.3776f
C3503 sar9b_0.net23 a_9870_27060# 0.01769f
C3504 sar9b_0.net46 single_9b_cdac_1.SW[2] 0.02228f
C3505 sar9b_0.net49 a_10098_19171# 0.02393f
C3506 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[7] 0.06019f
C3507 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C3508 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.CF[0] 0.12358f
C3509 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3510 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[0] 0.584f
C3511 th_dif_sw_0.th_sw_1.CK a_10482_3438# 0.1221f
C3512 VDPWR sar9b_0.net55 0.724f
C3513 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[2] 15.0435f
C3514 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[0] 0.27554f
C3515 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.07517f
C3516 sar9b_0.net43 a_6030_24396# 0.04681f
C3517 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] 1.50844f
C3518 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[0] 0.22444f
C3519 sar9b_0.clk_div_0.COUNT\[1\] a_3372_25734# 0.12822f
C3520 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 2.71729f
C3521 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] 0.17948f
C3522 a_5739_22488# sar9b_0.net60 0.01946f
C3523 a_7188_22119# a_7402_22441# 0.04522f
C3524 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.42509f
C3525 sar9b_0.net52 a_12047_26517# 0.22373f
C3526 a_6975_20813# sar9b_0.net10 0.03184f
C3527 sar9b_0.net27 a_12435_20806# 0.01148f
C3528 a_7470_22349# sar9b_0.net39 0.03069f
C3529 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C3530 sar9b_0.net41 a_10035_19474# 0.02751f
C3531 VDPWR a_11382_19478# 0.30104f
C3532 VDPWR a_10548_19053# 0.83308f
C3533 VDPWR a_4755_22138# 0.4525f
C3534 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.19266f
C3535 a_12182_18427# sar9b_0.net50 0.14036f
C3536 VDPWR a_9839_17527# 0.25186f
C3537 sar9b_0.net61 sar9b_0.net48 0.8171f
C3538 a_12182_18427# a_12618_18142# 0.16939f
C3539 th_dif_sw_0.CK single_9b_cdac_1.SW[1] 0.06557f
C3540 a_5443_19074# a_5811_19178# 0.08134f
C3541 sar9b_0.net7 sar9b_0.net73 1.54797f
C3542 single_9b_cdac_1.cdac_sw_9b_0.S[4] ua[0] 1.94611f
C3543 a_7890_26108# a_7692_26108# 0.06623f
C3544 VDPWR a_29134_26999# 1.81495f
C3545 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.26942f
C3546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C3547 sar9b_0.net40 a_6378_24802# 0.0119f
C3548 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C3549 sar9b_0.net50 single_9b_cdac_1.SW[8] 0.1731f
C3550 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.15428f
C3551 a_6534_27123# a_6880_26815# 0.07649f
C3552 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[8] 0.06897f
C3553 sar9b_0.net63 a_5682_23444# 0.04284f
C3554 VDPWR sar9b_0.net38 3.13581f
C3555 single_9b_cdac_1.CF[3] clk 0.109f
C3556 sar9b_0.net28 clk 0.52609f
C3557 single_9b_cdac_0.SW[6] uo_out[3] 0.30173f
C3558 sar9b_0._11_ sar9b_0.net65 0.09114f
C3559 a_13011_27234# a_13067_27662# 0.01136f
C3560 sar9b_0.net43 sar9b_0.net23 0.30643f
C3561 sar9b_0.net41 sar9b_0.net74 0.02251f
C3562 sar9b_0.net60 sar9b_0._10_ 0.38542f
C3563 a_7498_21109# sar9b_0.net10 0.03668f
C3564 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.0303f
C3565 sar9b_0.net36 a_10506_24506# 0.0206f
C3566 sar9b_0.net36 sar9b_0.net21 0.02863f
C3567 sar9b_0.net52 a_11430_24931# 0.16913f
C3568 uo_out[0] ui_in[0] 0.0743f
C3569 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[7] 2.07035f
C3570 a_10218_21842# sar9b_0.net38 0.02659f
C3571 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.19266f
C3572 sar9b_0.net1 sar9b_0.net38 0.03587f
C3573 a_8438_23755# a_8874_23470# 0.16939f
C3574 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.10626f
C3575 a_5439_24563# sar9b_0.net39 0.01949f
C3576 sar9b_0.net13 a_10742_25087# 0.02523f
C3577 a_10218_27466# a_11430_27595# 0.07766f
C3578 a_8166_27595# sar9b_0.net36 0.06865f
C3579 sar9b_0.net36 sar9b_0.net27 0.4102f
C3580 sar9b_0.net41 a_9942_20810# 0.01321f
C3581 a_8202_23174# sar9b_0.net11 0.26859f
C3582 sar9b_0.net33 sar9b_0.net42 0.01652f
C3583 a_48343_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.23864f
C3584 sar9b_0.net61 sar9b_0.net46 0.5339f
C3585 a_5010_28495# sar9b_0.net58 0.2625f
C3586 a_8595_17910# sar9b_0.net37 0.04816f
C3587 single_9b_cdac_1.CF[3] single_9b_cdac_1.SW[0] 0.2246f
C3588 sar9b_0.net61 sar9b_0.net50 0.03896f
C3589 sar9b_0.net59 sar9b_0.net20 0.0752f
C3590 single_9b_cdac_1.SW[3] sar9b_0.net61 0.02878f
C3591 a_8052_18123# sar9b_0.net5 0.06414f
C3592 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[7] 16.1938f
C3593 th_dif_sw_0.CKB dw_17224_1400# 0.01749f
C3594 a_11339_27039# sar9b_0.net45 0.10933f
C3595 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] 3.10218f
C3596 sar9b_0.net7 sar9b_0.net48 0.22803f
C3597 sar9b_0.net18 a_2847_27473# 0.03049f
C3598 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C3599 sar9b_0.net26 sar9b_0.net39 0.06931f
C3600 sar9b_0.net26 single_9b_cdac_1.CF[7] 0.18995f
C3601 tdc_0.OUTN a_16555_12412# 0.01287f
C3602 th_dif_sw_0.th_sw_1.CK a_21368_4076# 0.0478f
C3603 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C3604 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[7] 0.0313f
C3605 VDPWR a_9165_24988# 0.44778f
C3606 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.CF[2] 0.03547f
C3607 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.36334f
C3608 single_9b_cdac_1.CF[3] a_13011_20806# 0.35649f
C3609 sar9b_0.net52 sar9b_0.net54 0.82593f
C3610 a_10649_17131# single_9b_cdac_1.SW[0] 0.02173f
C3611 sar9b_0.net49 a_10182_20463# 0.2021f
C3612 a_3713_22522# a_4011_22488# 0.02614f
C3613 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A a_49926_15495# 0.01076f
C3614 sar9b_0.net35 a_6922_23534# 0.02301f
C3615 VDPWR a_9126_23599# 0.28311f
C3616 a_11658_23470# sar9b_0.net53 0.18176f
C3617 VDPWR sar9b_0.net6 2.96308f
C3618 a_4934_22432# a_5739_22488# 0.29207f
C3619 sar9b_0._18_ sar9b_0.net60 0.06258f
C3620 sar9b_0.net49 sar9b_0.net57 0.18506f
C3621 a_7306_19777# sar9b_0.net35 0.01601f
C3622 sar9b_0.net23 a_8340_26115# 0.02021f
C3623 sar9b_0._01_ sar9b_0.net60 0.26299f
C3624 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[2] 16.8504f
C3625 sar9b_0.net4 a_6030_24396# 0.01963f
C3626 sar9b_0.net41 sar9b_0.net8 0.02515f
C3627 sar9b_0.net1 sar9b_0.net6 0.06186f
C3628 sar9b_0.net7 sar9b_0.net50 0.20371f
C3629 sar9b_0.net59 sar9b_0.net44 0.32798f
C3630 a_8842_16874# a_8057_17131# 0.26257f
C3631 sar9b_0.net7 single_9b_cdac_1.SW[3] 0.03478f
C3632 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[3] 14.7603f
C3633 sar9b_0.net44 a_3156_27447# 0.236f
C3634 a_4125_25958# sar9b_0._03_ 0.1014f
C3635 sar9b_0.net8 a_11430_20935# 0.04729f
C3636 a_5938_22378# a_6540_22112# 0.01219f
C3637 VDPWR a_8970_20510# 0.9047f
C3638 sar9b_0.net11 sar9b_0.net37 0.02799f
C3639 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.6919f
C3640 a_5938_22378# sar9b_0.net39 0.0251f
C3641 a_10239_19235# a_9900_19047# 0.07649f
C3642 sar9b_0.net26 a_12435_20806# 0.0353f
C3643 sar9b_0.net46 a_6579_18832# 0.31908f
C3644 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 3.10218f
C3645 sar9b_0.net30 a_12064_22819# 0.2744f
C3646 VDPWR sar9b_0._14_ 0.55641f
C3647 a_43540_16877# single_9b_cdac_1.SW[4] 0.28324f
C3648 sar9b_0.net68 a_4044_24776# 0.041f
C3649 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.10499f
C3650 sar9b_0.net42 a_11178_24802# 0.01588f
C3651 a_11436_17742# sar9b_0.net61 0.18223f
C3652 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 3.27833f
C3653 a_6137_23791# sar9b_0.net11 0.11829f
C3654 VDPWR a_10218_21842# 0.36269f
C3655 sar9b_0.net52 sar9b_0.net74 0.7241f
C3656 VDPWR sar9b_0.net1 1.19391f
C3657 ua[3] dw_17224_1400# 1.4136f
C3658 a_4922_20857# sar9b_0._11_ 0.07006f
C3659 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C3660 a_3180_19448# a_3795_19512# 0.02106f
C3661 sar9b_0.net44 a_4330_27170# 0.07062f
C3662 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C3663 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0._03_ 0.03884f
C3664 tdc_0.OUTP a_16555_12124# 0.01017f
C3665 sar9b_0.net58 sar9b_0.net45 0.10292f
C3666 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[2] 4.15039f
C3667 single_9b_cdac_0.SW[2] sar9b_0.net27 0.06976f
C3668 a_11146_25483# sar9b_0.net74 0.0492f
C3669 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[5] 0.02056f
C3670 a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] 0.11932f
C3671 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.95338f
C3672 a_3946_27530# a_3438_27677# 0.19065f
C3673 a_8334_17021# sar9b_0.net27 0.06035f
C3674 a_11915_27039# sar9b_0.net30 0.22412f
C3675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 a_49221_26990# 0.14695f
C3676 sar9b_0.net31 sar9b_0.net52 0.77905f
C3677 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C3678 a_10254_2858# w_12795_1601# 0.14391f
C3679 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.22875f
C3680 a_8345_26455# sar9b_0.cyclic_flag_0.FINAL 0.12177f
C3681 a_7097_19795# sar9b_0.net40 0.16334f
C3682 a_8438_18958# sar9b_0.net48 0.14544f
C3683 sar9b_0.net24 a_9138_27163# 0.03746f
C3684 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3685 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.26942f
C3686 sar9b_0.net45 a_9323_27662# 0.10552f
C3687 sar9b_0.net53 sar9b_0.net39 0.01835f
C3688 single_9b_cdac_1.cdac_sw_9b_0.S[5] th_dif_sw_0.VCP 6.58553f
C3689 single_9b_cdac_0.cdac_sw_9b_0.S[8] ua[0] 16.2797f
C3690 a_7097_19795# sar9b_0.net51 0.02536f
C3691 sar9b_0.net26 sar9b_0.net36 0.0273f
C3692 sar9b_0.net70 a_3027_22138# 0.03062f
C3693 sar9b_0.net27 single_9b_cdac_1.CF[0] 0.02972f
C3694 sar9b_0.net64 sar9b_0.net4 0.04411f
C3695 a_3014_24136# a_2508_23444# 0.01366f
C3696 a_7638_19238# a_8303_18859# 0.19065f
C3697 single_9b_cdac_1.CF[5] clk 0.48018f
C3698 single_9b_cdac_0.SW[4] clk 0.1627f
C3699 sar9b_0.net60 a_5753_24250# 0.01748f
C3700 a_8098_23762# sar9b_0.net37 0.01305f
C3701 a_8883_27466# single_9b_cdac_0.SW[8] 0.0266f
C3702 sar9b_0.net19 uo_out[7] 0.03323f
C3703 VDPWR a_4083_28566# 0.47299f
C3704 a_10926_17021# a_10644_16791# 0.05462f
C3705 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[8] 0.80778f
C3706 a_4934_22432# sar9b_0._18_ 0.02193f
C3707 VDPWR a_2508_27440# 0.21708f
C3708 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 1.71649f
C3709 sar9b_0.net32 a_12531_28566# 0.02777f
C3710 sar9b_0.net54 a_6102_24806# 0.21862f
C3711 a_11842_23762# sar9b_0.net11 0.05371f
C3712 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.11216f
C3713 sar9b_0.net32 a_12870_23599# 0.0306f
C3714 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.19266f
C3715 sar9b_0.net59 a_4749_27652# 0.27144f
C3716 a_3695_23038# a_3725_23194# 0.0101f
C3717 a_10758_24459# a_11104_24151# 0.07649f
C3718 a_5289_22527# sar9b_0._12_ 0.0393f
C3719 a_10218_24802# sar9b_0.net57 0.2148f
C3720 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[0] 0.22459f
C3721 sar9b_0.net27 single_9b_cdac_1.SW[2] 0.12181f
C3722 a_10895_22855# sar9b_0.net53 0.2218f
C3723 a_3819_24136# a_2835_24136# 0.08669f
C3724 sar9b_0.net34 a_9593_26914# 0.02203f
C3725 a_10690_22806# a_10895_22855# 0.09983f
C3726 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.84061f
C3727 a_10506_23174# a_11466_23174# 0.03471f
C3728 a_12870_26263# a_13216_26469# 0.07649f
C3729 a_12182_26419# a_12047_26517# 0.35559f
C3730 sar9b_0.net33 a_11842_26426# 0.13675f
C3731 VDPWR sar9b_0.net29 1.26137f
C3732 a_9323_28371# uo_out[3] 0.04123f
C3733 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.6919f
C3734 a_7914_27466# a_8512_27801# 0.06623f
C3735 a_6636_20780# a_6834_20780# 0.06623f
C3736 sar9b_0.net60 uio_out[0] 0.09917f
C3737 a_3206_22432# a_3561_22527# 0.18757f
C3738 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.02618f
C3739 a_11466_23174# sar9b_0.net31 0.017f
C3740 a_9414_23127# sar9b_0.net54 0.18588f
C3741 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.01175f
C3742 a_3206_22432# sar9b_0.clknet_0_CLK 0.01173f
C3743 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C3744 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 2.82172f
C3745 a_8052_16791# sar9b_0.net6 0.02602f
C3746 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.11216f
C3747 sar9b_0.net35 sar9b_0._17_ 0.03063f
C3748 sar9b_0.net60 a_5506_26802# 0.02734f
C3749 tdc_0.OUTP single_9b_cdac_1.SW[2] 0.36499f
C3750 a_6954_27466# sar9b_0.net44 0.22029f
C3751 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[7] 0.06503f
C3752 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[6] 0.31534f
C3753 sar9b_0.net56 a_9359_20191# 0.01326f
C3754 a_3090_27163# sar9b_0.net19 0.05411f
C3755 VDPWR a_9472_18823# 0.21089f
C3756 a_11658_18142# a_12182_18427# 0.05022f
C3757 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._00_ 0.1706f
C3758 VDPWR a_5846_17626# 0.19864f
C3759 VDPWR a_5682_23444# 0.35048f
C3760 sar9b_0.net57 sar9b_0.net11 0.86992f
C3761 a_7347_24160# sar9b_0.net62 0.09083f
C3762 a_8386_22806# clk 0.03185f
C3763 sar9b_0.net27 single_9b_cdac_1.SW[8] 0.0444f
C3764 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.12358f
C3765 tdc_0.phase_detector_0.pd_out_0.B a_15052_11404# 0.18949f
C3766 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# 1.26208f
C3767 dw_12589_1395# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.26214f
C3768 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.42014f
C3769 sar9b_0._03_ sar9b_0.clknet_1_1__leaf_CLK 0.23577f
C3770 a_4934_22432# sar9b_0.net60 0.03501f
C3771 a_9472_18823# sar9b_0.net1 0.01552f
C3772 VDPWR a_9270_24566# 0.29709f
C3773 a_3014_24136# sar9b_0.net70 0.26822f
C3774 sar9b_0.net43 a_9323_27662# 0.04771f
C3775 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.17533f
C3776 a_11859_20574# sar9b_0.net51 0.08706f
C3777 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR 0.62555f
C3778 VDPWR a_11382_26138# 0.29139f
C3779 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.02638f
C3780 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.01152f
C3781 single_9b_cdac_1.CF[1] a_13011_20574# 0.01474f
C3782 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[7] 0.06019f
C3783 sar9b_0.net52 sar9b_0.net34 0.06265f
C3784 sar9b_0._09_ sar9b_0.net57 0.46567f
C3785 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[0] 0.7639f
C3786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3787 a_9996_16784# a_10194_16784# 0.06623f
C3788 single_9b_cdac_1.SW[5] th_dif_sw_0.VCN 0.09453f
C3789 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_50962_15501# 0.01076f
C3790 sar9b_0.net9 sar9b_0.net27 0.03863f
C3791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.07579f
C3792 VDPWR a_8052_16791# 0.86212f
C3793 sar9b_0.net36 sar9b_0.net53 0.06691f
C3794 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[7] 1.10355f
C3795 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.95338f
C3796 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[3] 14.7603f
C3797 a_10690_22806# sar9b_0.net36 0.01892f
C3798 a_6562_25094# a_6902_25087# 0.24088f
C3799 VDPWR a_11658_22138# 0.83163f
C3800 sar9b_0.net43 sar9b_0.net37 0.04982f
C3801 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.28523f
C3802 sar9b_0.net10 sar9b_0.net27 0.03534f
C3803 sar9b_0.net61 sar9b_0.net27 0.12915f
C3804 sar9b_0.net58 a_3754_26815# 0.14463f
C3805 sar9b_0.net48 a_5535_18149# 0.17429f
C3806 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.01175f
C3807 th_dif_sw_0.CKB tdc_0.OUTN 2.99096f
C3808 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.62443f
C3809 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38733f
C3810 sar9b_0.net58 a_3540_27045# 0.17959f
C3811 a_6307_27584# a_5460_28377# 0.01439f
C3812 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36044f
C3813 a_11658_18142# sar9b_0.net61 0.01086f
C3814 sar9b_0.net13 sar9b_0.net37 0.03945f
C3815 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.75853f
C3816 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C3817 a_2739_20140# a_3425_20244# 0.27693f
C3818 a_2918_20140# a_3166_20145# 0.05308f
C3819 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.SW[7] 0.17509f
C3820 a_5441_22522# a_5739_22488# 0.02614f
C3821 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C3822 sar9b_0.net38 a_8691_28566# 0.0583f
C3823 a_9802_26815# sar9b_0.net36 0.06626f
C3824 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] 0.17948f
C3825 a_10218_24802# a_11178_24802# 0.03432f
C3826 single_9b_cdac_1.SW[2] single_9b_cdac_1.SW[7] 0.2192f
C3827 VDPWR single_9b_cdac_0.SW[3] 2.47465f
C3828 sar9b_0.net56 a_4771_18260# 0.23559f
C3829 th_dif_sw_0.th_sw_1.CKB a_10482_3438# 0.0331f
C3830 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 2.82172f
C3831 a_11658_23470# a_12047_23853# 0.06034f
C3832 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C3833 a_8098_23762# sar9b_0.net57 0.06831f
C3834 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.02624f
C3835 tdc_0.OUTP sar9b_0.net61 0.10662f
C3836 sar9b_0.net43 a_9730_24138# 0.06642f
C3837 a_10858_17113# sar9b_0.net6 0.03245f
C3838 sar9b_0.net40 sar9b_0.net28 0.10374f
C3839 sar9b_0.net59 single_9b_cdac_0.SW[7] 0.07361f
C3840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C3841 VDPWR a_6678_27470# 0.2784f
C3842 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36301f
C3843 a_8554_26437# a_8622_26345# 0.35559f
C3844 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38715f
C3845 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[3] 12.6046f
C3846 a_8842_18206# sar9b_0.net73 0.04312f
C3847 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A 0.74663f
C3848 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.05472f
C3849 sar9b_0.net7 sar9b_0.net27 0.06127f
C3850 sar9b_0._07_ sar9b_0._10_ 0.0757f
C3851 a_4922_20857# a_5581_20992# 0.01403f
C3852 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.69086f
C3853 a_5628_19768# sar9b_0.net47 0.014f
C3854 sar9b_0.net58 a_4125_25958# 0.03759f
C3855 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.62443f
C3856 sar9b_0.net10 a_7470_22349# 0.07606f
C3857 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[7] 6.82494f
C3858 a_8874_19178# sar9b_0.net37 0.03852f
C3859 sar9b_0.net7 a_11658_18142# 0.21927f
C3860 a_5465_28246# a_5742_28392# 0.09983f
C3861 sar9b_0.net32 a_12435_24802# 0.03774f
C3862 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.08121f
C3863 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.05472f
C3864 sar9b_0.net23 sar9b_0.net38 0.02577f
C3865 sar9b_0.net35 clk 0.03859f
C3866 a_8340_26115# sar9b_0.net37 0.02741f
C3867 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[7] 3.98346f
C3868 a_12064_22819# clk 0.01615f
C3869 VDPWR a_10858_17113# 0.19951f
C3870 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.27795f
C3871 sar9b_0._08_ sar9b_0._10_ 0.25501f
C3872 a_10548_19053# a_10830_19068# 0.06034f
C3873 a_4755_22138# sar9b_0.net64 0.07292f
C3874 sar9b_0.net2 clk 0.03287f
C3875 sar9b_0.net58 sar9b_0._15_ 0.04426f
C3876 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.05472f
C3877 a_5846_26950# a_5322_27170# 0.04522f
C3878 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C3879 a_8591_22855# a_8726_22954# 0.35559f
C3880 single_9b_cdac_0.SW[1] a_13011_27234# 0.35197f
C3881 sar9b_0.net40 a_6282_27170# 0.0332f
C3882 a_6132_23451# a_6137_23791# 0.43491f
C3883 VDPWR a_4072_19474# 0.11411f
C3884 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.0303f
C3885 VDPWR sar9b_0.net71 0.30617f
C3886 a_8842_18206# sar9b_0.net48 0.06788f
C3887 sar9b_0.net58 sar9b_0.clk_div_0.COUNT\[2\] 0.06301f
C3888 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C3889 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C3890 a_11430_27595# single_9b_cdac_0.SW[5] 0.03357f
C3891 sar9b_0.net44 a_5846_26950# 0.05309f
C3892 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 3.27795f
C3893 a_9323_28371# single_9b_cdac_0.SW[8] 0.0233f
C3894 sar9b_0.net26 single_9b_cdac_1.SW[8] 0.03854f
C3895 VDPWR a_7193_22459# 0.22562f
C3896 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.0303f
C3897 sar9b_0._10_ sar9b_0.clknet_1_0__leaf_CLK 0.20402f
C3898 sar9b_0.net47 sar9b_0.net4 0.03459f
C3899 sar9b_0.net56 sar9b_0.net35 0.5676f
C3900 a_6744_23238# sar9b_0._17_ 0.03116f
C3901 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.37833f
C3902 a_7092_19455# a_6783_19481# 0.07766f
C3903 VDPWR a_12684_20379# 0.21989f
C3904 a_7539_28566# uo_out[5] 0.40403f
C3905 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.42509f
C3906 a_8019_17910# sar9b_0.net46 0.05518f
C3907 sar9b_0._06_ clk 0.01579f
C3908 sar9b_0._18_ sar9b_0._07_ 0.02201f
C3909 sar9b_0.net29 single_9b_cdac_0.SW[3] 0.06969f
C3910 sar9b_0.net21 a_7539_28566# 0.20381f
C3911 a_3369_24181# sar9b_0.clknet_1_1__leaf_CLK 0.06961f
C3912 a_8842_16874# sar9b_0.net46 0.19416f
C3913 a_9546_24506# sar9b_0.net12 0.21444f
C3914 a_11030_22954# sar9b_0.net2 0.01198f
C3915 sar9b_0.net9 sar9b_0.net26 0.02943f
C3916 a_6861_22828# sar9b_0.clk_div_0.COUNT\[2\] 0.04796f
C3917 tdc_0.OUTN single_9b_cdac_1.SW[0] 0.44367f
C3918 VDPWR a_6030_24396# 0.2481f
C3919 VDPWR a_8691_28566# 0.50803f
C3920 th_dif_sw_0.th_sw_1.CKB a_21368_4076# 0.06647f
C3921 sar9b_0._11_ sar9b_0._17_ 0.45057f
C3922 sar9b_0._01_ sar9b_0._07_ 0.14158f
C3923 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[0] 1.12533f
C3924 single_9b_cdac_1.cdac_sw_9b_0.S[6] ua[0] 1.67132f
C3925 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.94957f
C3926 VDPWR a_13216_26469# 0.21606f
C3927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.01003f
C3928 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] 0.12898f
C3929 sar9b_0.net26 sar9b_0.net61 0.01357f
C3930 sar9b_0.net26 sar9b_0.net10 0.0815f
C3931 sar9b_0._08_ sar9b_0._18_ 0.02837f
C3932 sar9b_0.net43 sar9b_0.net57 0.05729f
C3933 a_8052_18123# a_7743_18149# 0.07766f
C3934 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.363f
C3935 a_8842_18206# sar9b_0.net46 0.221f
C3936 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 2.82223f
C3937 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 ua[0] 0.14027f
C3938 sar9b_0.net27 a_13011_27234# 0.22439f
C3939 a_7404_16784# a_7602_16784# 0.06623f
C3940 sar9b_0._08_ sar9b_0._01_ 0.05213f
C3941 sar9b_0.net50 a_12618_19474# 0.26154f
C3942 a_6137_23791# sar9b_0.net4 0.01198f
C3943 sar9b_0.net35 a_7590_24931# 0.01235f
C3944 sar9b_0.net13 sar9b_0.net57 0.17396f
C3945 sar9b_0.net2 a_10803_18142# 0.0218f
C3946 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.10499f
C3947 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.SW[4] 0.01837f
C3948 a_8940_27039# a_9138_27163# 0.06623f
C3949 a_4210_22378# sar9b_0._12_ 0.04138f
C3950 sar9b_0.net41 sar9b_0.net73 0.0295f
C3951 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02618f
C3952 a_5151_28559# uo_out[7] 0.02535f
C3953 VDPWR sar9b_0._03_ 0.5857f
C3954 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.31534f
C3955 a_9942_27470# sar9b_0.net45 0.08179f
C3956 a_2603_17006# th_dif_sw_0.CKB 0.35268f
C3957 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[6] 0.26707f
C3958 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.03729f
C3959 sar9b_0.net63 sar9b_0.net58 0.25917f
C3960 a_10932_25713# a_10937_25582# 0.44532f
C3961 sar9b_0.net59 sar9b_0.net60 0.37207f
C3962 a_7936_25137# sar9b_0.net54 0.03507f
C3963 a_11722_25838# a_10932_25713# 0.1263f
C3964 a_10230_23234# sar9b_0.net11 0.04733f
C3965 sar9b_0.net7 a_9258_21842# 0.01005f
C3966 sar9b_0.net23 VDPWR 1.79675f
C3967 a_9258_21842# a_9442_21474# 0.44098f
C3968 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.42014f
C3969 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.A 0.02054f
C3970 VDPWR a_10742_25087# 0.19934f
C3971 a_8438_23755# sar9b_0.net54 0.02573f
C3972 uio_in[7] uio_in[6] 0.03102f
C3973 a_7638_19238# sar9b_0.net51 0.03553f
C3974 sar9b_0.net32 single_9b_cdac_1.CF[5] 0.011f
C3975 sar9b_0.net32 single_9b_cdac_0.SW[4] 0.02994f
C3976 sar9b_0._07_ a_3795_19512# 0.11659f
C3977 VDPWR a_5711_26851# 0.26739f
C3978 sar9b_0.net63 a_6861_22828# 0.16938f
C3979 sar9b_0.net7 sar9b_0.net26 0.07618f
C3980 a_7566_21017# sar9b_0.net51 0.02936f
C3981 sar9b_0._07_ sar9b_0.net60 0.56326f
C3982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.05472f
C3983 a_5441_22522# sar9b_0.net60 0.01343f
C3984 single_9b_cdac_1.CF[6] clk 0.13098f
C3985 a_7914_23470# clk 0.01168f
C3986 a_3206_22432# a_3027_22138# 0.54361f
C3987 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.1507f
C3988 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.84423f
C3989 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[6] 0.06019f
C3990 a_7978_22202# sar9b_0.net39 0.04787f
C3991 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C3992 sar9b_0.net41 sar9b_0.net48 0.33991f
C3993 a_59529_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.01076f
C3994 a_6132_23451# sar9b_0.net57 0.24363f
C3995 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.CF[5] 0.01608f
C3996 VDPWR a_10830_19068# 0.26619f
C3997 VDPWR sar9b_0.net64 0.46487f
C3998 a_3206_22432# sar9b_0.net65 0.02448f
C3999 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_1.CF[3] 0.01346f
C4000 a_12182_19759# sar9b_0.net50 0.14123f
C4001 sar9b_0._08_ sar9b_0.net60 0.18449f
C4002 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.81423f
C4003 sar9b_0.net40 a_13216_18477# 0.01664f
C4004 a_5126_20140# sar9b_0.net57 0.01075f
C4005 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.12431f
C4006 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62538f
C4007 a_12870_18271# a_13216_18477# 0.07649f
C4008 a_12182_18427# a_12047_18525# 0.35559f
C4009 sar9b_0.net58 sar9b_0.clknet_1_1__leaf_CLK 0.05967f
C4010 a_5931_20140# a_6130_20239# 0.29821f
C4011 a_5811_19178# a_6252_19074# 0.0184f
C4012 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP a_43540_26999# 0.04592f
C4013 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.11216f
C4014 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.22513f
C4015 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.06503f
C4016 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 3.27833f
C4017 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C4018 a_8031_26141# a_8340_26115# 0.07766f
C4019 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.31534f
C4020 sar9b_0._17_ sar9b_0.net39 0.02501f
C4021 a_6744_23238# clk 0.01136f
C4022 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.76578f
C4023 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.69086f
C4024 a_10859_26330# single_9b_cdac_0.SW[7] 0.37246f
C4025 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[0] 0.22459f
C4026 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.7611f
C4027 th_dif_sw_0.VCN ua[0] 0.86465f
C4028 sar9b_0.net63 a_6137_23791# 0.04828f
C4029 sar9b_0.net9 sar9b_0.net53 0.14548f
C4030 a_3994_19474# a_4072_19474# 0.01029f
C4031 sar9b_0.net60 a_5823_23477# 0.03124f
C4032 sar9b_0.net9 a_10690_22806# 0.03973f
C4033 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.71729f
C4034 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C4035 a_9359_20191# sar9b_0.net51 0.07207f
C4036 sar9b_0.net60 sar9b_0.clknet_1_0__leaf_CLK 0.04105f
C4037 VDPWR ui_in[0] 2.1737f
C4038 sar9b_0.net59 uio_out[0] 0.11978f
C4039 sar9b_0.net56 a_10218_20806# 0.21365f
C4040 a_10227_23490# sar9b_0.net54 0.18976f
C4041 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.95338f
C4042 sar9b_0.net10 sar9b_0.net53 0.31214f
C4043 sar9b_0._12_ a_5523_21528# 0.17627f
C4044 single_9b_cdac_1.CF[2] th_dif_sw_0.VCN 0.09453f
C4045 a_9126_23599# a_9472_23805# 0.07649f
C4046 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.84061f
C4047 sar9b_0.net13 a_11178_24802# 0.0805f
C4048 a_10402_27758# a_10742_27751# 0.24088f
C4049 a_8512_27801# sar9b_0.net36 0.04404f
C4050 sar9b_0.net41 single_9b_cdac_1.SW[3] 0.03054f
C4051 a_21684_3438# dw_17224_1400# 0.05479f
C4052 sar9b_0.net43 a_9942_27470# 0.17078f
C4053 a_5235_27466# sar9b_0.net36 0.073f
C4054 a_41357_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C4055 sar9b_0.net57 sar9b_0.net4 0.32464f
C4056 sar9b_0.net32 sar9b_0.net24 0.2487f
C4057 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.33229f
C4058 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.11907f
C4059 VDPWR a_17125_9355# 0.01057f
C4060 a_7338_24802# a_6378_24802# 0.03432f
C4061 a_33936_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.23864f
C4062 sar9b_0.net47 sar9b_0.net55 0.03364f
C4063 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 ua[0] 0.12069f
C4064 a_11722_25838# sar9b_0.net30 0.01802f
C4065 sar9b_0.net41 a_9154_20142# 0.02308f
C4066 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4067 a_11915_28371# uo_out[1] 0.04028f
C4068 a_16331_9671# th_dif_sw_0.VCP 0.10881f
C4069 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS w_12795_1601# 0.38264f
C4070 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4071 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.01198f
C4072 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[2\] 0.01818f
C4073 a_13011_24802# sar9b_0.net27 0.04101f
C4074 VDPWR a_7289_21127# 0.22771f
C4075 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C4076 single_9b_cdac_1.SW[4] sar9b_0.net27 0.46877f
C4077 a_4210_22378# a_4011_22488# 0.29821f
C4078 a_10926_17021# single_9b_cdac_1.SW[1] 0.02544f
C4079 a_7404_17715# sar9b_0.net35 0.03641f
C4080 VDPWR a_9472_23805# 0.20106f
C4081 sar9b_0.net58 sar9b_0.net38 0.14084f
C4082 a_8266_17113# a_8334_17021# 0.35559f
C4083 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[3] 0.06971f
C4084 a_4934_22432# sar9b_0._07_ 0.01085f
C4085 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.14695f
C4086 a_13011_17910# a_13216_18477# 0.01179f
C4087 sar9b_0.net14 a_12531_28566# 0.05077f
C4088 a_7306_19777# a_7374_19685# 0.35559f
C4089 a_2540_22432# sar9b_0._04_ 0.0164f
C4090 a_4934_22432# a_5441_22522# 0.21226f
C4091 a_7638_19238# a_7914_19178# 0.1263f
C4092 VDPWR a_11339_27039# 0.48115f
C4093 VDPWR a_3369_24181# 0.15274f
C4094 sar9b_0.net24 a_10995_28566# 0.21865f
C4095 sar9b_0.net1 a_9472_23805# 0.01959f
C4096 a_6954_27466# sar9b_0.net60 0.16181f
C4097 a_13011_25902# sar9b_0.net27 0.0399f
C4098 a_10662_17799# a_10410_17846# 0.27388f
C4099 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[2] 4.14971f
C4100 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.59531f
C4101 sar9b_0.net38 uo_out[4] 0.07167f
C4102 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 2.82172f
C4103 sar9b_0.net8 a_11776_21141# 0.3091f
C4104 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.12358f
C4105 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02589f
C4106 a_10402_25094# sar9b_0.net12 0.10692f
C4107 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.SW[0] 0.22983f
C4108 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C4109 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.84427f
C4110 a_8266_18445# a_8334_18353# 0.35559f
C4111 a_10548_19053# a_10098_19171# 0.03432f
C4112 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.SW[3] 0.019f
C4113 a_7188_22119# sar9b_0.net39 0.05015f
C4114 a_5581_20992# sar9b_0._17_ 0.04255f
C4115 a_6126_18353# a_6634_18206# 0.19065f
C4116 a_4467_24162# sar9b_0._15_ 0.11422f
C4117 sar9b_0.net41 a_11436_17742# 0.07436f
C4118 single_9b_cdac_1.CF[7] clk 0.16146f
C4119 sar9b_0.net63 sar9b_0.net57 0.63977f
C4120 single_9b_cdac_0.SW[7] a_30012_26990# 0.18991f
C4121 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[0] 0.01167f
C4122 a_11915_27039# a_11658_26134# 0.04032f
C4123 a_6346_23773# sar9b_0.net11 0.05901f
C4124 a_4467_24162# sar9b_0.clk_div_0.COUNT\[2\] 0.16437f
C4125 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C4126 a_3795_19512# a_3991_19768# 0.0388f
C4127 a_16185_13034# tdc_0.RDY 0.06167f
C4128 sar9b_0.net44 a_3156_26115# 0.23133f
C4129 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C4130 a_10098_19171# sar9b_0.net38 0.02641f
C4131 sar9b_0.net71 a_4072_19474# 0.10694f
C4132 a_8052_18123# sar9b_0.net73 0.05137f
C4133 sar9b_0.net36 a_9138_27163# 0.04377f
C4134 sar9b_0.net13 a_5580_24776# 0.01209f
C4135 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.28575f
C4136 VDPWR a_8202_23174# 0.87317f
C4137 a_8842_16874# sar9b_0.net27 0.08083f
C4138 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[0] 0.22459f
C4139 a_9730_24138# sar9b_0.net38 0.02314f
C4140 a_21368_4076# th_dif_sw_0.VCP 0.18144f
C4141 sar9b_0.net40 sar9b_0.net35 0.52689f
C4142 a_34814_17740# single_9b_cdac_1.SW[6] 0.18991f
C4143 single_9b_cdac_0.SW[0] single_9b_cdac_1.CF[0] 2.15297f
C4144 a_6444_19448# sar9b_0.net15 0.01357f
C4145 sar9b_0.clk_div_0.COUNT\[3\] a_4236_21738# 0.02104f
C4146 sar9b_0.net33 a_12870_26263# 0.07013f
C4147 a_10895_22855# clk 0.0165f
C4148 sar9b_0.net4 sar9b_0.clk_div_0.COUNT\[1\] 0.02438f
C4149 sar9b_0.net35 sar9b_0.net51 0.08262f
C4150 a_10402_27758# a_10607_27849# 0.09983f
C4151 sar9b_0.net27 a_12618_19474# 0.02681f
C4152 a_9165_24988# sar9b_0.net37 0.01216f
C4153 sar9b_0.net40 sar9b_0.net2 0.02933f
C4154 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[7] 0.05361f
C4155 single_9b_cdac_0.cdac_sw_9b_0.S[6] a_34814_26990# 0.22352f
C4156 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.42014f
C4157 a_8098_18810# a_8303_18859# 0.09983f
C4158 sar9b_0.net13 a_6378_24802# 0.08313f
C4159 a_15151_10456# tdc_0.phase_detector_0.INP 0.10793f
C4160 a_9126_23599# sar9b_0.net37 0.02665f
C4161 sar9b_0.net2 sar9b_0.net51 0.02425f
C4162 VDPWR sar9b_0.net58 3.35769f
C4163 sar9b_0.net34 single_9b_cdac_0.SW[8] 0.01408f
C4164 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.clk_div_0.COUNT\[1\] 0.12709f
C4165 sar9b_0.net6 sar9b_0.net37 0.05412f
C4166 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36301f
C4167 sar9b_0.net67 sar9b_0.clknet_1_0__leaf_CLK 0.18709f
C4168 a_11434_16874# a_10644_16791# 0.1263f
C4169 sar9b_0.net58 sar9b_0._14_ 0.12417f
C4170 a_8052_18123# sar9b_0.net48 0.02566f
C4171 VDPWR a_2706_27440# 0.37404f
C4172 sar9b_0.net32 sar9b_0._06_ 0.10957f
C4173 sar9b_0.net32 a_13216_23805# 0.28438f
C4174 sar9b_0.net26 a_13011_24802# 0.22283f
C4175 a_8074_20870# sar9b_0.net56 0.0467f
C4176 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.31534f
C4177 VDPWR a_9323_27662# 0.45921f
C4178 a_10402_25094# a_9942_24806# 0.26257f
C4179 VDPWR uo_out[4] 0.83671f
C4180 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C4181 sar9b_0.net10 a_6922_23534# 0.17349f
C4182 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.38397f
C4183 VDPWR sar9b_0.net47 2.56257f
C4184 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 1.71649f
C4185 a_4018_24235# a_3014_24136# 0.06302f
C4186 VDPWR a_6861_22828# 0.14773f
C4187 sar9b_0.net55 sar9b_0.net57 0.02755f
C4188 a_10895_22855# a_11030_22954# 0.35559f
C4189 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.75853f
C4190 single_9b_cdac_1.CF[4] th_dif_sw_0.VCN 0.09453f
C4191 a_8970_20510# sar9b_0.net37 0.02159f
C4192 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.17533f
C4193 a_8266_17113# sar9b_0.net61 0.04067f
C4194 th_dif_sw_0.CK a_9132_7271# 0.69795f
C4195 single_9b_cdac_1.CF[1] th_dif_sw_0.VCN 0.09453f
C4196 a_4332_23043# clk 0.4678f
C4197 sar9b_0._12_ sar9b_0.net39 0.48411f
C4198 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 a_39616_17740# 0.14695f
C4199 a_6252_19074# a_5844_18123# 0.01266f
C4200 a_3371_23106# sar9b_0.clk_div_0.COUNT\[2\] 0.10533f
C4201 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_53154_16877# 0.04592f
C4202 a_7306_19777# sar9b_0.net10 0.04467f
C4203 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.26942f
C4204 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02519f
C4205 a_45123_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.01076f
C4206 VDPWR a_2508_26108# 0.21993f
C4207 VDPWR sar9b_0.net37 2.42386f
C4208 a_7284_20787# a_6975_20813# 0.07766f
C4209 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.41793f
C4210 a_3206_22432# a_3454_22567# 0.05308f
C4211 sar9b_0.net2 a_10742_21091# 0.02055f
C4212 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.12431f
C4213 a_8266_18445# sar9b_0.net61 0.01651f
C4214 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 2.82165f
C4215 a_8052_18123# sar9b_0.net46 0.16885f
C4216 a_7743_16817# sar9b_0.net6 0.02026f
C4217 a_4755_22138# sar9b_0.net57 0.01782f
C4218 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.27832f
C4219 sar9b_0.net19 a_3754_26815# 0.0389f
C4220 sar9b_0.net36 clk 0.03715f
C4221 sar9b_0.net35 sar9b_0.net62 0.04291f
C4222 a_7138_27758# sar9b_0.net44 0.0155f
C4223 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.19143f
C4224 sar9b_0.net1 sar9b_0.net37 0.27714f
C4225 a_3540_27045# sar9b_0.net19 0.04938f
C4226 VDPWR a_10098_19171# 0.35321f
C4227 a_11842_18434# a_12182_18427# 0.24088f
C4228 VDPWR a_6137_23791# 0.21454f
C4229 sar9b_0.net38 a_10182_20463# 0.0163f
C4230 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.2428f
C4231 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02652f
C4232 a_8726_22954# clk 0.01799f
C4233 sar9b_0.net2 sar9b_0.net62 0.18559f
C4234 sar9b_0.net30 sar9b_0.net10 0.07137f
C4235 a_3922_20239# a_2918_20140# 0.06302f
C4236 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.84424f
C4237 a_5010_28495# a_5151_28559# 0.27388f
C4238 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 1.71649f
C4239 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[1\] 0.89565f
C4240 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.SW[6] 0.03532f
C4241 sar9b_0.net52 a_10482_25831# 0.33514f
C4242 clk tdc_0.phase_detector_0.INP 0.18819f
C4243 sar9b_0.net31 a_11382_22142# 0.03867f
C4244 VDPWR a_3370_26437# 0.20923f
C4245 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INN 0.0434f
C4246 VDPWR a_6642_19448# 0.3497f
C4247 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C4248 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] 3.14416f
C4249 a_5580_24776# sar9b_0._15_ 0.26726f
C4250 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.38397f
C4251 VDPWR a_9730_24138# 0.22331f
C4252 a_2508_27440# a_2706_27440# 0.06623f
C4253 a_11146_25483# a_10482_25831# 0.16939f
C4254 single_9b_cdac_1.CF[8] th_dif_sw_0.VCN 0.09453f
C4255 a_11658_19474# single_9b_cdac_1.SW[8] 0.01298f
C4256 a_11915_28371# single_9b_cdac_0.SW[5] 0.0323f
C4257 a_10166_3438# a_10482_3438# 0.62294f
C4258 sar9b_0.net36 single_9b_cdac_1.SW[0] 0.14f
C4259 a_7498_21109# a_7284_20787# 0.04522f
C4260 a_10644_16791# a_10335_16817# 0.07766f
C4261 sar9b_0.clk_div_0.COUNT\[2\] a_5580_24776# 0.02755f
C4262 VDPWR a_7602_18116# 0.3287f
C4263 a_10662_17799# a_11008_17491# 0.07649f
C4264 sar9b_0.net32 single_9b_cdac_1.CF[6] 0.03698f
C4265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C4266 VDPWR a_7743_16817# 0.26065f
C4267 sar9b_0.net60 sar9b_0.net54 0.10669f
C4268 sar9b_0.net41 sar9b_0.net27 0.03867f
C4269 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.12431f
C4270 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 ua[0] 0.15943f
C4271 sar9b_0.net70 sar9b_0._12_ 0.02802f
C4272 VDPWR a_11842_22430# 0.22622f
C4273 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.38397f
C4274 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] 1.14951f
C4275 a_7478_27751# sar9b_0.net45 0.02536f
C4276 a_7602_18116# sar9b_0.net1 0.03058f
C4277 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38715f
C4278 sar9b_0.net4 a_6378_24802# 0.2298f
C4279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.22875f
C4280 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.11216f
C4281 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.02638f
C4282 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.7611f
C4283 sar9b_0.net54 a_5753_24250# 0.09858f
C4284 a_2918_20140# a_3273_20185# 0.18752f
C4285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4286 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.42784f
C4287 sar9b_0.clk_div_0.COUNT\[1\] sar9b_0.clknet_1_1__leaf_CLK 1.13184f
C4288 a_10803_18142# sar9b_0.net36 0.02932f
C4289 VDPWR a_11842_23762# 0.2306f
C4290 a_5441_22522# sar9b_0._07_ 0.02011f
C4291 a_10402_25094# a_11430_24931# 0.07826f
C4292 sar9b_0.net26 a_12618_19474# 0.03006f
C4293 a_12531_28566# uo_out[0] 0.12656f
C4294 VDPWR a_3166_20145# 0.02403f
C4295 a_9165_24988# sar9b_0.net57 0.05719f
C4296 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C4297 sar9b_0.net40 a_6744_23238# 0.02487f
C4298 sar9b_0._08_ sar9b_0._07_ 0.02717f
C4299 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C4300 a_5506_26802# a_5846_26950# 0.24088f
C4301 sar9b_0.net43 a_10070_24286# 0.04223f
C4302 a_13011_16810# single_9b_cdac_1.SW[3] 0.03223f
C4303 sar9b_0._17_ a_6444_21738# 0.02137f
C4304 single_9b_cdac_0.cdac_sw_9b_0.S[0] clk 0.03331f
C4305 sar9b_0.net49 a_9359_20191# 0.18621f
C4306 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 ua[0] 0.12358f
C4307 sar9b_0.net43 a_7347_24160# 0.03385f
C4308 sar9b_0.net6 a_7404_18116# 0.28739f
C4309 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[1\] 0.02265f
C4310 sar9b_0.net72 a_4044_24776# 0.16551f
C4311 a_3371_23106# sar9b_0.clknet_1_1__leaf_CLK 0.02302f
C4312 single_9b_cdac_1.CF[3] th_dif_sw_0.VCN 0.09453f
C4313 sar9b_0.net9 a_7978_22202# 0.04916f
C4314 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.42509f
C4315 sar9b_0.net40 a_5748_24381# 0.02394f
C4316 a_10182_20463# a_8970_20510# 0.07766f
C4317 single_9b_cdac_0.SW[2] clk 0.13337f
C4318 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.A 0.26382f
C4319 sar9b_0.net10 a_7978_22202# 0.08861f
C4320 a_7978_22202# sar9b_0.net61 0.17441f
C4321 a_9472_18823# sar9b_0.net37 0.03442f
C4322 a_10218_20806# a_10742_21091# 0.05022f
C4323 sar9b_0.net7 a_11842_18434# 0.01552f
C4324 a_5460_28377# a_5674_28147# 0.05022f
C4325 VDPWR a_10182_20463# 0.26691f
C4326 VDPWR single_9b_cdac_1.SW[5] 2.51859f
C4327 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C4328 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4329 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.47485f
C4330 a_10482_3438# a_10254_2858# 0.11186f
C4331 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[7] 0.01887f
C4332 VDPWR sar9b_0.net57 1.46403f
C4333 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36037f
C4334 a_10644_16791# sar9b_0.net48 0.15925f
C4335 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.42509f
C4336 a_7914_23470# sar9b_0.net62 0.02516f
C4337 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[5] 18.8692f
C4338 VDPWR a_7404_18116# 0.19099f
C4339 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[7] 0.06503f
C4340 sar9b_0.net10 sar9b_0._17_ 0.01904f
C4341 VDPWR sar9b_0.net33 0.38773f
C4342 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] 1.55981f
C4343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR 0.62553f
C4344 sar9b_0.net7 a_9363_20826# 0.03016f
C4345 a_8386_22806# a_9162_23174# 0.3578f
C4346 single_9b_cdac_1.CF[0] clk 0.08196f
C4347 sar9b_0.net40 a_6880_26815# 0.01367f
C4348 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.12431f
C4349 a_5682_23444# a_6137_23791# 0.3578f
C4350 a_6132_23451# a_6346_23773# 0.04522f
C4351 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.42015f
C4352 ui_in[4] ui_in[3] 0.03102f
C4353 a_5506_17478# a_6534_17799# 0.07826f
C4354 a_9942_27470# sar9b_0.net38 0.01957f
C4355 sar9b_0.net51 a_5811_19178# 0.11557f
C4356 sar9b_0._16_ a_3372_25734# 0.26724f
C4357 VDPWR a_8031_26141# 0.26325f
C4358 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.28523f
C4359 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C4360 a_11776_27801# single_9b_cdac_0.SW[5] 0.01854f
C4361 sar9b_0.net52 sar9b_0.net27 0.01796f
C4362 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C4363 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.94957f
C4364 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 3.27803f
C4365 sar9b_0.net52 single_9b_cdac_0.SW[5] 0.12211f
C4366 sar9b_0.net11 a_13011_24570# 0.22279f
C4367 a_18214_3039# th_dif_sw_0.th_sw_1.CKB 0.42927f
C4368 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.11944f
C4369 sar9b_0.net22 uo_out[5] 0.01216f
C4370 a_9546_24506# a_9935_24187# 0.05462f
C4371 a_9270_24566# a_9730_24138# 0.26257f
C4372 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[0] 1.83507f
C4373 a_10194_16784# sar9b_0.net6 0.07207f
C4374 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.84061f
C4375 clk single_9b_cdac_1.SW[2] 0.17199f
C4376 a_10239_19235# sar9b_0.net48 0.22117f
C4377 sar9b_0.net41 sar9b_0.net26 0.02726f
C4378 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.03488f
C4379 sar9b_0.net43 a_11859_20574# 0.20839f
C4380 sar9b_0.net48 a_9634_17478# 0.1085f
C4381 single_9b_cdac_1.CF[8] sar9b_0.net13 0.01097f
C4382 sar9b_0.net32 single_9b_cdac_1.CF[7] 0.01485f
C4383 a_10402_25094# sar9b_0.net74 0.02019f
C4384 a_7914_27466# a_8115_28566# 0.01021f
C4385 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C4386 a_6540_22112# sar9b_0.net40 0.01639f
C4387 a_5083_21100# sar9b_0.net65 0.01754f
C4388 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[7] 6.17399f
C4389 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.22512f
C4390 a_5196_18116# a_5535_18149# 0.07649f
C4391 a_5844_18123# a_5394_18116# 0.03471f
C4392 a_8052_16791# a_7743_16817# 0.07766f
C4393 sar9b_0.net50 a_12047_19857# 0.22617f
C4394 a_6346_23773# sar9b_0.net4 0.01825f
C4395 sar9b_0.net40 sar9b_0.net39 0.04664f
C4396 single_9b_cdac_1.SW[0] a_9450_17846# 0.02044f
C4397 VDPWR a_4467_24162# 0.42883f
C4398 single_9b_cdac_1.SW[2] single_9b_cdac_1.SW[0] 0.98657f
C4399 sar9b_0.net42 sar9b_0.net2 0.15479f
C4400 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.42509f
C4401 a_9138_27163# a_9279_27227# 0.27388f
C4402 sar9b_0.net51 sar9b_0.net39 0.01895f
C4403 a_4467_24162# sar9b_0._14_ 0.11012f
C4404 sar9b_0.net56 a_9450_17846# 0.26827f
C4405 tdc_0.RDY a_5331_16810# 0.26021f
C4406 a_5465_28246# uo_out[7] 0.0105f
C4407 sar9b_0.net56 single_9b_cdac_1.SW[2] 0.31153f
C4408 a_7890_26108# sar9b_0.net59 0.30461f
C4409 clk a_16331_9671# 0.37638f
C4410 VDPWR a_10194_16784# 0.31773f
C4411 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C4412 sar9b_0.net52 a_7638_23474# 0.19487f
C4413 a_11658_22138# a_11842_22430# 0.44532f
C4414 a_10937_25582# a_11214_25728# 0.09983f
C4415 a_11338_19178# sar9b_0.net61 0.24596f
C4416 a_21368_4076# th_dif_sw_0.CKB 0.01417f
C4417 single_9b_cdac_1.SW[8] clk 0.08196f
C4418 VDPWR a_4496_20468# 0.33806f
C4419 a_11722_25838# a_11214_25728# 0.19065f
C4420 a_6767_25185# sar9b_0.net54 0.20328f
C4421 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.02149f
C4422 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.06503f
C4423 a_8982_21902# a_9647_21523# 0.19065f
C4424 a_9258_21842# a_9782_21622# 0.04522f
C4425 a_6534_17799# a_5322_17846# 0.07766f
C4426 VDPWR a_11178_24802# 0.33967f
C4427 sar9b_0.net9 a_7188_22119# 0.22374f
C4428 a_2835_24136# a_3262_24141# 0.04602f
C4429 a_8874_23470# sar9b_0.net54 0.09219f
C4430 a_10230_23234# sar9b_0.net38 0.01802f
C4431 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.01152f
C4432 a_9939_28566# uo_out[3] 0.40366f
C4433 a_8098_18810# sar9b_0.net51 0.0158f
C4434 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96978f
C4435 sar9b_0.net33 sar9b_0.net29 0.01075f
C4436 sar9b_0.net9 clk 0.02916f
C4437 a_7188_22119# sar9b_0.net10 0.01911f
C4438 sar9b_0.net47 a_7193_22459# 0.10511f
C4439 VDPWR a_16159_13315# 0.22342f
C4440 a_8074_20870# sar9b_0.net51 0.06285f
C4441 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.05105f
C4442 a_13011_19242# sar9b_0.net28 0.01241f
C4443 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[0] 0.02165f
C4444 a_2547_28132# uio_out[1] 0.03336f
C4445 a_9942_27470# VDPWR 0.30254f
C4446 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.17533f
C4447 a_5633_20244# a_5481_20185# 0.22338f
C4448 sar9b_0.net42 a_10758_24459# 0.01335f
C4449 VDPWR sar9b_0.clk_div_0.COUNT\[1\] 0.71891f
C4450 sar9b_0.net10 clk 0.1264f
C4451 tdc_0.RDY sar9b_0.net27 0.05081f
C4452 sar9b_0.net70 a_2892_23070# 0.01508f
C4453 sar9b_0.net49 sar9b_0.net2 0.02449f
C4454 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 0.19147f
C4455 VDPWR a_33936_26999# 1.81495f
C4456 sar9b_0._14_ sar9b_0.clk_div_0.COUNT\[1\] 0.03517f
C4457 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 3.10626f
C4458 a_5682_23444# sar9b_0.net57 0.06802f
C4459 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.22497f
C4460 VDPWR a_10410_17846# 0.32302f
C4461 single_9b_cdac_1.CF[5] th_dif_sw_0.VCN 0.09453f
C4462 single_9b_cdac_0.SW[4] th_dif_sw_0.VCN 0.09453f
C4463 a_8691_28566# uo_out[4] 0.37881f
C4464 a_10644_16791# a_11436_17742# 0.01113f
C4465 single_9b_cdac_0.SW[6] a_9323_28371# 0.38985f
C4466 a_6252_19074# a_6579_18832# 0.09203f
C4467 sar9b_0.net58 sar9b_0._03_ 0.03496f
C4468 a_11338_19178# sar9b_0.net7 0.0556f
C4469 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.12358f
C4470 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.06503f
C4471 sar9b_0.net62 sar9b_0.net39 0.02577f
C4472 sar9b_0.net52 a_8303_23853# 0.19552f
C4473 sar9b_0.net40 a_6902_25087# 0.0115f
C4474 sar9b_0.net12 a_9942_24806# 0.21789f
C4475 sar9b_0.net56 sar9b_0.net9 0.089f
C4476 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR 0.38716f
C4477 sar9b_0._10_ a_5196_19448# 0.10468f
C4478 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02813f
C4479 a_8303_18859# sar9b_0.net61 0.03127f
C4480 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.69086f
C4481 sar9b_0.net63 a_6346_23773# 0.03952f
C4482 a_5628_19768# a_5581_19664# 0.19021f
C4483 VDPWR a_3371_23106# 0.3848f
C4484 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.0303f
C4485 sar9b_0.net61 single_9b_cdac_1.SW[0] 0.03934f
C4486 sar9b_0.net41 sar9b_0.net53 0.28496f
C4487 sar9b_0.net33 a_11382_26138# 0.06166f
C4488 tdc_0.OUTP tdc_0.RDY 1.84081f
C4489 a_24332_26999# m2_23774_26966# 0.01541f
C4490 VDPWR a_6834_20780# 0.32839f
C4491 sar9b_0.net56 sar9b_0.net61 0.16507f
C4492 sar9b_0.net56 a_10402_21098# 0.01558f
C4493 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.26707f
C4494 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.26707f
C4495 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.38397f
C4496 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4497 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.75853f
C4498 sar9b_0.net58 a_5711_26851# 0.21873f
C4499 a_10402_27758# a_11178_27466# 0.3578f
C4500 VDPWR a_7443_21496# 0.44805f
C4501 a_8386_22806# sar9b_0.net11 0.15667f
C4502 VDPWR a_10803_19474# 0.44387f
C4503 a_21368_4076# ua[3] 0.65763f
C4504 sar9b_0.net45 single_9b_cdac_0.SW[4] 0.24467f
C4505 sar9b_0.net40 sar9b_0.net36 0.14787f
C4506 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C4507 a_4922_20857# a_5083_21100# 0.19021f
C4508 a_4136_25584# a_4365_25770# 0.18757f
C4509 a_8074_20870# sar9b_0.net62 0.01645f
C4510 VDPWR a_21177_7457# 1.54446f
C4511 a_5100_24375# a_5439_24563# 0.07649f
C4512 clk a_16527_10454# 0.20249f
C4513 a_13011_24802# single_9b_cdac_0.SW[0] 0.35451f
C4514 sar9b_0.net36 sar9b_0.net51 0.02568f
C4515 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.04988f
C4516 single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.26707f
C4517 sar9b_0._16_ a_3747_25724# 0.02266f
C4518 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.04988f
C4519 sar9b_0.net18 a_3438_27677# 0.04725f
C4520 sar9b_0.net41 a_9494_20290# 0.01451f
C4521 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 2.81139f
C4522 a_5581_19664# sar9b_0.net4 0.01002f
C4523 a_2547_28132# sar9b_0.net17 0.0815f
C4524 sar9b_0.net23 sar9b_0.net37 0.02446f
C4525 single_9b_cdac_0.cdac_sw_9b_0.S[4] th_dif_sw_0.VCN 13.5521f
C4526 a_3713_22522# sar9b_0.clknet_1_1__leaf_CLK 0.04145f
C4527 VDPWR a_10230_23234# 0.30161f
C4528 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[3] 0.02149f
C4529 VDPWR a_5580_24776# 0.24626f
C4530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[7] 0.42014f
C4531 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C4532 a_4210_22378# sar9b_0.clk_div_0.COUNT\[3\] 0.12081f
C4533 a_5711_26851# sar9b_0.net37 0.0259f
C4534 a_8595_17910# sar9b_0.net35 0.20113f
C4535 sar9b_0.net7 sar9b_0.net56 0.25867f
C4536 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C4537 single_9b_cdac_1.cdac_sw_9b_0.S[1] th_dif_sw_0.VCP 0.10984p
C4538 sar9b_0.net14 sar9b_0._06_ 0.04595f
C4539 sar9b_0.net38 a_10284_25707# 0.02385f
C4540 a_8098_18810# a_7914_19178# 0.44098f
C4541 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.04988f
C4542 sar9b_0.net51 a_5844_18123# 0.01122f
C4543 a_3206_22432# sar9b_0._12_ 0.04817f
C4544 a_7138_27758# sar9b_0.net60 0.0875f
C4545 VDPWR ua[0] 93.85329f
C4546 tdc_0.OUTP a_13011_16810# 0.01868f
C4547 sar9b_0.net36 a_10742_21091# 0.0132f
C4548 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.3196f
C4549 a_9802_26815# a_9593_26914# 0.24088f
C4550 VDPWR a_6378_24802# 0.83745f
C4551 single_9b_cdac_0.SW[8] uo_out[1] 0.10947f
C4552 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C4553 sar9b_0.net17 a_2451_27234# 0.0211f
C4554 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.22875f
C4555 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.84427f
C4556 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] 1.1512f
C4557 sar9b_0.net7 a_10803_18142# 0.01039f
C4558 sar9b_0.net49 a_10218_20806# 0.2026f
C4559 a_8512_27801# sar9b_0.cyclic_flag_0.FINAL 0.03823f
C4560 a_11430_24931# sar9b_0.net12 0.07831f
C4561 uo_out[4] ui_in[0] 0.06786f
C4562 VDPWR single_9b_cdac_1.CF[2] 3.12459f
C4563 sar9b_0.net55 a_7347_24160# 0.19384f
C4564 single_9b_cdac_0.cdac_sw_9b_0.S[2] ua[0] 1.2071f
C4565 sar9b_0.net24 sar9b_0.net45 0.03105f
C4566 sar9b_0._05_ a_4236_21738# 0.27985f
C4567 a_2508_20780# a_2918_20140# 0.05315f
C4568 sar9b_0.net68 sar9b_0.clk_div_0.COUNT\[2\] 0.49269f
C4569 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] 0.12898f
C4570 a_9930_20510# sar9b_0.net5 0.07266f
C4571 VDPWR sar9b_0.net19 0.3982f
C4572 sar9b_0.net52 sar9b_0.net53 0.37319f
C4573 sar9b_0._11_ a_6636_20780# 0.02384f
C4574 sar9b_0.net8 a_8694_20570# 0.05489f
C4575 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.SW[5] 0.03636f
C4576 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.84059f
C4577 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C4578 a_5823_23477# sar9b_0.net54 0.16953f
C4579 VDPWR a_13011_21906# 0.47029f
C4580 a_3545_26914# a_3822_27060# 0.09983f
C4581 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07517f
C4582 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.SW[8] 0.17126f
C4583 sar9b_0.net36 a_9588_27045# 0.07056f
C4584 sar9b_0.net35 sar9b_0.net11 0.02957f
C4585 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.22879f
C4586 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.06503f
C4587 sar9b_0.net65 a_4947_20140# 0.01364f
C4588 a_2451_27234# a_2892_27039# 0.01819f
C4589 a_7289_21127# sar9b_0.net47 0.10682f
C4590 sar9b_0.net2 sar9b_0.net11 0.02395f
C4591 sar9b_0.net73 a_11382_22142# 0.17249f
C4592 a_13011_19242# a_13216_18477# 0.01043f
C4593 sar9b_0.net12 sar9b_0.net54 0.03647f
C4594 th_dif_sw_0.CK sar9b_0.net73 0.16091f
C4595 a_10070_24286# sar9b_0.net38 0.01531f
C4596 a_3819_24136# a_4018_24235# 0.29821f
C4597 uio_in[1] uio_in[0] 0.03102f
C4598 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_21368_4076# 1.16499f
C4599 a_8622_26345# sar9b_0.cyclic_flag_0.FINAL 0.0786f
C4600 a_7374_19685# sar9b_0.net40 0.01327f
C4601 a_9126_19131# sar9b_0.net48 0.21244f
C4602 sar9b_0.net49 a_8982_21902# 0.22591f
C4603 sar9b_0.net33 a_13216_26469# 0.30861f
C4604 sar9b_0._09_ sar9b_0.net16 0.56465f
C4605 a_3946_26198# sar9b_0.net44 0.05662f
C4606 sar9b_0.net20 uo_out[5] 0.09694f
C4607 VDPWR a_11008_17491# 0.1898f
C4608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.22879f
C4609 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[6] 0.06019f
C4610 a_8303_18859# a_8438_18958# 0.35559f
C4611 sar9b_0.net20 sar9b_0.net21 0.32153f
C4612 single_9b_cdac_0.SW[4] a_12560_27128# 0.03746f
C4613 a_9450_17846# a_9174_17906# 0.1263f
C4614 a_11658_19474# a_12618_19474# 0.03432f
C4615 single_9b_cdac_0.SW[2] a_53154_26999# 0.28324f
C4616 single_9b_cdac_1.SW[2] a_9174_17906# 0.07801f
C4617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C4618 tdc_0.OUTP a_10644_16791# 0.07935f
C4619 a_10858_17113# a_10194_16784# 0.16939f
C4620 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C4621 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.10429f
C4622 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[3] 4.15032f
C4623 sar9b_0.net36 uo_out[7] 0.10138f
C4624 VDPWR a_10284_25707# 0.20062f
C4625 VDPWR a_3161_27787# 0.24214f
C4626 sar9b_0.net63 sar9b_0.net68 0.09062f
C4627 sar9b_0.net42 sar9b_0.net39 1.25124f
C4628 single_9b_cdac_1.SW[1] sar9b_0.net73 0.05555f
C4629 a_5182_22567# sar9b_0._12_ 0.01992f
C4630 sar9b_0.net35 a_7338_24802# 0.03288f
C4631 th_dif_sw_0.CK sar9b_0.net48 0.03264f
C4632 single_9b_cdac_1.CF[2] sar9b_0.net29 0.03358f
C4633 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] 3.10045f
C4634 a_11466_23174# sar9b_0.net53 0.28157f
C4635 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.84424f
C4636 sar9b_0._18_ a_3219_22860# 0.07732f
C4637 a_10690_22806# a_11466_23174# 0.3578f
C4638 a_5711_17527# sar9b_0.net46 0.26531f
C4639 th_dif_sw_0.CK th_dif_sw_0.th_sw_1.CK 0.01565f
C4640 a_3695_23038# sar9b_0.clk_div_0.COUNT\[2\] 0.21948f
C4641 sar9b_0.net23 a_8031_26141# 0.02315f
C4642 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.95338f
C4643 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C4644 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.01003f
C4645 sar9b_0.net43 sar9b_0.net24 0.02255f
C4646 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.7611f
C4647 sar9b_0.net74 sar9b_0.net12 0.05557f
C4648 sar9b_0.net60 a_4583_20468# 0.01054f
C4649 VDPWR a_2706_26108# 0.40591f
C4650 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.07579f
C4651 a_3206_22432# a_4011_22488# 0.29207f
C4652 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.23864f
C4653 sar9b_0.net44 sar9b_0.net21 0.03003f
C4654 a_16222_11316# tdc_0.phase_detector_0.INN 0.02415f
C4655 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP a_33936_26999# 0.04592f
C4656 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[0\] 0.03041f
C4657 sar9b_0.net64 sar9b_0.net57 0.02277f
C4658 sar9b_0.net31 sar9b_0.net12 0.61825f
C4659 a_6307_27584# sar9b_0.net40 0.10226f
C4660 VDPWR w_17430_1606# 0.44324f
C4661 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.75899f
C4662 sar9b_0.net68 sar9b_0.clknet_1_1__leaf_CLK 0.02176f
C4663 a_11658_19474# a_12182_19759# 0.05022f
C4664 sar9b_0.net49 sar9b_0.net39 0.01106f
C4665 clk tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.09743f
C4666 a_13011_20574# single_9b_cdac_1.CF[0] 0.36053f
C4667 VDPWR a_6346_23773# 0.20258f
C4668 VDPWR a_6534_17799# 0.26217f
C4669 sar9b_0.net15 a_6252_19074# 0.25177f
C4670 sar9b_0.net20 a_5460_28377# 0.09259f
C4671 a_5010_28495# a_5465_28246# 0.3578f
C4672 VDPWR a_3713_22522# 0.10433f
C4673 a_11915_27039# sar9b_0.net45 0.10003f
C4674 th_dif_sw_0.CK sar9b_0.net50 0.23424f
C4675 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[8] 0.01285f
C4676 sar9b_0.net48 single_9b_cdac_1.SW[1] 0.05838f
C4677 sar9b_0.net52 a_10932_25713# 0.17701f
C4678 sar9b_0.net58 a_2706_27440# 0.26179f
C4679 th_dif_sw_0.CK single_9b_cdac_1.SW[3] 0.69076f
C4680 single_9b_cdac_1.CF[1] sar9b_0.net6 0.01228f
C4681 VDPWR a_7097_19795# 0.22516f
C4682 sar9b_0.net40 single_9b_cdac_1.SW[8] 0.02686f
C4683 th_dif_sw_0.CK a_12618_18142# 0.06719f
C4684 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.15052f
C4685 a_4811_23656# sar9b_0.net72 0.2012f
C4686 VDPWR a_3922_20239# 0.38261f
C4687 VDPWR a_10070_24286# 0.20147f
C4688 a_11146_25483# a_10932_25713# 0.05022f
C4689 a_3156_27447# a_2847_27473# 0.07766f
C4690 a_11842_19766# single_9b_cdac_1.SW[8] 0.02175f
C4691 sar9b_0.net61 a_9174_17906# 0.04236f
C4692 a_10482_3438# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.63339f
C4693 sar9b_0.net45 sar9b_0._06_ 0.01013f
C4694 single_9b_cdac_1.SW[8] sar9b_0.net51 0.0423f
C4695 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C4696 VDPWR a_7347_24160# 0.44946f
C4697 single_9b_cdac_0.SW[7] uo_out[1] 0.04613f
C4698 sar9b_0.net59 sar9b_0.net34 0.14932f
C4699 a_7914_23470# sar9b_0.net11 0.07548f
C4700 single_9b_cdac_1.SW[4] clk 0.09021f
C4701 VDPWR a_8057_18463# 0.24516f
C4702 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[5] 17.8424f
C4703 a_3603_28156# uio_out[1] 0.013f
C4704 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.22879f
C4705 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C4706 single_9b_cdac_0.SW[3] ua[0] 0.16155f
C4707 VDPWR a_12870_22267# 0.25924f
C4708 a_6250_28502# a_5460_28377# 0.1263f
C4709 sar9b_0.net58 sar9b_0.net37 0.24097f
C4710 a_7914_27466# sar9b_0.net45 0.07701f
C4711 a_8057_18463# sar9b_0.net1 0.15171f
C4712 sar9b_0.net9 sar9b_0.net51 0.02854f
C4713 sar9b_0.net48 a_6126_18353# 0.22812f
C4714 a_6102_24806# a_6562_25094# 0.26257f
C4715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] 3.10215f
C4716 sar9b_0.net59 a_3156_26115# 0.17719f
C4717 a_5046_17906# sar9b_0.net46 0.41373f
C4718 sar9b_0.net40 sar9b_0.net10 0.35246f
C4719 sar9b_0.net40 sar9b_0.net61 0.03026f
C4720 VDPWR sar9b_0.net3 0.45768f
C4721 VDPWR single_9b_cdac_1.CF[4] 2.77384f
C4722 VDPWR single_9b_cdac_1.CF[1] 2.73909f
C4723 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.03729f
C4724 a_6484_22845# sar9b_0._02_ 0.01922f
C4725 a_2918_20140# a_3723_20140# 0.29221f
C4726 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[0] 0.02202f
C4727 sar9b_0.net10 sar9b_0.net51 0.09304f
C4728 sar9b_0.net61 sar9b_0.net51 0.06277f
C4729 single_9b_cdac_1.CF[6] th_dif_sw_0.VCN 0.09453f
C4730 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[1] 0.26555f
C4731 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.23119f
C4732 VDPWR a_12531_28566# 0.45349f
C4733 VDPWR a_12870_23599# 0.25929f
C4734 sar9b_0.net42 sar9b_0.net36 0.59867f
C4735 a_10742_25087# a_11178_24802# 0.16939f
C4736 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.10499f
C4737 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[8] 0.05858f
C4738 sar9b_0._06_ uo_out[0] 0.19708f
C4739 VDPWR a_3273_20185# 0.14496f
C4740 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.SW[7] 0.22983f
C4741 single_9b_cdac_1.cdac_sw_9b_0.S[6] a_33936_16877# 0.59531f
C4742 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36412f
C4743 sar9b_0.net6 a_11859_20574# 0.01121f
C4744 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31753_29911# 0.01076f
C4745 sar9b_0.net40 a_6538_24506# 0.01312f
C4746 sar9b_0.net43 sar9b_0.net35 0.06071f
C4747 a_5083_21100# sar9b_0._17_ 0.01853f
C4748 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C4749 a_9942_27470# sar9b_0.net23 0.02292f
C4750 a_3438_26345# sar9b_0.net59 0.22622f
C4751 a_10859_26330# sar9b_0.net74 0.1037f
C4752 a_11658_23470# sar9b_0.net11 0.24021f
C4753 single_9b_cdac_1.SW[8] a_13011_20574# 0.01361f
C4754 a_53154_16877# single_9b_cdac_1.SW[2] 0.28324f
C4755 VDPWR a_7478_27751# 0.20242f
C4756 sar9b_0.net13 sar9b_0.net35 0.02962f
C4757 sar9b_0.net43 sar9b_0.net2 1.88515f
C4758 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.62443f
C4759 a_10707_23470# sar9b_0.net38 0.01005f
C4760 a_3695_23038# sar9b_0.clknet_1_1__leaf_CLK 0.01667f
C4761 a_10239_19235# sar9b_0.net26 0.06761f
C4762 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] 1.15122f
C4763 sar9b_0._09_ sar9b_0._11_ 0.01658f
C4764 VDPWR a_11382_18146# 0.30035f
C4765 VDPWR dw_12589_1395# 1.90366f
C4766 sar9b_0.net46 a_3795_19512# 0.08659f
C4767 a_7914_23470# a_8098_23762# 0.44532f
C4768 VDPWR a_4236_21738# 0.23821f
C4769 VDPWR single_9b_cdac_1.CF[8] 2.63907f
C4770 a_6642_19448# sar9b_0.net47 0.33504f
C4771 sar9b_0.net7 sar9b_0.net40 0.02438f
C4772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.45521f
C4773 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.CF[7] 0.0174f
C4774 a_4947_20140# a_5931_20140# 0.08669f
C4775 a_10218_20806# a_11178_20806# 0.03432f
C4776 a_10402_21098# a_10742_21091# 0.24088f
C4777 a_5465_28246# sar9b_0.net45 0.02195f
C4778 a_5742_28392# a_5674_28147# 0.35559f
C4779 VDPWR a_11859_20574# 0.41872f
C4780 sar9b_0.net30 sar9b_0.net52 0.05789f
C4781 sar9b_0.net7 sar9b_0.net51 0.02342f
C4782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C4783 sar9b_0.net9 sar9b_0.net62 0.02856f
C4784 a_12491_27662# sar9b_0._06_ 0.04301f
C4785 sar9b_0.net42 a_10937_25582# 0.02311f
C4786 sar9b_0.net49 sar9b_0.net36 0.04379f
C4787 VDPWR a_12588_16784# 0.22693f
C4788 a_10553_18922# sar9b_0.net73 0.02068f
C4789 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] 1.14952f
C4790 a_10548_19053# a_10762_18823# 0.05022f
C4791 sar9b_0.net3 a_2508_27440# 0.02829f
C4792 sar9b_0.net45 a_7343_27849# 0.06174f
C4793 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# 0.18915f
C4794 sar9b_0.net10 sar9b_0.net62 0.15663f
C4795 sar9b_0.net61 sar9b_0.net62 0.26134f
C4796 a_6534_27123# a_5322_27170# 0.07766f
C4797 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.7611f
C4798 a_8726_22954# a_9162_23174# 0.16939f
C4799 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.02149f
C4800 sar9b_0.net43 a_10758_24459# 0.03693f
C4801 clk rst_n 0.03102f
C4802 a_5682_23444# a_6346_23773# 0.16939f
C4803 VDPWR a_5581_19664# 0.23366f
C4804 sar9b_0.net51 a_6579_18832# 0.26023f
C4805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.19266f
C4806 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.81428f
C4807 single_9b_cdac_1.cdac_sw_9b_0.S[8] th_dif_sw_0.VCP 0.85562f
C4808 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36044f
C4809 a_8019_17910# sar9b_0.net56 0.06841f
C4810 sar9b_0.net35 a_6132_23451# 0.01493f
C4811 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.31534f
C4812 uo_out[3] uo_out[2] 3.18986f
C4813 VDPWR a_7402_22441# 0.20328f
C4814 VDPWR a_5151_28559# 0.26391f
C4815 a_4755_22138# a_5289_22527# 0.35097f
C4816 single_9b_cdac_1.CF[4] sar9b_0.net29 0.03153f
C4817 a_11915_27039# a_12560_27128# 0.02698f
C4818 a_6538_24506# sar9b_0.net62 0.1665f
C4819 single_9b_cdac_1.CF[1] sar9b_0.net29 0.04096f
C4820 a_5580_24776# sar9b_0._03_ 0.1431f
C4821 a_8202_23174# sar9b_0.net57 0.01828f
C4822 a_7092_19455# a_7306_19777# 0.04522f
C4823 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.28523f
C4824 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 1.71649f
C4825 a_3747_25724# a_4136_25584# 0.06302f
C4826 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] 3.10217f
C4827 a_8303_23853# a_8438_23755# 0.35559f
C4828 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.38397f
C4829 sar9b_0.net7 a_10742_21091# 0.06412f
C4830 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26955f
C4831 a_11718_23127# a_12064_22819# 0.07649f
C4832 a_12560_27128# sar9b_0._06_ 0.0956f
C4833 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.75853f
C4834 a_10649_17131# sar9b_0.net6 0.09326f
C4835 sar9b_0.net56 a_8842_18206# 0.0572f
C4836 a_9935_24187# sar9b_0.net12 0.01643f
C4837 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.04988f
C4838 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.03484f
C4839 a_10553_18922# sar9b_0.net48 0.08167f
C4840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.69086f
C4841 sar9b_0.net11 sar9b_0.net39 0.01153f
C4842 single_9b_cdac_1.CF[7] sar9b_0.net11 0.03981f
C4843 a_2835_24136# sar9b_0.clknet_1_1__leaf_CLK 0.33556f
C4844 sar9b_0.net48 a_9974_17626# 0.13813f
C4845 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[7] 0.01285f
C4846 a_8512_27801# sar9b_0.net22 0.27285f
C4847 a_11430_24931# sar9b_0.net74 0.01382f
C4848 VDPWR single_9b_cdac_1.CF[3] 2.76152f
C4849 VDPWR sar9b_0.net28 1.71321f
C4850 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] 1.55946f
C4851 sar9b_0.net8 sar9b_0.net5 0.02967f
C4852 a_8052_18123# a_8266_18445# 0.04522f
C4853 VDPWR sar9b_0.net68 0.48583f
C4854 a_5844_18123# a_5849_18463# 0.44098f
C4855 a_5394_18116# a_5535_18149# 0.27388f
C4856 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36037f
C4857 VDPWR a_5812_21028# 0.2311f
C4858 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26427f
C4859 a_7602_16784# a_8057_17131# 0.3578f
C4860 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.42014f
C4861 sar9b_0._14_ sar9b_0.net68 0.7985f
C4862 sar9b_0.net31 a_11430_24931# 0.0265f
C4863 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.02638f
C4864 tdc_0.phase_detector_0.INN tdc_0.phase_detector_0.INP 1.21226f
C4865 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.05472f
C4866 tdc_0.OUTN a_6867_16810# 0.28739f
C4867 a_9279_27227# a_9588_27045# 0.07766f
C4868 a_9138_27163# a_9593_26914# 0.3578f
C4869 VDPWR a_10707_23470# 0.26572f
C4870 single_9b_cdac_1.CF[8] sar9b_0.net29 0.30185f
C4871 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C4872 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.01472f
C4873 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.11216f
C4874 VDPWR a_10816_21487# 0.20703f
C4875 a_10402_27758# sar9b_0.net45 0.09798f
C4876 a_21684_3438# a_21368_4076# 0.62294f
C4877 a_8345_26455# sar9b_0.net59 0.08274f
C4878 clk a_16357_9613# 0.01204f
C4879 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.7611f
C4880 VDPWR a_10649_17131# 0.21441f
C4881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.42784f
C4882 single_9b_cdac_1.CF[7] th_dif_sw_0.VCN 0.09453f
C4883 sar9b_0.clknet_1_0__leaf_CLK a_3425_20244# 0.0505f
C4884 sar9b_0._18_ sar9b_0.clknet_0_CLK 0.14719f
C4885 a_11658_22138# a_12870_22267# 0.07766f
C4886 sar9b_0.net47 sar9b_0.net57 0.03056f
C4887 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.26707f
C4888 a_3369_24181# sar9b_0.clk_div_0.COUNT\[1\] 0.0204f
C4889 sar9b_0.net1 a_10707_23470# 0.25386f
C4890 sar9b_0.net35 sar9b_0.clk_div_0.COUNT\[2\] 0.02371f
C4891 a_10895_22855# sar9b_0.net11 0.04486f
C4892 single_9b_cdac_0.SW[4] a_44418_26990# 0.18991f
C4893 a_9546_24506# a_10506_24506# 0.03504f
C4894 a_10816_21487# a_10218_21842# 0.06623f
C4895 a_9442_21474# a_9647_21523# 0.09983f
C4896 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[1] 17.5055f
C4897 VDPWR a_12435_24802# 0.45648f
C4898 a_13011_23238# sar9b_0.net27 0.04162f
C4899 a_3014_24136# a_3521_24240# 0.21226f
C4900 sar9b_0.net70 a_3262_24141# 0.13578f
C4901 a_9996_16784# sar9b_0.net36 0.27514f
C4902 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 1.56037f
C4903 a_7289_21127# a_6834_20780# 0.3578f
C4904 sar9b_0.net57 sar9b_0.net37 0.18597f
C4905 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_60565_29911# 0.01076f
C4906 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 ua[0] 0.12344f
C4907 VDPWR a_6282_27170# 0.35695f
C4908 a_25915_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.01076f
C4909 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[5] 0.11961f
C4910 a_15151_10456# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.09051f
C4911 VDPWR tdc_0.phase_detector_0.pd_out_0.B 1.26944f
C4912 sar9b_0.net41 clk 0.05496f
C4913 sar9b_0.clknet_1_0__leaf_CLK a_3027_21906# 0.01945f
C4914 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4915 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.10429f
C4916 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] 1.15121f
C4917 a_7404_16784# sar9b_0.net27 0.02142f
C4918 a_7188_22119# a_6879_22145# 0.07766f
C4919 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[6] 0.363f
C4920 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[3] 0.05403f
C4921 sar9b_0.net70 sar9b_0.net66 0.02815f
C4922 sar9b_0._08_ a_5196_19448# 0.06291f
C4923 a_11178_20806# sar9b_0.net39 0.01531f
C4924 a_6137_23791# sar9b_0.net57 0.07535f
C4925 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C4926 VDPWR a_10762_18823# 0.20297f
C4927 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C4928 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.26427f
C4929 th_dif_sw_0.CK sar9b_0.net27 0.02592f
C4930 sar9b_0.net43 a_5748_24381# 0.02206f
C4931 a_4467_24162# sar9b_0.net58 0.09475f
C4932 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[8] 0.36652f
C4933 th_dif_sw_0.CK a_11658_18142# 0.06562f
C4934 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C4935 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.3196f
C4936 sar9b_0.net13 a_5748_24381# 0.24967f
C4937 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] 0.12898f
C4938 a_8554_26437# a_8340_26115# 0.04522f
C4939 VDPWR a_13011_24570# 0.48259f
C4940 single_9b_cdac_1.CF[3] sar9b_0.net29 0.47519f
C4941 sar9b_0.net29 sar9b_0.net28 1.82558f
C4942 sar9b_0.net41 sar9b_0.net56 0.06968f
C4943 VDPWR a_3695_23038# 0.22559f
C4944 VDPWR a_5289_22527# 0.14221f
C4945 single_9b_cdac_1.SW[6] clk 0.08446f
C4946 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.06503f
C4947 a_7602_18116# a_7404_18116# 0.06623f
C4948 sar9b_0.net63 sar9b_0.net35 0.03292f
C4949 sar9b_0.net60 sar9b_0.clknet_0_CLK 0.01871f
C4950 single_9b_cdac_1.cdac_sw_9b_0.S[2] a_54032_17740# 0.22367f
C4951 a_10506_23174# sar9b_0.net74 0.05564f
C4952 a_24332_26999# VDPWR 1.81495f
C4953 a_18214_3039# ua[3] 0.12559f
C4954 sar9b_0.net36 sar9b_0.net11 0.02201f
C4955 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C4956 single_9b_cdac_0.cdac_sw_9b_0.S[4] a_44418_26990# 0.22513f
C4957 tdc_0.OUTP th_dif_sw_0.CK 0.05462f
C4958 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[3] 0.01573f
C4959 a_6954_27466# a_7138_27758# 0.44532f
C4960 a_11430_27595# a_11178_27466# 0.27388f
C4961 sar9b_0._18_ a_4812_21738# 0.01257f
C4962 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.22875f
C4963 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.22497f
C4964 a_8726_22954# sar9b_0.net11 0.06796f
C4965 a_55773_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C4966 a_7926_23234# sar9b_0.net54 0.22246f
C4967 VDPWR dw_17224_1400# 1.89831f
C4968 single_9b_cdac_1.SW[1] sar9b_0.net27 0.17807f
C4969 sar9b_0.net31 sar9b_0.net74 0.23142f
C4970 sar9b_0.net9 sar9b_0.net42 0.01827f
C4971 a_5581_20992# sar9b_0._09_ 0.10212f
C4972 a_10742_21091# a_10607_21189# 0.35559f
C4973 a_4365_25770# a_4293_25852# 0.22517f
C4974 a_10218_27466# sar9b_0.net59 0.16798f
C4975 a_5298_24499# a_5748_24381# 0.03432f
C4976 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[0] 0.02174f
C4977 a_7743_18149# sar9b_0.net5 0.0249f
C4978 clk tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.09625f
C4979 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.45521f
C4980 a_8057_17131# sar9b_0.net5 0.05766f
C4981 VDPWR a_7638_19238# 0.30428f
C4982 a_7338_24802# a_6902_25087# 0.16939f
C4983 sar9b_0.net24 sar9b_0.net38 0.18f
C4984 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4985 sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# 0.24895f
C4986 a_4136_25584# a_4698_25851# 0.05308f
C4987 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[0\] 0.02059f
C4988 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.45521f
C4989 sar9b_0.net42 sar9b_0.net10 0.04131f
C4990 sar9b_0.net42 sar9b_0.net61 0.08366f
C4991 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36446f
C4992 single_9b_cdac_0.SW[8] uo_out[2] 0.10257f
C4993 a_8340_26115# a_8940_27039# 0.0165f
C4994 th_dif_sw_0.CK th_dif_sw_0.th_sw_1.CKB 0.09539f
C4995 a_5748_24381# a_6132_23451# 0.15019f
C4996 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 0.19143f
C4997 VDPWR a_7566_21017# 0.26799f
C4998 a_7404_17715# a_8019_17910# 0.02256f
C4999 a_4210_22378# sar9b_0.clknet_1_1__leaf_CLK 0.09811f
C5000 single_9b_cdac_1.cdac_sw_9b_0.S[2] ua[0] 1.21558f
C5001 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C5002 a_6861_22828# sar9b_0.clk_div_0.COUNT\[1\] 0.05496f
C5003 tdc_0.OUTP single_9b_cdac_1.SW[1] 0.10358f
C5004 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.02149f
C5005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A a_30717_15495# 0.01076f
C5006 sar9b_0.net40 single_9b_cdac_1.SW[4] 0.1589f
C5007 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] 3.10215f
C5008 VDPWR single_9b_cdac_1.CF[5] 2.58659f
C5009 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.36512f
C5010 VDPWR single_9b_cdac_0.SW[4] 2.61739f
C5011 a_10227_23490# sar9b_0.net53 0.38452f
C5012 sar9b_0.net60 sar9b_0.net21 0.08339f
C5013 sar9b_0.net38 a_10623_25895# 0.02019f
C5014 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.SW[4] 0.22983f
C5015 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.11216f
C5016 a_9930_20510# a_10528_20155# 0.06623f
C5017 sar9b_0.net43 sar9b_0.net39 0.08882f
C5018 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C5019 a_8438_18958# a_7914_19178# 0.04522f
C5020 a_4947_20140# a_5633_20244# 0.27693f
C5021 a_5126_20140# a_5374_20145# 0.05308f
C5022 a_6636_20780# sar9b_0.net10 0.29165f
C5023 sar9b_0.net52 clk 0.01379f
C5024 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.19147f
C5025 VDPWR a_13216_18477# 0.21525f
C5026 a_8166_27595# sar9b_0.net60 0.17093f
C5027 a_8694_20570# a_9154_20142# 0.26257f
C5028 a_8970_20510# a_9359_20191# 0.05462f
C5029 th_dif_sw_0.CKB tdc_0.RDY 0.6441f
C5030 VDPWR a_2835_24136# 0.52652f
C5031 sar9b_0.net36 sar9b_0.net45 0.56715f
C5032 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.12358f
C5033 a_10378_27170# a_9588_27045# 0.1263f
C5034 a_10926_17021# a_11434_16874# 0.19065f
C5035 sar9b_0.net35 sar9b_0.net55 0.02784f
C5036 sar9b_0.net29 a_13011_24570# 0.02017f
C5037 a_5938_22378# a_5739_22488# 0.29821f
C5038 a_3219_22860# sar9b_0._07_ 0.20806f
C5039 single_9b_cdac_1.CF[3] single_9b_cdac_0.SW[3] 1.96064f
C5040 sar9b_0.net28 single_9b_cdac_0.SW[3] 0.05131f
C5041 VDPWR a_9359_20191# 0.26316f
C5042 sar9b_0.net49 sar9b_0.net61 0.13664f
C5043 sar9b_0.net49 a_10402_21098# 0.10002f
C5044 sar9b_0.net7 sar9b_0.net42 0.12319f
C5045 a_6744_23238# sar9b_0.clk_div_0.COUNT\[2\] 0.03621f
C5046 a_11776_25137# sar9b_0.net12 0.07772f
C5047 sar9b_0.net25 uo_out[1] 0.06669f
C5048 a_6834_20780# sar9b_0.net47 0.26333f
C5049 sar9b_0.net8 a_9942_20810# 0.03985f
C5050 sar9b_0._11_ sar9b_0.net4 0.03423f
C5051 a_10607_25185# sar9b_0.net36 0.02216f
C5052 sar9b_0.net40 sar9b_0.net15 0.04777f
C5053 single_9b_cdac_0.SW[0] a_62748_26999# 0.28324f
C5054 sar9b_0.net27 a_12618_26134# 0.03607f
C5055 sar9b_0.net1 a_9359_20191# 0.01823f
C5056 sar9b_0.net47 a_7443_21496# 0.31185f
C5057 a_30012_17740# single_9b_cdac_1.SW[7] 0.18991f
C5058 a_8595_17910# single_9b_cdac_1.SW[2] 0.09011f
C5059 sar9b_0.net15 sar9b_0.net51 0.14145f
C5060 sar9b_0.net43 a_10895_22855# 0.02011f
C5061 a_9996_16784# a_9450_17846# 0.0165f
C5062 a_10528_20155# sar9b_0.net5 0.02721f
C5063 a_6252_20780# sar9b_0._01_ 0.14179f
C5064 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.38397f
C5065 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.75849f
C5066 VDPWR a_2508_20780# 1.55529f
C5067 a_7890_26108# a_8345_26455# 0.3578f
C5068 a_5298_24499# sar9b_0.net39 0.01755f
C5069 sar9b_0.net36 a_9870_27060# 0.04885f
C5070 VDPWR w_12795_1601# 0.45037f
C5071 single_9b_cdac_0.cdac_sw_9b_0.S[0] th_dif_sw_0.VCN 0.21769p
C5072 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[7] 0.21737f
C5073 a_18214_3039# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.33121f
C5074 a_3231_27227# a_3545_26914# 0.07826f
C5075 sar9b_0.net4 a_5811_19178# 0.07105f
C5076 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[4] 4.15222f
C5077 a_2892_27039# a_3090_27163# 0.06623f
C5078 VDPWR a_8386_22806# 0.24182f
C5079 sar9b_0.net63 sar9b_0._16_ 0.23068f
C5080 a_7193_22459# a_7402_22441# 0.24088f
C5081 sar9b_0.net60 a_5460_28377# 0.02635f
C5082 a_3603_28156# sar9b_0.net18 0.02874f
C5083 sar9b_0.net24 VDPWR 0.56782f
C5084 a_9130_26198# sar9b_0.cyclic_flag_0.FINAL 0.05175f
C5085 sar9b_0.net7 sar9b_0.net49 0.47708f
C5086 a_7882_19538# sar9b_0.net40 0.04062f
C5087 a_9900_19047# sar9b_0.net48 0.04064f
C5088 sar9b_0.net2 sar9b_0.net38 0.03026f
C5089 single_9b_cdac_0.SW[2] th_dif_sw_0.VCN 0.09453f
C5090 sar9b_0.net49 a_9442_21474# 0.10581f
C5091 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[7] 0.03585f
C5092 single_9b_cdac_1.SW[4] a_13011_17910# 0.07172f
C5093 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[2] 16.7662f
C5094 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.62443f
C5095 a_11466_23174# clk 0.02108f
C5096 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 2.82172f
C5097 a_7882_19538# sar9b_0.net51 0.01799f
C5098 sar9b_0._07_ sar9b_0.net46 0.15475f
C5099 VDPWR a_11859_17910# 0.40675f
C5100 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.28033f
C5101 single_9b_cdac_1.CF[5] sar9b_0.net29 0.09978f
C5102 single_9b_cdac_0.SW[4] sar9b_0.net29 0.07482f
C5103 sar9b_0.net63 a_6744_23238# 0.07362f
C5104 sar9b_0.net13 a_6902_25087# 0.05284f
C5105 sar9b_0.net26 single_9b_cdac_1.SW[1] 0.02116f
C5106 a_8098_18810# a_8874_19178# 0.3578f
C5107 sar9b_0.net60 a_5962_24151# 0.02401f
C5108 sar9b_0.net40 a_12618_19474# 0.06297f
C5109 VDPWR a_4771_18260# 0.42657f
C5110 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.28813f
C5111 a_11658_19474# a_12047_19857# 0.06034f
C5112 a_11842_19766# a_12618_19474# 0.3578f
C5113 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C5114 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C5115 sar9b_0.net67 sar9b_0.clknet_0_CLK 0.0173f
C5116 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[8] 0.24288f
C5117 a_10858_17113# a_10649_17131# 0.24088f
C5118 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07579f
C5119 VDPWR a_10623_25895# 0.25685f
C5120 a_4125_25958# sar9b_0.net39 0.02409f
C5121 sar9b_0._08_ sar9b_0.net46 0.2868f
C5122 VDPWR a_3370_27769# 0.20008f
C5123 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.28813f
C5124 single_9b_cdac_1.CF[0] th_dif_sw_0.VCN 0.09453f
C5125 sar9b_0.net58 sar9b_0.net19 0.19557f
C5126 a_6252_20780# sar9b_0.net60 0.02523f
C5127 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.19266f
C5128 sar9b_0.net3 ui_in[0] 0.05952f
C5129 sar9b_0.net43 sar9b_0.net36 0.11895f
C5130 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 3.27824f
C5131 single_9b_cdac_1.SW[8] a_13216_19809# 0.01788f
C5132 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.3196f
C5133 single_9b_cdac_1.SW[3] a_49221_17740# 0.18991f
C5134 a_5753_24250# a_5962_24151# 0.24088f
C5135 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.62443f
C5136 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] 3.10226f
C5137 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C5138 a_8595_17910# sar9b_0.net61 0.0485f
C5139 a_9546_24506# sar9b_0.net53 0.19966f
C5140 sar9b_0.clk_div_0.COUNT\[2\] a_2508_23444# 0.03301f
C5141 sar9b_0._16_ sar9b_0.clknet_1_1__leaf_CLK 0.07072f
C5142 sar9b_0.net13 sar9b_0.net36 0.024f
C5143 sar9b_0._18_ sar9b_0.net65 0.08636f
C5144 a_11030_22954# a_11466_23174# 0.16939f
C5145 sar9b_0.net4 sar9b_0.net39 0.0209f
C5146 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] 1.15113f
C5147 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] 1.56115f
C5148 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26218f
C5149 sar9b_0._15_ sar9b_0.net39 0.09291f
C5150 sar9b_0.net56 a_8052_18123# 0.21417f
C5151 sar9b_0.net35 sar9b_0.net6 0.53411f
C5152 single_9b_cdac_0.SW[6] uo_out[1] 0.04587f
C5153 a_4211_19474# sar9b_0.net46 0.02075f
C5154 single_9b_cdac_0.SW[7] uo_out[2] 0.69613f
C5155 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.12367f
C5156 VDPWR a_3161_26455# 0.25277f
C5157 a_5439_24563# a_5753_24250# 0.07826f
C5158 th_dif_sw_0.VCN single_9b_cdac_1.SW[2] 0.09468f
C5159 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net39 0.06168f
C5160 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[1\] 0.01596f
C5161 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.42014f
C5162 sar9b_0.net2 sar9b_0.net6 0.19883f
C5163 single_9b_cdac_1.SW[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.24456f
C5164 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.19147f
C5165 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 a_34814_26990# 0.14695f
C5166 a_16527_10454# tdc_0.phase_detector_0.INN 0.10585f
C5167 sar9b_0.net53 a_11382_22142# 0.2367f
C5168 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[0] 0.0313f
C5169 a_5235_27466# a_5322_27170# 0.01145f
C5170 sar9b_0.net19 sar9b_0.net37 0.21509f
C5171 a_7602_16784# sar9b_0.net46 0.25599f
C5172 a_10662_17799# sar9b_0.net36 0.03369f
C5173 sar9b_0.net60 a_6534_27123# 0.01098f
C5174 a_7882_19538# sar9b_0.net62 0.20424f
C5175 sar9b_0.net73 a_6634_18206# 0.17082f
C5176 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A a_64331_15495# 0.01076f
C5177 sar9b_0.net40 a_12182_19759# 0.06762f
C5178 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.84059f
C5179 a_11842_19766# a_12182_19759# 0.24088f
C5180 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.42014f
C5181 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 2.71729f
C5182 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07517f
C5183 sar9b_0.net32 a_11915_28371# 0.04795f
C5184 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.0313f
C5185 a_9414_23127# clk 0.01589f
C5186 sar9b_0.net20 a_5742_28392# 0.07038f
C5187 VDPWR a_4210_22378# 0.37875f
C5188 a_7539_28566# uo_out[6] 0.08058f
C5189 sar9b_0.net58 a_3161_27787# 0.10647f
C5190 sar9b_0.net52 a_11214_25728# 0.27195f
C5191 sar9b_0.net31 a_12182_22423# 0.02073f
C5192 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.10429f
C5193 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.81428f
C5194 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C5195 VDPWR sar9b_0.net35 1.86196f
C5196 th_dif_sw_0.CK a_12047_18525# 0.04966f
C5197 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07517f
C5198 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.23119f
C5199 VDPWR sar9b_0.net16 1.35456f
C5200 sar9b_0.net13 a_10937_25582# 0.03829f
C5201 a_2706_27440# a_3161_27787# 0.3578f
C5202 a_11146_25483# a_11214_25728# 0.35559f
C5203 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A a_54737_29917# 0.01076f
C5204 a_12870_19603# single_9b_cdac_1.SW[8] 0.01567f
C5205 VDPWR a_12064_22819# 0.1986f
C5206 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] 0.17948f
C5207 a_10378_27170# sar9b_0.net42 0.16789f
C5208 a_16331_9671# th_dif_sw_0.VCN 0.0647f
C5209 sar9b_0.net56 a_7284_20787# 0.21387f
C5210 uio_in[6] uio_in[5] 0.03102f
C5211 sar9b_0.net13 a_11722_25838# 0.05888f
C5212 sar9b_0.net5 sar9b_0.net73 1.10057f
C5213 VDPWR sar9b_0.net2 1.0982f
C5214 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[3] 0.02002f
C5215 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.3196f
C5216 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[7] 0.02149f
C5217 single_9b_cdac_0.SW[4] single_9b_cdac_0.SW[3] 12.7151f
C5218 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[7] 0.31534f
C5219 single_9b_cdac_1.SW[8] th_dif_sw_0.VCN 0.09453f
C5220 sar9b_0.net35 sar9b_0.net1 0.20023f
C5221 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31753_15501# 0.01076f
C5222 sar9b_0.net10 sar9b_0.net11 0.2401f
C5223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[7] 0.0313f
C5224 a_10926_17021# sar9b_0.net48 0.19705f
C5225 a_5748_24381# sar9b_0.net55 0.0128f
C5226 VDPWR tdc_0.OUTN 0.62093f
C5227 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.3186f
C5228 sar9b_0.net41 sar9b_0.net40 0.06786f
C5229 sar9b_0.net38 a_10218_20806# 0.01292f
C5230 a_5938_22378# sar9b_0.net60 0.01049f
C5231 VDPWR a_13216_22473# 0.20771f
C5232 a_6250_28502# a_5742_28392# 0.19065f
C5233 sar9b_0.net48 a_6634_18206# 0.28205f
C5234 sar9b_0.net59 a_2847_26141# 0.17414f
C5235 VDPWR a_11915_27039# 0.44729f
C5236 sar9b_0.net41 sar9b_0.net51 0.02663f
C5237 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.26707f
C5238 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0303f
C5239 sar9b_0.net63 sar9b_0.net39 0.2717f
C5240 a_6307_27584# sar9b_0.net45 0.3888f
C5241 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C5242 a_12491_27662# single_9b_cdac_0.SW[2] 0.03543f
C5243 sar9b_0.net1 tdc_0.OUTN 0.04134f
C5244 sar9b_0.net40 a_6879_22145# 0.02015f
C5245 sar9b_0.net49 a_10607_21189# 0.22001f
C5246 VDPWR sar9b_0._06_ 0.47072f
C5247 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C5248 a_53154_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.23864f
C5249 VDPWR a_13216_23805# 0.20771f
C5250 a_11430_24931# a_11776_25137# 0.07649f
C5251 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 1.55978f
C5252 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.17533f
C5253 th_dif_sw_0.CK th_dif_sw_0.VCP 0.0144f
C5254 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.84426f
C5255 VDPWR a_3723_20140# 0.08905f
C5256 sar9b_0.net55 a_5811_19178# 0.26511f
C5257 single_9b_cdac_0.SW[5] sar9b_0.net25 0.1111f
C5258 VDPWR a_10758_24459# 0.26555f
C5259 a_4332_23043# sar9b_0.clk_div_0.COUNT\[2\] 0.1269f
C5260 sar9b_0.net48 sar9b_0.net5 0.3854f
C5261 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.11216f
C5262 a_5506_26802# a_6534_27123# 0.07826f
C5263 a_3946_26198# sar9b_0.net59 0.24509f
C5264 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.01175f
C5265 VDPWR a_7914_27466# 0.35464f
C5266 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.03484f
C5267 a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK 1.86751f
C5268 a_9130_26198# sar9b_0.net41 0.17586f
C5269 a_2508_26108# a_2706_26108# 0.06623f
C5270 single_9b_cdac_1.SW[5] ua[0] 0.13353f
C5271 a_4922_20857# sar9b_0._18_ 0.14576f
C5272 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26427f
C5273 sar9b_0.net72 sar9b_0.clk_div_0.COUNT\[2\] 0.29657f
C5274 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C5275 sar9b_0.net52 a_11658_26134# 0.18819f
C5276 a_10553_18922# sar9b_0.net26 0.13039f
C5277 a_5581_20992# a_5761_21100# 0.01239f
C5278 a_7914_23470# a_9126_23599# 0.07766f
C5279 a_9930_20510# a_9154_20142# 0.3578f
C5280 a_4812_28371# uo_out[7] 0.0141f
C5281 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.07579f
C5282 VDPWR a_5523_21528# 0.22726f
C5283 a_5235_27466# a_4749_27652# 0.13237f
C5284 sar9b_0._07_ sar9b_0.clknet_0_CLK 0.16508f
C5285 sar9b_0.net39 sar9b_0.clknet_1_1__leaf_CLK 0.01422f
C5286 a_7097_19795# sar9b_0.net47 0.13999f
C5287 a_5126_20140# a_6130_20239# 0.06302f
C5288 a_10402_21098# a_11178_20806# 0.3578f
C5289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5290 sar9b_0.net46 sar9b_0.net5 1.36216f
C5291 a_3438_26345# a_3156_26115# 0.05462f
C5292 a_3370_26437# a_2706_26108# 0.16939f
C5293 sar9b_0._09_ a_5481_20185# 0.02188f
C5294 sar9b_0.net50 sar9b_0.net5 0.49397f
C5295 a_10830_19068# a_10762_18823# 0.35559f
C5296 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C5297 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[1] 0.01285f
C5298 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_15265_9613# 0.16728f
C5299 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] 1.17995f
C5300 sar9b_0.net41 a_13011_17910# 0.2244f
C5301 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.05472f
C5302 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 a_63626_17740# 0.14695f
C5303 sar9b_0.net55 sar9b_0.net39 0.04945f
C5304 sar9b_0.net70 sar9b_0._05_ 0.12818f
C5305 a_6137_23791# a_6346_23773# 0.24088f
C5306 a_10402_27758# sar9b_0.net38 0.02612f
C5307 VDPWR a_8554_26437# 0.21407f
C5308 sar9b_0.net32 sar9b_0.net52 0.06191f
C5309 a_3371_23106# sar9b_0.clk_div_0.COUNT\[1\] 0.10763f
C5310 sar9b_0.net29 a_13216_22473# 0.01568f
C5311 sar9b_0.net5 a_9154_20142# 0.01312f
C5312 VDPWR single_9b_cdac_1.CF[6] 2.73682f
C5313 VDPWR a_7914_23470# 0.85718f
C5314 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.03488f
C5315 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.SW[4] 0.1516f
C5316 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.06503f
C5317 VDPWR a_10218_20806# 0.83839f
C5318 VDPWR a_5465_28246# 0.21298f
C5319 VDPWR a_3946_27530# 0.29317f
C5320 a_4934_22432# a_5938_22378# 0.06302f
C5321 sar9b_0.clknet_1_0__leaf_CLK sar9b_0.clknet_0_CLK 0.03854f
C5322 VDPWR sar9b_0._16_ 0.84748f
C5323 sar9b_0.net41 a_9647_21523# 0.0288f
C5324 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.01472f
C5325 a_6642_19448# a_7097_19795# 0.3578f
C5326 sar9b_0._14_ sar9b_0._16_ 0.12248f
C5327 sar9b_0.net59 single_9b_cdac_0.SW[5] 0.02001f
C5328 a_6130_20239# sar9b_0.net4 0.03123f
C5329 sar9b_0.net63 sar9b_0.net72 0.26712f
C5330 a_10548_19053# sar9b_0.net39 0.01144f
C5331 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP a_24332_16877# 0.04592f
C5332 sar9b_0._06_ sar9b_0.net29 0.03732f
C5333 a_4755_22138# sar9b_0.net39 0.1069f
C5334 a_4125_25958# a_4136_25584# 0.54361f
C5335 sar9b_0.net29 a_13216_23805# 0.01558f
C5336 a_9730_24138# a_10070_24286# 0.24088f
C5337 sar9b_0.net7 a_11178_20806# 0.04419f
C5338 a_10218_21842# a_10218_20806# 0.01915f
C5339 a_10662_17799# a_9450_17846# 0.07766f
C5340 VDPWR a_7343_27849# 0.26147f
C5341 a_10662_17799# single_9b_cdac_1.SW[2] 0.03662f
C5342 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.45521f
C5343 sar9b_0.net2 a_9270_24566# 0.03939f
C5344 a_3819_24136# a_3521_24240# 0.02614f
C5345 VDPWR a_6744_23238# 0.16029f
C5346 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.19129f
C5347 a_13011_17910# single_9b_cdac_1.SW[6] 0.35507f
C5348 sar9b_0.net70 sar9b_0.clknet_1_1__leaf_CLK 0.27895f
C5349 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.12431f
C5350 a_13011_19242# single_9b_cdac_1.SW[8] 0.01098f
C5351 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[5] 8.69008f
C5352 sar9b_0.net38 sar9b_0.net39 0.02578f
C5353 a_7602_18116# a_8057_18463# 0.3578f
C5354 a_12064_22819# a_11658_22138# 0.0165f
C5355 a_5535_18149# a_5849_18463# 0.07826f
C5356 a_5844_18123# a_6058_18445# 0.04522f
C5357 a_21684_3438# a_18214_3039# 0.11186f
C5358 VDPWR sar9b_0._11_ 0.2748f
C5359 VDPWR a_8940_27039# 0.24411f
C5360 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C5361 VDPWR a_5748_24381# 0.75977f
C5362 sar9b_0.net43 sar9b_0.net9 0.0248f
C5363 VDPWR a_2603_17006# 0.51948f
C5364 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.25152f
C5365 a_9588_27045# a_9593_26914# 0.44532f
C5366 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_65367_15501# 0.01076f
C5367 sar9b_0.net67 a_3027_22138# 0.0723f
C5368 VDPWR a_11658_23470# 0.84308f
C5369 sar9b_0.net56 a_9634_17478# 0.02665f
C5370 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.03729f
C5371 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07579f
C5372 VDPWR a_8982_21902# 0.33673f
C5373 single_9b_cdac_1.cdac_sw_9b_0.S[7] a_29134_16877# 0.59531f
C5374 sar9b_0.net67 sar9b_0.net65 0.11461f
C5375 sar9b_0.net43 sar9b_0.net10 0.02603f
C5376 sar9b_0.net44 a_3545_26914# 0.05842f
C5377 a_11382_22142# a_12047_22521# 0.19065f
C5378 a_11842_22430# a_12870_22267# 0.07826f
C5379 a_9939_28566# a_9323_28371# 0.03551f
C5380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.01175f
C5381 sar9b_0.net72 sar9b_0.clknet_1_1__leaf_CLK 0.02825f
C5382 VDPWR a_16222_11316# 0.52162f
C5383 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.08121f
C5384 sar9b_0.net58 a_5151_28559# 0.19397f
C5385 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 1.50841f
C5386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.84427f
C5387 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[5] 4.15352f
C5388 VDPWR a_5374_20145# 0.01375f
C5389 a_10035_19474# sar9b_0.net48 0.35551f
C5390 a_9647_21523# a_9782_21622# 0.35559f
C5391 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C5392 a_8982_21902# sar9b_0.net1 0.01917f
C5393 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C5394 a_53154_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.23864f
C5395 VDPWR a_5811_19178# 0.21566f
C5396 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[6] 17.8424f
C5397 sar9b_0.net47 a_5581_19664# 0.07464f
C5398 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.01751f
C5399 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.CF[0] 0.10499f
C5400 VDPWR a_6880_26815# 0.20981f
C5401 sar9b_0.net43 a_6538_24506# 0.03826f
C5402 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.SW[8] 0.15864f
C5403 a_7092_19455# sar9b_0.net40 0.0376f
C5404 sar9b_0.net52 sar9b_0.net62 0.03789f
C5405 a_9132_7271# th_dif_sw_0.th_sw_1.CK 2.28032f
C5406 sar9b_0.net47 a_7402_22441# 0.15391f
C5407 a_7092_19455# sar9b_0.net51 0.02272f
C5408 single_9b_cdac_1.CF[6] sar9b_0.net29 0.19274f
C5409 a_10402_27758# VDPWR 0.22246f
C5410 sar9b_0.net13 a_6538_24506# 0.03555f
C5411 a_7602_16784# sar9b_0.net27 0.05862f
C5412 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.81423f
C5413 sar9b_0.net6 sar9b_0.net39 0.02562f
C5414 a_10662_17799# sar9b_0.net61 0.05961f
C5415 sar9b_0.net58 sar9b_0.net68 0.02945f
C5416 a_11842_23762# a_12870_23599# 0.07826f
C5417 a_6346_23773# sar9b_0.net57 0.03377f
C5418 VDPWR a_33936_16877# 1.81495f
C5419 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[5] 0.31534f
C5420 sar9b_0._06_ single_9b_cdac_0.SW[3] 0.08528f
C5421 sar9b_0.net23 sar9b_0.net24 0.18313f
C5422 a_3166_20145# a_3273_20185# 0.14439f
C5423 sar9b_0.net43 sar9b_0.net7 0.59584f
C5424 th_dif_sw_0.CK a_11842_18434# 0.11252f
C5425 single_9b_cdac_0.SW[8] clk 0.42402f
C5426 a_7289_21127# a_7566_21017# 0.09983f
C5427 VDPWR a_2508_23444# 1.56828f
C5428 a_8874_19178# sar9b_0.net61 0.01101f
C5429 th_dif_sw_0.CK a_10166_3438# 0.0136f
C5430 sar9b_0.net8 sar9b_0.net73 0.02045f
C5431 sar9b_0.net40 a_6102_24806# 0.01823f
C5432 VDPWR a_6540_22112# 0.20318f
C5433 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.SW[8] 0.1495f
C5434 sar9b_0.net16 a_4072_19474# 0.04195f
C5435 sar9b_0.net16 sar9b_0.net71 0.48375f
C5436 a_6954_27466# sar9b_0.net21 0.03499f
C5437 sar9b_0.net35 a_7193_22459# 0.01725f
C5438 a_6880_17491# sar9b_0.net5 0.27459f
C5439 clk ena 0.03102f
C5440 VDPWR sar9b_0.net39 1.30812f
C5441 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 3.10626f
C5442 VDPWR single_9b_cdac_1.CF[7] 2.59279f
C5443 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.03433f
C5444 a_11718_23127# sar9b_0.net10 0.07252f
C5445 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.36044f
C5446 a_6954_27466# a_8166_27595# 0.07766f
C5447 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.CF[3] 0.105f
C5448 sar9b_0.net58 a_6282_27170# 0.26031f
C5449 sar9b_0.net36 sar9b_0.net38 0.92018f
C5450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 ua[0] 0.11944f
C5451 a_11178_27466# a_11776_27801# 0.06623f
C5452 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[8] 0.363f
C5453 single_9b_cdac_0.cdac_sw_9b_0.S[7] a_30012_26990# 0.22513f
C5454 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22497f
C5455 sar9b_0.net1 sar9b_0.net39 0.02611f
C5456 a_10227_23490# clk 0.01166f
C5457 a_7284_20787# sar9b_0.net51 0.07994f
C5458 sar9b_0.net6 a_12435_20806# 0.19538f
C5459 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] 0.17948f
C5460 a_7092_19455# sar9b_0.net62 0.03046f
C5461 a_11008_17491# a_10410_17846# 0.06623f
C5462 a_11339_27039# single_9b_cdac_0.SW[4] 0.03465f
C5463 VDPWR a_8098_18810# 0.26718f
C5464 a_6767_25185# a_6562_25094# 0.09983f
C5465 a_7936_25137# a_7590_24931# 0.07649f
C5466 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0._02_ 0.06001f
C5467 a_4136_25584# sar9b_0.clknet_1_1__leaf_CLK 0.10289f
C5468 sar9b_0._07_ a_5443_19074# 0.02952f
C5469 sar9b_0.net42 a_11430_20935# 0.01027f
C5470 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 a_25210_26990# 0.14695f
C5471 a_10378_27170# sar9b_0.net45 0.05318f
C5472 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.02632f
C5473 VDPWR a_8074_20870# 0.30584f
C5474 a_3369_24181# a_2835_24136# 0.35097f
C5475 a_11658_26134# a_12182_26419# 0.05022f
C5476 a_10218_27466# sar9b_0.net34 0.05477f
C5477 a_13011_16810# sar9b_0.net40 0.21779f
C5478 a_10926_17021# sar9b_0.net27 0.03167f
C5479 VDPWR a_10895_22855# 0.26689f
C5480 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[3] 0.02012f
C5481 a_6282_27170# sar9b_0.net37 0.06133f
C5482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.12358f
C5483 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.26707f
C5484 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[8] 1.41793f
C5485 VDPWR a_12435_20806# 0.43957f
C5486 single_9b_cdac_1.CF[2] ua[0] 3.58697f
C5487 a_9900_19047# sar9b_0.net26 0.04584f
C5488 sar9b_0.net10 sar9b_0.clk_div_0.COUNT\[2\] 0.03438f
C5489 a_5126_20140# a_5481_20185# 0.18752f
C5490 single_9b_cdac_1.SW[4] th_dif_sw_0.VCN 0.09453f
C5491 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.45521f
C5492 VDPWR sar9b_0.net70 0.75523f
C5493 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.84042f
C5494 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[5] 0.06019f
C5495 sar9b_0.net41 sar9b_0.net49 0.52224f
C5496 sar9b_0.net36 sar9b_0.net6 0.05014f
C5497 a_10378_27170# a_9870_27060# 0.19065f
C5498 sar9b_0.net41 a_9162_23174# 0.01093f
C5499 a_10926_17021# tdc_0.OUTP 0.06343f
C5500 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22367f
C5501 th_dif_sw_0.CK th_dif_sw_0.CKB 0.08006f
C5502 sar9b_0.net27 sar9b_0.net5 0.07039f
C5503 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07517f
C5504 VDPWR a_6902_25087# 0.2038f
C5505 sar9b_0._18_ sar9b_0._17_ 0.19231f
C5506 a_8115_28566# sar9b_0.net22 0.0346f
C5507 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02666f
C5508 sar9b_0.net49 a_11430_20935# 0.17358f
C5509 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.62443f
C5510 sar9b_0.net26 sar9b_0.net12 0.02943f
C5511 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.10429f
C5512 sar9b_0.net8 sar9b_0.net50 0.34359f
C5513 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[6] 0.0313f
C5514 a_7284_20787# sar9b_0.net62 0.023f
C5515 sar9b_0._01_ sar9b_0._17_ 0.03752f
C5516 sar9b_0.net32 a_12182_26419# 0.01466f
C5517 a_6678_27470# a_7343_27849# 0.19065f
C5518 a_10762_18823# a_10098_19171# 0.16939f
C5519 VDPWR a_4332_23043# 1.38139f
C5520 a_8052_18123# a_7914_19178# 0.26288f
C5521 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.10499f
C5522 a_12618_19474# a_13216_19809# 0.06623f
C5523 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.SW[7] 0.22983f
C5524 a_10742_27751# single_9b_cdac_0.SW[7] 0.02243f
C5525 single_9b_cdac_1.CF[7] sar9b_0.net29 0.04004f
C5526 sar9b_0.net32 uo_out[3] 0.13894f
C5527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.10499f
C5528 a_13011_21906# single_9b_cdac_1.CF[2] 0.08337f
C5529 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.31534f
C5530 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.69086f
C5531 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.26942f
C5532 sar9b_0.net8 a_9154_20142# 0.01901f
C5533 VDPWR sar9b_0.net72 0.65198f
C5534 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.07852f
C5535 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.38397f
C5536 a_6414_23681# sar9b_0.net54 0.20382f
C5537 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.02632f
C5538 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C5539 VDPWR a_5581_20992# 0.1971f
C5540 sar9b_0.net72 sar9b_0._14_ 1.15565f
C5541 VDPWR sar9b_0.net36 1.87634f
C5542 sar9b_0.net6 a_5844_18123# 0.23512f
C5543 a_3822_27060# a_3754_26815# 0.35559f
C5544 a_10830_19068# sar9b_0.net2 0.018f
C5545 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 1.71649f
C5546 a_7743_18149# sar9b_0.net73 0.09002f
C5547 a_11915_28371# sar9b_0.net14 0.20706f
C5548 sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# 0.26938f
C5549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C5550 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.27833f
C5551 a_3540_27045# a_3822_27060# 0.06034f
C5552 a_4812_28371# a_5010_28495# 0.06623f
C5553 single_9b_cdac_1.SW[5] sar9b_0.net28 0.01641f
C5554 VDPWR a_8726_22954# 0.22795f
C5555 sar9b_0.net65 sar9b_0.clknet_1_0__leaf_CLK 0.03848f
C5556 a_3090_27163# a_3231_27227# 0.27388f
C5557 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP a_57946_16877# 0.04592f
C5558 a_7566_21017# sar9b_0.net47 0.24689f
C5559 sar9b_0.net63 sar9b_0.net10 0.04452f
C5560 sar9b_0.net1 sar9b_0.net36 0.01195f
C5561 a_13011_16810# a_13011_17910# 0.0246f
C5562 VDPWR tdc_0.phase_detector_0.INP 0.59622f
C5563 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.11216f
C5564 sar9b_0.net60 a_5742_28392# 0.06229f
C5565 sar9b_0._01_ a_5633_20244# 0.01113f
C5566 sar9b_0.net42 sar9b_0.net52 0.15052f
C5567 a_9802_26815# sar9b_0.net59 0.17205f
C5568 a_13011_23238# clk 0.0315f
C5569 sar9b_0.net49 a_9782_21622# 0.15031f
C5570 single_9b_cdac_1.cdac_sw_9b_0.S[3] ua[0] 1.59889f
C5571 single_9b_cdac_0.SW[7] clk 1.04996f
C5572 a_11146_25483# sar9b_0.net42 0.01506f
C5573 single_9b_cdac_0.SW[6] uo_out[2] 0.04371f
C5574 sar9b_0._04_ sar9b_0.net69 0.13306f
C5575 sar9b_0.net45 sar9b_0.cyclic_flag_0.FINAL 0.18011f
C5576 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] 0.17948f
C5577 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 1.55946f
C5578 a_8438_18958# a_8874_19178# 0.16939f
C5579 sar9b_0.net40 a_12047_19857# 0.04975f
C5580 sar9b_0.net60 sar9b_0._17_ 0.04099f
C5581 VDPWR a_5844_18123# 0.83758f
C5582 ui_in[3] ui_in[2] 0.03102f
C5583 a_9174_17906# a_9634_17478# 0.26257f
C5584 a_9450_17846# a_9839_17527# 0.05462f
C5585 sar9b_0.net67 a_3454_22567# 0.1221f
C5586 a_11842_19766# a_12047_19857# 0.09983f
C5587 a_12870_19603# a_12618_19474# 0.27388f
C5588 a_2931_28566# uio_out[1] 0.4065f
C5589 a_8202_23174# a_8386_22806# 0.43491f
C5590 single_9b_cdac_1.SW[2] a_9839_17527# 0.06063f
C5591 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38317f
C5592 sar9b_0.net56 a_9126_19131# 0.02432f
C5593 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.11216f
C5594 sar9b_0.net55 a_6444_21738# 0.02142f
C5595 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[5] 1.06635f
C5596 VDPWR a_10937_25582# 0.2119f
C5597 a_7743_18149# sar9b_0.net48 0.03022f
C5598 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26218f
C5599 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.42784f
C5600 a_5711_17527# sar9b_0.net56 0.06214f
C5601 VDPWR a_11722_25838# 0.30045f
C5602 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INN 0.06563f
C5603 th_dif_sw_0.th_sw_1.CK ua[4] 0.42268f
C5604 a_7289_21127# sar9b_0.net35 0.02113f
C5605 a_5739_22488# sar9b_0._12_ 0.0684f
C5606 a_6282_17846# sar9b_0.net46 0.32729f
C5607 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.0115f
C5608 a_8334_17021# sar9b_0.net6 0.03019f
C5609 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.37833f
C5610 VDPWR a_6130_20239# 0.38534f
C5611 sar9b_0.net64 a_5523_21528# 0.03232f
C5612 sar9b_0.net12 sar9b_0.net53 0.44449f
C5613 sar9b_0.net23 a_8554_26437# 0.01362f
C5614 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[3] 0.02029f
C5615 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.95338f
C5616 sar9b_0.net41 a_10227_18142# 0.01117f
C5617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.03484f
C5618 th_dif_sw_0.CK single_9b_cdac_1.SW[0] 0.05143f
C5619 a_3206_22432# sar9b_0.clknet_1_1__leaf_CLK 0.06142f
C5620 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5621 a_5748_24381# a_6030_24396# 0.06034f
C5622 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[0] 4.151f
C5623 a_7743_18149# sar9b_0.net46 0.17277f
C5624 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.06503f
C5625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[8] 0.01887f
C5626 VDPWR a_4136_25584# 0.84755f
C5627 a_8057_17131# sar9b_0.net46 0.08295f
C5628 a_11466_23174# sar9b_0.net42 0.01972f
C5629 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.22879f
C5630 sar9b_0.net26 sar9b_0.net5 0.02305f
C5631 single_9b_cdac_1.SW[1] clk 0.99126f
C5632 a_6286_22804# sar9b_0._02_ 0.01706f
C5633 a_4018_24235# sar9b_0.clk_div_0.COUNT\[2\] 0.15815f
C5634 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.SW[6] 0.22497f
C5635 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.27794f
C5636 a_4922_20857# sar9b_0._08_ 0.02439f
C5637 VDPWR single_9b_cdac_0.SW[2] 2.53031f
C5638 sar9b_0.net40 sar9b_0.net44 0.06639f
C5639 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.70254f
C5640 a_5010_28495# a_5674_28147# 0.16939f
C5641 sar9b_0.net58 a_3370_27769# 0.14413f
C5642 sar9b_0.net31 a_12618_22138# 0.06744f
C5643 VDPWR a_8334_17021# 0.2535f
C5644 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.42509f
C5645 a_3747_25724# a_3855_25792# 0.29821f
C5646 a_8386_22806# sar9b_0.net37 0.03128f
C5647 sar9b_0.net55 a_6538_24506# 0.0859f
C5648 VDPWR a_7374_19685# 0.26931f
C5649 single_9b_cdac_0.SW[7] a_10607_27849# 0.02998f
C5650 a_10548_19053# sar9b_0.net61 0.01669f
C5651 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C5652 a_3156_27447# a_3438_27677# 0.05462f
C5653 a_10803_18142# th_dif_sw_0.CK 0.095f
C5654 a_2706_27440# a_3370_27769# 0.16939f
C5655 a_2547_28132# sar9b_0.net60 0.23163f
C5656 sar9b_0.net17 a_2931_28566# 0.22067f
C5657 sar9b_0.net24 sar9b_0.net37 0.25988f
C5658 sar9b_0.net61 a_9839_17527# 0.01999f
C5659 a_16357_9613# th_dif_sw_0.VCN 0.10892f
C5660 sar9b_0.net41 sar9b_0.net11 0.07372f
C5661 sar9b_0.net13 a_13011_25902# 0.2478f
C5662 sar9b_0.net6 single_9b_cdac_1.SW[2] 0.15073f
C5663 single_9b_cdac_1.CF[4] ua[0] 3.57685f
C5664 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22543f
C5665 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.19143f
C5666 sar9b_0.net9 sar9b_0.net38 0.32278f
C5667 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[0] 19.2136f
C5668 a_10194_16784# a_10649_17131# 0.3578f
C5669 single_9b_cdac_1.CF[1] ua[0] 3.57763f
C5670 VDPWR a_8334_18353# 0.25378f
C5671 a_7638_23474# sar9b_0.net54 0.09716f
C5672 a_14897_9355# a_14871_9671# 0.06748f
C5673 sar9b_0.net56 a_5046_17906# 0.13749f
C5674 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.12898f
C5675 VDPWR single_9b_cdac_1.CF[0] 2.72978f
C5676 sar9b_0._12_ sar9b_0.net69 0.23206f
C5677 a_11434_16874# sar9b_0.net48 0.19635f
C5678 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[6] 0.42014f
C5679 sar9b_0.net13 sar9b_0.cyclic_flag_0.FINAL 0.03185f
C5680 sar9b_0.net10 sar9b_0.net38 0.02721f
C5681 sar9b_0.net38 a_10402_21098# 0.0282f
C5682 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[2] 0.07133f
C5683 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[2] 16.4998f
C5684 a_8334_18353# sar9b_0.net1 0.01172f
C5685 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.12431f
C5686 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[6] 0.02149f
C5687 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.19266f
C5688 sar9b_0.net68 sar9b_0.clk_div_0.COUNT\[1\] 0.35672f
C5689 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C5690 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.28523f
C5691 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5692 sar9b_0.net60 clk 0.04516f
C5693 a_7193_22459# sar9b_0.net39 0.17464f
C5694 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.22875f
C5695 sar9b_0.net31 sar9b_0.net27 0.03712f
C5696 a_12182_18427# sar9b_0.net6 0.02363f
C5697 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.04592f
C5698 sar9b_0.net54 a_5962_24151# 0.14491f
C5699 sar9b_0.net31 single_9b_cdac_0.SW[5] 0.01126f
C5700 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.62443f
C5701 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5702 VDPWR a_9450_17846# 0.85429f
C5703 sar9b_0.net3 sar9b_0.net19 0.0315f
C5704 VDPWR single_9b_cdac_1.SW[2] 2.86879f
C5705 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.17156f
C5706 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 3.10626f
C5707 a_10803_18142# single_9b_cdac_1.SW[1] 0.0113f
C5708 sar9b_0._18_ sar9b_0._12_ 0.02191f
C5709 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[4] 0.31534f
C5710 a_13011_21906# single_9b_cdac_1.CF[4] 0.35507f
C5711 sar9b_0.net55 a_6579_18832# 0.01696f
C5712 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[5] 1.95851f
C5713 sar9b_0.net6 single_9b_cdac_1.SW[8] 0.1227f
C5714 a_10548_19053# sar9b_0.net7 0.21355f
C5715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.02545f
C5716 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.36006f
C5717 single_9b_cdac_1.CF[8] ua[0] 5.00726f
C5718 sar9b_0.net35 sar9b_0.net58 0.03409f
C5719 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.24288f
C5720 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.SW[3] 0.14997f
C5721 a_5439_24563# sar9b_0.net54 0.16847f
C5722 a_9132_7271# th_dif_sw_0.th_sw_1.CKB 0.01594f
C5723 a_3156_26115# a_2847_26141# 0.07766f
C5724 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C5725 single_9b_cdac_1.cdac_sw_9b_0.S[7] th_dif_sw_0.VCP 1.61586f
C5726 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.B 0.38171f
C5727 VDPWR a_6307_27584# 0.36193f
C5728 a_8303_23853# sar9b_0.net54 0.0633f
C5729 sar9b_0.net52 a_11842_26426# 0.09411f
C5730 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[2] 0.01481f
C5731 sar9b_0.net52 a_10218_24802# 0.16549f
C5732 VDPWR a_12182_18427# 0.20217f
C5733 sar9b_0.net12 a_10932_25713# 0.01703f
C5734 sar9b_0.net7 sar9b_0.net38 0.02694f
C5735 a_9442_21474# sar9b_0.net38 0.01689f
C5736 single_9b_cdac_1.SW[6] th_dif_sw_0.VCN 0.09453f
C5737 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.10626f
C5738 a_9930_20510# a_9494_20290# 0.16939f
C5739 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL 0.2316f
C5740 single_9b_cdac_0.SW[2] sar9b_0.net29 0.33939f
C5741 sar9b_0.net20 uo_out[7] 0.0338f
C5742 VDPWR a_6444_21738# 0.29205f
C5743 a_6678_27470# sar9b_0.net36 0.05745f
C5744 sar9b_0.net47 sar9b_0.net35 0.11331f
C5745 VDPWR a_16331_9671# 0.67026f
C5746 VDPWR a_10482_3438# 0.07094f
C5747 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.SW[5] 0.22549f
C5748 sar9b_0.net61 sar9b_0.net6 0.4224f
C5749 sar9b_0.net39 sar9b_0._03_ 0.13967f
C5750 a_11430_20935# a_11178_20806# 0.27388f
C5751 sar9b_0.net8 sar9b_0.net27 0.0426f
C5752 VDPWR single_9b_cdac_1.SW[8] 2.60138f
C5753 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 ua[0] 0.12358f
C5754 a_3370_26437# a_3161_26455# 0.24088f
C5755 a_3946_26198# a_3156_26115# 0.1263f
C5756 sar9b_0.net35 sar9b_0.net37 0.35869f
C5757 sar9b_0.net4 a_5535_18149# 0.03052f
C5758 a_10553_18922# a_11338_19178# 0.26257f
C5759 a_10335_16817# sar9b_0.net48 0.17419f
C5760 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.CF[4] 0.01514f
C5761 a_11915_28371# uo_out[0] 0.38176f
C5762 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01175f
C5763 sar9b_0.net29 single_9b_cdac_1.CF[0] 0.10817f
C5764 sar9b_0.net2 sar9b_0.net37 0.03346f
C5765 a_9162_23174# a_9414_23127# 0.27388f
C5766 a_38738_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.23864f
C5767 VDPWR sar9b_0.net9 1.21348f
C5768 a_6282_17846# a_6880_17491# 0.06623f
C5769 sar9b_0.net52 sar9b_0.net11 0.15337f
C5770 sar9b_0.net20 a_8115_28566# 0.21703f
C5771 a_3695_23038# sar9b_0.clk_div_0.COUNT\[1\] 0.07641f
C5772 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38702f
C5773 sar9b_0.net60 sar9b_0._12_ 0.23194f
C5774 sar9b_0.net5 a_9494_20290# 0.0262f
C5775 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.02632f
C5776 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.42784f
C5777 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.7611f
C5778 VDPWR sar9b_0.net10 3.17323f
C5779 VDPWR sar9b_0.net61 2.29778f
C5780 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.12358f
C5781 VDPWR a_10402_21098# 0.21902f
C5782 a_4755_22138# a_5182_22567# 0.04602f
C5783 sar9b_0.net9 a_10218_21842# 0.02303f
C5784 single_9b_cdac_1.CF[3] ua[0] 3.58897f
C5785 a_11382_23474# sar9b_0.net74 0.18434f
C5786 sar9b_0.net9 sar9b_0.net1 0.02842f
C5787 a_3438_26345# a_3946_26198# 0.19065f
C5788 a_6642_19448# sar9b_0.net35 0.01573f
C5789 sar9b_0.net45 a_9593_26914# 0.02056f
C5790 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.01003f
C5791 a_8386_22806# sar9b_0.net57 0.03019f
C5792 sar9b_0.net63 a_2940_25096# 0.02555f
C5793 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5794 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C5795 sar9b_0.net15 sar9b_0.net4 0.47161f
C5796 a_5235_27466# sar9b_0.net59 0.05706f
C5797 a_8595_17910# a_8052_18123# 0.0131f
C5798 a_4125_25958# a_4293_25852# 0.27693f
C5799 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.14972f
C5800 sar9b_0.net1 sar9b_0.net10 0.02729f
C5801 sar9b_0.net1 sar9b_0.net61 0.02364f
C5802 VDPWR a_3206_22432# 0.86795f
C5803 a_2739_20140# a_2918_20140# 0.54426f
C5804 single_9b_cdac_1.CF[3] single_9b_cdac_1.CF[2] 14.3503f
C5805 sar9b_0.net48 sar9b_0.net73 0.46206f
C5806 single_9b_cdac_1.CF[2] sar9b_0.net28 0.04267f
C5807 a_8266_17113# a_7602_16784# 0.16939f
C5808 a_8334_17021# a_8052_16791# 0.05462f
C5809 sar9b_0.net2 a_9730_24138# 0.07985f
C5810 VDPWR a_6538_24506# 0.27686f
C5811 a_3371_23106# a_3695_23038# 0.15159f
C5812 sar9b_0.net38 a_7539_28566# 0.05709f
C5813 single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.10499f
C5814 VDPWR uio_out[1] 1.23314f
C5815 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.27843f
C5816 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.71729f
C5817 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.07579f
C5818 single_9b_cdac_0.SW[0] a_63626_26990# 0.18991f
C5819 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.28813f
C5820 sar9b_0.net57 a_4771_18260# 0.29258f
C5821 single_9b_cdac_1.SW[0] a_9974_17626# 0.0138f
C5822 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.17268f
C5823 sar9b_0.net31 sar9b_0.net26 0.03062f
C5824 VDPWR a_9279_27227# 0.27846f
C5825 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07517f
C5826 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.24495f
C5827 a_13011_21906# single_9b_cdac_1.CF[3] 0.02875f
C5828 a_48343_26999# single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.59531f
C5829 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[3] 14.7461f
C5830 a_9593_26914# a_9870_27060# 0.09983f
C5831 tdc_0.OUTN a_7743_16817# 0.05748f
C5832 sar9b_0.net30 sar9b_0.net12 0.09512f
C5833 sar9b_0.net43 sar9b_0.net41 0.34712f
C5834 VDPWR sar9b_0.net7 1.0007f
C5835 a_5484_23444# sar9b_0.net11 0.29424f
C5836 VDPWR a_21368_4076# 0.07949f
C5837 VDPWR a_9442_21474# 0.23612f
C5838 a_8622_26345# sar9b_0.net59 0.24081f
C5839 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.95338f
C5840 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.69086f
C5841 sar9b_0.net52 a_8098_23762# 0.0833f
C5842 sar9b_0.net29 single_9b_cdac_1.SW[8] 0.04274f
C5843 a_12182_22423# a_12618_22138# 0.16939f
C5844 sar9b_0.net41 sar9b_0.net13 0.0247f
C5845 VDPWR a_16527_10454# 0.3789f
C5846 sar9b_0.net46 sar9b_0.net73 0.14249f
C5847 sar9b_0.net58 a_3946_27530# 0.24636f
C5848 sar9b_0.net58 a_5465_28246# 0.07923f
C5849 sar9b_0.net52 sar9b_0.net45 0.18401f
C5850 a_14897_9355# clk 0.02917f
C5851 sar9b_0.net50 sar9b_0.net73 0.28503f
C5852 sar9b_0.net53 sar9b_0.net54 0.39148f
C5853 VDPWR a_5481_20185# 0.14537f
C5854 a_11466_23174# sar9b_0.net11 0.0513f
C5855 a_9730_24138# a_10758_24459# 0.07826f
C5856 sar9b_0.net32 single_9b_cdac_0.SW[7] 0.02288f
C5857 single_9b_cdac_1.SW[3] sar9b_0.net73 0.09966f
C5858 a_9442_21474# a_10218_21842# 0.3578f
C5859 a_9442_21474# sar9b_0.net1 0.02634f
C5860 uio_in[0] ui_in[7] 0.03102f
C5861 a_2835_24136# sar9b_0.clk_div_0.COUNT\[1\] 0.02455f
C5862 VDPWR a_6579_18832# 0.41927f
C5863 a_10607_25185# sar9b_0.net52 0.19466f
C5864 sar9b_0._09_ a_4947_20140# 0.01531f
C5865 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[4] 0.02164f
C5866 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C5867 sar9b_0.net23 sar9b_0.net36 0.02152f
C5868 sar9b_0.net41 a_10662_17799# 0.06166f
C5869 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 2.82222f
C5870 sar9b_0.net38 a_10607_21189# 0.01344f
C5871 sar9b_0.net22 sar9b_0.net45 0.14216f
C5872 a_11859_21906# sar9b_0.net26 0.01146f
C5873 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.24288f
C5874 a_10742_25087# sar9b_0.net36 0.01344f
C5875 a_11430_27595# VDPWR 0.26904f
C5876 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.SW[8] 0.22497f
C5877 a_8057_17131# sar9b_0.net27 0.01567f
C5878 a_8874_23470# clk 0.01286f
C5879 a_2892_23070# sar9b_0.net69 0.01085f
C5880 sar9b_0.net8 sar9b_0.net26 0.0267f
C5881 a_4934_22432# sar9b_0._12_ 0.06662f
C5882 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[0] 0.06503f
C5883 a_12182_23755# a_12618_23470# 0.16939f
C5884 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[8] 1.08672f
C5885 a_10378_27170# sar9b_0.net38 0.01469f
C5886 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[5] 0.06503f
C5887 a_4749_27652# uo_out[7] 0.01802f
C5888 sar9b_0.net43 a_9593_26914# 0.01648f
C5889 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 1.55985f
C5890 sar9b_0.net54 a_6562_25094# 0.07487f
C5891 VDPWR sar9b_0.net17 0.77016f
C5892 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C5893 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.26942f
C5894 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[6] 14.2348f
C5895 sar9b_0.net59 a_9138_27163# 0.3052f
C5896 sar9b_0.net35 sar9b_0.net57 0.03434f
C5897 sar9b_0.net40 th_dif_sw_0.CK 0.08068f
C5898 a_6484_22845# sar9b_0._17_ 0.03367f
C5899 a_6861_22828# a_6744_23238# 0.3009f
C5900 sar9b_0._07_ sar9b_0._17_ 0.02418f
C5901 sar9b_0.net48 sar9b_0.net46 0.56511f
C5902 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.26427f
C5903 th_dif_sw_0.CK a_12870_18271# 0.06999f
C5904 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 a_58824_17740# 0.14695f
C5905 sar9b_0.net48 sar9b_0.net50 0.03024f
C5906 sar9b_0.net16 sar9b_0.net57 0.01547f
C5907 sar9b_0.net35 a_7404_18116# 0.01538f
C5908 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02632f
C5909 a_7289_21127# a_8074_20870# 0.26257f
C5910 a_10830_19068# sar9b_0.net36 0.02201f
C5911 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.12358f
C5912 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 1.71649f
C5913 a_6783_19481# a_6444_19448# 0.07649f
C5914 a_2892_23070# sar9b_0._18_ 0.28345f
C5915 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5916 VDPWR a_5182_22567# 0.0129f
C5917 a_10506_23174# sar9b_0.net53 0.17591f
C5918 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[4] 0.01525f
C5919 VDPWR a_7539_28566# 0.41703f
C5920 sar9b_0._08_ sar9b_0._17_ 0.25385f
C5921 a_10506_23174# a_10690_22806# 0.44098f
C5922 a_10239_19235# sar9b_0.net49 0.02293f
C5923 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[1] 0.0147f
C5924 sar9b_0.net74 sar9b_0.net53 0.63719f
C5925 a_9942_27470# sar9b_0.net24 0.01062f
C5926 a_10690_22806# sar9b_0.net74 0.04092f
C5927 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.0303f
C5928 a_7138_27758# sar9b_0.net21 0.0211f
C5929 sar9b_0.net20 uo_out[6] 0.34847f
C5930 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.07579f
C5931 VDPWR a_13011_27234# 0.41846f
C5932 ui_in[0] ui_in[1] 0.03102f
C5933 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 1.71649f
C5934 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 a_44418_26990# 0.14695f
C5935 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.02666f
C5936 a_7138_27758# a_8166_27595# 0.07826f
C5937 VDPWR a_3822_27060# 0.26946f
C5938 sar9b_0.net31 sar9b_0.net53 0.91386f
C5939 a_9414_23127# sar9b_0.net11 0.06993f
C5940 a_8940_27039# sar9b_0.net37 0.05651f
C5941 a_10690_22806# sar9b_0.net31 0.01488f
C5942 a_8591_22855# sar9b_0.net54 0.22373f
C5943 VDPWR a_2892_27039# 0.25024f
C5944 a_6307_27584# a_6678_27470# 0.04761f
C5945 VDPWR a_4018_24235# 0.3802f
C5946 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.CF[0] 0.10499f
C5947 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5948 sar9b_0.net61 a_8052_16791# 0.07136f
C5949 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.19266f
C5950 a_12491_27662# sar9b_0.net52 0.01099f
C5951 sar9b_0.net67 sar9b_0._12_ 0.06679f
C5952 sar9b_0._07_ a_5633_20244# 0.0155f
C5953 sar9b_0.net40 single_9b_cdac_1.SW[1] 0.10842f
C5954 a_10742_27751# sar9b_0.net59 0.14619f
C5955 th_dif_sw_0.th_sw_1.CKB ua[4] 0.08416f
C5956 a_8982_21902# sar9b_0.net37 0.02238f
C5957 a_8266_18445# sar9b_0.net5 0.04964f
C5958 a_10858_17113# single_9b_cdac_1.SW[2] 0.02538f
C5959 sar9b_0.net56 a_8694_20570# 0.01417f
C5960 sar9b_0.net43 sar9b_0.net52 0.08027f
C5961 VDPWR a_8438_18958# 0.21428f
C5962 sar9b_0.net47 a_5811_19178# 0.01123f
C5963 sar9b_0.net10 a_11658_22138# 0.24856f
C5964 single_9b_cdac_1.CF[5] ua[0] 3.57763f
C5965 single_9b_cdac_0.SW[4] ua[0] 0.17308f
C5966 a_4293_25852# sar9b_0.clknet_1_1__leaf_CLK 0.04421f
C5967 single_9b_cdac_0.SW[3] a_49221_26990# 0.18991f
C5968 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[4] 0.26707f
C5969 a_6250_28502# uo_out[6] 0.02897f
C5970 a_4136_25584# sar9b_0._03_ 0.29527f
C5971 a_12618_18142# sar9b_0.net50 0.26153f
C5972 a_3603_28156# sar9b_0.net60 0.28939f
C5973 sar9b_0.net55 sar9b_0.net15 0.43777f
C5974 sar9b_0.net13 sar9b_0.net52 1.35209f
C5975 a_3369_24181# sar9b_0.net70 0.01723f
C5976 sar9b_0.net17 a_2508_27440# 0.01561f
C5977 a_16159_13315# a_16185_12837# 0.01114f
C5978 a_11842_26426# a_12182_26419# 0.24088f
C5979 a_11658_26134# a_12618_26134# 0.03432f
C5980 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.01751f
C5981 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[2] 0.02195f
C5982 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[0] 0.06019f
C5983 a_6880_26815# sar9b_0.net37 0.04911f
C5984 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.81428f
C5985 sar9b_0.net69 a_3372_25734# 0.14523f
C5986 VDPWR a_10607_21189# 0.26776f
C5987 sar9b_0.net30 a_12047_26517# 0.02505f
C5988 a_9126_19131# a_7914_19178# 0.07766f
C5989 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.17533f
C5990 sar9b_0.net58 sar9b_0.net39 0.55587f
C5991 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.69086f
C5992 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[3] 12.1694f
C5993 single_9b_cdac_1.CF[4] sar9b_0.net28 0.36381f
C5994 sar9b_0.net52 a_12560_27128# 0.08336f
C5995 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.24443f
C5996 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[3] 0.05125f
C5997 single_9b_cdac_1.CF[1] sar9b_0.net28 0.04257f
C5998 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.38397f
C5999 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01156f
C6000 VDPWR a_10378_27170# 0.30084f
C6001 sar9b_0.net16 a_4496_20468# 0.03603f
C6002 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.75815f
C6003 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[0\] 0.86907f
C6004 sar9b_0.net40 sar9b_0.net60 0.49844f
C6005 sar9b_0.net41 a_9760_22819# 0.28794f
C6006 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 1.71649f
C6007 a_11434_16874# tdc_0.OUTP 0.04839f
C6008 sar9b_0.net43 a_5100_24375# 0.27992f
C6009 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.24311f
C6010 single_9b_cdac_1.cdac_sw_9b_0.S[1] a_57946_16877# 0.59531f
C6011 a_7188_22119# a_6738_22112# 0.03529f
C6012 sar9b_0.net32 a_12618_26134# 0.01453f
C6013 sar9b_0.net47 sar9b_0.net39 0.20215f
C6014 single_9b_cdac_0.SW[6] clk 0.22166f
C6015 a_6484_22845# clk 0.01293f
C6016 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[6] 0.01475f
C6017 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 1.71649f
C6018 sar9b_0.net35 sar9b_0.clk_div_0.COUNT\[1\] 0.03758f
C6019 a_11658_23470# a_11842_23762# 0.44532f
C6020 sar9b_0.net40 a_5753_24250# 0.01091f
C6021 single_9b_cdac_0.cdac_sw_9b_0.S[4] ua[0] 1.93763f
C6022 a_13011_27234# sar9b_0.net29 0.01376f
C6023 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.7611f
C6024 a_7914_23470# sar9b_0.net57 0.22944f
C6025 sar9b_0.net26 a_12182_22423# 0.0187f
C6026 VDPWR a_2940_25096# 0.20267f
C6027 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.06503f
C6028 sar9b_0.net37 sar9b_0.net39 0.18921f
C6029 single_9b_cdac_1.SW[4] sar9b_0.net6 0.02588f
C6030 sar9b_0._14_ a_2940_25096# 0.01562f
C6031 a_2893_24992# a_3364_25120# 0.01114f
C6032 a_6922_23534# sar9b_0.net54 0.26015f
C6033 a_16159_13315# tdc_0.OUTN 0.01845f
C6034 a_3545_26914# a_4330_27170# 0.26257f
C6035 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6036 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[3] 0.01497f
C6037 single_9b_cdac_1.CF[8] sar9b_0.net28 0.04086f
C6038 sar9b_0.net74 a_10932_25713# 0.06691f
C6039 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._04_ 0.01564f
C6040 sar9b_0.net9 a_7193_22459# 0.01552f
C6041 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] 3.10215f
C6042 a_10227_18142# a_9634_17478# 0.01011f
C6043 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.11216f
C6044 sar9b_0.net26 a_12182_23755# 0.01551f
C6045 VDPWR tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.45583f
C6046 a_5010_28495# sar9b_0.net20 0.08006f
C6047 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.42784f
C6048 a_3231_27227# a_3540_27045# 0.07766f
C6049 a_8074_20870# sar9b_0.net47 0.22159f
C6050 a_10335_16817# sar9b_0.net27 0.02939f
C6051 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 2.71729f
C6052 a_5100_24375# a_5298_24499# 0.06623f
C6053 sar9b_0.net10 a_7193_22459# 0.01351f
C6054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.01152f
C6055 a_8098_18810# sar9b_0.net37 0.01309f
C6056 a_6834_20780# sar9b_0.net35 0.03194f
C6057 VDPWR a_13011_24802# 0.4961f
C6058 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.02778f
C6059 w_17430_1606# dw_17224_1400# 9.71413f
C6060 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 a_30012_17740# 0.14695f
C6061 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.SW[3] 0.15108f
C6062 sar9b_0._13_ a_4811_23656# 0.11957f
C6063 VDPWR single_9b_cdac_1.SW[4] 2.6945f
C6064 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] 1.15132f
C6065 sar9b_0.net35 a_7443_21496# 0.01956f
C6066 sar9b_0._11_ sar9b_0.net57 0.0163f
C6067 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.07517f
C6068 VDPWR a_5535_18149# 0.2712f
C6069 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07517f
C6070 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C6071 a_8202_23174# a_8726_22954# 0.04522f
C6072 a_7926_23234# a_8591_22855# 0.19065f
C6073 sar9b_0.net13 a_6102_24806# 0.23362f
C6074 sar9b_0.net59 a_10607_27849# 0.21965f
C6075 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.22875f
C6076 a_4811_23656# a_5002_23764# 0.01358f
C6077 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.SW[4] 0.17175f
C6078 a_8982_21902# sar9b_0.net57 0.05351f
C6079 sar9b_0.net2 a_10803_19474# 0.02668f
C6080 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.03729f
C6081 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.10503f
C6082 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.22549f
C6083 sar9b_0.net58 sar9b_0.net72 0.01694f
C6084 VDPWR a_13011_25902# 0.47442f
C6085 a_4947_20140# a_5126_20140# 0.54426f
C6086 a_5374_20145# sar9b_0.net57 0.01527f
C6087 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.95338f
C6088 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.62443f
C6089 sar9b_0.net58 sar9b_0.net36 0.27889f
C6090 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[5] 0.0187f
C6091 a_6030_24396# a_6538_24506# 0.19065f
C6092 sar9b_0._07_ sar9b_0._12_ 0.03077f
C6093 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.27554f
C6094 a_9935_24187# sar9b_0.net53 0.2035f
C6095 a_11466_23174# a_11718_23127# 0.27388f
C6096 a_6880_17491# sar9b_0.net46 0.03742f
C6097 a_5441_22522# sar9b_0._12_ 0.04735f
C6098 VDPWR sar9b_0.cyclic_flag_0.FINAL 0.90593f
C6099 single_9b_cdac_1.CF[3] sar9b_0.net28 0.03461f
C6100 a_8842_16874# sar9b_0.net6 0.05357f
C6101 VDPWR sar9b_0.net15 0.41783f
C6102 sar9b_0.net64 a_6444_21738# 0.1416f
C6103 a_13011_27234# single_9b_cdac_0.SW[3] 0.01848f
C6104 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C6105 sar9b_0.net36 a_9323_27662# 0.03315f
C6106 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.03729f
C6107 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_53154_26999# 0.04592f
C6108 a_5100_24375# sar9b_0._15_ 0.06016f
C6109 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C6110 sar9b_0.net53 a_12182_22423# 0.14409f
C6111 VDPWR a_4293_25852# 0.10504f
C6112 sar9b_0.net42 single_9b_cdac_0.SW[7] 0.0472f
C6113 sar9b_0.net36 sar9b_0.net37 0.0292f
C6114 sar9b_0.net30 sar9b_0.net74 0.03698f
C6115 sar9b_0.net48 sar9b_0.net27 0.34189f
C6116 sar9b_0.net60 uo_out[7] 0.02565f
C6117 VDPWR a_8019_17910# 0.39892f
C6118 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.75849f
C6119 sar9b_0.net20 sar9b_0.net45 0.05044f
C6120 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._12_ 0.12298f
C6121 sar9b_0.net53 a_12182_23755# 0.14448f
C6122 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[4] 9.91576f
C6123 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[4] 1.90123f
C6124 sar9b_0.net31 a_12047_22521# 0.04699f
C6125 VDPWR a_8842_16874# 0.29337f
C6126 sar9b_0.net41 a_9839_17527# 0.06481f
C6127 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.05472f
C6128 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07517f
C6129 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[5] 0.02038f
C6130 sar9b_0._16_ sar9b_0.clk_div_0.COUNT\[1\] 0.1686f
C6131 a_3855_25792# a_4125_25958# 0.08669f
C6132 a_8726_22954# sar9b_0.net37 0.01269f
C6133 VDPWR a_7882_19538# 0.30688f
C6134 a_10284_25707# a_10623_25895# 0.07649f
C6135 a_13011_24802# sar9b_0.net29 0.01443f
C6136 sar9b_0.net31 sar9b_0.net30 0.08627f
C6137 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[7] 0.01475f
C6138 sar9b_0.net42 a_11382_22142# 0.01996f
C6139 a_3161_27787# a_3370_27769# 0.24088f
C6140 a_10098_19171# sar9b_0.net36 0.0123f
C6141 a_8019_17910# sar9b_0.net1 0.01265f
C6142 sar9b_0._11_ a_4496_20468# 0.09559f
C6143 a_10470_21795# a_9258_21842# 0.07766f
C6144 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.6919f
C6145 sar9b_0.net74 a_11104_24151# 0.01447f
C6146 sar9b_0.net57 sar9b_0.net39 0.68049f
C6147 VDPWR a_8842_18206# 0.30615f
C6148 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95338f
C6149 sar9b_0.net41 sar9b_0.net38 0.17261f
C6150 VDPWR a_12618_19474# 0.35538f
C6151 a_17125_9355# a_16331_9671# 0.06748f
C6152 a_6744_23238# sar9b_0.clk_div_0.COUNT\[1\] 0.02511f
C6153 VDPWR a_5046_27230# 0.28883f
C6154 tdc_0.OUTP sar9b_0.net48 0.1166f
C6155 sar9b_0.net40 a_6767_25185# 0.02519f
C6156 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.02624f
C6157 a_6250_28502# sar9b_0.net45 0.03629f
C6158 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.SW[2] 0.22543f
C6159 a_8842_18206# sar9b_0.net1 0.03616f
C6160 sar9b_0.net52 a_12870_26263# 0.17285f
C6161 VDPWR a_4812_28371# 0.19653f
C6162 sar9b_0.net27 sar9b_0.net46 0.77693f
C6163 a_13011_25902# sar9b_0.net29 0.01649f
C6164 clk single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.02119f
C6165 VDPWR sar9b_0.net18 1.35357f
C6166 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.19266f
C6167 sar9b_0.net27 sar9b_0.net50 0.03263f
C6168 ua[4] th_dif_sw_0.VCP 3.30291f
C6169 a_6102_24806# sar9b_0.net4 0.02847f
C6170 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.3196f
C6171 single_9b_cdac_1.SW[3] sar9b_0.net27 0.02529f
C6172 a_12182_19759# sar9b_0.net6 0.02207f
C6173 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C6174 sar9b_0.net32 sar9b_0.net25 0.11681f
C6175 a_24332_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.23864f
C6176 sar9b_0.net58 a_4136_25584# 0.04102f
C6177 sar9b_0.net27 a_12618_18142# 0.02447f
C6178 a_13011_21906# a_13216_22473# 0.01179f
C6179 a_11658_18142# sar9b_0.net50 0.17638f
C6180 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[5] 0.01577f
C6181 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[4] 0.0154f
C6182 sar9b_0.net44 sar9b_0.net45 0.33602f
C6183 single_9b_cdac_1.SW[3] a_11658_18142# 0.02689f
C6184 sar9b_0.net63 a_5100_24375# 0.0166f
C6185 a_11658_18142# a_12618_18142# 0.03432f
C6186 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[4] 0.06503f
C6187 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.69086f
C6188 a_10830_19068# sar9b_0.net7 0.01607f
C6189 sar9b_0.net49 th_dif_sw_0.CK 0.01033f
C6190 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.84082f
C6191 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR 0.38397f
C6192 uio_out[0] uo_out[7] 2.91188f
C6193 uio_out[1] ui_in[0] 1.11045f
C6194 a_11008_17491# sar9b_0.net2 0.03502f
C6195 sar9b_0.net63 a_5484_23444# 0.04251f
C6196 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.31809f
C6197 single_9b_cdac_0.SW[8] th_dif_sw_0.VCN 0.15316f
C6198 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.CKB 4.72443f
C6199 a_7338_24802# a_7936_25137# 0.06623f
C6200 a_13011_27234# a_13216_26469# 0.01043f
C6201 sar9b_0.net38 a_9593_26914# 0.0231f
C6202 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] 0.28871f
C6203 a_2706_26108# a_3161_26455# 0.3578f
C6204 tdc_0.OUTP single_9b_cdac_1.SW[3] 0.04678f
C6205 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.8438f
C6206 sar9b_0.net26 sar9b_0.net73 0.02035f
C6207 a_7289_21127# sar9b_0.net10 0.01176f
C6208 sar9b_0.net5 single_9b_cdac_1.SW[0] 0.03107f
C6209 VDPWR a_5083_21100# 0.18914f
C6210 VDPWR a_12182_19759# 0.20727f
C6211 sar9b_0.net41 sar9b_0.net6 0.02799f
C6212 single_9b_cdac_0.SW[5] uo_out[1] 0.07247f
C6213 a_8098_23762# a_8438_23755# 0.24088f
C6214 sar9b_0.net56 sar9b_0.net5 1.07927f
C6215 a_9942_27470# a_10402_27758# 0.26257f
C6216 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.59531f
C6217 a_7374_19685# sar9b_0.net47 0.29639f
C6218 VDPWR a_16357_9613# 0.18873f
C6219 a_11178_20806# a_11776_21141# 0.06623f
C6220 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.3601f
C6221 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.22875f
C6222 a_4083_28566# a_4812_28371# 0.01209f
C6223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.42509f
C6224 sar9b_0.net57 a_4332_23043# 0.0332f
C6225 single_9b_cdac_1.CF[6] ua[0] 3.57763f
C6226 sar9b_0.net18 a_4083_28566# 0.2051f
C6227 a_3603_28156# sar9b_0.net59 0.32304f
C6228 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[0\] 0.08053f
C6229 a_11915_28371# VDPWR 0.45787f
C6230 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C6231 a_5938_22378# sar9b_0.clk_div_0.COUNT\[0\] 0.11986f
C6232 sar9b_0.net8 a_11658_19474# 0.2065f
C6233 dw_12589_1395# w_12795_1601# 9.86148f
C6234 sar9b_0.net18 a_2508_27440# 0.28434f
C6235 a_3603_28156# a_3156_27447# 0.02744f
C6236 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.81434f
C6237 sar9b_0.net45 single_9b_cdac_0.SW[8] 0.08609f
C6238 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[1] 4.14969f
C6239 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 2.82223f
C6240 a_9414_23127# a_9760_22819# 0.07649f
C6241 a_2508_23444# sar9b_0.clk_div_0.COUNT\[1\] 0.06012f
C6242 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[3] 0.02744f
C6243 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[2] 0.02038f
C6244 single_9b_cdac_1.CF[5] sar9b_0.net28 0.03576f
C6245 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.28523f
C6246 sar9b_0.net63 a_7483_23174# 0.01409f
C6247 VDPWR sar9b_0.net41 1.4128f
C6248 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0313f
C6249 a_11436_17742# sar9b_0.net27 0.04295f
C6250 sar9b_0.net26 sar9b_0.net48 0.4034f
C6251 a_9363_20826# sar9b_0.net8 0.03842f
C6252 sar9b_0.net52 sar9b_0.net38 0.0649f
C6253 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.04988f
C6254 sar9b_0.net28 a_13216_18477# 0.28248f
C6255 VDPWR a_11430_20935# 0.27331f
C6256 VDPWR a_5674_28147# 0.19864f
C6257 sar9b_0.net64 a_5182_22567# 0.12016f
C6258 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.36013f
C6259 sar9b_0.clk_div_0.COUNT\[1\] sar9b_0.net39 0.0203f
C6260 a_7097_19795# sar9b_0.net35 0.01811f
C6261 sar9b_0.net41 sar9b_0.net1 0.90489f
C6262 VDPWR a_6879_22145# 0.27369f
C6263 a_43540_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.23864f
C6264 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.42509f
C6265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.26942f
C6266 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 2.82172f
C6267 sar9b_0.net17 ui_in[0] 0.02606f
C6268 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[7] 0.06912f
C6269 sar9b_0.net40 sar9b_0.net59 0.03006f
C6270 VDPWR a_38738_16877# 1.81495f
C6271 a_3922_20239# sar9b_0.net16 0.1201f
C6272 a_8019_17910# a_8052_16791# 0.03036f
C6273 a_10662_17799# a_9634_17478# 0.07826f
C6274 sar9b_0.net35 a_7347_24160# 0.03326f
C6275 a_7188_22119# sar9b_0.net54 0.01061f
C6276 sar9b_0.net32 single_9b_cdac_0.SW[6] 0.05164f
C6277 m2_23774_26966# single_9b_cdac_0.SW[8] 0.02037f
C6278 a_2918_20140# sar9b_0._00_ 0.27567f
C6279 a_8842_16874# a_8052_16791# 0.1263f
C6280 a_8266_17113# a_8057_17131# 0.24088f
C6281 sar9b_0.net2 a_10070_24286# 0.0649f
C6282 a_3855_25792# sar9b_0.clknet_1_1__leaf_CLK 0.07223f
C6283 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 3.10626f
C6284 single_9b_cdac_0.SW[8] uo_out[0] 0.10191f
C6285 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.05472f
C6286 sar9b_0.net38 sar9b_0.net22 0.04437f
C6287 single_9b_cdac_1.SW[2] sar9b_0.net37 0.07696f
C6288 VDPWR tdc_0.phase_detector_0.pd_out_0.A 1.77491f
C6289 sar9b_0.net54 clk 0.11407f
C6290 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.3196f
C6291 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.31534f
C6292 sar9b_0.net12 a_11658_26134# 0.21062f
C6293 VDPWR a_2739_20140# 0.47557f
C6294 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.SW[2] 0.15027f
C6295 a_8202_23174# sar9b_0.net61 0.01019f
C6296 a_5748_24381# a_6378_24802# 0.01007f
C6297 VDPWR single_9b_cdac_1.SW[6] 2.4631f
C6298 a_6738_22112# sar9b_0.net40 0.02168f
C6299 a_5849_18463# a_6126_18353# 0.09983f
C6300 sar9b_0.net26 sar9b_0.net50 0.09003f
C6301 a_18214_3039# VDPWR 0.51112f
C6302 single_9b_cdac_1.cdac_sw_9b_0.S[5] ua[0] 1.57219f
C6303 sar9b_0.net60 uo_out[6] 0.01362f
C6304 VDPWR a_9593_26914# 0.22537f
C6305 sar9b_0.net53 sar9b_0.net73 0.13314f
C6306 a_10227_18142# th_dif_sw_0.CK 0.35616f
C6307 sar9b_0.net42 a_10402_25094# 0.01861f
C6308 sar9b_0.net52 a_9165_24988# 0.35265f
C6309 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.42509f
C6310 VDPWR a_9782_21622# 0.20774f
C6311 a_9130_26198# sar9b_0.net59 0.27842f
C6312 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.81434f
C6313 a_4467_24162# sar9b_0.net72 0.02699f
C6314 sar9b_0.net52 a_9126_23599# 0.20232f
C6315 sar9b_0.net13 a_7936_25137# 0.0469f
C6316 a_12870_22267# a_13216_22473# 0.07649f
C6317 single_9b_cdac_0.SW[6] a_10995_28566# 0.01025f
C6318 a_12182_22423# a_12047_22521# 0.35559f
C6319 VDPWR tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.45581f
C6320 a_3922_20239# a_3723_20140# 0.29821f
C6321 single_9b_cdac_1.SW[3] a_48343_16877# 0.28324f
C6322 a_3540_27045# sar9b_0.net44 0.27099f
C6323 a_9782_21622# a_10218_21842# 0.16939f
C6324 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.10429f
C6325 single_9b_cdac_1.cdac_sw_9b_0.S[0] a_62748_16877# 0.59531f
C6326 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 ua[0] 0.12344f
C6327 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.17533f
C6328 a_3946_27530# a_3161_27787# 0.26257f
C6329 sar9b_0.net70 sar9b_0.clk_div_0.COUNT\[1\] 0.23038f
C6330 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6331 sar9b_0.net9 sar9b_0.net47 0.32405f
C6332 a_10194_16784# sar9b_0.net36 0.05607f
C6333 sar9b_0.net32 sar9b_0.net12 0.03166f
C6334 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] 0.12898f
C6335 a_10553_18922# sar9b_0.net42 0.018f
C6336 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.02618f
C6337 sar9b_0._09_ sar9b_0._10_ 0.14294f
C6338 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C6339 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C6340 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C6341 sar9b_0.net30 a_12182_23755# 0.02293f
C6342 sar9b_0.net47 sar9b_0.net10 1.99512f
C6343 sar9b_0.net47 sar9b_0.net61 0.15705f
C6344 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.02778f
C6345 a_10506_23174# clk 0.01873f
C6346 sar9b_0.net74 clk 0.07221f
C6347 sar9b_0.net9 sar9b_0.net37 0.08996f
C6348 a_4332_23043# sar9b_0.clk_div_0.COUNT\[1\] 0.81462f
C6349 sar9b_0.net66 sar9b_0.net69 0.14538f
C6350 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[6] 0.02149f
C6351 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.07517f
C6352 a_11776_27801# VDPWR 0.20399f
C6353 single_9b_cdac_0.SW[1] sar9b_0.net27 0.088f
C6354 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.08121f
C6355 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[5] 0.01299f
C6356 single_9b_cdac_0.SW[7] th_dif_sw_0.VCN 0.0955f
C6357 a_12531_28566# sar9b_0._06_ 0.02926f
C6358 a_2828_22432# sar9b_0._05_ 0.01634f
C6359 a_5331_16810# sar9b_0.net27 0.05702f
C6360 a_12182_23755# a_12047_23853# 0.35559f
C6361 a_12870_23599# a_13216_23805# 0.07649f
C6362 sar9b_0.net70 a_3371_23106# 0.01159f
C6363 a_13011_25902# a_13216_26469# 0.01179f
C6364 sar9b_0.net27 a_12618_22138# 0.02584f
C6365 VDPWR sar9b_0.net52 3.91808f
C6366 sar9b_0.net61 sar9b_0.net37 0.52176f
C6367 sar9b_0.net54 a_7590_24931# 0.20557f
C6368 sar9b_0.net10 sar9b_0.net37 0.02841f
C6369 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36542f
C6370 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.03729f
C6371 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.969f
C6372 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62573f
C6373 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.18989f
C6374 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.12898f
C6375 a_62748_16877# single_9b_cdac_1.SW[0] 0.28324f
C6376 sar9b_0.net31 clk 0.0477f
C6377 sar9b_0.net72 sar9b_0.clk_div_0.COUNT\[1\] 0.04678f
C6378 a_10166_3438# ua[4] 0.65763f
C6379 sar9b_0.net59 a_9588_27045# 0.18035f
C6380 VDPWR a_11146_25483# 0.19884f
C6381 sar9b_0._02_ sar9b_0._17_ 0.15132f
C6382 single_9b_cdac_1.CF[7] ua[0] 3.57763f
C6383 sar9b_0.net21 uo_out[5] 0.07619f
C6384 a_12588_16784# sar9b_0.net2 0.14533f
C6385 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[0] 0.56248f
C6386 sar9b_0._18_ sar9b_0.net66 0.0125f
C6387 sar9b_0.net27 a_12618_23470# 0.02584f
C6388 sar9b_0.net36 a_10410_17846# 0.02317f
C6389 single_9b_cdac_0.SW[5] a_13164_28398# 0.01688f
C6390 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.42784f
C6391 VDPWR sar9b_0.net22 0.53629f
C6392 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[2] 0.02011f
C6393 sar9b_0.net16 a_5581_19664# 0.01792f
C6394 a_10506_23174# a_11030_22954# 0.04522f
C6395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.12431f
C6396 a_10230_23234# a_10895_22855# 0.19065f
C6397 sar9b_0.net41 a_9270_24566# 0.01466f
C6398 a_11030_22954# sar9b_0.net74 0.01098f
C6399 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.28523f
C6400 sar9b_0.net35 a_7402_22441# 0.01975f
C6401 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[5] 1.26495f
C6402 a_7404_17715# sar9b_0.net5 0.05199f
C6403 single_9b_cdac_0.SW[7] sar9b_0.net45 0.21976f
C6404 sar9b_0._09_ sar9b_0._18_ 0.1776f
C6405 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[7] 1.64863f
C6406 sar9b_0.net56 a_9942_20810# 0.04264f
C6407 a_7478_27751# a_7914_27466# 0.16939f
C6408 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96893f
C6409 a_9279_27227# sar9b_0.net37 0.07713f
C6410 sar9b_0._09_ sar9b_0._01_ 0.03554f
C6411 sar9b_0.net19 sar9b_0.net39 0.0141f
C6412 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[4] 0.06951f
C6413 a_62748_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.23864f
C6414 VDPWR a_3231_27227# 0.28136f
C6415 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[2] 0.22004f
C6416 VDPWR a_5100_24375# 0.1934f
C6417 sar9b_0.net59 uo_out[7] 0.02838f
C6418 a_25210_26990# single_9b_cdac_0.SW[8] 0.18991f
C6419 a_11178_27466# sar9b_0.net59 0.26568f
C6420 a_9442_21474# sar9b_0.net37 0.01287f
C6421 sar9b_0.net23 sar9b_0.cyclic_flag_0.FINAL 0.03316f
C6422 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C6423 sar9b_0.net10 a_11842_22430# 0.03989f
C6424 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36041f
C6425 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38733f
C6426 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.26942f
C6427 VDPWR a_5484_23444# 0.19999f
C6428 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.27833f
C6429 sar9b_0.net36 a_10803_19474# 0.21894f
C6430 a_5010_28495# sar9b_0.net60 0.06731f
C6431 sar9b_0.net58 sar9b_0.net17 0.01182f
C6432 VDPWR a_7692_26108# 0.20712f
C6433 a_12047_18525# sar9b_0.net50 0.22675f
C6434 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[4] 0.02215f
C6435 a_7926_23234# clk 0.01904f
C6436 single_9b_cdac_1.SW[1] th_dif_sw_0.VCN 0.0955f
C6437 single_9b_cdac_1.SW[3] a_12047_18525# 0.01367f
C6438 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[6] 0.02011f
C6439 VDPWR a_4947_20140# 0.39022f
C6440 a_29134_16877# single_9b_cdac_1.SW[7] 0.28324f
C6441 sar9b_0.net17 a_2706_27440# 0.02173f
C6442 VDPWR a_7092_19455# 0.85935f
C6443 a_11658_26134# a_12047_26517# 0.06034f
C6444 a_11842_26426# a_12618_26134# 0.3578f
C6445 uio_in[5] uio_in[4] 0.03102f
C6446 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCP 1.0224f
C6447 VDPWR a_11466_23174# 0.34557f
C6448 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C6449 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.11216f
C6450 single_9b_cdac_0.SW[7] uo_out[0] 0.04546f
C6451 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[3] 1.26495f
C6452 a_9930_20510# sar9b_0.net51 0.07643f
C6453 VDPWR a_8052_18123# 0.76662f
C6454 sar9b_0.net60 sar9b_0.net11 0.10348f
C6455 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.07517f
C6456 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[8] 0.04036f
C6457 VDPWR tdc_0.RDY 0.57898f
C6458 a_10230_23234# sar9b_0.net36 0.01418f
C6459 uo_out[2] uo_out[1] 3.05143f
C6460 sar9b_0.net56 sar9b_0.net8 0.13034f
C6461 a_6378_24802# a_6902_25087# 0.05022f
C6462 VDPWR a_3855_25792# 0.09015f
C6463 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.26684f
C6464 sar9b_0._09_ a_3795_19512# 0.09292f
C6465 a_9154_20142# a_9494_20290# 0.24088f
C6466 a_10254_2858# ua[4] 0.12559f
C6467 sar9b_0.net58 a_3822_27060# 0.22673f
C6468 a_8052_18123# sar9b_0.net1 0.02679f
C6469 sar9b_0._09_ a_3180_19448# 0.26014f
C6470 sar9b_0.net17 a_2508_26108# 0.28355f
C6471 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.3196f
C6472 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.71729f
C6473 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.3196f
C6474 sar9b_0._09_ sar9b_0.net60 0.06706f
C6475 a_4018_24235# sar9b_0.net58 0.01775f
C6476 sar9b_0.net32 a_9323_28371# 0.22468f
C6477 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[6] 0.02343f
C6478 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.01608f
C6479 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.22983f
C6480 sar9b_0.net8 a_13011_20806# 0.22594f
C6481 sar9b_0.net40 sar9b_0.net5 0.02461f
C6482 VDPWR a_6102_24806# 0.29526f
C6483 a_7478_27751# a_7343_27849# 0.35559f
C6484 sar9b_0.net32 a_12047_26517# 0.01148f
C6485 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.04592f
C6486 VDPWR a_24332_16877# 1.81495f
C6487 a_10218_24802# a_10402_25094# 0.44532f
C6488 a_3521_24240# sar9b_0.clknet_1_1__leaf_CLK 0.04554f
C6489 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.SW[6] 0.14966f
C6490 sar9b_0._02_ clk 0.01536f
C6491 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6492 sar9b_0.net9 sar9b_0.net57 0.06836f
C6493 sar9b_0.net5 sar9b_0.net51 1.21471f
C6494 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] 1.15121f
C6495 a_11658_23470# a_12870_23599# 0.07766f
C6496 sar9b_0.net26 a_12618_22138# 0.02736f
C6497 VDPWR a_5196_24776# 0.23838f
C6498 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.CF[5] 0.12358f
C6499 sar9b_0.net43 a_9546_24506# 0.06524f
C6500 a_10194_16784# a_9450_17846# 0.01861f
C6501 a_5046_27230# a_5711_26851# 0.19065f
C6502 sar9b_0.net38 uo_out[3] 0.26142f
C6503 VDPWR a_7284_20787# 0.86664f
C6504 sar9b_0.net61 sar9b_0.net57 0.18181f
C6505 sar9b_0.net10 sar9b_0.net57 0.09558f
C6506 sar9b_0.net52 a_9270_24566# 0.02178f
C6507 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C6508 sar9b_0.net49 a_8694_20570# 0.22589f
C6509 a_8345_26455# a_8622_26345# 0.09983f
C6510 tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTN 0.19342f
C6511 a_3561_22527# a_3027_22138# 0.35097f
C6512 sar9b_0.net52 a_11382_26138# 0.24197f
C6513 a_10762_18823# sar9b_0.net2 0.01126f
C6514 a_8266_18445# sar9b_0.net73 0.05509f
C6515 sar9b_0.net46 a_5196_18116# 0.01474f
C6516 sar9b_0.net74 a_11214_25728# 0.06877f
C6517 a_11382_19478# a_12047_19857# 0.19065f
C6518 a_3561_22527# sar9b_0.net65 0.0125f
C6519 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.03729f
C6520 sar9b_0.net26 a_12618_23470# 0.02755f
C6521 sar9b_0.net36 sar9b_0.net19 0.07564f
C6522 sar9b_0.net65 sar9b_0.clknet_0_CLK 0.2446f
C6523 VDPWR a_9414_23127# 0.27453f
C6524 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.84424f
C6525 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.05472f
C6526 sar9b_0.net60 sar9b_0.net45 1.09005f
C6527 a_5151_28559# a_5465_28246# 0.07826f
C6528 sar9b_0.net31 a_11214_25728# 0.01178f
C6529 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.11216f
C6530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.28813f
C6531 sar9b_0.net42 sar9b_0.net59 0.13366f
C6532 VDPWR a_43540_26999# 1.81495f
C6533 VDPWR a_13011_16810# 0.4276f
C6534 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.02513f
C6535 a_6879_22145# a_7193_22459# 0.07826f
C6536 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.42784f
C6537 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C6538 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.69086f
C6539 a_49926_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.01076f
C6540 sar9b_0.net1 a_9414_23127# 0.02489f
C6541 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[8] 4.16545f
C6542 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR 0.38716f
C6543 sar9b_0.net26 sar9b_0.net27 0.67638f
C6544 a_10239_19235# a_10548_19053# 0.07766f
C6545 a_8874_19178# a_9126_19131# 0.27388f
C6546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C6547 sar9b_0.net5 a_13011_20574# 0.2669f
C6548 a_9634_17478# a_9839_17527# 0.09983f
C6549 a_9450_17846# a_10410_17846# 0.03493f
C6550 ui_in[0] rst_n 0.03102f
C6551 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[3] 0.02091f
C6552 single_9b_cdac_1.CF[6] sar9b_0.net28 0.04016f
C6553 single_9b_cdac_1.SW[2] a_10410_17846# 0.06269f
C6554 a_5484_23444# a_5682_23444# 0.06623f
C6555 sar9b_0.net20 sar9b_0.net38 0.02978f
C6556 a_5506_17478# a_5711_17527# 0.09983f
C6557 a_9442_21474# sar9b_0.net57 0.0155f
C6558 a_65367_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C6559 a_8266_18445# sar9b_0.net48 0.02071f
C6560 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.19266f
C6561 sar9b_0.net14 sar9b_0.net25 0.2521f
C6562 a_6282_17846# sar9b_0.net56 0.06691f
C6563 a_13216_23805# a_13011_24570# 0.01043f
C6564 a_5126_20140# sar9b_0._10_ 0.06232f
C6565 sar9b_0.net68 sar9b_0._16_ 0.0172f
C6566 sar9b_0.net63 a_2893_24992# 0.0883f
C6567 a_5628_19768# sar9b_0._10_ 0.06416f
C6568 single_9b_cdac_0.cdac_sw_9b_0.S[0] ua[0] 1.19231f
C6569 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[7] 0.02091f
C6570 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[7] 0.01994f
C6571 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96841f
C6572 sar9b_0._12_ sar9b_0._02_ 0.12883f
C6573 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[5] 0.42014f
C6574 a_8303_23853# a_7638_23474# 0.19065f
C6575 a_10816_21487# a_10218_20806# 0.0165f
C6576 a_10644_16791# sar9b_0.net6 0.22613f
C6577 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C6578 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.17533f
C6579 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[0] 0.26707f
C6580 sar9b_0.net23 sar9b_0.net41 0.03354f
C6581 a_8266_17113# sar9b_0.net46 0.13705f
C6582 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] 1.15113f
C6583 a_6250_28502# sar9b_0.net38 0.16677f
C6584 single_9b_cdac_0.SW[2] ua[0] 0.15413f
C6585 sar9b_0.net40 sar9b_0.net54 0.09214f
C6586 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.3196f
C6587 VDPWR a_12182_26419# 0.20236f
C6588 sar9b_0._04_ a_3027_21906# 0.24347f
C6589 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 2.82223f
C6590 sar9b_0.net53 a_12618_22138# 0.26166f
C6591 a_54032_17740# single_9b_cdac_1.SW[2] 0.18991f
C6592 a_8266_18445# sar9b_0.net46 0.14299f
C6593 VDPWR a_62748_26999# 1.81495f
C6594 sar9b_0.net6 a_12047_19857# 0.01561f
C6595 a_11466_23174# a_11658_22138# 0.01821f
C6596 VDPWR uo_out[3] 0.80535f
C6597 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.07579f
C6598 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[2] 2.01677f
C6599 sar9b_0.net65 a_4812_21738# 0.15545f
C6600 a_5812_21028# sar9b_0._11_ 0.06033f
C6601 a_6867_16810# a_7404_16784# 0.01177f
C6602 a_5711_17527# sar9b_0.net4 0.01409f
C6603 sar9b_0.net31 a_11658_26134# 0.02303f
C6604 sar9b_0.net5 a_7914_19178# 0.20518f
C6605 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.02513f
C6606 sar9b_0.net42 sar9b_0.net12 0.02691f
C6607 a_11382_18146# sar9b_0.net39 0.01041f
C6608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 a_25210_17740# 0.14695f
C6609 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.02618f
C6610 a_10607_25185# a_10402_25094# 0.09983f
C6611 single_9b_cdac_1.CF[0] ua[0] 3.29077f
C6612 a_11915_27039# single_9b_cdac_0.SW[4] 0.38596f
C6613 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[7] 3.85504f
C6614 sar9b_0.net40 a_10035_19474# 0.05886f
C6615 sar9b_0.net53 a_12618_23470# 0.26167f
C6616 VDPWR a_10644_16791# 0.84151f
C6617 sar9b_0.net43 sar9b_0.net60 0.02362f
C6618 a_10482_25831# a_10932_25713# 0.03432f
C6619 single_9b_cdac_1.CF[1] a_12435_20806# 0.35667f
C6620 sar9b_0.net53 a_10506_24506# 0.24393f
C6621 single_9b_cdac_0.SW[4] sar9b_0._06_ 0.22289f
C6622 sar9b_0.net61 a_10410_17846# 0.05361f
C6623 sar9b_0._01_ a_5126_20140# 0.2535f
C6624 single_9b_cdac_1.CF[2] single_9b_cdac_1.CF[0] 0.03575f
C6625 a_5506_17478# a_5046_17906# 0.26257f
C6626 a_5711_17527# a_5322_17846# 0.05462f
C6627 sar9b_0.net13 sar9b_0.net60 0.03465f
C6628 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22526f
C6629 sar9b_0.net49 a_9900_19047# 0.01024f
C6630 single_9b_cdac_1.CF[6] a_13011_24570# 0.35426f
C6631 VDPWR a_12047_19857# 0.26705f
C6632 th_dif_sw_0.th_sw_1.CK a_10166_3438# 0.04891f
C6633 a_14897_9355# th_dif_sw_0.VCN 0.05461f
C6634 sar9b_0.net53 sar9b_0.net27 0.03024f
C6635 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.28523f
C6636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A a_35519_15495# 0.01076f
C6637 sar9b_0.net43 a_5753_24250# 0.01111f
C6638 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[3] 0.26707f
C6639 single_9b_cdac_1.SW[2] ua[0] 0.14772f
C6640 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.03729f
C6641 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.84042f
C6642 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C6643 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.24371f
C6644 VDPWR sar9b_0.net20 0.27201f
C6645 sar9b_0.net13 a_5753_24250# 0.07055f
C6646 a_6834_20780# sar9b_0.net10 0.0738f
C6647 single_9b_cdac_0.SW[5] uo_out[2] 0.04146f
C6648 a_7402_22441# sar9b_0.net39 0.03886f
C6649 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.17533f
C6650 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.11216f
C6651 VDPWR a_3521_24240# 0.10938f
C6652 sar9b_0.net54 sar9b_0.net62 0.89973f
C6653 single_9b_cdac_1.CF[2] single_9b_cdac_1.SW[2] 1.79549f
C6654 VDPWR a_10239_19235# 0.26788f
C6655 sar9b_0.net38 single_9b_cdac_0.SW[8] 0.02501f
C6656 a_11842_18434# sar9b_0.net50 0.09528f
C6657 sar9b_0.net47 sar9b_0.net15 0.02183f
C6658 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] 1.56015f
C6659 a_11658_19474# sar9b_0.net50 0.19816f
C6660 sar9b_0.net10 a_7443_21496# 0.02366f
C6661 VDPWR a_9634_17478# 0.21868f
C6662 single_9b_cdac_1.SW[3] a_11842_18434# 0.10099f
C6663 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C6664 sar9b_0.net63 sar9b_0._13_ 0.05991f
C6665 a_11658_18142# a_12047_18525# 0.06034f
C6666 sar9b_0.net22 a_8691_28566# 0.2096f
C6667 a_11842_18434# a_12618_18142# 0.3578f
C6668 a_5298_24499# sar9b_0.net60 0.011f
C6669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.SW[0] 0.14962f
C6670 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38397f
C6671 sar9b_0._01_ sar9b_0.net4 0.03109f
C6672 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C6673 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.75899f
C6674 sar9b_0.cyclic_flag_0.FINAL sar9b_0.net37 0.17246f
C6675 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[6] 0.24288f
C6676 a_6282_27170# a_6880_26815# 0.06623f
C6677 a_11859_17910# sar9b_0.net2 0.11023f
C6678 a_5046_17906# sar9b_0.net4 0.01394f
C6679 sar9b_0._18_ sar9b_0.clk_div_0.COUNT\[2\] 0.71169f
C6680 VDPWR a_6250_28502# 0.29018f
C6681 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[3] 0.02038f
C6682 single_9b_cdac_1.CF[7] sar9b_0.net28 0.03957f
C6683 sar9b_0.net9 a_10230_23234# 0.03894f
C6684 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A 0.74663f
C6685 single_9b_cdac_1.SW[8] ua[0] 0.13942f
C6686 VDPWR a_5322_27170# 0.86299f
C6687 sar9b_0.net60 a_5126_20140# 0.02835f
C6688 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.26427f
C6689 a_5298_24499# a_5753_24250# 0.3578f
C6690 sar9b_0.net68 sar9b_0.net39 0.01595f
C6691 sar9b_0.net52 a_10742_25087# 0.12673f
C6692 ua[1] VGND 0.14595f
C6693 ua[2] VGND 0.14595f
C6694 ua[5] VGND 0.14595f
C6695 ua[6] VGND 0.14595f
C6696 ua[7] VGND 0.14595f
C6697 ena VGND 0.06982f
C6698 rst_n VGND 0.04231f
C6699 ui_in[1] VGND 0.04231f
C6700 ui_in[2] VGND 0.04231f
C6701 ui_in[3] VGND 0.04231f
C6702 ui_in[4] VGND 0.04231f
C6703 ui_in[5] VGND 0.04231f
C6704 ui_in[6] VGND 0.04231f
C6705 ui_in[7] VGND 0.04231f
C6706 uio_in[0] VGND 0.04231f
C6707 uio_in[1] VGND 0.04231f
C6708 uio_in[2] VGND 0.04231f
C6709 uio_in[3] VGND 0.04231f
C6710 uio_in[4] VGND 0.04231f
C6711 uio_in[5] VGND 0.04231f
C6712 uio_in[6] VGND 0.04231f
C6713 uio_in[7] VGND 0.04264f
C6714 ua[3] VGND 13.5574f
C6715 ua[4] VGND 13.4686f
C6716 clk VGND 28.193f
C6717 ui_in[0] VGND 17.1737f
C6718 uo_out[7] VGND 5.41879f
C6719 uo_out[1] VGND 4.49964f
C6720 uo_out[0] VGND 6.32256f
C6721 uo_out[2] VGND 4.375f
C6722 uo_out[3] VGND 4.4898f
C6723 uo_out[4] VGND 4.97269f
C6724 uo_out[6] VGND 5.39467f
C6725 uo_out[5] VGND 5.08381f
C6726 uio_out[0] VGND 5.71643f
C6727 uio_out[1] VGND 7.50245f
C6728 ua[0] VGND 0.11733p
C6729 VDPWR VGND 0.97985p
C6730 m2_23774_17236# VGND 0.24462f
C6731 m2_23774_26966# VGND 0.24462f
C6732 a_18214_3039# VGND 1.49705f $ **FLOATING
C6733 a_21684_3438# VGND 4.00493f $ **FLOATING
C6734 a_21368_4076# VGND 15.5335f $ **FLOATING
C6735 a_10254_2858# VGND 1.4958f $ **FLOATING
C6736 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VGND 3.32878f $ **FLOATING
C6737 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VGND 3.32496f $ **FLOATING
C6738 a_10482_3438# VGND 4.00493f $ **FLOATING
C6739 a_10166_3438# VGND 16.0184f $ **FLOATING
C6740 th_dif_sw_0.th_sw_1.CKB VGND 8.08199f $ **FLOATING
C6741 th_dif_sw_0.th_sw_1.CK VGND 9.07818f $ **FLOATING
C6742 a_21177_7457# VGND 2.80515f $ **FLOATING
C6743 a_9132_7271# VGND 2.80492f $ **FLOATING
C6744 a_17125_9355# VGND 0.09476f $ **FLOATING
C6745 a_14897_9355# VGND 0.09476f $ **FLOATING
C6746 th_dif_sw_0.VCP VGND 55.6678f $ **FLOATING
C6747 th_dif_sw_0.VCN VGND 67.3957f $ **FLOATING
C6748 a_16357_9613# VGND 0.05938f $ **FLOATING
C6749 a_15265_9613# VGND 0.05938f $ **FLOATING
C6750 a_16331_9671# VGND 0.82151f $ **FLOATING
C6751 a_14871_9671# VGND 0.82187f $ **FLOATING
C6752 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VGND 0.66688f $ **FLOATING
C6753 a_16881_10256# VGND 0.01123f $ **FLOATING
C6754 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VGND 0.66603f $ **FLOATING
C6755 a_15197_10290# VGND 0.01123f $ **FLOATING
C6756 a_16527_10454# VGND 0.18095f $ **FLOATING
C6757 a_15151_10456# VGND 0.18103f $ **FLOATING
C6758 a_16222_11316# VGND 0.04271f $ **FLOATING
C6759 a_15400_11316# VGND 0.04271f $ **FLOATING
C6760 tdc_0.phase_detector_0.INP VGND 1.24598f $ **FLOATING
C6761 tdc_0.phase_detector_0.INN VGND 1.87249f $ **FLOATING
C6762 a_16970_11404# VGND 0.20846f $ **FLOATING
C6763 a_15052_11404# VGND 0.20846f $ **FLOATING
C6764 tdc_0.phase_detector_0.pd_out_0.A VGND 2.40659f $ **FLOATING
C6765 tdc_0.phase_detector_0.pd_out_0.B VGND 1.65957f $ **FLOATING
C6766 a_16159_13315# VGND 0.26136f $ **FLOATING
C6767 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6768 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.41378f $ **FLOATING
C6769 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6770 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.45426f $ **FLOATING
C6771 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6772 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND 1.60512f $ **FLOATING
C6773 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND 1.57322f $ **FLOATING
C6774 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.39423f $ **FLOATING
C6775 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6776 a_63626_17740# VGND 0.89497f $ **FLOATING
C6777 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND 2.68117f $ **FLOATING
C6778 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6779 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6780 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6781 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6783 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND 3.19276f $ **FLOATING
C6784 a_62748_16877# VGND 0.16243f $ **FLOATING
C6785 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6787 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND 4.52812f $ **FLOATING
C6788 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND 94.0914f $ **FLOATING
C6789 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6790 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND 6.36367f $ **FLOATING
C6792 a_58824_17740# VGND 0.89548f $ **FLOATING
C6793 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND 2.66663f $ **FLOATING
C6794 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6795 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.405f $ **FLOATING
C6796 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6797 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44881f $ **FLOATING
C6798 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6799 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND 3.16257f $ **FLOATING
C6800 a_57946_16877# VGND 0.16243f $ **FLOATING
C6801 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND 1.58431f $ **FLOATING
C6802 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND 1.56057f $ **FLOATING
C6803 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND 4.51086f $ **FLOATING
C6804 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND 47.9165f $ **FLOATING
C6805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37225f $ **FLOATING
C6806 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6807 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND 6.34714f $ **FLOATING
C6808 a_54032_17740# VGND 0.89543f $ **FLOATING
C6809 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND 2.66664f $ **FLOATING
C6810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40542f $ **FLOATING
C6812 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6813 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44912f $ **FLOATING
C6814 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6815 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND 3.16256f $ **FLOATING
C6816 a_53154_16877# VGND 0.16243f $ **FLOATING
C6817 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND 1.58193f $ **FLOATING
C6818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND 1.56099f $ **FLOATING
C6819 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND 4.51373f $ **FLOATING
C6820 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND 30.3253f $ **FLOATING
C6821 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37352f $ **FLOATING
C6822 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6823 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND 6.34762f $ **FLOATING
C6824 a_49221_17740# VGND 0.89502f $ **FLOATING
C6825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND 2.66535f $ **FLOATING
C6826 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6827 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40525f $ **FLOATING
C6828 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6829 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44899f $ **FLOATING
C6830 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6831 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND 3.16312f $ **FLOATING
C6832 a_48343_16877# VGND 0.16243f $ **FLOATING
C6833 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND 1.58513f $ **FLOATING
C6834 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND 1.56081f $ **FLOATING
C6835 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND 4.51233f $ **FLOATING
C6836 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND 21.4947f $ **FLOATING
C6837 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37301f $ **FLOATING
C6838 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6839 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND 6.3477f $ **FLOATING
C6840 a_44418_17740# VGND 0.89497f $ **FLOATING
C6841 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND 2.665f $ **FLOATING
C6842 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6843 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6844 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6845 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6846 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6847 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND 3.16281f $ **FLOATING
C6848 a_43540_16877# VGND 0.16243f $ **FLOATING
C6849 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6850 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6851 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND 4.51195f $ **FLOATING
C6852 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND 20.61f $ **FLOATING
C6853 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6854 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6856 a_39616_17740# VGND 0.89497f $ **FLOATING
C6857 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND 2.66616f $ **FLOATING
C6858 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6859 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6860 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6861 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6862 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6863 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6864 a_38738_16877# VGND 0.16243f $ **FLOATING
C6865 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6866 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6867 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND 4.51201f $ **FLOATING
C6868 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND 16.1449f $ **FLOATING
C6869 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6870 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6871 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6872 a_34814_17740# VGND 0.89548f $ **FLOATING
C6873 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND 2.66683f $ **FLOATING
C6874 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6875 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6876 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6877 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6878 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6879 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6880 a_33936_16877# VGND 0.16243f $ **FLOATING
C6881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6882 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND 4.51252f $ **FLOATING
C6884 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND 15.6371f $ **FLOATING
C6885 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6886 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6888 a_30012_17740# VGND 0.89497f $ **FLOATING
C6889 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND 2.66498f $ **FLOATING
C6890 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6891 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6892 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6893 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6894 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6895 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6896 a_29134_16877# VGND 0.16243f $ **FLOATING
C6897 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6898 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6899 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND 4.51193f $ **FLOATING
C6900 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND 14.5496f $ **FLOATING
C6901 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6902 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6903 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND 6.34748f $ **FLOATING
C6904 a_25210_17740# VGND 0.89548f $ **FLOATING
C6905 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND 2.68106f $ **FLOATING
C6906 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND 3.16216f $ **FLOATING
C6907 a_24332_16877# VGND 0.16243f $ **FLOATING
C6908 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND 4.71828f $ **FLOATING
C6909 single_9b_cdac_1.SW[5] VGND 6.60196f $ **FLOATING
C6910 a_13011_16810# VGND 0.63654f $ **FLOATING
C6911 tdc_0.OUTP VGND 3.42864f $ **FLOATING
C6912 a_12588_16784# VGND 0.3641f $ **FLOATING
C6913 a_11434_16874# VGND 0.16615f $ **FLOATING
C6914 a_10926_17021# VGND 0.17322f $ **FLOATING
C6915 a_10858_17113# VGND 0.13557f $ **FLOATING
C6916 a_10649_17131# VGND 0.93597f $ **FLOATING
C6917 a_10335_16817# VGND 0.30597f $ **FLOATING
C6918 a_10194_16784# VGND 0.35867f $ **FLOATING
C6919 a_10644_16791# VGND 0.61756f $ **FLOATING
C6920 a_9996_16784# VGND 0.3018f $ **FLOATING
C6921 a_8842_16874# VGND 0.13599f $ **FLOATING
C6922 a_8334_17021# VGND 0.17338f $ **FLOATING
C6923 a_8266_17113# VGND 0.13376f $ **FLOATING
C6924 a_8057_17131# VGND 0.92848f $ **FLOATING
C6925 a_7743_16817# VGND 0.30616f $ **FLOATING
C6926 a_7602_16784# VGND 0.36252f $ **FLOATING
C6927 a_8052_16791# VGND 0.6075f $ **FLOATING
C6928 a_7404_16784# VGND 0.30035f $ **FLOATING
C6929 a_6867_16810# VGND 0.38007f $ **FLOATING
C6930 tdc_0.OUTN VGND 5.01507f $ **FLOATING
C6931 a_5331_16810# VGND 0.38321f $ **FLOATING
C6932 tdc_0.RDY VGND 6.15869f $ **FLOATING
C6933 th_dif_sw_0.CKB VGND 16.3637f $ **FLOATING
C6934 a_2603_17006# VGND 0.67873f $ **FLOATING
C6935 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND 13.6188f $ **FLOATING
C6936 single_9b_cdac_1.SW[6] VGND 6.72589f $ **FLOATING
C6937 a_13011_17910# VGND 0.63061f $ **FLOATING
C6938 single_9b_cdac_1.SW[4] VGND 6.88153f $ **FLOATING
C6939 a_11859_17910# VGND 0.6882f $ **FLOATING
C6940 a_11436_17742# VGND 0.33062f $ **FLOATING
C6941 a_11008_17491# VGND 0.27893f $ **FLOATING
C6942 a_10662_17799# VGND 0.29366f $ **FLOATING
C6943 a_10410_17846# VGND 0.34331f $ **FLOATING
C6944 a_9974_17626# VGND 0.1176f $ **FLOATING
C6945 a_9839_17527# VGND 0.15642f $ **FLOATING
C6946 a_9634_17478# VGND 0.88707f $ **FLOATING
C6947 a_9174_17906# VGND 0.1327f $ **FLOATING
C6948 a_9450_17846# VGND 0.59308f $ **FLOATING
C6949 single_9b_cdac_1.SW[0] VGND 15.1733f $ **FLOATING
C6950 single_9b_cdac_1.SW[2] VGND 7.72854f $ **FLOATING
C6951 a_8595_17910# VGND 0.5964f $ **FLOATING
C6952 a_8019_17910# VGND 0.60315f $ **FLOATING
C6953 a_7404_17715# VGND 0.24299f $ **FLOATING
C6954 a_6880_17491# VGND 0.29519f $ **FLOATING
C6955 a_6534_17799# VGND 0.31348f $ **FLOATING
C6956 a_6282_17846# VGND 0.36418f $ **FLOATING
C6957 a_5846_17626# VGND 0.1724f $ **FLOATING
C6958 a_5711_17527# VGND 0.19862f $ **FLOATING
C6959 a_5506_17478# VGND 0.95291f $ **FLOATING
C6960 a_5046_17906# VGND 0.14415f $ **FLOATING
C6961 a_5322_17846# VGND 0.6425f $ **FLOATING
C6962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND 6.37641f $ **FLOATING
C6963 a_12047_18525# VGND 0.1897f $ **FLOATING
C6964 a_13216_18477# VGND 0.28599f $ **FLOATING
C6965 a_12618_18142# VGND 0.35255f $ **FLOATING
C6966 a_12870_18271# VGND 0.29854f $ **FLOATING
C6967 a_12182_18427# VGND 0.1325f $ **FLOATING
C6968 a_11842_18434# VGND 0.9417f $ **FLOATING
C6969 a_11658_18142# VGND 0.67802f $ **FLOATING
C6970 a_11382_18146# VGND 0.1608f $ **FLOATING
C6971 single_9b_cdac_1.SW[3] VGND 8.35662f $ **FLOATING
C6972 th_dif_sw_0.CK VGND 10.2695f $ **FLOATING
C6973 a_10803_18142# VGND 0.61263f $ **FLOATING
C6974 a_10227_18142# VGND 0.62055f $ **FLOATING
C6975 a_8842_18206# VGND 0.12267f $ **FLOATING
C6976 a_8334_18353# VGND 0.15504f $ **FLOATING
C6977 a_8266_18445# VGND 0.11469f $ **FLOATING
C6978 a_8057_18463# VGND 0.88109f $ **FLOATING
C6979 a_7743_18149# VGND 0.29328f $ **FLOATING
C6980 a_7602_18116# VGND 0.33292f $ **FLOATING
C6981 a_8052_18123# VGND 0.56532f $ **FLOATING
C6982 a_7404_18116# VGND 0.27413f $ **FLOATING
C6983 a_6634_18206# VGND 0.15117f $ **FLOATING
C6984 a_6126_18353# VGND 0.19104f $ **FLOATING
C6985 a_6058_18445# VGND 0.16799f $ **FLOATING
C6986 a_5849_18463# VGND 0.98369f $ **FLOATING
C6987 a_5535_18149# VGND 0.31139f $ **FLOATING
C6988 a_5394_18116# VGND 0.39633f $ **FLOATING
C6989 a_5844_18123# VGND 0.62179f $ **FLOATING
C6990 a_5196_18116# VGND 0.28271f $ **FLOATING
C6991 a_4771_18260# VGND 0.50939f $ **FLOATING
C6992 single_9b_cdac_1.SW[7] VGND 6.05886f $ **FLOATING
C6993 a_13011_19242# VGND 0.63648f $ **FLOATING
C6994 a_11338_19178# VGND 0.17146f $ **FLOATING
C6995 a_10762_18823# VGND 0.12318f $ **FLOATING
C6996 a_10830_19068# VGND 0.1661f $ **FLOATING
C6997 a_10553_18922# VGND 0.91659f $ **FLOATING
C6998 a_10548_19053# VGND 0.59692f $ **FLOATING
C6999 a_10239_19235# VGND 0.2919f $ **FLOATING
C7000 a_10098_19171# VGND 0.34247f $ **FLOATING
C7001 a_9900_19047# VGND 0.28365f $ **FLOATING
C7002 a_9472_18823# VGND 0.27623f $ **FLOATING
C7003 a_9126_19131# VGND 0.29177f $ **FLOATING
C7004 a_8874_19178# VGND 0.34094f $ **FLOATING
C7005 a_8438_18958# VGND 0.13218f $ **FLOATING
C7006 a_8303_18859# VGND 0.17139f $ **FLOATING
C7007 a_8098_18810# VGND 0.9231f $ **FLOATING
C7008 a_7638_19238# VGND 0.13759f $ **FLOATING
C7009 a_7914_19178# VGND 0.58482f $ **FLOATING
C7010 a_6579_18832# VGND 0.45588f $ **FLOATING
C7011 a_6252_19074# VGND 0.32141f $ **FLOATING
C7012 a_5811_19178# VGND 0.27961f $ **FLOATING
C7013 a_5443_19074# VGND 0.44526f $ **FLOATING
C7014 a_12047_19857# VGND 0.19066f $ **FLOATING
C7015 a_13216_19809# VGND 0.29524f $ **FLOATING
C7016 a_12618_19474# VGND 0.35239f $ **FLOATING
C7017 a_12870_19603# VGND 0.29287f $ **FLOATING
C7018 a_12182_19759# VGND 0.13111f $ **FLOATING
C7019 a_11842_19766# VGND 0.96526f $ **FLOATING
C7020 a_11658_19474# VGND 0.62067f $ **FLOATING
C7021 a_11382_19478# VGND 0.17055f $ **FLOATING
C7022 single_9b_cdac_1.SW[1] VGND 7.77706f $ **FLOATING
C7023 sar9b_0.net48 VGND 3.00596f $ **FLOATING
C7024 a_10803_19474# VGND 0.61976f $ **FLOATING
C7025 a_10035_19474# VGND 0.62781f $ **FLOATING
C7026 a_7882_19538# VGND 0.1244f $ **FLOATING
C7027 a_7374_19685# VGND 0.15921f $ **FLOATING
C7028 a_7306_19777# VGND 0.1167f $ **FLOATING
C7029 a_5761_19487# VGND 0.01222f $ **FLOATING
C7030 a_7097_19795# VGND 0.88857f $ **FLOATING
C7031 a_6783_19481# VGND 0.29276f $ **FLOATING
C7032 a_6642_19448# VGND 0.34651f $ **FLOATING
C7033 a_5628_19768# VGND 0.01308f $ **FLOATING
C7034 a_7092_19455# VGND 0.59664f $ **FLOATING
C7035 a_6444_19448# VGND 0.28777f $ **FLOATING
C7036 a_5581_19664# VGND 0.29099f $ **FLOATING
C7037 a_5196_19448# VGND 0.34938f $ **FLOATING
C7038 a_4072_19474# VGND 0.47181f $ **FLOATING
C7039 a_3795_19512# VGND 0.2312f $ **FLOATING
C7040 sar9b_0.net46 VGND 3.29711f $ **FLOATING
C7041 sar9b_0.net71 VGND 0.32339f $ **FLOATING
C7042 a_3180_19448# VGND 0.35853f $ **FLOATING
C7043 sar9b_0.net50 VGND 1.2487f $ **FLOATING
C7044 a_13011_20574# VGND 0.61397f $ **FLOATING
C7045 sar9b_0.net5 VGND 1.48438f $ **FLOATING
C7046 a_12684_20379# VGND 0.25006f $ **FLOATING
C7047 single_9b_cdac_1.SW[8] VGND 6.02413f $ **FLOATING
C7048 a_11859_20574# VGND 0.71415f $ **FLOATING
C7049 a_10528_20155# VGND 0.29045f $ **FLOATING
C7050 a_10182_20463# VGND 0.30322f $ **FLOATING
C7051 a_9930_20510# VGND 0.34846f $ **FLOATING
C7052 a_9494_20290# VGND 0.13056f $ **FLOATING
C7053 a_9359_20191# VGND 0.16916f $ **FLOATING
C7054 a_9154_20142# VGND 0.92156f $ **FLOATING
C7055 a_8694_20570# VGND 0.13812f $ **FLOATING
C7056 a_8970_20510# VGND 0.66102f $ **FLOATING
C7057 sar9b_0.net15 VGND 0.46616f $ **FLOATING
C7058 a_6130_20239# VGND 0.46131f $ **FLOATING
C7059 a_5931_20140# VGND 0.28737f $ **FLOATING
C7060 a_5481_20185# VGND 0.15828f $ **FLOATING
C7061 a_5633_20244# VGND 0.20547f $ **FLOATING
C7062 a_5374_20145# VGND 0.01758f $ **FLOATING
C7063 a_4496_20468# VGND 0.17016f $ **FLOATING
C7064 sar9b_0._10_ VGND 0.37869f $ **FLOATING
C7065 a_5126_20140# VGND 0.71166f $ **FLOATING
C7066 a_4947_20140# VGND 1.23378f $ **FLOATING
C7067 sar9b_0.net16 VGND 1.53593f $ **FLOATING
C7068 a_3922_20239# VGND 0.41543f $ **FLOATING
C7069 a_3723_20140# VGND 0.24243f $ **FLOATING
C7070 a_3273_20185# VGND 0.15798f $ **FLOATING
C7071 a_3425_20244# VGND 0.18716f $ **FLOATING
C7072 a_3166_20145# VGND 0.02072f $ **FLOATING
C7073 sar9b_0._00_ VGND 0.34642f $ **FLOATING
C7074 a_2918_20140# VGND 0.66229f $ **FLOATING
C7075 a_2739_20140# VGND 1.25389f $ **FLOATING
C7076 a_10607_21189# VGND 0.16031f $ **FLOATING
C7077 a_13011_20806# VGND 0.62155f $ **FLOATING
C7078 a_12435_20806# VGND 0.63677f $ **FLOATING
C7079 sar9b_0.net6 VGND 1.99773f $ **FLOATING
C7080 a_11776_21141# VGND 0.31771f $ **FLOATING
C7081 a_11178_20806# VGND 0.34832f $ **FLOATING
C7082 a_11430_20935# VGND 0.29503f $ **FLOATING
C7083 a_10742_21091# VGND 0.11828f $ **FLOATING
C7084 a_10402_21098# VGND 0.89532f $ **FLOATING
C7085 a_10218_20806# VGND 0.58532f $ **FLOATING
C7086 a_9942_20810# VGND 0.14176f $ **FLOATING
C7087 a_9363_20826# VGND 0.45753f $ **FLOATING
C7088 sar9b_0.net56 VGND 1.44734f $ **FLOATING
C7089 a_8074_20870# VGND 0.14861f $ **FLOATING
C7090 a_7566_21017# VGND 0.17208f $ **FLOATING
C7091 a_7498_21109# VGND 0.13435f $ **FLOATING
C7092 a_5183_20819# VGND 0.01178f $ **FLOATING
C7093 a_7289_21127# VGND 0.92471f $ **FLOATING
C7094 a_6975_20813# VGND 0.30878f $ **FLOATING
C7095 a_6834_20780# VGND 0.37224f $ **FLOATING
C7096 sar9b_0._01_ VGND 0.97665f $ **FLOATING
C7097 a_7284_20787# VGND 0.60133f $ **FLOATING
C7098 a_6636_20780# VGND 0.29286f $ **FLOATING
C7099 sar9b_0._11_ VGND 0.67367f $ **FLOATING
C7100 a_6252_20780# VGND 0.39203f $ **FLOATING
C7101 a_5812_21028# VGND 0.3166f $ **FLOATING
C7102 sar9b_0._08_ VGND 0.57215f $ **FLOATING
C7103 sar9b_0._09_ VGND 0.59924f $ **FLOATING
C7104 a_5581_20992# VGND 0.30562f $ **FLOATING
C7105 a_4922_20857# VGND 0.24594f $ **FLOATING
C7106 a_2508_20780# VGND 2.7729f $ **FLOATING
C7107 a_13011_21906# VGND 0.63044f $ **FLOATING
C7108 a_11859_21906# VGND 0.72107f $ **FLOATING
C7109 sar9b_0.net7 VGND 1.24263f $ **FLOATING
C7110 a_10816_21487# VGND 0.30071f $ **FLOATING
C7111 a_10470_21795# VGND 0.3024f $ **FLOATING
C7112 a_10218_21842# VGND 0.34969f $ **FLOATING
C7113 a_9782_21622# VGND 0.13363f $ **FLOATING
C7114 a_9647_21523# VGND 0.17263f $ **FLOATING
C7115 a_9442_21474# VGND 0.92619f $ **FLOATING
C7116 a_8982_21902# VGND 0.13981f $ **FLOATING
C7117 a_9258_21842# VGND 0.60132f $ **FLOATING
C7118 sar9b_0.net49 VGND 2.18775f $ **FLOATING
C7119 sar9b_0.net8 VGND 3.73402f $ **FLOATING
C7120 a_7443_21496# VGND 0.49853f $ **FLOATING
C7121 sar9b_0.net51 VGND 2.5769f $ **FLOATING
C7122 a_6444_21738# VGND 0.39129f $ **FLOATING
C7123 a_5523_21528# VGND 0.30787f $ **FLOATING
C7124 a_4812_21738# VGND 0.38426f $ **FLOATING
C7125 a_4236_21738# VGND 0.35329f $ **FLOATING
C7126 a_3027_21906# VGND 0.35644f $ **FLOATING
C7127 a_12047_22521# VGND 0.20349f $ **FLOATING
C7128 a_13216_22473# VGND 0.29599f $ **FLOATING
C7129 a_12618_22138# VGND 0.36248f $ **FLOATING
C7130 a_12870_22267# VGND 0.30878f $ **FLOATING
C7131 a_12182_22423# VGND 0.1466f $ **FLOATING
C7132 a_11842_22430# VGND 0.97398f $ **FLOATING
C7133 a_11658_22138# VGND 0.64577f $ **FLOATING
C7134 a_11382_22142# VGND 0.15492f $ **FLOATING
C7135 sar9b_0.net73 VGND 2.09299f $ **FLOATING
C7136 sar9b_0.net61 VGND 3.33314f $ **FLOATING
C7137 a_7978_22202# VGND 0.12351f $ **FLOATING
C7138 a_7470_22349# VGND 0.15862f $ **FLOATING
C7139 a_7402_22441# VGND 0.11773f $ **FLOATING
C7140 a_7193_22459# VGND 0.888f $ **FLOATING
C7141 a_6879_22145# VGND 0.29152f $ **FLOATING
C7142 sar9b_0.net47 VGND 2.48893f $ **FLOATING
C7143 a_6738_22112# VGND 0.33464f $ **FLOATING
C7144 a_5739_22488# VGND 0.25938f $ **FLOATING
C7145 a_5182_22567# VGND 0.01826f $ **FLOATING
C7146 a_7188_22119# VGND 0.58869f $ **FLOATING
C7147 a_6540_22112# VGND 0.2837f $ **FLOATING
C7148 a_5938_22378# VGND 0.43981f $ **FLOATING
C7149 a_5289_22527# VGND 0.1531f $ **FLOATING
C7150 a_5441_22522# VGND 0.18149f $ **FLOATING
C7151 sar9b_0.net64 VGND 1.22538f $ **FLOATING
C7152 a_4934_22432# VGND 0.65617f $ **FLOATING
C7153 a_4755_22138# VGND 1.27206f $ **FLOATING
C7154 sar9b_0.clk_div_0.COUNT\[3\] VGND 0.68828f $ **FLOATING
C7155 a_4011_22488# VGND 0.2324f $ **FLOATING
C7156 a_3454_22567# VGND 0.01679f $ **FLOATING
C7157 a_4210_22378# VGND 0.40953f $ **FLOATING
C7158 a_3561_22527# VGND 0.15284f $ **FLOATING
C7159 a_3713_22522# VGND 0.18104f $ **FLOATING
C7160 sar9b_0.net67 VGND 0.81321f $ **FLOATING
C7161 a_3206_22432# VGND 0.66139f $ **FLOATING
C7162 sar9b_0._05_ VGND 0.79927f $ **FLOATING
C7163 sar9b_0._04_ VGND 0.78117f $ **FLOATING
C7164 a_3027_22138# VGND 1.2701f $ **FLOATING
C7165 sar9b_0.clknet_1_0__leaf_CLK VGND 1.92116f $ **FLOATING
C7166 a_13011_23238# VGND 0.6362f $ **FLOATING
C7167 a_12064_22819# VGND 0.32582f $ **FLOATING
C7168 a_11718_23127# VGND 0.32104f $ **FLOATING
C7169 a_11466_23174# VGND 0.37219f $ **FLOATING
C7170 a_11030_22954# VGND 0.1247f $ **FLOATING
C7171 a_10895_22855# VGND 0.16542f $ **FLOATING
C7172 a_10690_22806# VGND 0.91522f $ **FLOATING
C7173 a_10230_23234# VGND 0.13716f $ **FLOATING
C7174 a_10506_23174# VGND 0.64615f $ **FLOATING
C7175 sar9b_0.net9 VGND 2.28378f $ **FLOATING
C7176 a_9760_22819# VGND 0.28806f $ **FLOATING
C7177 a_9414_23127# VGND 0.2958f $ **FLOATING
C7178 a_9162_23174# VGND 0.35069f $ **FLOATING
C7179 a_8726_22954# VGND 0.12072f $ **FLOATING
C7180 a_8591_22855# VGND 0.15931f $ **FLOATING
C7181 a_8386_22806# VGND 0.90687f $ **FLOATING
C7182 a_7926_23234# VGND 0.13601f $ **FLOATING
C7183 a_8202_23174# VGND 0.60825f $ **FLOATING
C7184 a_7597_23174# VGND 0.01081f $ **FLOATING
C7185 sar9b_0._17_ VGND 0.54536f $ **FLOATING
C7186 a_6744_23238# VGND 0.27119f $ **FLOATING
C7187 sar9b_0._02_ VGND 0.50023f $ **FLOATING
C7188 a_6861_22828# VGND 0.22749f $ **FLOATING
C7189 a_6484_22845# VGND 0.38938f $ **FLOATING
C7190 sar9b_0._12_ VGND 2.03947f $ **FLOATING
C7191 a_4332_23043# VGND 2.49415f $ **FLOATING
C7192 sar9b_0.clk_div_0.COUNT\[0\] VGND 0.5303f $ **FLOATING
C7193 sar9b_0._07_ VGND 3.63856f $ **FLOATING
C7194 sar9b_0.net66 VGND 0.36733f $ **FLOATING
C7195 sar9b_0.net65 VGND 1.04893f $ **FLOATING
C7196 a_3695_23038# VGND 0.27588f $ **FLOATING
C7197 a_3219_22860# VGND 0.23516f $ **FLOATING
C7198 a_3371_23106# VGND 0.25044f $ **FLOATING
C7199 sar9b_0._18_ VGND 0.52436f $ **FLOATING
C7200 a_2892_23070# VGND 0.3304f $ **FLOATING
C7201 a_12047_23853# VGND 0.20399f $ **FLOATING
C7202 a_13216_23805# VGND 0.29598f $ **FLOATING
C7203 a_12618_23470# VGND 0.36236f $ **FLOATING
C7204 a_12870_23599# VGND 0.3087f $ **FLOATING
C7205 a_12182_23755# VGND 0.14911f $ **FLOATING
C7206 a_11842_23762# VGND 0.97787f $ **FLOATING
C7207 a_11658_23470# VGND 0.66469f $ **FLOATING
C7208 a_11382_23474# VGND 0.15995f $ **FLOATING
C7209 a_10707_23470# VGND 0.36843f $ **FLOATING
C7210 sar9b_0.net1 VGND 2.40289f $ **FLOATING
C7211 a_10227_23490# VGND 0.467f $ **FLOATING
C7212 a_8303_23853# VGND 0.16637f $ **FLOATING
C7213 a_9472_23805# VGND 0.29613f $ **FLOATING
C7214 a_8874_23470# VGND 0.35331f $ **FLOATING
C7215 a_9126_23599# VGND 0.29994f $ **FLOATING
C7216 a_8438_23755# VGND 0.13265f $ **FLOATING
C7217 a_8098_23762# VGND 0.9183f $ **FLOATING
C7218 a_7914_23470# VGND 0.6159f $ **FLOATING
C7219 a_7638_23474# VGND 0.11866f $ **FLOATING
C7220 sar9b_0.net10 VGND 1.74489f $ **FLOATING
C7221 a_6922_23534# VGND 0.11783f $ **FLOATING
C7222 a_6414_23681# VGND 0.16683f $ **FLOATING
C7223 a_6346_23773# VGND 0.12324f $ **FLOATING
C7224 a_6137_23791# VGND 0.93229f $ **FLOATING
C7225 a_5823_23477# VGND 0.31555f $ **FLOATING
C7226 a_5682_23444# VGND 0.37293f $ **FLOATING
C7227 a_6132_23451# VGND 0.58878f $ **FLOATING
C7228 a_5484_23444# VGND 0.29255f $ **FLOATING
C7229 a_4811_23656# VGND 0.28975f $ **FLOATING
C7230 sar9b_0.clknet_0_CLK VGND 2.22837f $ **FLOATING
C7231 a_2508_23444# VGND 2.77512f $ **FLOATING
C7232 a_13011_24570# VGND 0.62981f $ **FLOATING
C7233 sar9b_0.net11 VGND 3.57213f $ **FLOATING
C7234 a_11104_24151# VGND 0.30915f $ **FLOATING
C7235 a_10758_24459# VGND 0.303f $ **FLOATING
C7236 a_10506_24506# VGND 0.35537f $ **FLOATING
C7237 a_10070_24286# VGND 0.13107f $ **FLOATING
C7238 a_9935_24187# VGND 0.16193f $ **FLOATING
C7239 a_9730_24138# VGND 0.91556f $ **FLOATING
C7240 a_9270_24566# VGND 0.1136f $ **FLOATING
C7241 a_9546_24506# VGND 0.60387f $ **FLOATING
C7242 sar9b_0.net2 VGND 1.31622f $ **FLOATING
C7243 a_8940_24402# VGND 0.33197f $ **FLOATING
C7244 a_7347_24160# VGND 0.51748f $ **FLOATING
C7245 sar9b_0.net55 VGND 1.13897f $ **FLOATING
C7246 sar9b_0.net62 VGND 1.27467f $ **FLOATING
C7247 a_6538_24506# VGND 0.1602f $ **FLOATING
C7248 a_5962_24151# VGND 0.17011f $ **FLOATING
C7249 a_6030_24396# VGND 0.20052f $ **FLOATING
C7250 a_5753_24250# VGND 0.95497f $ **FLOATING
C7251 a_5748_24381# VGND 0.60642f $ **FLOATING
C7252 a_5439_24563# VGND 0.30942f $ **FLOATING
C7253 a_4467_24162# VGND 0.1655f $ **FLOATING
C7254 sar9b_0._13_ VGND 0.30005f $ **FLOATING
C7255 a_5298_24499# VGND 0.38655f $ **FLOATING
C7256 a_5100_24375# VGND 0.29673f $ **FLOATING
C7257 a_4018_24235# VGND 0.41892f $ **FLOATING
C7258 a_3819_24136# VGND 0.2435f $ **FLOATING
C7259 a_3369_24181# VGND 0.15303f $ **FLOATING
C7260 a_3521_24240# VGND 0.18898f $ **FLOATING
C7261 a_3262_24141# VGND 0.02073f $ **FLOATING
C7262 sar9b_0.net70 VGND 0.58889f $ **FLOATING
C7263 a_3014_24136# VGND 0.63058f $ **FLOATING
C7264 a_2835_24136# VGND 1.26692f $ **FLOATING
C7265 a_10607_25185# VGND 0.16691f $ **FLOATING
C7266 a_13011_24802# VGND 0.62905f $ **FLOATING
C7267 sar9b_0.net26 VGND 2.14803f $ **FLOATING
C7268 a_12435_24802# VGND 0.64526f $ **FLOATING
C7269 a_11776_25137# VGND 0.32738f $ **FLOATING
C7270 a_11178_24802# VGND 0.35816f $ **FLOATING
C7271 a_11430_24931# VGND 0.30602f $ **FLOATING
C7272 a_10742_25087# VGND 0.13219f $ **FLOATING
C7273 a_10402_25094# VGND 0.91973f $ **FLOATING
C7274 a_10218_24802# VGND 0.5916f $ **FLOATING
C7275 sar9b_0.net57 VGND 2.74111f $ **FLOATING
C7276 a_9942_24806# VGND 0.1549f $ **FLOATING
C7277 sar9b_0.net53 VGND 2.57915f $ **FLOATING
C7278 a_6767_25185# VGND 0.17399f $ **FLOATING
C7279 a_9165_24988# VGND 0.47483f $ **FLOATING
C7280 a_7936_25137# VGND 0.3013f $ **FLOATING
C7281 a_7338_24802# VGND 0.35928f $ **FLOATING
C7282 a_7590_24931# VGND 0.30299f $ **FLOATING
C7283 a_6902_25087# VGND 0.1354f $ **FLOATING
C7284 a_6562_25094# VGND 0.92936f $ **FLOATING
C7285 a_6378_24802# VGND 0.661f $ **FLOATING
C7286 sar9b_0.net4 VGND 1.56917f $ **FLOATING
C7287 a_6102_24806# VGND 0.15486f $ **FLOATING
C7288 sar9b_0.net54 VGND 2.72635f $ **FLOATING
C7289 sar9b_0._15_ VGND 0.7538f $ **FLOATING
C7290 a_5580_24776# VGND 0.35113f $ **FLOATING
C7291 sar9b_0.clk_div_0.COUNT\[2\] VGND 0.9962f $ **FLOATING
C7292 a_5196_24776# VGND 0.33541f $ **FLOATING
C7293 a_4044_24776# VGND 0.344f $ **FLOATING
C7294 sar9b_0.net68 VGND 0.89917f $ **FLOATING
C7295 sar9b_0._14_ VGND 0.97587f $ **FLOATING
C7296 a_2893_24992# VGND 0.22912f $ **FLOATING
C7297 sar9b_0.net72 VGND 1.71102f $ **FLOATING
C7298 sar9b_0.net63 VGND 1.46347f $ **FLOATING
C7299 a_13011_25902# VGND 0.63761f $ **FLOATING
C7300 a_11722_25838# VGND 0.17423f $ **FLOATING
C7301 sar9b_0.net13 VGND 1.83091f $ **FLOATING
C7302 a_11146_25483# VGND 0.13526f $ **FLOATING
C7303 a_11214_25728# VGND 0.17226f $ **FLOATING
C7304 a_10937_25582# VGND 0.93944f $ **FLOATING
C7305 a_10932_25713# VGND 0.63975f $ **FLOATING
C7306 a_10623_25895# VGND 0.30445f $ **FLOATING
C7307 a_10482_25831# VGND 0.35993f $ **FLOATING
C7308 a_10284_25707# VGND 0.30192f $ **FLOATING
C7309 sar9b_0.clknet_1_1__leaf_CLK VGND 1.99526f $ **FLOATING
C7310 a_4698_25851# VGND 0.02231f $ **FLOATING
C7311 sar9b_0._03_ VGND 0.34487f $ **FLOATING
C7312 a_4293_25852# VGND 0.18854f $ **FLOATING
C7313 a_4365_25770# VGND 0.16167f $ **FLOATING
C7314 a_4136_25584# VGND 0.6886f $ **FLOATING
C7315 sar9b_0.clk_div_0.COUNT\[1\] VGND 1.70819f $ **FLOATING
C7316 sar9b_0.net69 VGND 1.15997f $ **FLOATING
C7317 a_4125_25958# VGND 1.27131f $ **FLOATING
C7318 a_3855_25792# VGND 0.24272f $ **FLOATING
C7319 a_3747_25724# VGND 0.41638f $ **FLOATING
C7320 sar9b_0._16_ VGND 0.40855f $ **FLOATING
C7321 a_3372_25734# VGND 0.33769f $ **FLOATING
C7322 a_12047_26517# VGND 0.19151f $ **FLOATING
C7323 a_13216_26469# VGND 0.28884f $ **FLOATING
C7324 a_12618_26134# VGND 0.35065f $ **FLOATING
C7325 a_12870_26263# VGND 0.29813f $ **FLOATING
C7326 a_12182_26419# VGND 0.13385f $ **FLOATING
C7327 a_11842_26426# VGND 0.96869f $ **FLOATING
C7328 a_11658_26134# VGND 0.62093f $ **FLOATING
C7329 sar9b_0.net12 VGND 1.66742f $ **FLOATING
C7330 a_11382_26138# VGND 0.14597f $ **FLOATING
C7331 sar9b_0.net74 VGND 1.58493f $ **FLOATING
C7332 sar9b_0.net33 VGND 1.05333f $ **FLOATING
C7333 a_10859_26330# VGND 0.61787f $ **FLOATING
C7334 sar9b_0.net41 VGND 2.17416f $ **FLOATING
C7335 a_9130_26198# VGND 0.15692f $ **FLOATING
C7336 a_8622_26345# VGND 0.17118f $ **FLOATING
C7337 a_8554_26437# VGND 0.13269f $ **FLOATING
C7338 a_8345_26455# VGND 0.92555f $ **FLOATING
C7339 a_8031_26141# VGND 0.30485f $ **FLOATING
C7340 a_7890_26108# VGND 0.35529f $ **FLOATING
C7341 a_8340_26115# VGND 0.61091f $ **FLOATING
C7342 a_7692_26108# VGND 0.30296f $ **FLOATING
C7343 sar9b_0.net35 VGND 2.44446f $ **FLOATING
C7344 a_3946_26198# VGND 0.15782f $ **FLOATING
C7345 a_3438_26345# VGND 0.17121f $ **FLOATING
C7346 a_3370_26437# VGND 0.13251f $ **FLOATING
C7347 a_3161_26455# VGND 0.9217f $ **FLOATING
C7348 a_2847_26141# VGND 0.3046f $ **FLOATING
C7349 a_2706_26108# VGND 0.36022f $ **FLOATING
C7350 a_3156_26115# VGND 0.59376f $ **FLOATING
C7351 a_2508_26108# VGND 0.30075f $ **FLOATING
C7352 a_63626_26990# VGND 0.89497f $ **FLOATING
C7353 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND 2.68117f $ **FLOATING
C7354 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND 3.19275f $ **FLOATING
C7355 a_62748_26999# VGND 0.16243f $ **FLOATING
C7356 single_9b_cdac_0.SW[0] VGND 11.0253f $ **FLOATING
C7357 a_58824_26990# VGND 0.89548f $ **FLOATING
C7358 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND 2.66663f $ **FLOATING
C7359 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND 6.36459f $ **FLOATING
C7360 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.39423f $ **FLOATING
C7361 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7362 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.45426f $ **FLOATING
C7363 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7364 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND 1.57322f $ **FLOATING
C7365 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND 1.60512f $ **FLOATING
C7366 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND 94.5927f $ **FLOATING
C7367 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND 3.16256f $ **FLOATING
C7368 a_57946_26999# VGND 0.16243f $ **FLOATING
C7369 a_54032_26990# VGND 0.89543f $ **FLOATING
C7370 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND 2.66664f $ **FLOATING
C7371 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND 6.34807f $ **FLOATING
C7372 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7374 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7375 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7376 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND 4.52773f $ **FLOATING
C7377 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7378 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.41378f $ **FLOATING
C7380 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7381 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND 47.9165f $ **FLOATING
C7382 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND 3.16255f $ **FLOATING
C7383 a_53154_26999# VGND 0.16243f $ **FLOATING
C7384 a_49221_26990# VGND 0.89502f $ **FLOATING
C7385 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND 2.66535f $ **FLOATING
C7386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND 6.34853f $ **FLOATING
C7387 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37221f $ **FLOATING
C7388 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7389 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44881f $ **FLOATING
C7390 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7391 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND 4.51045f $ **FLOATING
C7392 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND 1.56057f $ **FLOATING
C7393 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7394 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7395 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND 1.58431f $ **FLOATING
C7396 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND 30.3253f $ **FLOATING
C7397 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND 3.16311f $ **FLOATING
C7398 a_48343_26999# VGND 0.16243f $ **FLOATING
C7399 a_44418_26990# VGND 0.89497f $ **FLOATING
C7400 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND 2.665f $ **FLOATING
C7401 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND 6.34862f $ **FLOATING
C7402 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37348f $ **FLOATING
C7403 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7404 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44912f $ **FLOATING
C7405 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7406 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND 4.51335f $ **FLOATING
C7407 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND 1.56099f $ **FLOATING
C7408 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.405f $ **FLOATING
C7410 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND 1.58193f $ **FLOATING
C7411 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND 21.4947f $ **FLOATING
C7412 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND 3.16279f $ **FLOATING
C7413 a_43540_26999# VGND 0.16243f $ **FLOATING
C7414 a_39616_26990# VGND 0.89497f $ **FLOATING
C7415 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND 2.66616f $ **FLOATING
C7416 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND 6.34842f $ **FLOATING
C7417 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37296f $ **FLOATING
C7418 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7419 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44899f $ **FLOATING
C7420 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7421 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND 4.51193f $ **FLOATING
C7422 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND 1.56081f $ **FLOATING
C7423 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7424 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40542f $ **FLOATING
C7425 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND 1.58513f $ **FLOATING
C7426 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND 20.61f $ **FLOATING
C7427 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7428 a_38738_26999# VGND 0.16243f $ **FLOATING
C7429 a_34814_26990# VGND 0.89548f $ **FLOATING
C7430 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND 2.66683f $ **FLOATING
C7431 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND 6.34843f $ **FLOATING
C7432 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7433 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7434 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7435 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7436 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND 4.51156f $ **FLOATING
C7437 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7438 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7439 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40525f $ **FLOATING
C7440 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7441 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND 16.1449f $ **FLOATING
C7442 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7443 a_33936_26999# VGND 0.16243f $ **FLOATING
C7444 a_30012_26990# VGND 0.89497f $ **FLOATING
C7445 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND 2.66498f $ **FLOATING
C7446 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND 6.34843f $ **FLOATING
C7447 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7448 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7449 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7450 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND 4.51162f $ **FLOATING
C7452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7453 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7454 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7455 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7456 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND 15.6371f $ **FLOATING
C7457 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7458 a_29134_26999# VGND 0.16243f $ **FLOATING
C7459 single_9b_cdac_0.SW[7] VGND 7.22415f $ **FLOATING
C7460 a_25210_26990# VGND 0.89548f $ **FLOATING
C7461 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND 2.68106f $ **FLOATING
C7462 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND 6.3484f $ **FLOATING
C7463 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7464 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7465 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7467 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND 4.51212f $ **FLOATING
C7468 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7469 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7470 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7471 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7472 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND 14.5496f $ **FLOATING
C7473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND 3.17698f $ **FLOATING
C7474 a_24332_26999# VGND 0.16243f $ **FLOATING
C7475 single_9b_cdac_0.SW[1] VGND 7.88723f $ **FLOATING
C7476 a_12647_27128# VGND 0.01049f $ **FLOATING
C7477 a_12560_27128# VGND 0.18115f $ **FLOATING
C7478 a_13011_27234# VGND 0.59986f $ **FLOATING
C7479 sar9b_0.net27 VGND 1.75655f $ **FLOATING
C7480 single_9b_cdac_0.SW[4] VGND 7.53235f $ **FLOATING
C7481 single_9b_cdac_0.SW[5] VGND 7.99262f $ **FLOATING
C7482 sar9b_0.net52 VGND 3.396f $ **FLOATING
C7483 sar9b_0.net30 VGND 0.98276f $ **FLOATING
C7484 a_11915_27039# VGND 0.68615f $ **FLOATING
C7485 sar9b_0.net31 VGND 0.75736f $ **FLOATING
C7486 a_11339_27039# VGND 0.62214f $ **FLOATING
C7487 sar9b_0.net42 VGND 1.35212f $ **FLOATING
C7488 a_10378_27170# VGND 0.13252f $ **FLOATING
C7489 a_9802_26815# VGND 0.11561f $ **FLOATING
C7490 a_9870_27060# VGND 0.16016f $ **FLOATING
C7491 a_9593_26914# VGND 0.89305f $ **FLOATING
C7492 a_9588_27045# VGND 0.60592f $ **FLOATING
C7493 a_9279_27227# VGND 0.28615f $ **FLOATING
C7494 a_9138_27163# VGND 0.33078f $ **FLOATING
C7495 a_8940_27039# VGND 0.28409f $ **FLOATING
C7496 a_6880_26815# VGND 0.30246f $ **FLOATING
C7497 a_6534_27123# VGND 0.29776f $ **FLOATING
C7498 a_6282_27170# VGND 0.35829f $ **FLOATING
C7499 a_5846_26950# VGND 0.15475f $ **FLOATING
C7500 a_5711_26851# VGND 0.20102f $ **FLOATING
C7501 a_5506_26802# VGND 0.94424f $ **FLOATING
C7502 a_5046_27230# VGND 0.11169f $ **FLOATING
C7503 a_5322_27170# VGND 0.61739f $ **FLOATING
C7504 sar9b_0.net39 VGND 5.04702f $ **FLOATING
C7505 sar9b_0.net37 VGND 3.30771f $ **FLOATING
C7506 a_4330_27170# VGND 0.1075f $ **FLOATING
C7507 a_3754_26815# VGND 0.11452f $ **FLOATING
C7508 a_3822_27060# VGND 0.15534f $ **FLOATING
C7509 a_3545_26914# VGND 0.88258f $ **FLOATING
C7510 a_3540_27045# VGND 0.57229f $ **FLOATING
C7511 a_3231_27227# VGND 0.28633f $ **FLOATING
C7512 a_3090_27163# VGND 0.3281f $ **FLOATING
C7513 a_2892_27039# VGND 0.27715f $ **FLOATING
C7514 a_2451_27234# VGND 0.36326f $ **FLOATING
C7515 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND 6.37207f $ **FLOATING
C7516 single_9b_cdac_0.SW[2] VGND 7.79108f $ **FLOATING
C7517 single_9b_cdac_0.SW[3] VGND 7.69147f $ **FLOATING
C7518 a_10607_27849# VGND 0.17037f $ **FLOATING
C7519 sar9b_0.net28 VGND 2.13028f $ **FLOATING
C7520 a_13067_27662# VGND 0.62659f $ **FLOATING
C7521 sar9b_0.net29 VGND 1.17448f $ **FLOATING
C7522 a_12491_27662# VGND 0.63745f $ **FLOATING
C7523 a_11776_27801# VGND 0.33209f $ **FLOATING
C7524 a_11178_27466# VGND 0.37061f $ **FLOATING
C7525 a_11430_27595# VGND 0.30882f $ **FLOATING
C7526 a_10742_27751# VGND 0.13782f $ **FLOATING
C7527 a_10402_27758# VGND 0.92755f $ **FLOATING
C7528 a_10218_27466# VGND 0.65521f $ **FLOATING
C7529 a_9942_27470# VGND 0.15547f $ **FLOATING
C7530 sar9b_0.net43 VGND 2.18762f $ **FLOATING
C7531 single_9b_cdac_0.SW[8] VGND 9.42114f $ **FLOATING
C7532 a_7343_27849# VGND 0.16308f $ **FLOATING
C7533 sar9b_0.net34 VGND 0.84365f $ **FLOATING
C7534 a_9323_27662# VGND 0.63074f $ **FLOATING
C7535 a_8883_27466# VGND 0.45025f $ **FLOATING
C7536 sar9b_0.cyclic_flag_0.FINAL VGND 1.13968f $ **FLOATING
C7537 a_8512_27801# VGND 0.28448f $ **FLOATING
C7538 a_7914_27466# VGND 0.34106f $ **FLOATING
C7539 a_8166_27595# VGND 0.29361f $ **FLOATING
C7540 a_7478_27751# VGND 0.12296f $ **FLOATING
C7541 a_7138_27758# VGND 0.91809f $ **FLOATING
C7542 a_6954_27466# VGND 0.61234f $ **FLOATING
C7543 a_6678_27470# VGND 0.11676f $ **FLOATING
C7544 sar9b_0.net40 VGND 4.42282f $ **FLOATING
C7545 a_6307_27584# VGND 0.41924f $ **FLOATING
C7546 a_5235_27466# VGND 0.61697f $ **FLOATING
C7547 sar9b_0.net19 VGND 1.72645f $ **FLOATING
C7548 a_4749_27652# VGND 0.44592f $ **FLOATING
C7549 sar9b_0.net36 VGND 3.44267f $ **FLOATING
C7550 sar9b_0.net44 VGND 1.32306f $ **FLOATING
C7551 a_3946_27530# VGND 0.1577f $ **FLOATING
C7552 a_3438_27677# VGND 0.1683f $ **FLOATING
C7553 a_3370_27769# VGND 0.13183f $ **FLOATING
C7554 a_3161_27787# VGND 0.91973f $ **FLOATING
C7555 a_2847_27473# VGND 0.30295f $ **FLOATING
C7556 a_2706_27440# VGND 0.35511f $ **FLOATING
C7557 a_3156_27447# VGND 0.60874f $ **FLOATING
C7558 a_2508_27440# VGND 0.29951f $ **FLOATING
C7559 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7560 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7561 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7562 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7563 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND 4.51154f $ **FLOATING
C7564 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7565 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7567 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7568 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND 13.6188f $ **FLOATING
C7569 sar9b_0._06_ VGND 0.51759f $ **FLOATING
C7570 a_13164_28398# VGND 0.35538f $ **FLOATING
C7571 a_12531_28566# VGND 0.66182f $ **FLOATING
C7572 sar9b_0.net25 VGND 0.48263f $ **FLOATING
C7573 sar9b_0.net14 VGND 0.57635f $ **FLOATING
C7574 a_11915_28371# VGND 0.69798f $ **FLOATING
C7575 a_10995_28566# VGND 0.63419f $ **FLOATING
C7576 sar9b_0.net24 VGND 1.19162f $ **FLOATING
C7577 a_9939_28566# VGND 0.66415f $ **FLOATING
C7578 sar9b_0.net23 VGND 0.45975f $ **FLOATING
C7579 single_9b_cdac_0.SW[6] VGND 7.61708f $ **FLOATING
C7580 sar9b_0.net32 VGND 2.57466f $ **FLOATING
C7581 a_9323_28371# VGND 0.65565f $ **FLOATING
C7582 a_8691_28566# VGND 0.6426f $ **FLOATING
C7583 sar9b_0.net22 VGND 0.37611f $ **FLOATING
C7584 a_8115_28566# VGND 0.63526f $ **FLOATING
C7585 a_7539_28566# VGND 0.63297f $ **FLOATING
C7586 sar9b_0.net21 VGND 0.59997f $ **FLOATING
C7587 sar9b_0.net38 VGND 1.58614f $ **FLOATING
C7588 a_6250_28502# VGND 0.14552f $ **FLOATING
C7589 sar9b_0.net45 VGND 1.28036f $ **FLOATING
C7590 a_5674_28147# VGND 0.15778f $ **FLOATING
C7591 a_5742_28392# VGND 0.21088f $ **FLOATING
C7592 a_5465_28246# VGND 0.95941f $ **FLOATING
C7593 a_5460_28377# VGND 0.66988f $ **FLOATING
C7594 a_5151_28559# VGND 0.30729f $ **FLOATING
C7595 sar9b_0.net58 VGND 3.01825f $ **FLOATING
C7596 sar9b_0.net20 VGND 1.32881f $ **FLOATING
C7597 a_5010_28495# VGND 0.36594f $ **FLOATING
C7598 a_4812_28371# VGND 0.29879f $ **FLOATING
C7599 sar9b_0.net59 VGND 2.86651f $ **FLOATING
C7600 a_4083_28566# VGND 0.64865f $ **FLOATING
C7601 sar9b_0.net18 VGND 0.41648f $ **FLOATING
C7602 a_3603_28156# VGND 0.47335f $ **FLOATING
C7603 sar9b_0.net60 VGND 3.34485f $ **FLOATING
C7604 a_2931_28566# VGND 0.64119f $ **FLOATING
C7605 sar9b_0.net17 VGND 0.6804f $ **FLOATING
C7606 a_2547_28132# VGND 0.43769f $ **FLOATING
C7607 sar9b_0.net3 VGND 0.60828f $ **FLOATING
C7608 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND 4.71478f $ **FLOATING
C7609 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7611 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7612 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7613 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7614 single_9b_cdac_1.CF[0] VGND 15.8339f $ **FLOATING
C7615 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7616 single_9b_cdac_1.CF[1] VGND 11.5306f $ **FLOATING
C7617 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7618 single_9b_cdac_1.CF[2] VGND 11.2901f $ **FLOATING
C7619 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7620 single_9b_cdac_1.CF[3] VGND 10.9802f $ **FLOATING
C7621 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7622 single_9b_cdac_1.CF[4] VGND 10.9973f $ **FLOATING
C7623 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7624 single_9b_cdac_1.CF[5] VGND 10.4191f $ **FLOATING
C7625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7626 single_9b_cdac_1.CF[6] VGND 10.1217f $ **FLOATING
C7627 single_9b_cdac_1.CF[7] VGND 10.1149f $ **FLOATING
C7628 single_9b_cdac_1.CF[8] VGND 8.83586f $ **FLOATING
C7629 dw_17224_1400# VGND 27.9938f $ **FLOATING
C7630 dw_12589_1395# VGND 28.2006f $ **FLOATING
.ends
