magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< nwell >>
rect -211 -348 211 348
<< pmos >>
rect -15 -200 15 200
<< pdiff >>
rect -73 188 -15 200
rect -73 -188 -61 188
rect -27 -188 -15 188
rect -73 -200 -15 -188
rect 15 188 73 200
rect 15 -188 27 188
rect 61 -188 73 188
rect 15 -200 73 -188
<< pdiffc >>
rect -61 -188 -27 188
rect 27 -188 61 188
<< nsubdiff >>
rect -175 278 -79 312
rect 79 278 175 312
rect -175 216 -141 278
rect 141 216 175 278
rect -175 -278 -141 -216
rect 141 -278 175 -216
rect -175 -312 -79 -278
rect 79 -312 175 -278
<< nsubdiffcont >>
rect -79 278 79 312
rect -175 -216 -141 216
rect 141 -216 175 216
rect -79 -312 79 -278
<< poly >>
rect -15 200 15 226
rect -15 -226 15 -200
<< locali >>
rect -175 278 -79 312
rect 79 278 175 312
rect -175 216 -141 278
rect 141 216 175 278
rect -61 188 -27 204
rect -61 -204 -27 -188
rect 27 188 61 204
rect 27 -204 61 -188
rect -175 -278 -141 -216
rect 141 -278 175 -216
rect -175 -312 -79 -278
rect 79 -312 175 -278
<< viali >>
rect -61 -188 -27 188
rect 27 -188 61 188
<< metal1 >>
rect -67 188 -21 200
rect -67 -188 -61 188
rect -27 -188 -21 188
rect -67 -200 -21 -188
rect 21 188 67 200
rect 21 -188 27 188
rect 61 -188 67 188
rect 21 -200 67 -188
<< properties >>
string FIXED_BBOX -158 -295 158 295
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
