magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< nwell >>
rect -211 -223 211 223
<< pmos >>
rect -15 -75 15 75
<< pdiff >>
rect -73 63 -15 75
rect -73 -63 -61 63
rect -27 -63 -15 63
rect -73 -75 -15 -63
rect 15 63 73 75
rect 15 -63 27 63
rect 61 -63 73 63
rect 15 -75 73 -63
<< pdiffc >>
rect -61 -63 -27 63
rect 27 -63 61 63
<< nsubdiff >>
rect -175 153 -79 187
rect 79 153 175 187
rect -175 91 -141 153
rect 141 91 175 153
rect -175 -153 -141 -91
rect 141 -153 175 -91
rect -175 -187 -79 -153
rect 79 -187 175 -153
<< nsubdiffcont >>
rect -79 153 79 187
rect -175 -91 -141 91
rect 141 -91 175 91
rect -79 -187 79 -153
<< poly >>
rect -15 75 15 101
rect -15 -101 15 -75
<< locali >>
rect -175 153 -79 187
rect 79 153 175 187
rect -175 91 -141 153
rect 141 91 175 153
rect -61 63 -27 79
rect -61 -79 -27 -63
rect 27 63 61 79
rect 27 -79 61 -63
rect -175 -153 -141 -91
rect 141 -153 175 -91
rect -175 -187 -79 -153
rect 79 -187 175 -153
<< viali >>
rect -61 -63 -27 63
rect 27 -63 61 63
<< metal1 >>
rect -67 63 -21 75
rect -67 -63 -61 63
rect -27 -63 -21 63
rect -67 -75 -21 -63
rect 21 63 67 75
rect 21 -63 27 63
rect 61 -63 67 63
rect 21 -75 67 -63
<< properties >>
string FIXED_BBOX -158 -170 158 170
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.75 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
