magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< error_p >>
rect -29 -407 29 -401
rect -29 -441 -17 -407
rect -29 -447 29 -441
<< pwell >>
rect -201 -569 201 569
<< nmos >>
rect -15 -369 15 431
<< ndiff >>
rect -73 388 -15 431
rect -73 354 -61 388
rect -27 354 -15 388
rect -73 320 -15 354
rect -73 286 -61 320
rect -27 286 -15 320
rect -73 252 -15 286
rect -73 218 -61 252
rect -27 218 -15 252
rect -73 184 -15 218
rect -73 150 -61 184
rect -27 150 -15 184
rect -73 116 -15 150
rect -73 82 -61 116
rect -27 82 -15 116
rect -73 48 -15 82
rect -73 14 -61 48
rect -27 14 -15 48
rect -73 -20 -15 14
rect -73 -54 -61 -20
rect -27 -54 -15 -20
rect -73 -88 -15 -54
rect -73 -122 -61 -88
rect -27 -122 -15 -88
rect -73 -156 -15 -122
rect -73 -190 -61 -156
rect -27 -190 -15 -156
rect -73 -224 -15 -190
rect -73 -258 -61 -224
rect -27 -258 -15 -224
rect -73 -292 -15 -258
rect -73 -326 -61 -292
rect -27 -326 -15 -292
rect -73 -369 -15 -326
rect 15 388 73 431
rect 15 354 27 388
rect 61 354 73 388
rect 15 320 73 354
rect 15 286 27 320
rect 61 286 73 320
rect 15 252 73 286
rect 15 218 27 252
rect 61 218 73 252
rect 15 184 73 218
rect 15 150 27 184
rect 61 150 73 184
rect 15 116 73 150
rect 15 82 27 116
rect 61 82 73 116
rect 15 48 73 82
rect 15 14 27 48
rect 61 14 73 48
rect 15 -20 73 14
rect 15 -54 27 -20
rect 61 -54 73 -20
rect 15 -88 73 -54
rect 15 -122 27 -88
rect 61 -122 73 -88
rect 15 -156 73 -122
rect 15 -190 27 -156
rect 61 -190 73 -156
rect 15 -224 73 -190
rect 15 -258 27 -224
rect 61 -258 73 -224
rect 15 -292 73 -258
rect 15 -326 27 -292
rect 61 -326 73 -292
rect 15 -369 73 -326
<< ndiffc >>
rect -61 354 -27 388
rect -61 286 -27 320
rect -61 218 -27 252
rect -61 150 -27 184
rect -61 82 -27 116
rect -61 14 -27 48
rect -61 -54 -27 -20
rect -61 -122 -27 -88
rect -61 -190 -27 -156
rect -61 -258 -27 -224
rect -61 -326 -27 -292
rect 27 354 61 388
rect 27 286 61 320
rect 27 218 61 252
rect 27 150 61 184
rect 27 82 61 116
rect 27 14 61 48
rect 27 -54 61 -20
rect 27 -122 61 -88
rect 27 -190 61 -156
rect 27 -258 61 -224
rect 27 -326 61 -292
<< psubdiff >>
rect -175 509 -51 543
rect -17 509 17 543
rect 51 509 175 543
rect -175 -509 -141 509
rect 141 425 175 509
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -509 175 -425
rect -175 -543 -51 -509
rect -17 -543 17 -509
rect 51 -543 175 -509
<< psubdiffcont >>
rect -51 509 -17 543
rect 17 509 51 543
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect -51 -543 -17 -509
rect 17 -543 51 -509
<< poly >>
rect -15 431 15 457
rect -15 -391 15 -369
rect -33 -407 33 -391
rect -33 -441 -17 -407
rect 17 -441 33 -407
rect -33 -457 33 -441
<< polycont >>
rect -17 -441 17 -407
<< locali >>
rect -175 509 -51 543
rect -17 509 17 543
rect 51 509 175 543
rect -175 -509 -141 509
rect -61 408 -27 435
rect -61 336 -27 354
rect -61 264 -27 286
rect -61 192 -27 218
rect -61 120 -27 150
rect -61 48 -27 82
rect -61 -20 -27 14
rect -61 -88 -27 -58
rect -61 -156 -27 -130
rect -61 -224 -27 -202
rect -61 -292 -27 -274
rect -61 -373 -27 -346
rect 27 408 61 435
rect 27 336 61 354
rect 27 264 61 286
rect 27 192 61 218
rect 27 120 61 150
rect 27 48 61 82
rect 27 -20 61 14
rect 27 -88 61 -58
rect 27 -156 61 -130
rect 27 -224 61 -202
rect 27 -292 61 -274
rect 27 -373 61 -346
rect 141 425 175 509
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect -33 -441 -17 -407
rect 17 -441 33 -407
rect 141 -509 175 -425
rect -175 -543 -51 -509
rect -17 -543 17 -509
rect 51 -543 175 -509
<< viali >>
rect -61 388 -27 408
rect -61 374 -27 388
rect -61 320 -27 336
rect -61 302 -27 320
rect -61 252 -27 264
rect -61 230 -27 252
rect -61 184 -27 192
rect -61 158 -27 184
rect -61 116 -27 120
rect -61 86 -27 116
rect -61 14 -27 48
rect -61 -54 -27 -24
rect -61 -58 -27 -54
rect -61 -122 -27 -96
rect -61 -130 -27 -122
rect -61 -190 -27 -168
rect -61 -202 -27 -190
rect -61 -258 -27 -240
rect -61 -274 -27 -258
rect -61 -326 -27 -312
rect -61 -346 -27 -326
rect 27 388 61 408
rect 27 374 61 388
rect 27 320 61 336
rect 27 302 61 320
rect 27 252 61 264
rect 27 230 61 252
rect 27 184 61 192
rect 27 158 61 184
rect 27 116 61 120
rect 27 86 61 116
rect 27 14 61 48
rect 27 -54 61 -24
rect 27 -58 61 -54
rect 27 -122 61 -96
rect 27 -130 61 -122
rect 27 -190 61 -168
rect 27 -202 61 -190
rect 27 -258 61 -240
rect 27 -274 61 -258
rect 27 -326 61 -312
rect 27 -346 61 -326
rect -17 -441 17 -407
<< metal1 >>
rect -67 408 -21 431
rect -67 374 -61 408
rect -27 374 -21 408
rect -67 336 -21 374
rect -67 302 -61 336
rect -27 302 -21 336
rect -67 264 -21 302
rect -67 230 -61 264
rect -27 230 -21 264
rect -67 192 -21 230
rect -67 158 -61 192
rect -27 158 -21 192
rect -67 120 -21 158
rect -67 86 -61 120
rect -27 86 -21 120
rect -67 48 -21 86
rect -67 14 -61 48
rect -27 14 -21 48
rect -67 -24 -21 14
rect -67 -58 -61 -24
rect -27 -58 -21 -24
rect -67 -96 -21 -58
rect -67 -130 -61 -96
rect -27 -130 -21 -96
rect -67 -168 -21 -130
rect -67 -202 -61 -168
rect -27 -202 -21 -168
rect -67 -240 -21 -202
rect -67 -274 -61 -240
rect -27 -274 -21 -240
rect -67 -312 -21 -274
rect -67 -346 -61 -312
rect -27 -346 -21 -312
rect -67 -369 -21 -346
rect 21 408 67 431
rect 21 374 27 408
rect 61 374 67 408
rect 21 336 67 374
rect 21 302 27 336
rect 61 302 67 336
rect 21 264 67 302
rect 21 230 27 264
rect 61 230 67 264
rect 21 192 67 230
rect 21 158 27 192
rect 61 158 67 192
rect 21 120 67 158
rect 21 86 27 120
rect 61 86 67 120
rect 21 48 67 86
rect 21 14 27 48
rect 61 14 67 48
rect 21 -24 67 14
rect 21 -58 27 -24
rect 61 -58 67 -24
rect 21 -96 67 -58
rect 21 -130 27 -96
rect 61 -130 67 -96
rect 21 -168 67 -130
rect 21 -202 27 -168
rect 61 -202 67 -168
rect 21 -240 67 -202
rect 21 -274 27 -240
rect 61 -274 67 -240
rect 21 -312 67 -274
rect 21 -346 27 -312
rect 61 -346 67 -312
rect 21 -369 67 -346
rect -29 -407 29 -401
rect -29 -441 -17 -407
rect 17 -441 29 -407
rect -29 -447 29 -441
<< properties >>
string FIXED_BBOX -158 -526 158 526
<< end >>
