magic
tech sky130A
magscale 1 2
timestamp 1749307785
<< error_p >>
rect -29 156 29 162
rect -29 122 -17 156
rect -29 116 29 122
rect -29 -122 29 -116
rect -29 -156 -17 -122
rect -29 -162 29 -156
<< nwell >>
rect -211 -294 211 294
<< pmos >>
rect -15 -75 15 75
<< pdiff >>
rect -73 63 -15 75
rect -73 -63 -61 63
rect -27 -63 -15 63
rect -73 -75 -15 -63
rect 15 63 73 75
rect 15 -63 27 63
rect 61 -63 73 63
rect 15 -75 73 -63
<< pdiffc >>
rect -61 -63 -27 63
rect 27 -63 61 63
<< nsubdiff >>
rect -175 224 -79 258
rect 79 224 175 258
rect -175 162 -141 224
rect 141 162 175 224
rect -175 -224 -141 -162
rect 141 -224 175 -162
rect -175 -258 -79 -224
rect 79 -258 175 -224
<< nsubdiffcont >>
rect -79 224 79 258
rect -175 -162 -141 162
rect 141 -162 175 162
rect -79 -258 79 -224
<< poly >>
rect -33 156 33 172
rect -33 122 -17 156
rect 17 122 33 156
rect -33 106 33 122
rect -15 75 15 106
rect -15 -106 15 -75
rect -33 -122 33 -106
rect -33 -156 -17 -122
rect 17 -156 33 -122
rect -33 -172 33 -156
<< polycont >>
rect -17 122 17 156
rect -17 -156 17 -122
<< locali >>
rect -175 224 -79 258
rect 79 224 175 258
rect -175 162 -141 224
rect 141 162 175 224
rect -33 122 -17 156
rect 17 122 33 156
rect -61 63 -27 79
rect -61 -79 -27 -63
rect 27 63 61 79
rect 27 -79 61 -63
rect -33 -156 -17 -122
rect 17 -156 33 -122
rect -175 -224 -141 -162
rect 141 -224 175 -162
rect -175 -258 -79 -224
rect 79 -258 175 -224
<< viali >>
rect -17 122 17 156
rect -61 -63 -27 63
rect 27 -63 61 63
rect -17 -156 17 -122
<< metal1 >>
rect -29 156 29 162
rect -29 122 -17 156
rect 17 122 29 156
rect -29 116 29 122
rect -67 63 -21 75
rect -67 -63 -61 63
rect -27 -63 -21 63
rect -67 -75 -21 -63
rect 21 63 67 75
rect 21 -63 27 63
rect 61 -63 67 63
rect 21 -75 67 -63
rect -29 -122 29 -116
rect -29 -156 -17 -122
rect 17 -156 29 -122
rect -29 -162 29 -156
<< properties >>
string FIXED_BBOX -158 -241 158 241
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.75 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
