magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal3 >>
rect -2704 4312 -1532 4360
rect -2704 4248 -1616 4312
rect -1552 4248 -1532 4312
rect -2704 4232 -1532 4248
rect -2704 4168 -1616 4232
rect -1552 4168 -1532 4232
rect -2704 4152 -1532 4168
rect -2704 4088 -1616 4152
rect -1552 4088 -1532 4152
rect -2704 4072 -1532 4088
rect -2704 4008 -1616 4072
rect -1552 4008 -1532 4072
rect -2704 3992 -1532 4008
rect -2704 3928 -1616 3992
rect -1552 3928 -1532 3992
rect -2704 3912 -1532 3928
rect -2704 3848 -1616 3912
rect -1552 3848 -1532 3912
rect -2704 3832 -1532 3848
rect -2704 3768 -1616 3832
rect -1552 3768 -1532 3832
rect -2704 3752 -1532 3768
rect -2704 3688 -1616 3752
rect -1552 3688 -1532 3752
rect -2704 3672 -1532 3688
rect -2704 3608 -1616 3672
rect -1552 3608 -1532 3672
rect -2704 3592 -1532 3608
rect -2704 3528 -1616 3592
rect -1552 3528 -1532 3592
rect -2704 3480 -1532 3528
rect -1292 4312 -120 4360
rect -1292 4248 -204 4312
rect -140 4248 -120 4312
rect -1292 4232 -120 4248
rect -1292 4168 -204 4232
rect -140 4168 -120 4232
rect -1292 4152 -120 4168
rect -1292 4088 -204 4152
rect -140 4088 -120 4152
rect -1292 4072 -120 4088
rect -1292 4008 -204 4072
rect -140 4008 -120 4072
rect -1292 3992 -120 4008
rect -1292 3928 -204 3992
rect -140 3928 -120 3992
rect -1292 3912 -120 3928
rect -1292 3848 -204 3912
rect -140 3848 -120 3912
rect -1292 3832 -120 3848
rect -1292 3768 -204 3832
rect -140 3768 -120 3832
rect -1292 3752 -120 3768
rect -1292 3688 -204 3752
rect -140 3688 -120 3752
rect -1292 3672 -120 3688
rect -1292 3608 -204 3672
rect -140 3608 -120 3672
rect -1292 3592 -120 3608
rect -1292 3528 -204 3592
rect -140 3528 -120 3592
rect -1292 3480 -120 3528
rect 120 4312 1292 4360
rect 120 4248 1208 4312
rect 1272 4248 1292 4312
rect 120 4232 1292 4248
rect 120 4168 1208 4232
rect 1272 4168 1292 4232
rect 120 4152 1292 4168
rect 120 4088 1208 4152
rect 1272 4088 1292 4152
rect 120 4072 1292 4088
rect 120 4008 1208 4072
rect 1272 4008 1292 4072
rect 120 3992 1292 4008
rect 120 3928 1208 3992
rect 1272 3928 1292 3992
rect 120 3912 1292 3928
rect 120 3848 1208 3912
rect 1272 3848 1292 3912
rect 120 3832 1292 3848
rect 120 3768 1208 3832
rect 1272 3768 1292 3832
rect 120 3752 1292 3768
rect 120 3688 1208 3752
rect 1272 3688 1292 3752
rect 120 3672 1292 3688
rect 120 3608 1208 3672
rect 1272 3608 1292 3672
rect 120 3592 1292 3608
rect 120 3528 1208 3592
rect 1272 3528 1292 3592
rect 120 3480 1292 3528
rect 1532 4312 2704 4360
rect 1532 4248 2620 4312
rect 2684 4248 2704 4312
rect 1532 4232 2704 4248
rect 1532 4168 2620 4232
rect 2684 4168 2704 4232
rect 1532 4152 2704 4168
rect 1532 4088 2620 4152
rect 2684 4088 2704 4152
rect 1532 4072 2704 4088
rect 1532 4008 2620 4072
rect 2684 4008 2704 4072
rect 1532 3992 2704 4008
rect 1532 3928 2620 3992
rect 2684 3928 2704 3992
rect 1532 3912 2704 3928
rect 1532 3848 2620 3912
rect 2684 3848 2704 3912
rect 1532 3832 2704 3848
rect 1532 3768 2620 3832
rect 2684 3768 2704 3832
rect 1532 3752 2704 3768
rect 1532 3688 2620 3752
rect 2684 3688 2704 3752
rect 1532 3672 2704 3688
rect 1532 3608 2620 3672
rect 2684 3608 2704 3672
rect 1532 3592 2704 3608
rect 1532 3528 2620 3592
rect 2684 3528 2704 3592
rect 1532 3480 2704 3528
rect -2704 3192 -1532 3240
rect -2704 3128 -1616 3192
rect -1552 3128 -1532 3192
rect -2704 3112 -1532 3128
rect -2704 3048 -1616 3112
rect -1552 3048 -1532 3112
rect -2704 3032 -1532 3048
rect -2704 2968 -1616 3032
rect -1552 2968 -1532 3032
rect -2704 2952 -1532 2968
rect -2704 2888 -1616 2952
rect -1552 2888 -1532 2952
rect -2704 2872 -1532 2888
rect -2704 2808 -1616 2872
rect -1552 2808 -1532 2872
rect -2704 2792 -1532 2808
rect -2704 2728 -1616 2792
rect -1552 2728 -1532 2792
rect -2704 2712 -1532 2728
rect -2704 2648 -1616 2712
rect -1552 2648 -1532 2712
rect -2704 2632 -1532 2648
rect -2704 2568 -1616 2632
rect -1552 2568 -1532 2632
rect -2704 2552 -1532 2568
rect -2704 2488 -1616 2552
rect -1552 2488 -1532 2552
rect -2704 2472 -1532 2488
rect -2704 2408 -1616 2472
rect -1552 2408 -1532 2472
rect -2704 2360 -1532 2408
rect -1292 3192 -120 3240
rect -1292 3128 -204 3192
rect -140 3128 -120 3192
rect -1292 3112 -120 3128
rect -1292 3048 -204 3112
rect -140 3048 -120 3112
rect -1292 3032 -120 3048
rect -1292 2968 -204 3032
rect -140 2968 -120 3032
rect -1292 2952 -120 2968
rect -1292 2888 -204 2952
rect -140 2888 -120 2952
rect -1292 2872 -120 2888
rect -1292 2808 -204 2872
rect -140 2808 -120 2872
rect -1292 2792 -120 2808
rect -1292 2728 -204 2792
rect -140 2728 -120 2792
rect -1292 2712 -120 2728
rect -1292 2648 -204 2712
rect -140 2648 -120 2712
rect -1292 2632 -120 2648
rect -1292 2568 -204 2632
rect -140 2568 -120 2632
rect -1292 2552 -120 2568
rect -1292 2488 -204 2552
rect -140 2488 -120 2552
rect -1292 2472 -120 2488
rect -1292 2408 -204 2472
rect -140 2408 -120 2472
rect -1292 2360 -120 2408
rect 120 3192 1292 3240
rect 120 3128 1208 3192
rect 1272 3128 1292 3192
rect 120 3112 1292 3128
rect 120 3048 1208 3112
rect 1272 3048 1292 3112
rect 120 3032 1292 3048
rect 120 2968 1208 3032
rect 1272 2968 1292 3032
rect 120 2952 1292 2968
rect 120 2888 1208 2952
rect 1272 2888 1292 2952
rect 120 2872 1292 2888
rect 120 2808 1208 2872
rect 1272 2808 1292 2872
rect 120 2792 1292 2808
rect 120 2728 1208 2792
rect 1272 2728 1292 2792
rect 120 2712 1292 2728
rect 120 2648 1208 2712
rect 1272 2648 1292 2712
rect 120 2632 1292 2648
rect 120 2568 1208 2632
rect 1272 2568 1292 2632
rect 120 2552 1292 2568
rect 120 2488 1208 2552
rect 1272 2488 1292 2552
rect 120 2472 1292 2488
rect 120 2408 1208 2472
rect 1272 2408 1292 2472
rect 120 2360 1292 2408
rect 1532 3192 2704 3240
rect 1532 3128 2620 3192
rect 2684 3128 2704 3192
rect 1532 3112 2704 3128
rect 1532 3048 2620 3112
rect 2684 3048 2704 3112
rect 1532 3032 2704 3048
rect 1532 2968 2620 3032
rect 2684 2968 2704 3032
rect 1532 2952 2704 2968
rect 1532 2888 2620 2952
rect 2684 2888 2704 2952
rect 1532 2872 2704 2888
rect 1532 2808 2620 2872
rect 2684 2808 2704 2872
rect 1532 2792 2704 2808
rect 1532 2728 2620 2792
rect 2684 2728 2704 2792
rect 1532 2712 2704 2728
rect 1532 2648 2620 2712
rect 2684 2648 2704 2712
rect 1532 2632 2704 2648
rect 1532 2568 2620 2632
rect 2684 2568 2704 2632
rect 1532 2552 2704 2568
rect 1532 2488 2620 2552
rect 2684 2488 2704 2552
rect 1532 2472 2704 2488
rect 1532 2408 2620 2472
rect 2684 2408 2704 2472
rect 1532 2360 2704 2408
rect -2704 2072 -1532 2120
rect -2704 2008 -1616 2072
rect -1552 2008 -1532 2072
rect -2704 1992 -1532 2008
rect -2704 1928 -1616 1992
rect -1552 1928 -1532 1992
rect -2704 1912 -1532 1928
rect -2704 1848 -1616 1912
rect -1552 1848 -1532 1912
rect -2704 1832 -1532 1848
rect -2704 1768 -1616 1832
rect -1552 1768 -1532 1832
rect -2704 1752 -1532 1768
rect -2704 1688 -1616 1752
rect -1552 1688 -1532 1752
rect -2704 1672 -1532 1688
rect -2704 1608 -1616 1672
rect -1552 1608 -1532 1672
rect -2704 1592 -1532 1608
rect -2704 1528 -1616 1592
rect -1552 1528 -1532 1592
rect -2704 1512 -1532 1528
rect -2704 1448 -1616 1512
rect -1552 1448 -1532 1512
rect -2704 1432 -1532 1448
rect -2704 1368 -1616 1432
rect -1552 1368 -1532 1432
rect -2704 1352 -1532 1368
rect -2704 1288 -1616 1352
rect -1552 1288 -1532 1352
rect -2704 1240 -1532 1288
rect -1292 2072 -120 2120
rect -1292 2008 -204 2072
rect -140 2008 -120 2072
rect -1292 1992 -120 2008
rect -1292 1928 -204 1992
rect -140 1928 -120 1992
rect -1292 1912 -120 1928
rect -1292 1848 -204 1912
rect -140 1848 -120 1912
rect -1292 1832 -120 1848
rect -1292 1768 -204 1832
rect -140 1768 -120 1832
rect -1292 1752 -120 1768
rect -1292 1688 -204 1752
rect -140 1688 -120 1752
rect -1292 1672 -120 1688
rect -1292 1608 -204 1672
rect -140 1608 -120 1672
rect -1292 1592 -120 1608
rect -1292 1528 -204 1592
rect -140 1528 -120 1592
rect -1292 1512 -120 1528
rect -1292 1448 -204 1512
rect -140 1448 -120 1512
rect -1292 1432 -120 1448
rect -1292 1368 -204 1432
rect -140 1368 -120 1432
rect -1292 1352 -120 1368
rect -1292 1288 -204 1352
rect -140 1288 -120 1352
rect -1292 1240 -120 1288
rect 120 2072 1292 2120
rect 120 2008 1208 2072
rect 1272 2008 1292 2072
rect 120 1992 1292 2008
rect 120 1928 1208 1992
rect 1272 1928 1292 1992
rect 120 1912 1292 1928
rect 120 1848 1208 1912
rect 1272 1848 1292 1912
rect 120 1832 1292 1848
rect 120 1768 1208 1832
rect 1272 1768 1292 1832
rect 120 1752 1292 1768
rect 120 1688 1208 1752
rect 1272 1688 1292 1752
rect 120 1672 1292 1688
rect 120 1608 1208 1672
rect 1272 1608 1292 1672
rect 120 1592 1292 1608
rect 120 1528 1208 1592
rect 1272 1528 1292 1592
rect 120 1512 1292 1528
rect 120 1448 1208 1512
rect 1272 1448 1292 1512
rect 120 1432 1292 1448
rect 120 1368 1208 1432
rect 1272 1368 1292 1432
rect 120 1352 1292 1368
rect 120 1288 1208 1352
rect 1272 1288 1292 1352
rect 120 1240 1292 1288
rect 1532 2072 2704 2120
rect 1532 2008 2620 2072
rect 2684 2008 2704 2072
rect 1532 1992 2704 2008
rect 1532 1928 2620 1992
rect 2684 1928 2704 1992
rect 1532 1912 2704 1928
rect 1532 1848 2620 1912
rect 2684 1848 2704 1912
rect 1532 1832 2704 1848
rect 1532 1768 2620 1832
rect 2684 1768 2704 1832
rect 1532 1752 2704 1768
rect 1532 1688 2620 1752
rect 2684 1688 2704 1752
rect 1532 1672 2704 1688
rect 1532 1608 2620 1672
rect 2684 1608 2704 1672
rect 1532 1592 2704 1608
rect 1532 1528 2620 1592
rect 2684 1528 2704 1592
rect 1532 1512 2704 1528
rect 1532 1448 2620 1512
rect 2684 1448 2704 1512
rect 1532 1432 2704 1448
rect 1532 1368 2620 1432
rect 2684 1368 2704 1432
rect 1532 1352 2704 1368
rect 1532 1288 2620 1352
rect 2684 1288 2704 1352
rect 1532 1240 2704 1288
rect -2704 952 -1532 1000
rect -2704 888 -1616 952
rect -1552 888 -1532 952
rect -2704 872 -1532 888
rect -2704 808 -1616 872
rect -1552 808 -1532 872
rect -2704 792 -1532 808
rect -2704 728 -1616 792
rect -1552 728 -1532 792
rect -2704 712 -1532 728
rect -2704 648 -1616 712
rect -1552 648 -1532 712
rect -2704 632 -1532 648
rect -2704 568 -1616 632
rect -1552 568 -1532 632
rect -2704 552 -1532 568
rect -2704 488 -1616 552
rect -1552 488 -1532 552
rect -2704 472 -1532 488
rect -2704 408 -1616 472
rect -1552 408 -1532 472
rect -2704 392 -1532 408
rect -2704 328 -1616 392
rect -1552 328 -1532 392
rect -2704 312 -1532 328
rect -2704 248 -1616 312
rect -1552 248 -1532 312
rect -2704 232 -1532 248
rect -2704 168 -1616 232
rect -1552 168 -1532 232
rect -2704 120 -1532 168
rect -1292 952 -120 1000
rect -1292 888 -204 952
rect -140 888 -120 952
rect -1292 872 -120 888
rect -1292 808 -204 872
rect -140 808 -120 872
rect -1292 792 -120 808
rect -1292 728 -204 792
rect -140 728 -120 792
rect -1292 712 -120 728
rect -1292 648 -204 712
rect -140 648 -120 712
rect -1292 632 -120 648
rect -1292 568 -204 632
rect -140 568 -120 632
rect -1292 552 -120 568
rect -1292 488 -204 552
rect -140 488 -120 552
rect -1292 472 -120 488
rect -1292 408 -204 472
rect -140 408 -120 472
rect -1292 392 -120 408
rect -1292 328 -204 392
rect -140 328 -120 392
rect -1292 312 -120 328
rect -1292 248 -204 312
rect -140 248 -120 312
rect -1292 232 -120 248
rect -1292 168 -204 232
rect -140 168 -120 232
rect -1292 120 -120 168
rect 120 952 1292 1000
rect 120 888 1208 952
rect 1272 888 1292 952
rect 120 872 1292 888
rect 120 808 1208 872
rect 1272 808 1292 872
rect 120 792 1292 808
rect 120 728 1208 792
rect 1272 728 1292 792
rect 120 712 1292 728
rect 120 648 1208 712
rect 1272 648 1292 712
rect 120 632 1292 648
rect 120 568 1208 632
rect 1272 568 1292 632
rect 120 552 1292 568
rect 120 488 1208 552
rect 1272 488 1292 552
rect 120 472 1292 488
rect 120 408 1208 472
rect 1272 408 1292 472
rect 120 392 1292 408
rect 120 328 1208 392
rect 1272 328 1292 392
rect 120 312 1292 328
rect 120 248 1208 312
rect 1272 248 1292 312
rect 120 232 1292 248
rect 120 168 1208 232
rect 1272 168 1292 232
rect 120 120 1292 168
rect 1532 952 2704 1000
rect 1532 888 2620 952
rect 2684 888 2704 952
rect 1532 872 2704 888
rect 1532 808 2620 872
rect 2684 808 2704 872
rect 1532 792 2704 808
rect 1532 728 2620 792
rect 2684 728 2704 792
rect 1532 712 2704 728
rect 1532 648 2620 712
rect 2684 648 2704 712
rect 1532 632 2704 648
rect 1532 568 2620 632
rect 2684 568 2704 632
rect 1532 552 2704 568
rect 1532 488 2620 552
rect 2684 488 2704 552
rect 1532 472 2704 488
rect 1532 408 2620 472
rect 2684 408 2704 472
rect 1532 392 2704 408
rect 1532 328 2620 392
rect 2684 328 2704 392
rect 1532 312 2704 328
rect 1532 248 2620 312
rect 2684 248 2704 312
rect 1532 232 2704 248
rect 1532 168 2620 232
rect 2684 168 2704 232
rect 1532 120 2704 168
rect -2704 -168 -1532 -120
rect -2704 -232 -1616 -168
rect -1552 -232 -1532 -168
rect -2704 -248 -1532 -232
rect -2704 -312 -1616 -248
rect -1552 -312 -1532 -248
rect -2704 -328 -1532 -312
rect -2704 -392 -1616 -328
rect -1552 -392 -1532 -328
rect -2704 -408 -1532 -392
rect -2704 -472 -1616 -408
rect -1552 -472 -1532 -408
rect -2704 -488 -1532 -472
rect -2704 -552 -1616 -488
rect -1552 -552 -1532 -488
rect -2704 -568 -1532 -552
rect -2704 -632 -1616 -568
rect -1552 -632 -1532 -568
rect -2704 -648 -1532 -632
rect -2704 -712 -1616 -648
rect -1552 -712 -1532 -648
rect -2704 -728 -1532 -712
rect -2704 -792 -1616 -728
rect -1552 -792 -1532 -728
rect -2704 -808 -1532 -792
rect -2704 -872 -1616 -808
rect -1552 -872 -1532 -808
rect -2704 -888 -1532 -872
rect -2704 -952 -1616 -888
rect -1552 -952 -1532 -888
rect -2704 -1000 -1532 -952
rect -1292 -168 -120 -120
rect -1292 -232 -204 -168
rect -140 -232 -120 -168
rect -1292 -248 -120 -232
rect -1292 -312 -204 -248
rect -140 -312 -120 -248
rect -1292 -328 -120 -312
rect -1292 -392 -204 -328
rect -140 -392 -120 -328
rect -1292 -408 -120 -392
rect -1292 -472 -204 -408
rect -140 -472 -120 -408
rect -1292 -488 -120 -472
rect -1292 -552 -204 -488
rect -140 -552 -120 -488
rect -1292 -568 -120 -552
rect -1292 -632 -204 -568
rect -140 -632 -120 -568
rect -1292 -648 -120 -632
rect -1292 -712 -204 -648
rect -140 -712 -120 -648
rect -1292 -728 -120 -712
rect -1292 -792 -204 -728
rect -140 -792 -120 -728
rect -1292 -808 -120 -792
rect -1292 -872 -204 -808
rect -140 -872 -120 -808
rect -1292 -888 -120 -872
rect -1292 -952 -204 -888
rect -140 -952 -120 -888
rect -1292 -1000 -120 -952
rect 120 -168 1292 -120
rect 120 -232 1208 -168
rect 1272 -232 1292 -168
rect 120 -248 1292 -232
rect 120 -312 1208 -248
rect 1272 -312 1292 -248
rect 120 -328 1292 -312
rect 120 -392 1208 -328
rect 1272 -392 1292 -328
rect 120 -408 1292 -392
rect 120 -472 1208 -408
rect 1272 -472 1292 -408
rect 120 -488 1292 -472
rect 120 -552 1208 -488
rect 1272 -552 1292 -488
rect 120 -568 1292 -552
rect 120 -632 1208 -568
rect 1272 -632 1292 -568
rect 120 -648 1292 -632
rect 120 -712 1208 -648
rect 1272 -712 1292 -648
rect 120 -728 1292 -712
rect 120 -792 1208 -728
rect 1272 -792 1292 -728
rect 120 -808 1292 -792
rect 120 -872 1208 -808
rect 1272 -872 1292 -808
rect 120 -888 1292 -872
rect 120 -952 1208 -888
rect 1272 -952 1292 -888
rect 120 -1000 1292 -952
rect 1532 -168 2704 -120
rect 1532 -232 2620 -168
rect 2684 -232 2704 -168
rect 1532 -248 2704 -232
rect 1532 -312 2620 -248
rect 2684 -312 2704 -248
rect 1532 -328 2704 -312
rect 1532 -392 2620 -328
rect 2684 -392 2704 -328
rect 1532 -408 2704 -392
rect 1532 -472 2620 -408
rect 2684 -472 2704 -408
rect 1532 -488 2704 -472
rect 1532 -552 2620 -488
rect 2684 -552 2704 -488
rect 1532 -568 2704 -552
rect 1532 -632 2620 -568
rect 2684 -632 2704 -568
rect 1532 -648 2704 -632
rect 1532 -712 2620 -648
rect 2684 -712 2704 -648
rect 1532 -728 2704 -712
rect 1532 -792 2620 -728
rect 2684 -792 2704 -728
rect 1532 -808 2704 -792
rect 1532 -872 2620 -808
rect 2684 -872 2704 -808
rect 1532 -888 2704 -872
rect 1532 -952 2620 -888
rect 2684 -952 2704 -888
rect 1532 -1000 2704 -952
rect -2704 -1288 -1532 -1240
rect -2704 -1352 -1616 -1288
rect -1552 -1352 -1532 -1288
rect -2704 -1368 -1532 -1352
rect -2704 -1432 -1616 -1368
rect -1552 -1432 -1532 -1368
rect -2704 -1448 -1532 -1432
rect -2704 -1512 -1616 -1448
rect -1552 -1512 -1532 -1448
rect -2704 -1528 -1532 -1512
rect -2704 -1592 -1616 -1528
rect -1552 -1592 -1532 -1528
rect -2704 -1608 -1532 -1592
rect -2704 -1672 -1616 -1608
rect -1552 -1672 -1532 -1608
rect -2704 -1688 -1532 -1672
rect -2704 -1752 -1616 -1688
rect -1552 -1752 -1532 -1688
rect -2704 -1768 -1532 -1752
rect -2704 -1832 -1616 -1768
rect -1552 -1832 -1532 -1768
rect -2704 -1848 -1532 -1832
rect -2704 -1912 -1616 -1848
rect -1552 -1912 -1532 -1848
rect -2704 -1928 -1532 -1912
rect -2704 -1992 -1616 -1928
rect -1552 -1992 -1532 -1928
rect -2704 -2008 -1532 -1992
rect -2704 -2072 -1616 -2008
rect -1552 -2072 -1532 -2008
rect -2704 -2120 -1532 -2072
rect -1292 -1288 -120 -1240
rect -1292 -1352 -204 -1288
rect -140 -1352 -120 -1288
rect -1292 -1368 -120 -1352
rect -1292 -1432 -204 -1368
rect -140 -1432 -120 -1368
rect -1292 -1448 -120 -1432
rect -1292 -1512 -204 -1448
rect -140 -1512 -120 -1448
rect -1292 -1528 -120 -1512
rect -1292 -1592 -204 -1528
rect -140 -1592 -120 -1528
rect -1292 -1608 -120 -1592
rect -1292 -1672 -204 -1608
rect -140 -1672 -120 -1608
rect -1292 -1688 -120 -1672
rect -1292 -1752 -204 -1688
rect -140 -1752 -120 -1688
rect -1292 -1768 -120 -1752
rect -1292 -1832 -204 -1768
rect -140 -1832 -120 -1768
rect -1292 -1848 -120 -1832
rect -1292 -1912 -204 -1848
rect -140 -1912 -120 -1848
rect -1292 -1928 -120 -1912
rect -1292 -1992 -204 -1928
rect -140 -1992 -120 -1928
rect -1292 -2008 -120 -1992
rect -1292 -2072 -204 -2008
rect -140 -2072 -120 -2008
rect -1292 -2120 -120 -2072
rect 120 -1288 1292 -1240
rect 120 -1352 1208 -1288
rect 1272 -1352 1292 -1288
rect 120 -1368 1292 -1352
rect 120 -1432 1208 -1368
rect 1272 -1432 1292 -1368
rect 120 -1448 1292 -1432
rect 120 -1512 1208 -1448
rect 1272 -1512 1292 -1448
rect 120 -1528 1292 -1512
rect 120 -1592 1208 -1528
rect 1272 -1592 1292 -1528
rect 120 -1608 1292 -1592
rect 120 -1672 1208 -1608
rect 1272 -1672 1292 -1608
rect 120 -1688 1292 -1672
rect 120 -1752 1208 -1688
rect 1272 -1752 1292 -1688
rect 120 -1768 1292 -1752
rect 120 -1832 1208 -1768
rect 1272 -1832 1292 -1768
rect 120 -1848 1292 -1832
rect 120 -1912 1208 -1848
rect 1272 -1912 1292 -1848
rect 120 -1928 1292 -1912
rect 120 -1992 1208 -1928
rect 1272 -1992 1292 -1928
rect 120 -2008 1292 -1992
rect 120 -2072 1208 -2008
rect 1272 -2072 1292 -2008
rect 120 -2120 1292 -2072
rect 1532 -1288 2704 -1240
rect 1532 -1352 2620 -1288
rect 2684 -1352 2704 -1288
rect 1532 -1368 2704 -1352
rect 1532 -1432 2620 -1368
rect 2684 -1432 2704 -1368
rect 1532 -1448 2704 -1432
rect 1532 -1512 2620 -1448
rect 2684 -1512 2704 -1448
rect 1532 -1528 2704 -1512
rect 1532 -1592 2620 -1528
rect 2684 -1592 2704 -1528
rect 1532 -1608 2704 -1592
rect 1532 -1672 2620 -1608
rect 2684 -1672 2704 -1608
rect 1532 -1688 2704 -1672
rect 1532 -1752 2620 -1688
rect 2684 -1752 2704 -1688
rect 1532 -1768 2704 -1752
rect 1532 -1832 2620 -1768
rect 2684 -1832 2704 -1768
rect 1532 -1848 2704 -1832
rect 1532 -1912 2620 -1848
rect 2684 -1912 2704 -1848
rect 1532 -1928 2704 -1912
rect 1532 -1992 2620 -1928
rect 2684 -1992 2704 -1928
rect 1532 -2008 2704 -1992
rect 1532 -2072 2620 -2008
rect 2684 -2072 2704 -2008
rect 1532 -2120 2704 -2072
rect -2704 -2408 -1532 -2360
rect -2704 -2472 -1616 -2408
rect -1552 -2472 -1532 -2408
rect -2704 -2488 -1532 -2472
rect -2704 -2552 -1616 -2488
rect -1552 -2552 -1532 -2488
rect -2704 -2568 -1532 -2552
rect -2704 -2632 -1616 -2568
rect -1552 -2632 -1532 -2568
rect -2704 -2648 -1532 -2632
rect -2704 -2712 -1616 -2648
rect -1552 -2712 -1532 -2648
rect -2704 -2728 -1532 -2712
rect -2704 -2792 -1616 -2728
rect -1552 -2792 -1532 -2728
rect -2704 -2808 -1532 -2792
rect -2704 -2872 -1616 -2808
rect -1552 -2872 -1532 -2808
rect -2704 -2888 -1532 -2872
rect -2704 -2952 -1616 -2888
rect -1552 -2952 -1532 -2888
rect -2704 -2968 -1532 -2952
rect -2704 -3032 -1616 -2968
rect -1552 -3032 -1532 -2968
rect -2704 -3048 -1532 -3032
rect -2704 -3112 -1616 -3048
rect -1552 -3112 -1532 -3048
rect -2704 -3128 -1532 -3112
rect -2704 -3192 -1616 -3128
rect -1552 -3192 -1532 -3128
rect -2704 -3240 -1532 -3192
rect -1292 -2408 -120 -2360
rect -1292 -2472 -204 -2408
rect -140 -2472 -120 -2408
rect -1292 -2488 -120 -2472
rect -1292 -2552 -204 -2488
rect -140 -2552 -120 -2488
rect -1292 -2568 -120 -2552
rect -1292 -2632 -204 -2568
rect -140 -2632 -120 -2568
rect -1292 -2648 -120 -2632
rect -1292 -2712 -204 -2648
rect -140 -2712 -120 -2648
rect -1292 -2728 -120 -2712
rect -1292 -2792 -204 -2728
rect -140 -2792 -120 -2728
rect -1292 -2808 -120 -2792
rect -1292 -2872 -204 -2808
rect -140 -2872 -120 -2808
rect -1292 -2888 -120 -2872
rect -1292 -2952 -204 -2888
rect -140 -2952 -120 -2888
rect -1292 -2968 -120 -2952
rect -1292 -3032 -204 -2968
rect -140 -3032 -120 -2968
rect -1292 -3048 -120 -3032
rect -1292 -3112 -204 -3048
rect -140 -3112 -120 -3048
rect -1292 -3128 -120 -3112
rect -1292 -3192 -204 -3128
rect -140 -3192 -120 -3128
rect -1292 -3240 -120 -3192
rect 120 -2408 1292 -2360
rect 120 -2472 1208 -2408
rect 1272 -2472 1292 -2408
rect 120 -2488 1292 -2472
rect 120 -2552 1208 -2488
rect 1272 -2552 1292 -2488
rect 120 -2568 1292 -2552
rect 120 -2632 1208 -2568
rect 1272 -2632 1292 -2568
rect 120 -2648 1292 -2632
rect 120 -2712 1208 -2648
rect 1272 -2712 1292 -2648
rect 120 -2728 1292 -2712
rect 120 -2792 1208 -2728
rect 1272 -2792 1292 -2728
rect 120 -2808 1292 -2792
rect 120 -2872 1208 -2808
rect 1272 -2872 1292 -2808
rect 120 -2888 1292 -2872
rect 120 -2952 1208 -2888
rect 1272 -2952 1292 -2888
rect 120 -2968 1292 -2952
rect 120 -3032 1208 -2968
rect 1272 -3032 1292 -2968
rect 120 -3048 1292 -3032
rect 120 -3112 1208 -3048
rect 1272 -3112 1292 -3048
rect 120 -3128 1292 -3112
rect 120 -3192 1208 -3128
rect 1272 -3192 1292 -3128
rect 120 -3240 1292 -3192
rect 1532 -2408 2704 -2360
rect 1532 -2472 2620 -2408
rect 2684 -2472 2704 -2408
rect 1532 -2488 2704 -2472
rect 1532 -2552 2620 -2488
rect 2684 -2552 2704 -2488
rect 1532 -2568 2704 -2552
rect 1532 -2632 2620 -2568
rect 2684 -2632 2704 -2568
rect 1532 -2648 2704 -2632
rect 1532 -2712 2620 -2648
rect 2684 -2712 2704 -2648
rect 1532 -2728 2704 -2712
rect 1532 -2792 2620 -2728
rect 2684 -2792 2704 -2728
rect 1532 -2808 2704 -2792
rect 1532 -2872 2620 -2808
rect 2684 -2872 2704 -2808
rect 1532 -2888 2704 -2872
rect 1532 -2952 2620 -2888
rect 2684 -2952 2704 -2888
rect 1532 -2968 2704 -2952
rect 1532 -3032 2620 -2968
rect 2684 -3032 2704 -2968
rect 1532 -3048 2704 -3032
rect 1532 -3112 2620 -3048
rect 2684 -3112 2704 -3048
rect 1532 -3128 2704 -3112
rect 1532 -3192 2620 -3128
rect 2684 -3192 2704 -3128
rect 1532 -3240 2704 -3192
rect -2704 -3528 -1532 -3480
rect -2704 -3592 -1616 -3528
rect -1552 -3592 -1532 -3528
rect -2704 -3608 -1532 -3592
rect -2704 -3672 -1616 -3608
rect -1552 -3672 -1532 -3608
rect -2704 -3688 -1532 -3672
rect -2704 -3752 -1616 -3688
rect -1552 -3752 -1532 -3688
rect -2704 -3768 -1532 -3752
rect -2704 -3832 -1616 -3768
rect -1552 -3832 -1532 -3768
rect -2704 -3848 -1532 -3832
rect -2704 -3912 -1616 -3848
rect -1552 -3912 -1532 -3848
rect -2704 -3928 -1532 -3912
rect -2704 -3992 -1616 -3928
rect -1552 -3992 -1532 -3928
rect -2704 -4008 -1532 -3992
rect -2704 -4072 -1616 -4008
rect -1552 -4072 -1532 -4008
rect -2704 -4088 -1532 -4072
rect -2704 -4152 -1616 -4088
rect -1552 -4152 -1532 -4088
rect -2704 -4168 -1532 -4152
rect -2704 -4232 -1616 -4168
rect -1552 -4232 -1532 -4168
rect -2704 -4248 -1532 -4232
rect -2704 -4312 -1616 -4248
rect -1552 -4312 -1532 -4248
rect -2704 -4360 -1532 -4312
rect -1292 -3528 -120 -3480
rect -1292 -3592 -204 -3528
rect -140 -3592 -120 -3528
rect -1292 -3608 -120 -3592
rect -1292 -3672 -204 -3608
rect -140 -3672 -120 -3608
rect -1292 -3688 -120 -3672
rect -1292 -3752 -204 -3688
rect -140 -3752 -120 -3688
rect -1292 -3768 -120 -3752
rect -1292 -3832 -204 -3768
rect -140 -3832 -120 -3768
rect -1292 -3848 -120 -3832
rect -1292 -3912 -204 -3848
rect -140 -3912 -120 -3848
rect -1292 -3928 -120 -3912
rect -1292 -3992 -204 -3928
rect -140 -3992 -120 -3928
rect -1292 -4008 -120 -3992
rect -1292 -4072 -204 -4008
rect -140 -4072 -120 -4008
rect -1292 -4088 -120 -4072
rect -1292 -4152 -204 -4088
rect -140 -4152 -120 -4088
rect -1292 -4168 -120 -4152
rect -1292 -4232 -204 -4168
rect -140 -4232 -120 -4168
rect -1292 -4248 -120 -4232
rect -1292 -4312 -204 -4248
rect -140 -4312 -120 -4248
rect -1292 -4360 -120 -4312
rect 120 -3528 1292 -3480
rect 120 -3592 1208 -3528
rect 1272 -3592 1292 -3528
rect 120 -3608 1292 -3592
rect 120 -3672 1208 -3608
rect 1272 -3672 1292 -3608
rect 120 -3688 1292 -3672
rect 120 -3752 1208 -3688
rect 1272 -3752 1292 -3688
rect 120 -3768 1292 -3752
rect 120 -3832 1208 -3768
rect 1272 -3832 1292 -3768
rect 120 -3848 1292 -3832
rect 120 -3912 1208 -3848
rect 1272 -3912 1292 -3848
rect 120 -3928 1292 -3912
rect 120 -3992 1208 -3928
rect 1272 -3992 1292 -3928
rect 120 -4008 1292 -3992
rect 120 -4072 1208 -4008
rect 1272 -4072 1292 -4008
rect 120 -4088 1292 -4072
rect 120 -4152 1208 -4088
rect 1272 -4152 1292 -4088
rect 120 -4168 1292 -4152
rect 120 -4232 1208 -4168
rect 1272 -4232 1292 -4168
rect 120 -4248 1292 -4232
rect 120 -4312 1208 -4248
rect 1272 -4312 1292 -4248
rect 120 -4360 1292 -4312
rect 1532 -3528 2704 -3480
rect 1532 -3592 2620 -3528
rect 2684 -3592 2704 -3528
rect 1532 -3608 2704 -3592
rect 1532 -3672 2620 -3608
rect 2684 -3672 2704 -3608
rect 1532 -3688 2704 -3672
rect 1532 -3752 2620 -3688
rect 2684 -3752 2704 -3688
rect 1532 -3768 2704 -3752
rect 1532 -3832 2620 -3768
rect 2684 -3832 2704 -3768
rect 1532 -3848 2704 -3832
rect 1532 -3912 2620 -3848
rect 2684 -3912 2704 -3848
rect 1532 -3928 2704 -3912
rect 1532 -3992 2620 -3928
rect 2684 -3992 2704 -3928
rect 1532 -4008 2704 -3992
rect 1532 -4072 2620 -4008
rect 2684 -4072 2704 -4008
rect 1532 -4088 2704 -4072
rect 1532 -4152 2620 -4088
rect 2684 -4152 2704 -4088
rect 1532 -4168 2704 -4152
rect 1532 -4232 2620 -4168
rect 2684 -4232 2704 -4168
rect 1532 -4248 2704 -4232
rect 1532 -4312 2620 -4248
rect 2684 -4312 2704 -4248
rect 1532 -4360 2704 -4312
<< via3 >>
rect -1616 4248 -1552 4312
rect -1616 4168 -1552 4232
rect -1616 4088 -1552 4152
rect -1616 4008 -1552 4072
rect -1616 3928 -1552 3992
rect -1616 3848 -1552 3912
rect -1616 3768 -1552 3832
rect -1616 3688 -1552 3752
rect -1616 3608 -1552 3672
rect -1616 3528 -1552 3592
rect -204 4248 -140 4312
rect -204 4168 -140 4232
rect -204 4088 -140 4152
rect -204 4008 -140 4072
rect -204 3928 -140 3992
rect -204 3848 -140 3912
rect -204 3768 -140 3832
rect -204 3688 -140 3752
rect -204 3608 -140 3672
rect -204 3528 -140 3592
rect 1208 4248 1272 4312
rect 1208 4168 1272 4232
rect 1208 4088 1272 4152
rect 1208 4008 1272 4072
rect 1208 3928 1272 3992
rect 1208 3848 1272 3912
rect 1208 3768 1272 3832
rect 1208 3688 1272 3752
rect 1208 3608 1272 3672
rect 1208 3528 1272 3592
rect 2620 4248 2684 4312
rect 2620 4168 2684 4232
rect 2620 4088 2684 4152
rect 2620 4008 2684 4072
rect 2620 3928 2684 3992
rect 2620 3848 2684 3912
rect 2620 3768 2684 3832
rect 2620 3688 2684 3752
rect 2620 3608 2684 3672
rect 2620 3528 2684 3592
rect -1616 3128 -1552 3192
rect -1616 3048 -1552 3112
rect -1616 2968 -1552 3032
rect -1616 2888 -1552 2952
rect -1616 2808 -1552 2872
rect -1616 2728 -1552 2792
rect -1616 2648 -1552 2712
rect -1616 2568 -1552 2632
rect -1616 2488 -1552 2552
rect -1616 2408 -1552 2472
rect -204 3128 -140 3192
rect -204 3048 -140 3112
rect -204 2968 -140 3032
rect -204 2888 -140 2952
rect -204 2808 -140 2872
rect -204 2728 -140 2792
rect -204 2648 -140 2712
rect -204 2568 -140 2632
rect -204 2488 -140 2552
rect -204 2408 -140 2472
rect 1208 3128 1272 3192
rect 1208 3048 1272 3112
rect 1208 2968 1272 3032
rect 1208 2888 1272 2952
rect 1208 2808 1272 2872
rect 1208 2728 1272 2792
rect 1208 2648 1272 2712
rect 1208 2568 1272 2632
rect 1208 2488 1272 2552
rect 1208 2408 1272 2472
rect 2620 3128 2684 3192
rect 2620 3048 2684 3112
rect 2620 2968 2684 3032
rect 2620 2888 2684 2952
rect 2620 2808 2684 2872
rect 2620 2728 2684 2792
rect 2620 2648 2684 2712
rect 2620 2568 2684 2632
rect 2620 2488 2684 2552
rect 2620 2408 2684 2472
rect -1616 2008 -1552 2072
rect -1616 1928 -1552 1992
rect -1616 1848 -1552 1912
rect -1616 1768 -1552 1832
rect -1616 1688 -1552 1752
rect -1616 1608 -1552 1672
rect -1616 1528 -1552 1592
rect -1616 1448 -1552 1512
rect -1616 1368 -1552 1432
rect -1616 1288 -1552 1352
rect -204 2008 -140 2072
rect -204 1928 -140 1992
rect -204 1848 -140 1912
rect -204 1768 -140 1832
rect -204 1688 -140 1752
rect -204 1608 -140 1672
rect -204 1528 -140 1592
rect -204 1448 -140 1512
rect -204 1368 -140 1432
rect -204 1288 -140 1352
rect 1208 2008 1272 2072
rect 1208 1928 1272 1992
rect 1208 1848 1272 1912
rect 1208 1768 1272 1832
rect 1208 1688 1272 1752
rect 1208 1608 1272 1672
rect 1208 1528 1272 1592
rect 1208 1448 1272 1512
rect 1208 1368 1272 1432
rect 1208 1288 1272 1352
rect 2620 2008 2684 2072
rect 2620 1928 2684 1992
rect 2620 1848 2684 1912
rect 2620 1768 2684 1832
rect 2620 1688 2684 1752
rect 2620 1608 2684 1672
rect 2620 1528 2684 1592
rect 2620 1448 2684 1512
rect 2620 1368 2684 1432
rect 2620 1288 2684 1352
rect -1616 888 -1552 952
rect -1616 808 -1552 872
rect -1616 728 -1552 792
rect -1616 648 -1552 712
rect -1616 568 -1552 632
rect -1616 488 -1552 552
rect -1616 408 -1552 472
rect -1616 328 -1552 392
rect -1616 248 -1552 312
rect -1616 168 -1552 232
rect -204 888 -140 952
rect -204 808 -140 872
rect -204 728 -140 792
rect -204 648 -140 712
rect -204 568 -140 632
rect -204 488 -140 552
rect -204 408 -140 472
rect -204 328 -140 392
rect -204 248 -140 312
rect -204 168 -140 232
rect 1208 888 1272 952
rect 1208 808 1272 872
rect 1208 728 1272 792
rect 1208 648 1272 712
rect 1208 568 1272 632
rect 1208 488 1272 552
rect 1208 408 1272 472
rect 1208 328 1272 392
rect 1208 248 1272 312
rect 1208 168 1272 232
rect 2620 888 2684 952
rect 2620 808 2684 872
rect 2620 728 2684 792
rect 2620 648 2684 712
rect 2620 568 2684 632
rect 2620 488 2684 552
rect 2620 408 2684 472
rect 2620 328 2684 392
rect 2620 248 2684 312
rect 2620 168 2684 232
rect -1616 -232 -1552 -168
rect -1616 -312 -1552 -248
rect -1616 -392 -1552 -328
rect -1616 -472 -1552 -408
rect -1616 -552 -1552 -488
rect -1616 -632 -1552 -568
rect -1616 -712 -1552 -648
rect -1616 -792 -1552 -728
rect -1616 -872 -1552 -808
rect -1616 -952 -1552 -888
rect -204 -232 -140 -168
rect -204 -312 -140 -248
rect -204 -392 -140 -328
rect -204 -472 -140 -408
rect -204 -552 -140 -488
rect -204 -632 -140 -568
rect -204 -712 -140 -648
rect -204 -792 -140 -728
rect -204 -872 -140 -808
rect -204 -952 -140 -888
rect 1208 -232 1272 -168
rect 1208 -312 1272 -248
rect 1208 -392 1272 -328
rect 1208 -472 1272 -408
rect 1208 -552 1272 -488
rect 1208 -632 1272 -568
rect 1208 -712 1272 -648
rect 1208 -792 1272 -728
rect 1208 -872 1272 -808
rect 1208 -952 1272 -888
rect 2620 -232 2684 -168
rect 2620 -312 2684 -248
rect 2620 -392 2684 -328
rect 2620 -472 2684 -408
rect 2620 -552 2684 -488
rect 2620 -632 2684 -568
rect 2620 -712 2684 -648
rect 2620 -792 2684 -728
rect 2620 -872 2684 -808
rect 2620 -952 2684 -888
rect -1616 -1352 -1552 -1288
rect -1616 -1432 -1552 -1368
rect -1616 -1512 -1552 -1448
rect -1616 -1592 -1552 -1528
rect -1616 -1672 -1552 -1608
rect -1616 -1752 -1552 -1688
rect -1616 -1832 -1552 -1768
rect -1616 -1912 -1552 -1848
rect -1616 -1992 -1552 -1928
rect -1616 -2072 -1552 -2008
rect -204 -1352 -140 -1288
rect -204 -1432 -140 -1368
rect -204 -1512 -140 -1448
rect -204 -1592 -140 -1528
rect -204 -1672 -140 -1608
rect -204 -1752 -140 -1688
rect -204 -1832 -140 -1768
rect -204 -1912 -140 -1848
rect -204 -1992 -140 -1928
rect -204 -2072 -140 -2008
rect 1208 -1352 1272 -1288
rect 1208 -1432 1272 -1368
rect 1208 -1512 1272 -1448
rect 1208 -1592 1272 -1528
rect 1208 -1672 1272 -1608
rect 1208 -1752 1272 -1688
rect 1208 -1832 1272 -1768
rect 1208 -1912 1272 -1848
rect 1208 -1992 1272 -1928
rect 1208 -2072 1272 -2008
rect 2620 -1352 2684 -1288
rect 2620 -1432 2684 -1368
rect 2620 -1512 2684 -1448
rect 2620 -1592 2684 -1528
rect 2620 -1672 2684 -1608
rect 2620 -1752 2684 -1688
rect 2620 -1832 2684 -1768
rect 2620 -1912 2684 -1848
rect 2620 -1992 2684 -1928
rect 2620 -2072 2684 -2008
rect -1616 -2472 -1552 -2408
rect -1616 -2552 -1552 -2488
rect -1616 -2632 -1552 -2568
rect -1616 -2712 -1552 -2648
rect -1616 -2792 -1552 -2728
rect -1616 -2872 -1552 -2808
rect -1616 -2952 -1552 -2888
rect -1616 -3032 -1552 -2968
rect -1616 -3112 -1552 -3048
rect -1616 -3192 -1552 -3128
rect -204 -2472 -140 -2408
rect -204 -2552 -140 -2488
rect -204 -2632 -140 -2568
rect -204 -2712 -140 -2648
rect -204 -2792 -140 -2728
rect -204 -2872 -140 -2808
rect -204 -2952 -140 -2888
rect -204 -3032 -140 -2968
rect -204 -3112 -140 -3048
rect -204 -3192 -140 -3128
rect 1208 -2472 1272 -2408
rect 1208 -2552 1272 -2488
rect 1208 -2632 1272 -2568
rect 1208 -2712 1272 -2648
rect 1208 -2792 1272 -2728
rect 1208 -2872 1272 -2808
rect 1208 -2952 1272 -2888
rect 1208 -3032 1272 -2968
rect 1208 -3112 1272 -3048
rect 1208 -3192 1272 -3128
rect 2620 -2472 2684 -2408
rect 2620 -2552 2684 -2488
rect 2620 -2632 2684 -2568
rect 2620 -2712 2684 -2648
rect 2620 -2792 2684 -2728
rect 2620 -2872 2684 -2808
rect 2620 -2952 2684 -2888
rect 2620 -3032 2684 -2968
rect 2620 -3112 2684 -3048
rect 2620 -3192 2684 -3128
rect -1616 -3592 -1552 -3528
rect -1616 -3672 -1552 -3608
rect -1616 -3752 -1552 -3688
rect -1616 -3832 -1552 -3768
rect -1616 -3912 -1552 -3848
rect -1616 -3992 -1552 -3928
rect -1616 -4072 -1552 -4008
rect -1616 -4152 -1552 -4088
rect -1616 -4232 -1552 -4168
rect -1616 -4312 -1552 -4248
rect -204 -3592 -140 -3528
rect -204 -3672 -140 -3608
rect -204 -3752 -140 -3688
rect -204 -3832 -140 -3768
rect -204 -3912 -140 -3848
rect -204 -3992 -140 -3928
rect -204 -4072 -140 -4008
rect -204 -4152 -140 -4088
rect -204 -4232 -140 -4168
rect -204 -4312 -140 -4248
rect 1208 -3592 1272 -3528
rect 1208 -3672 1272 -3608
rect 1208 -3752 1272 -3688
rect 1208 -3832 1272 -3768
rect 1208 -3912 1272 -3848
rect 1208 -3992 1272 -3928
rect 1208 -4072 1272 -4008
rect 1208 -4152 1272 -4088
rect 1208 -4232 1272 -4168
rect 1208 -4312 1272 -4248
rect 2620 -3592 2684 -3528
rect 2620 -3672 2684 -3608
rect 2620 -3752 2684 -3688
rect 2620 -3832 2684 -3768
rect 2620 -3912 2684 -3848
rect 2620 -3992 2684 -3928
rect 2620 -4072 2684 -4008
rect 2620 -4152 2684 -4088
rect 2620 -4232 2684 -4168
rect 2620 -4312 2684 -4248
<< mimcap >>
rect -2664 4272 -1864 4320
rect -2664 3568 -2616 4272
rect -1912 3568 -1864 4272
rect -2664 3520 -1864 3568
rect -1252 4272 -452 4320
rect -1252 3568 -1204 4272
rect -500 3568 -452 4272
rect -1252 3520 -452 3568
rect 160 4272 960 4320
rect 160 3568 208 4272
rect 912 3568 960 4272
rect 160 3520 960 3568
rect 1572 4272 2372 4320
rect 1572 3568 1620 4272
rect 2324 3568 2372 4272
rect 1572 3520 2372 3568
rect -2664 3152 -1864 3200
rect -2664 2448 -2616 3152
rect -1912 2448 -1864 3152
rect -2664 2400 -1864 2448
rect -1252 3152 -452 3200
rect -1252 2448 -1204 3152
rect -500 2448 -452 3152
rect -1252 2400 -452 2448
rect 160 3152 960 3200
rect 160 2448 208 3152
rect 912 2448 960 3152
rect 160 2400 960 2448
rect 1572 3152 2372 3200
rect 1572 2448 1620 3152
rect 2324 2448 2372 3152
rect 1572 2400 2372 2448
rect -2664 2032 -1864 2080
rect -2664 1328 -2616 2032
rect -1912 1328 -1864 2032
rect -2664 1280 -1864 1328
rect -1252 2032 -452 2080
rect -1252 1328 -1204 2032
rect -500 1328 -452 2032
rect -1252 1280 -452 1328
rect 160 2032 960 2080
rect 160 1328 208 2032
rect 912 1328 960 2032
rect 160 1280 960 1328
rect 1572 2032 2372 2080
rect 1572 1328 1620 2032
rect 2324 1328 2372 2032
rect 1572 1280 2372 1328
rect -2664 912 -1864 960
rect -2664 208 -2616 912
rect -1912 208 -1864 912
rect -2664 160 -1864 208
rect -1252 912 -452 960
rect -1252 208 -1204 912
rect -500 208 -452 912
rect -1252 160 -452 208
rect 160 912 960 960
rect 160 208 208 912
rect 912 208 960 912
rect 160 160 960 208
rect 1572 912 2372 960
rect 1572 208 1620 912
rect 2324 208 2372 912
rect 1572 160 2372 208
rect -2664 -208 -1864 -160
rect -2664 -912 -2616 -208
rect -1912 -912 -1864 -208
rect -2664 -960 -1864 -912
rect -1252 -208 -452 -160
rect -1252 -912 -1204 -208
rect -500 -912 -452 -208
rect -1252 -960 -452 -912
rect 160 -208 960 -160
rect 160 -912 208 -208
rect 912 -912 960 -208
rect 160 -960 960 -912
rect 1572 -208 2372 -160
rect 1572 -912 1620 -208
rect 2324 -912 2372 -208
rect 1572 -960 2372 -912
rect -2664 -1328 -1864 -1280
rect -2664 -2032 -2616 -1328
rect -1912 -2032 -1864 -1328
rect -2664 -2080 -1864 -2032
rect -1252 -1328 -452 -1280
rect -1252 -2032 -1204 -1328
rect -500 -2032 -452 -1328
rect -1252 -2080 -452 -2032
rect 160 -1328 960 -1280
rect 160 -2032 208 -1328
rect 912 -2032 960 -1328
rect 160 -2080 960 -2032
rect 1572 -1328 2372 -1280
rect 1572 -2032 1620 -1328
rect 2324 -2032 2372 -1328
rect 1572 -2080 2372 -2032
rect -2664 -2448 -1864 -2400
rect -2664 -3152 -2616 -2448
rect -1912 -3152 -1864 -2448
rect -2664 -3200 -1864 -3152
rect -1252 -2448 -452 -2400
rect -1252 -3152 -1204 -2448
rect -500 -3152 -452 -2448
rect -1252 -3200 -452 -3152
rect 160 -2448 960 -2400
rect 160 -3152 208 -2448
rect 912 -3152 960 -2448
rect 160 -3200 960 -3152
rect 1572 -2448 2372 -2400
rect 1572 -3152 1620 -2448
rect 2324 -3152 2372 -2448
rect 1572 -3200 2372 -3152
rect -2664 -3568 -1864 -3520
rect -2664 -4272 -2616 -3568
rect -1912 -4272 -1864 -3568
rect -2664 -4320 -1864 -4272
rect -1252 -3568 -452 -3520
rect -1252 -4272 -1204 -3568
rect -500 -4272 -452 -3568
rect -1252 -4320 -452 -4272
rect 160 -3568 960 -3520
rect 160 -4272 208 -3568
rect 912 -4272 960 -3568
rect 160 -4320 960 -4272
rect 1572 -3568 2372 -3520
rect 1572 -4272 1620 -3568
rect 2324 -4272 2372 -3568
rect 1572 -4320 2372 -4272
<< mimcapcontact >>
rect -2616 3568 -1912 4272
rect -1204 3568 -500 4272
rect 208 3568 912 4272
rect 1620 3568 2324 4272
rect -2616 2448 -1912 3152
rect -1204 2448 -500 3152
rect 208 2448 912 3152
rect 1620 2448 2324 3152
rect -2616 1328 -1912 2032
rect -1204 1328 -500 2032
rect 208 1328 912 2032
rect 1620 1328 2324 2032
rect -2616 208 -1912 912
rect -1204 208 -500 912
rect 208 208 912 912
rect 1620 208 2324 912
rect -2616 -912 -1912 -208
rect -1204 -912 -500 -208
rect 208 -912 912 -208
rect 1620 -912 2324 -208
rect -2616 -2032 -1912 -1328
rect -1204 -2032 -500 -1328
rect 208 -2032 912 -1328
rect 1620 -2032 2324 -1328
rect -2616 -3152 -1912 -2448
rect -1204 -3152 -500 -2448
rect 208 -3152 912 -2448
rect 1620 -3152 2324 -2448
rect -2616 -4272 -1912 -3568
rect -1204 -4272 -500 -3568
rect 208 -4272 912 -3568
rect 1620 -4272 2324 -3568
<< metal4 >>
rect -2316 4281 -2212 4480
rect -1636 4312 -1532 4480
rect -2625 4272 -1903 4281
rect -2625 3568 -2616 4272
rect -1912 3568 -1903 4272
rect -2625 3559 -1903 3568
rect -1636 4248 -1616 4312
rect -1552 4248 -1532 4312
rect -904 4281 -800 4480
rect -224 4312 -120 4480
rect -1636 4232 -1532 4248
rect -1636 4168 -1616 4232
rect -1552 4168 -1532 4232
rect -1636 4152 -1532 4168
rect -1636 4088 -1616 4152
rect -1552 4088 -1532 4152
rect -1636 4072 -1532 4088
rect -1636 4008 -1616 4072
rect -1552 4008 -1532 4072
rect -1636 3992 -1532 4008
rect -1636 3928 -1616 3992
rect -1552 3928 -1532 3992
rect -1636 3912 -1532 3928
rect -1636 3848 -1616 3912
rect -1552 3848 -1532 3912
rect -1636 3832 -1532 3848
rect -1636 3768 -1616 3832
rect -1552 3768 -1532 3832
rect -1636 3752 -1532 3768
rect -1636 3688 -1616 3752
rect -1552 3688 -1532 3752
rect -1636 3672 -1532 3688
rect -1636 3608 -1616 3672
rect -1552 3608 -1532 3672
rect -1636 3592 -1532 3608
rect -2316 3161 -2212 3559
rect -1636 3528 -1616 3592
rect -1552 3528 -1532 3592
rect -1213 4272 -491 4281
rect -1213 3568 -1204 4272
rect -500 3568 -491 4272
rect -1213 3559 -491 3568
rect -224 4248 -204 4312
rect -140 4248 -120 4312
rect 508 4281 612 4480
rect 1188 4312 1292 4480
rect -224 4232 -120 4248
rect -224 4168 -204 4232
rect -140 4168 -120 4232
rect -224 4152 -120 4168
rect -224 4088 -204 4152
rect -140 4088 -120 4152
rect -224 4072 -120 4088
rect -224 4008 -204 4072
rect -140 4008 -120 4072
rect -224 3992 -120 4008
rect -224 3928 -204 3992
rect -140 3928 -120 3992
rect -224 3912 -120 3928
rect -224 3848 -204 3912
rect -140 3848 -120 3912
rect -224 3832 -120 3848
rect -224 3768 -204 3832
rect -140 3768 -120 3832
rect -224 3752 -120 3768
rect -224 3688 -204 3752
rect -140 3688 -120 3752
rect -224 3672 -120 3688
rect -224 3608 -204 3672
rect -140 3608 -120 3672
rect -224 3592 -120 3608
rect -1636 3192 -1532 3528
rect -2625 3152 -1903 3161
rect -2625 2448 -2616 3152
rect -1912 2448 -1903 3152
rect -2625 2439 -1903 2448
rect -1636 3128 -1616 3192
rect -1552 3128 -1532 3192
rect -904 3161 -800 3559
rect -224 3528 -204 3592
rect -140 3528 -120 3592
rect 199 4272 921 4281
rect 199 3568 208 4272
rect 912 3568 921 4272
rect 199 3559 921 3568
rect 1188 4248 1208 4312
rect 1272 4248 1292 4312
rect 1920 4281 2024 4480
rect 2600 4312 2704 4480
rect 1188 4232 1292 4248
rect 1188 4168 1208 4232
rect 1272 4168 1292 4232
rect 1188 4152 1292 4168
rect 1188 4088 1208 4152
rect 1272 4088 1292 4152
rect 1188 4072 1292 4088
rect 1188 4008 1208 4072
rect 1272 4008 1292 4072
rect 1188 3992 1292 4008
rect 1188 3928 1208 3992
rect 1272 3928 1292 3992
rect 1188 3912 1292 3928
rect 1188 3848 1208 3912
rect 1272 3848 1292 3912
rect 1188 3832 1292 3848
rect 1188 3768 1208 3832
rect 1272 3768 1292 3832
rect 1188 3752 1292 3768
rect 1188 3688 1208 3752
rect 1272 3688 1292 3752
rect 1188 3672 1292 3688
rect 1188 3608 1208 3672
rect 1272 3608 1292 3672
rect 1188 3592 1292 3608
rect -224 3192 -120 3528
rect -1636 3112 -1532 3128
rect -1636 3048 -1616 3112
rect -1552 3048 -1532 3112
rect -1636 3032 -1532 3048
rect -1636 2968 -1616 3032
rect -1552 2968 -1532 3032
rect -1636 2952 -1532 2968
rect -1636 2888 -1616 2952
rect -1552 2888 -1532 2952
rect -1636 2872 -1532 2888
rect -1636 2808 -1616 2872
rect -1552 2808 -1532 2872
rect -1636 2792 -1532 2808
rect -1636 2728 -1616 2792
rect -1552 2728 -1532 2792
rect -1636 2712 -1532 2728
rect -1636 2648 -1616 2712
rect -1552 2648 -1532 2712
rect -1636 2632 -1532 2648
rect -1636 2568 -1616 2632
rect -1552 2568 -1532 2632
rect -1636 2552 -1532 2568
rect -1636 2488 -1616 2552
rect -1552 2488 -1532 2552
rect -1636 2472 -1532 2488
rect -2316 2041 -2212 2439
rect -1636 2408 -1616 2472
rect -1552 2408 -1532 2472
rect -1213 3152 -491 3161
rect -1213 2448 -1204 3152
rect -500 2448 -491 3152
rect -1213 2439 -491 2448
rect -224 3128 -204 3192
rect -140 3128 -120 3192
rect 508 3161 612 3559
rect 1188 3528 1208 3592
rect 1272 3528 1292 3592
rect 1611 4272 2333 4281
rect 1611 3568 1620 4272
rect 2324 3568 2333 4272
rect 1611 3559 2333 3568
rect 2600 4248 2620 4312
rect 2684 4248 2704 4312
rect 2600 4232 2704 4248
rect 2600 4168 2620 4232
rect 2684 4168 2704 4232
rect 2600 4152 2704 4168
rect 2600 4088 2620 4152
rect 2684 4088 2704 4152
rect 2600 4072 2704 4088
rect 2600 4008 2620 4072
rect 2684 4008 2704 4072
rect 2600 3992 2704 4008
rect 2600 3928 2620 3992
rect 2684 3928 2704 3992
rect 2600 3912 2704 3928
rect 2600 3848 2620 3912
rect 2684 3848 2704 3912
rect 2600 3832 2704 3848
rect 2600 3768 2620 3832
rect 2684 3768 2704 3832
rect 2600 3752 2704 3768
rect 2600 3688 2620 3752
rect 2684 3688 2704 3752
rect 2600 3672 2704 3688
rect 2600 3608 2620 3672
rect 2684 3608 2704 3672
rect 2600 3592 2704 3608
rect 1188 3192 1292 3528
rect -224 3112 -120 3128
rect -224 3048 -204 3112
rect -140 3048 -120 3112
rect -224 3032 -120 3048
rect -224 2968 -204 3032
rect -140 2968 -120 3032
rect -224 2952 -120 2968
rect -224 2888 -204 2952
rect -140 2888 -120 2952
rect -224 2872 -120 2888
rect -224 2808 -204 2872
rect -140 2808 -120 2872
rect -224 2792 -120 2808
rect -224 2728 -204 2792
rect -140 2728 -120 2792
rect -224 2712 -120 2728
rect -224 2648 -204 2712
rect -140 2648 -120 2712
rect -224 2632 -120 2648
rect -224 2568 -204 2632
rect -140 2568 -120 2632
rect -224 2552 -120 2568
rect -224 2488 -204 2552
rect -140 2488 -120 2552
rect -224 2472 -120 2488
rect -1636 2072 -1532 2408
rect -2625 2032 -1903 2041
rect -2625 1328 -2616 2032
rect -1912 1328 -1903 2032
rect -2625 1319 -1903 1328
rect -1636 2008 -1616 2072
rect -1552 2008 -1532 2072
rect -904 2041 -800 2439
rect -224 2408 -204 2472
rect -140 2408 -120 2472
rect 199 3152 921 3161
rect 199 2448 208 3152
rect 912 2448 921 3152
rect 199 2439 921 2448
rect 1188 3128 1208 3192
rect 1272 3128 1292 3192
rect 1920 3161 2024 3559
rect 2600 3528 2620 3592
rect 2684 3528 2704 3592
rect 2600 3192 2704 3528
rect 1188 3112 1292 3128
rect 1188 3048 1208 3112
rect 1272 3048 1292 3112
rect 1188 3032 1292 3048
rect 1188 2968 1208 3032
rect 1272 2968 1292 3032
rect 1188 2952 1292 2968
rect 1188 2888 1208 2952
rect 1272 2888 1292 2952
rect 1188 2872 1292 2888
rect 1188 2808 1208 2872
rect 1272 2808 1292 2872
rect 1188 2792 1292 2808
rect 1188 2728 1208 2792
rect 1272 2728 1292 2792
rect 1188 2712 1292 2728
rect 1188 2648 1208 2712
rect 1272 2648 1292 2712
rect 1188 2632 1292 2648
rect 1188 2568 1208 2632
rect 1272 2568 1292 2632
rect 1188 2552 1292 2568
rect 1188 2488 1208 2552
rect 1272 2488 1292 2552
rect 1188 2472 1292 2488
rect -224 2072 -120 2408
rect -1636 1992 -1532 2008
rect -1636 1928 -1616 1992
rect -1552 1928 -1532 1992
rect -1636 1912 -1532 1928
rect -1636 1848 -1616 1912
rect -1552 1848 -1532 1912
rect -1636 1832 -1532 1848
rect -1636 1768 -1616 1832
rect -1552 1768 -1532 1832
rect -1636 1752 -1532 1768
rect -1636 1688 -1616 1752
rect -1552 1688 -1532 1752
rect -1636 1672 -1532 1688
rect -1636 1608 -1616 1672
rect -1552 1608 -1532 1672
rect -1636 1592 -1532 1608
rect -1636 1528 -1616 1592
rect -1552 1528 -1532 1592
rect -1636 1512 -1532 1528
rect -1636 1448 -1616 1512
rect -1552 1448 -1532 1512
rect -1636 1432 -1532 1448
rect -1636 1368 -1616 1432
rect -1552 1368 -1532 1432
rect -1636 1352 -1532 1368
rect -2316 921 -2212 1319
rect -1636 1288 -1616 1352
rect -1552 1288 -1532 1352
rect -1213 2032 -491 2041
rect -1213 1328 -1204 2032
rect -500 1328 -491 2032
rect -1213 1319 -491 1328
rect -224 2008 -204 2072
rect -140 2008 -120 2072
rect 508 2041 612 2439
rect 1188 2408 1208 2472
rect 1272 2408 1292 2472
rect 1611 3152 2333 3161
rect 1611 2448 1620 3152
rect 2324 2448 2333 3152
rect 1611 2439 2333 2448
rect 2600 3128 2620 3192
rect 2684 3128 2704 3192
rect 2600 3112 2704 3128
rect 2600 3048 2620 3112
rect 2684 3048 2704 3112
rect 2600 3032 2704 3048
rect 2600 2968 2620 3032
rect 2684 2968 2704 3032
rect 2600 2952 2704 2968
rect 2600 2888 2620 2952
rect 2684 2888 2704 2952
rect 2600 2872 2704 2888
rect 2600 2808 2620 2872
rect 2684 2808 2704 2872
rect 2600 2792 2704 2808
rect 2600 2728 2620 2792
rect 2684 2728 2704 2792
rect 2600 2712 2704 2728
rect 2600 2648 2620 2712
rect 2684 2648 2704 2712
rect 2600 2632 2704 2648
rect 2600 2568 2620 2632
rect 2684 2568 2704 2632
rect 2600 2552 2704 2568
rect 2600 2488 2620 2552
rect 2684 2488 2704 2552
rect 2600 2472 2704 2488
rect 1188 2072 1292 2408
rect -224 1992 -120 2008
rect -224 1928 -204 1992
rect -140 1928 -120 1992
rect -224 1912 -120 1928
rect -224 1848 -204 1912
rect -140 1848 -120 1912
rect -224 1832 -120 1848
rect -224 1768 -204 1832
rect -140 1768 -120 1832
rect -224 1752 -120 1768
rect -224 1688 -204 1752
rect -140 1688 -120 1752
rect -224 1672 -120 1688
rect -224 1608 -204 1672
rect -140 1608 -120 1672
rect -224 1592 -120 1608
rect -224 1528 -204 1592
rect -140 1528 -120 1592
rect -224 1512 -120 1528
rect -224 1448 -204 1512
rect -140 1448 -120 1512
rect -224 1432 -120 1448
rect -224 1368 -204 1432
rect -140 1368 -120 1432
rect -224 1352 -120 1368
rect -1636 952 -1532 1288
rect -2625 912 -1903 921
rect -2625 208 -2616 912
rect -1912 208 -1903 912
rect -2625 199 -1903 208
rect -1636 888 -1616 952
rect -1552 888 -1532 952
rect -904 921 -800 1319
rect -224 1288 -204 1352
rect -140 1288 -120 1352
rect 199 2032 921 2041
rect 199 1328 208 2032
rect 912 1328 921 2032
rect 199 1319 921 1328
rect 1188 2008 1208 2072
rect 1272 2008 1292 2072
rect 1920 2041 2024 2439
rect 2600 2408 2620 2472
rect 2684 2408 2704 2472
rect 2600 2072 2704 2408
rect 1188 1992 1292 2008
rect 1188 1928 1208 1992
rect 1272 1928 1292 1992
rect 1188 1912 1292 1928
rect 1188 1848 1208 1912
rect 1272 1848 1292 1912
rect 1188 1832 1292 1848
rect 1188 1768 1208 1832
rect 1272 1768 1292 1832
rect 1188 1752 1292 1768
rect 1188 1688 1208 1752
rect 1272 1688 1292 1752
rect 1188 1672 1292 1688
rect 1188 1608 1208 1672
rect 1272 1608 1292 1672
rect 1188 1592 1292 1608
rect 1188 1528 1208 1592
rect 1272 1528 1292 1592
rect 1188 1512 1292 1528
rect 1188 1448 1208 1512
rect 1272 1448 1292 1512
rect 1188 1432 1292 1448
rect 1188 1368 1208 1432
rect 1272 1368 1292 1432
rect 1188 1352 1292 1368
rect -224 952 -120 1288
rect -1636 872 -1532 888
rect -1636 808 -1616 872
rect -1552 808 -1532 872
rect -1636 792 -1532 808
rect -1636 728 -1616 792
rect -1552 728 -1532 792
rect -1636 712 -1532 728
rect -1636 648 -1616 712
rect -1552 648 -1532 712
rect -1636 632 -1532 648
rect -1636 568 -1616 632
rect -1552 568 -1532 632
rect -1636 552 -1532 568
rect -1636 488 -1616 552
rect -1552 488 -1532 552
rect -1636 472 -1532 488
rect -1636 408 -1616 472
rect -1552 408 -1532 472
rect -1636 392 -1532 408
rect -1636 328 -1616 392
rect -1552 328 -1532 392
rect -1636 312 -1532 328
rect -1636 248 -1616 312
rect -1552 248 -1532 312
rect -1636 232 -1532 248
rect -2316 -199 -2212 199
rect -1636 168 -1616 232
rect -1552 168 -1532 232
rect -1213 912 -491 921
rect -1213 208 -1204 912
rect -500 208 -491 912
rect -1213 199 -491 208
rect -224 888 -204 952
rect -140 888 -120 952
rect 508 921 612 1319
rect 1188 1288 1208 1352
rect 1272 1288 1292 1352
rect 1611 2032 2333 2041
rect 1611 1328 1620 2032
rect 2324 1328 2333 2032
rect 1611 1319 2333 1328
rect 2600 2008 2620 2072
rect 2684 2008 2704 2072
rect 2600 1992 2704 2008
rect 2600 1928 2620 1992
rect 2684 1928 2704 1992
rect 2600 1912 2704 1928
rect 2600 1848 2620 1912
rect 2684 1848 2704 1912
rect 2600 1832 2704 1848
rect 2600 1768 2620 1832
rect 2684 1768 2704 1832
rect 2600 1752 2704 1768
rect 2600 1688 2620 1752
rect 2684 1688 2704 1752
rect 2600 1672 2704 1688
rect 2600 1608 2620 1672
rect 2684 1608 2704 1672
rect 2600 1592 2704 1608
rect 2600 1528 2620 1592
rect 2684 1528 2704 1592
rect 2600 1512 2704 1528
rect 2600 1448 2620 1512
rect 2684 1448 2704 1512
rect 2600 1432 2704 1448
rect 2600 1368 2620 1432
rect 2684 1368 2704 1432
rect 2600 1352 2704 1368
rect 1188 952 1292 1288
rect -224 872 -120 888
rect -224 808 -204 872
rect -140 808 -120 872
rect -224 792 -120 808
rect -224 728 -204 792
rect -140 728 -120 792
rect -224 712 -120 728
rect -224 648 -204 712
rect -140 648 -120 712
rect -224 632 -120 648
rect -224 568 -204 632
rect -140 568 -120 632
rect -224 552 -120 568
rect -224 488 -204 552
rect -140 488 -120 552
rect -224 472 -120 488
rect -224 408 -204 472
rect -140 408 -120 472
rect -224 392 -120 408
rect -224 328 -204 392
rect -140 328 -120 392
rect -224 312 -120 328
rect -224 248 -204 312
rect -140 248 -120 312
rect -224 232 -120 248
rect -1636 -168 -1532 168
rect -2625 -208 -1903 -199
rect -2625 -912 -2616 -208
rect -1912 -912 -1903 -208
rect -2625 -921 -1903 -912
rect -1636 -232 -1616 -168
rect -1552 -232 -1532 -168
rect -904 -199 -800 199
rect -224 168 -204 232
rect -140 168 -120 232
rect 199 912 921 921
rect 199 208 208 912
rect 912 208 921 912
rect 199 199 921 208
rect 1188 888 1208 952
rect 1272 888 1292 952
rect 1920 921 2024 1319
rect 2600 1288 2620 1352
rect 2684 1288 2704 1352
rect 2600 952 2704 1288
rect 1188 872 1292 888
rect 1188 808 1208 872
rect 1272 808 1292 872
rect 1188 792 1292 808
rect 1188 728 1208 792
rect 1272 728 1292 792
rect 1188 712 1292 728
rect 1188 648 1208 712
rect 1272 648 1292 712
rect 1188 632 1292 648
rect 1188 568 1208 632
rect 1272 568 1292 632
rect 1188 552 1292 568
rect 1188 488 1208 552
rect 1272 488 1292 552
rect 1188 472 1292 488
rect 1188 408 1208 472
rect 1272 408 1292 472
rect 1188 392 1292 408
rect 1188 328 1208 392
rect 1272 328 1292 392
rect 1188 312 1292 328
rect 1188 248 1208 312
rect 1272 248 1292 312
rect 1188 232 1292 248
rect -224 -168 -120 168
rect -1636 -248 -1532 -232
rect -1636 -312 -1616 -248
rect -1552 -312 -1532 -248
rect -1636 -328 -1532 -312
rect -1636 -392 -1616 -328
rect -1552 -392 -1532 -328
rect -1636 -408 -1532 -392
rect -1636 -472 -1616 -408
rect -1552 -472 -1532 -408
rect -1636 -488 -1532 -472
rect -1636 -552 -1616 -488
rect -1552 -552 -1532 -488
rect -1636 -568 -1532 -552
rect -1636 -632 -1616 -568
rect -1552 -632 -1532 -568
rect -1636 -648 -1532 -632
rect -1636 -712 -1616 -648
rect -1552 -712 -1532 -648
rect -1636 -728 -1532 -712
rect -1636 -792 -1616 -728
rect -1552 -792 -1532 -728
rect -1636 -808 -1532 -792
rect -1636 -872 -1616 -808
rect -1552 -872 -1532 -808
rect -1636 -888 -1532 -872
rect -2316 -1319 -2212 -921
rect -1636 -952 -1616 -888
rect -1552 -952 -1532 -888
rect -1213 -208 -491 -199
rect -1213 -912 -1204 -208
rect -500 -912 -491 -208
rect -1213 -921 -491 -912
rect -224 -232 -204 -168
rect -140 -232 -120 -168
rect 508 -199 612 199
rect 1188 168 1208 232
rect 1272 168 1292 232
rect 1611 912 2333 921
rect 1611 208 1620 912
rect 2324 208 2333 912
rect 1611 199 2333 208
rect 2600 888 2620 952
rect 2684 888 2704 952
rect 2600 872 2704 888
rect 2600 808 2620 872
rect 2684 808 2704 872
rect 2600 792 2704 808
rect 2600 728 2620 792
rect 2684 728 2704 792
rect 2600 712 2704 728
rect 2600 648 2620 712
rect 2684 648 2704 712
rect 2600 632 2704 648
rect 2600 568 2620 632
rect 2684 568 2704 632
rect 2600 552 2704 568
rect 2600 488 2620 552
rect 2684 488 2704 552
rect 2600 472 2704 488
rect 2600 408 2620 472
rect 2684 408 2704 472
rect 2600 392 2704 408
rect 2600 328 2620 392
rect 2684 328 2704 392
rect 2600 312 2704 328
rect 2600 248 2620 312
rect 2684 248 2704 312
rect 2600 232 2704 248
rect 1188 -168 1292 168
rect -224 -248 -120 -232
rect -224 -312 -204 -248
rect -140 -312 -120 -248
rect -224 -328 -120 -312
rect -224 -392 -204 -328
rect -140 -392 -120 -328
rect -224 -408 -120 -392
rect -224 -472 -204 -408
rect -140 -472 -120 -408
rect -224 -488 -120 -472
rect -224 -552 -204 -488
rect -140 -552 -120 -488
rect -224 -568 -120 -552
rect -224 -632 -204 -568
rect -140 -632 -120 -568
rect -224 -648 -120 -632
rect -224 -712 -204 -648
rect -140 -712 -120 -648
rect -224 -728 -120 -712
rect -224 -792 -204 -728
rect -140 -792 -120 -728
rect -224 -808 -120 -792
rect -224 -872 -204 -808
rect -140 -872 -120 -808
rect -224 -888 -120 -872
rect -1636 -1288 -1532 -952
rect -2625 -1328 -1903 -1319
rect -2625 -2032 -2616 -1328
rect -1912 -2032 -1903 -1328
rect -2625 -2041 -1903 -2032
rect -1636 -1352 -1616 -1288
rect -1552 -1352 -1532 -1288
rect -904 -1319 -800 -921
rect -224 -952 -204 -888
rect -140 -952 -120 -888
rect 199 -208 921 -199
rect 199 -912 208 -208
rect 912 -912 921 -208
rect 199 -921 921 -912
rect 1188 -232 1208 -168
rect 1272 -232 1292 -168
rect 1920 -199 2024 199
rect 2600 168 2620 232
rect 2684 168 2704 232
rect 2600 -168 2704 168
rect 1188 -248 1292 -232
rect 1188 -312 1208 -248
rect 1272 -312 1292 -248
rect 1188 -328 1292 -312
rect 1188 -392 1208 -328
rect 1272 -392 1292 -328
rect 1188 -408 1292 -392
rect 1188 -472 1208 -408
rect 1272 -472 1292 -408
rect 1188 -488 1292 -472
rect 1188 -552 1208 -488
rect 1272 -552 1292 -488
rect 1188 -568 1292 -552
rect 1188 -632 1208 -568
rect 1272 -632 1292 -568
rect 1188 -648 1292 -632
rect 1188 -712 1208 -648
rect 1272 -712 1292 -648
rect 1188 -728 1292 -712
rect 1188 -792 1208 -728
rect 1272 -792 1292 -728
rect 1188 -808 1292 -792
rect 1188 -872 1208 -808
rect 1272 -872 1292 -808
rect 1188 -888 1292 -872
rect -224 -1288 -120 -952
rect -1636 -1368 -1532 -1352
rect -1636 -1432 -1616 -1368
rect -1552 -1432 -1532 -1368
rect -1636 -1448 -1532 -1432
rect -1636 -1512 -1616 -1448
rect -1552 -1512 -1532 -1448
rect -1636 -1528 -1532 -1512
rect -1636 -1592 -1616 -1528
rect -1552 -1592 -1532 -1528
rect -1636 -1608 -1532 -1592
rect -1636 -1672 -1616 -1608
rect -1552 -1672 -1532 -1608
rect -1636 -1688 -1532 -1672
rect -1636 -1752 -1616 -1688
rect -1552 -1752 -1532 -1688
rect -1636 -1768 -1532 -1752
rect -1636 -1832 -1616 -1768
rect -1552 -1832 -1532 -1768
rect -1636 -1848 -1532 -1832
rect -1636 -1912 -1616 -1848
rect -1552 -1912 -1532 -1848
rect -1636 -1928 -1532 -1912
rect -1636 -1992 -1616 -1928
rect -1552 -1992 -1532 -1928
rect -1636 -2008 -1532 -1992
rect -2316 -2439 -2212 -2041
rect -1636 -2072 -1616 -2008
rect -1552 -2072 -1532 -2008
rect -1213 -1328 -491 -1319
rect -1213 -2032 -1204 -1328
rect -500 -2032 -491 -1328
rect -1213 -2041 -491 -2032
rect -224 -1352 -204 -1288
rect -140 -1352 -120 -1288
rect 508 -1319 612 -921
rect 1188 -952 1208 -888
rect 1272 -952 1292 -888
rect 1611 -208 2333 -199
rect 1611 -912 1620 -208
rect 2324 -912 2333 -208
rect 1611 -921 2333 -912
rect 2600 -232 2620 -168
rect 2684 -232 2704 -168
rect 2600 -248 2704 -232
rect 2600 -312 2620 -248
rect 2684 -312 2704 -248
rect 2600 -328 2704 -312
rect 2600 -392 2620 -328
rect 2684 -392 2704 -328
rect 2600 -408 2704 -392
rect 2600 -472 2620 -408
rect 2684 -472 2704 -408
rect 2600 -488 2704 -472
rect 2600 -552 2620 -488
rect 2684 -552 2704 -488
rect 2600 -568 2704 -552
rect 2600 -632 2620 -568
rect 2684 -632 2704 -568
rect 2600 -648 2704 -632
rect 2600 -712 2620 -648
rect 2684 -712 2704 -648
rect 2600 -728 2704 -712
rect 2600 -792 2620 -728
rect 2684 -792 2704 -728
rect 2600 -808 2704 -792
rect 2600 -872 2620 -808
rect 2684 -872 2704 -808
rect 2600 -888 2704 -872
rect 1188 -1288 1292 -952
rect -224 -1368 -120 -1352
rect -224 -1432 -204 -1368
rect -140 -1432 -120 -1368
rect -224 -1448 -120 -1432
rect -224 -1512 -204 -1448
rect -140 -1512 -120 -1448
rect -224 -1528 -120 -1512
rect -224 -1592 -204 -1528
rect -140 -1592 -120 -1528
rect -224 -1608 -120 -1592
rect -224 -1672 -204 -1608
rect -140 -1672 -120 -1608
rect -224 -1688 -120 -1672
rect -224 -1752 -204 -1688
rect -140 -1752 -120 -1688
rect -224 -1768 -120 -1752
rect -224 -1832 -204 -1768
rect -140 -1832 -120 -1768
rect -224 -1848 -120 -1832
rect -224 -1912 -204 -1848
rect -140 -1912 -120 -1848
rect -224 -1928 -120 -1912
rect -224 -1992 -204 -1928
rect -140 -1992 -120 -1928
rect -224 -2008 -120 -1992
rect -1636 -2408 -1532 -2072
rect -2625 -2448 -1903 -2439
rect -2625 -3152 -2616 -2448
rect -1912 -3152 -1903 -2448
rect -2625 -3161 -1903 -3152
rect -1636 -2472 -1616 -2408
rect -1552 -2472 -1532 -2408
rect -904 -2439 -800 -2041
rect -224 -2072 -204 -2008
rect -140 -2072 -120 -2008
rect 199 -1328 921 -1319
rect 199 -2032 208 -1328
rect 912 -2032 921 -1328
rect 199 -2041 921 -2032
rect 1188 -1352 1208 -1288
rect 1272 -1352 1292 -1288
rect 1920 -1319 2024 -921
rect 2600 -952 2620 -888
rect 2684 -952 2704 -888
rect 2600 -1288 2704 -952
rect 1188 -1368 1292 -1352
rect 1188 -1432 1208 -1368
rect 1272 -1432 1292 -1368
rect 1188 -1448 1292 -1432
rect 1188 -1512 1208 -1448
rect 1272 -1512 1292 -1448
rect 1188 -1528 1292 -1512
rect 1188 -1592 1208 -1528
rect 1272 -1592 1292 -1528
rect 1188 -1608 1292 -1592
rect 1188 -1672 1208 -1608
rect 1272 -1672 1292 -1608
rect 1188 -1688 1292 -1672
rect 1188 -1752 1208 -1688
rect 1272 -1752 1292 -1688
rect 1188 -1768 1292 -1752
rect 1188 -1832 1208 -1768
rect 1272 -1832 1292 -1768
rect 1188 -1848 1292 -1832
rect 1188 -1912 1208 -1848
rect 1272 -1912 1292 -1848
rect 1188 -1928 1292 -1912
rect 1188 -1992 1208 -1928
rect 1272 -1992 1292 -1928
rect 1188 -2008 1292 -1992
rect -224 -2408 -120 -2072
rect -1636 -2488 -1532 -2472
rect -1636 -2552 -1616 -2488
rect -1552 -2552 -1532 -2488
rect -1636 -2568 -1532 -2552
rect -1636 -2632 -1616 -2568
rect -1552 -2632 -1532 -2568
rect -1636 -2648 -1532 -2632
rect -1636 -2712 -1616 -2648
rect -1552 -2712 -1532 -2648
rect -1636 -2728 -1532 -2712
rect -1636 -2792 -1616 -2728
rect -1552 -2792 -1532 -2728
rect -1636 -2808 -1532 -2792
rect -1636 -2872 -1616 -2808
rect -1552 -2872 -1532 -2808
rect -1636 -2888 -1532 -2872
rect -1636 -2952 -1616 -2888
rect -1552 -2952 -1532 -2888
rect -1636 -2968 -1532 -2952
rect -1636 -3032 -1616 -2968
rect -1552 -3032 -1532 -2968
rect -1636 -3048 -1532 -3032
rect -1636 -3112 -1616 -3048
rect -1552 -3112 -1532 -3048
rect -1636 -3128 -1532 -3112
rect -2316 -3559 -2212 -3161
rect -1636 -3192 -1616 -3128
rect -1552 -3192 -1532 -3128
rect -1213 -2448 -491 -2439
rect -1213 -3152 -1204 -2448
rect -500 -3152 -491 -2448
rect -1213 -3161 -491 -3152
rect -224 -2472 -204 -2408
rect -140 -2472 -120 -2408
rect 508 -2439 612 -2041
rect 1188 -2072 1208 -2008
rect 1272 -2072 1292 -2008
rect 1611 -1328 2333 -1319
rect 1611 -2032 1620 -1328
rect 2324 -2032 2333 -1328
rect 1611 -2041 2333 -2032
rect 2600 -1352 2620 -1288
rect 2684 -1352 2704 -1288
rect 2600 -1368 2704 -1352
rect 2600 -1432 2620 -1368
rect 2684 -1432 2704 -1368
rect 2600 -1448 2704 -1432
rect 2600 -1512 2620 -1448
rect 2684 -1512 2704 -1448
rect 2600 -1528 2704 -1512
rect 2600 -1592 2620 -1528
rect 2684 -1592 2704 -1528
rect 2600 -1608 2704 -1592
rect 2600 -1672 2620 -1608
rect 2684 -1672 2704 -1608
rect 2600 -1688 2704 -1672
rect 2600 -1752 2620 -1688
rect 2684 -1752 2704 -1688
rect 2600 -1768 2704 -1752
rect 2600 -1832 2620 -1768
rect 2684 -1832 2704 -1768
rect 2600 -1848 2704 -1832
rect 2600 -1912 2620 -1848
rect 2684 -1912 2704 -1848
rect 2600 -1928 2704 -1912
rect 2600 -1992 2620 -1928
rect 2684 -1992 2704 -1928
rect 2600 -2008 2704 -1992
rect 1188 -2408 1292 -2072
rect -224 -2488 -120 -2472
rect -224 -2552 -204 -2488
rect -140 -2552 -120 -2488
rect -224 -2568 -120 -2552
rect -224 -2632 -204 -2568
rect -140 -2632 -120 -2568
rect -224 -2648 -120 -2632
rect -224 -2712 -204 -2648
rect -140 -2712 -120 -2648
rect -224 -2728 -120 -2712
rect -224 -2792 -204 -2728
rect -140 -2792 -120 -2728
rect -224 -2808 -120 -2792
rect -224 -2872 -204 -2808
rect -140 -2872 -120 -2808
rect -224 -2888 -120 -2872
rect -224 -2952 -204 -2888
rect -140 -2952 -120 -2888
rect -224 -2968 -120 -2952
rect -224 -3032 -204 -2968
rect -140 -3032 -120 -2968
rect -224 -3048 -120 -3032
rect -224 -3112 -204 -3048
rect -140 -3112 -120 -3048
rect -224 -3128 -120 -3112
rect -1636 -3528 -1532 -3192
rect -2625 -3568 -1903 -3559
rect -2625 -4272 -2616 -3568
rect -1912 -4272 -1903 -3568
rect -2625 -4281 -1903 -4272
rect -1636 -3592 -1616 -3528
rect -1552 -3592 -1532 -3528
rect -904 -3559 -800 -3161
rect -224 -3192 -204 -3128
rect -140 -3192 -120 -3128
rect 199 -2448 921 -2439
rect 199 -3152 208 -2448
rect 912 -3152 921 -2448
rect 199 -3161 921 -3152
rect 1188 -2472 1208 -2408
rect 1272 -2472 1292 -2408
rect 1920 -2439 2024 -2041
rect 2600 -2072 2620 -2008
rect 2684 -2072 2704 -2008
rect 2600 -2408 2704 -2072
rect 1188 -2488 1292 -2472
rect 1188 -2552 1208 -2488
rect 1272 -2552 1292 -2488
rect 1188 -2568 1292 -2552
rect 1188 -2632 1208 -2568
rect 1272 -2632 1292 -2568
rect 1188 -2648 1292 -2632
rect 1188 -2712 1208 -2648
rect 1272 -2712 1292 -2648
rect 1188 -2728 1292 -2712
rect 1188 -2792 1208 -2728
rect 1272 -2792 1292 -2728
rect 1188 -2808 1292 -2792
rect 1188 -2872 1208 -2808
rect 1272 -2872 1292 -2808
rect 1188 -2888 1292 -2872
rect 1188 -2952 1208 -2888
rect 1272 -2952 1292 -2888
rect 1188 -2968 1292 -2952
rect 1188 -3032 1208 -2968
rect 1272 -3032 1292 -2968
rect 1188 -3048 1292 -3032
rect 1188 -3112 1208 -3048
rect 1272 -3112 1292 -3048
rect 1188 -3128 1292 -3112
rect -224 -3528 -120 -3192
rect -1636 -3608 -1532 -3592
rect -1636 -3672 -1616 -3608
rect -1552 -3672 -1532 -3608
rect -1636 -3688 -1532 -3672
rect -1636 -3752 -1616 -3688
rect -1552 -3752 -1532 -3688
rect -1636 -3768 -1532 -3752
rect -1636 -3832 -1616 -3768
rect -1552 -3832 -1532 -3768
rect -1636 -3848 -1532 -3832
rect -1636 -3912 -1616 -3848
rect -1552 -3912 -1532 -3848
rect -1636 -3928 -1532 -3912
rect -1636 -3992 -1616 -3928
rect -1552 -3992 -1532 -3928
rect -1636 -4008 -1532 -3992
rect -1636 -4072 -1616 -4008
rect -1552 -4072 -1532 -4008
rect -1636 -4088 -1532 -4072
rect -1636 -4152 -1616 -4088
rect -1552 -4152 -1532 -4088
rect -1636 -4168 -1532 -4152
rect -1636 -4232 -1616 -4168
rect -1552 -4232 -1532 -4168
rect -1636 -4248 -1532 -4232
rect -2316 -4480 -2212 -4281
rect -1636 -4312 -1616 -4248
rect -1552 -4312 -1532 -4248
rect -1213 -3568 -491 -3559
rect -1213 -4272 -1204 -3568
rect -500 -4272 -491 -3568
rect -1213 -4281 -491 -4272
rect -224 -3592 -204 -3528
rect -140 -3592 -120 -3528
rect 508 -3559 612 -3161
rect 1188 -3192 1208 -3128
rect 1272 -3192 1292 -3128
rect 1611 -2448 2333 -2439
rect 1611 -3152 1620 -2448
rect 2324 -3152 2333 -2448
rect 1611 -3161 2333 -3152
rect 2600 -2472 2620 -2408
rect 2684 -2472 2704 -2408
rect 2600 -2488 2704 -2472
rect 2600 -2552 2620 -2488
rect 2684 -2552 2704 -2488
rect 2600 -2568 2704 -2552
rect 2600 -2632 2620 -2568
rect 2684 -2632 2704 -2568
rect 2600 -2648 2704 -2632
rect 2600 -2712 2620 -2648
rect 2684 -2712 2704 -2648
rect 2600 -2728 2704 -2712
rect 2600 -2792 2620 -2728
rect 2684 -2792 2704 -2728
rect 2600 -2808 2704 -2792
rect 2600 -2872 2620 -2808
rect 2684 -2872 2704 -2808
rect 2600 -2888 2704 -2872
rect 2600 -2952 2620 -2888
rect 2684 -2952 2704 -2888
rect 2600 -2968 2704 -2952
rect 2600 -3032 2620 -2968
rect 2684 -3032 2704 -2968
rect 2600 -3048 2704 -3032
rect 2600 -3112 2620 -3048
rect 2684 -3112 2704 -3048
rect 2600 -3128 2704 -3112
rect 1188 -3528 1292 -3192
rect -224 -3608 -120 -3592
rect -224 -3672 -204 -3608
rect -140 -3672 -120 -3608
rect -224 -3688 -120 -3672
rect -224 -3752 -204 -3688
rect -140 -3752 -120 -3688
rect -224 -3768 -120 -3752
rect -224 -3832 -204 -3768
rect -140 -3832 -120 -3768
rect -224 -3848 -120 -3832
rect -224 -3912 -204 -3848
rect -140 -3912 -120 -3848
rect -224 -3928 -120 -3912
rect -224 -3992 -204 -3928
rect -140 -3992 -120 -3928
rect -224 -4008 -120 -3992
rect -224 -4072 -204 -4008
rect -140 -4072 -120 -4008
rect -224 -4088 -120 -4072
rect -224 -4152 -204 -4088
rect -140 -4152 -120 -4088
rect -224 -4168 -120 -4152
rect -224 -4232 -204 -4168
rect -140 -4232 -120 -4168
rect -224 -4248 -120 -4232
rect -1636 -4480 -1532 -4312
rect -904 -4480 -800 -4281
rect -224 -4312 -204 -4248
rect -140 -4312 -120 -4248
rect 199 -3568 921 -3559
rect 199 -4272 208 -3568
rect 912 -4272 921 -3568
rect 199 -4281 921 -4272
rect 1188 -3592 1208 -3528
rect 1272 -3592 1292 -3528
rect 1920 -3559 2024 -3161
rect 2600 -3192 2620 -3128
rect 2684 -3192 2704 -3128
rect 2600 -3528 2704 -3192
rect 1188 -3608 1292 -3592
rect 1188 -3672 1208 -3608
rect 1272 -3672 1292 -3608
rect 1188 -3688 1292 -3672
rect 1188 -3752 1208 -3688
rect 1272 -3752 1292 -3688
rect 1188 -3768 1292 -3752
rect 1188 -3832 1208 -3768
rect 1272 -3832 1292 -3768
rect 1188 -3848 1292 -3832
rect 1188 -3912 1208 -3848
rect 1272 -3912 1292 -3848
rect 1188 -3928 1292 -3912
rect 1188 -3992 1208 -3928
rect 1272 -3992 1292 -3928
rect 1188 -4008 1292 -3992
rect 1188 -4072 1208 -4008
rect 1272 -4072 1292 -4008
rect 1188 -4088 1292 -4072
rect 1188 -4152 1208 -4088
rect 1272 -4152 1292 -4088
rect 1188 -4168 1292 -4152
rect 1188 -4232 1208 -4168
rect 1272 -4232 1292 -4168
rect 1188 -4248 1292 -4232
rect -224 -4480 -120 -4312
rect 508 -4480 612 -4281
rect 1188 -4312 1208 -4248
rect 1272 -4312 1292 -4248
rect 1611 -3568 2333 -3559
rect 1611 -4272 1620 -3568
rect 2324 -4272 2333 -3568
rect 1611 -4281 2333 -4272
rect 2600 -3592 2620 -3528
rect 2684 -3592 2704 -3528
rect 2600 -3608 2704 -3592
rect 2600 -3672 2620 -3608
rect 2684 -3672 2704 -3608
rect 2600 -3688 2704 -3672
rect 2600 -3752 2620 -3688
rect 2684 -3752 2704 -3688
rect 2600 -3768 2704 -3752
rect 2600 -3832 2620 -3768
rect 2684 -3832 2704 -3768
rect 2600 -3848 2704 -3832
rect 2600 -3912 2620 -3848
rect 2684 -3912 2704 -3848
rect 2600 -3928 2704 -3912
rect 2600 -3992 2620 -3928
rect 2684 -3992 2704 -3928
rect 2600 -4008 2704 -3992
rect 2600 -4072 2620 -4008
rect 2684 -4072 2704 -4008
rect 2600 -4088 2704 -4072
rect 2600 -4152 2620 -4088
rect 2684 -4152 2704 -4088
rect 2600 -4168 2704 -4152
rect 2600 -4232 2620 -4168
rect 2684 -4232 2704 -4168
rect 2600 -4248 2704 -4232
rect 1188 -4480 1292 -4312
rect 1920 -4480 2024 -4281
rect 2600 -4312 2620 -4248
rect 2684 -4312 2704 -4248
rect 2600 -4480 2704 -4312
<< properties >>
string FIXED_BBOX 1532 3480 2412 4360
<< end >>
