magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< pwell >>
rect -236 -1405 236 1405
<< nmos >>
rect -50 1105 50 1205
rect -50 895 50 995
rect -50 685 50 785
rect -50 475 50 575
rect -50 265 50 365
rect -50 55 50 155
rect -50 -155 50 -55
rect -50 -365 50 -265
rect -50 -575 50 -475
rect -50 -785 50 -685
rect -50 -995 50 -895
rect -50 -1205 50 -1105
<< ndiff >>
rect -108 1172 -50 1205
rect -108 1138 -96 1172
rect -62 1138 -50 1172
rect -108 1105 -50 1138
rect 50 1172 108 1205
rect 50 1138 62 1172
rect 96 1138 108 1172
rect 50 1105 108 1138
rect -108 962 -50 995
rect -108 928 -96 962
rect -62 928 -50 962
rect -108 895 -50 928
rect 50 962 108 995
rect 50 928 62 962
rect 96 928 108 962
rect 50 895 108 928
rect -108 752 -50 785
rect -108 718 -96 752
rect -62 718 -50 752
rect -108 685 -50 718
rect 50 752 108 785
rect 50 718 62 752
rect 96 718 108 752
rect 50 685 108 718
rect -108 542 -50 575
rect -108 508 -96 542
rect -62 508 -50 542
rect -108 475 -50 508
rect 50 542 108 575
rect 50 508 62 542
rect 96 508 108 542
rect 50 475 108 508
rect -108 332 -50 365
rect -108 298 -96 332
rect -62 298 -50 332
rect -108 265 -50 298
rect 50 332 108 365
rect 50 298 62 332
rect 96 298 108 332
rect 50 265 108 298
rect -108 122 -50 155
rect -108 88 -96 122
rect -62 88 -50 122
rect -108 55 -50 88
rect 50 122 108 155
rect 50 88 62 122
rect 96 88 108 122
rect 50 55 108 88
rect -108 -88 -50 -55
rect -108 -122 -96 -88
rect -62 -122 -50 -88
rect -108 -155 -50 -122
rect 50 -88 108 -55
rect 50 -122 62 -88
rect 96 -122 108 -88
rect 50 -155 108 -122
rect -108 -298 -50 -265
rect -108 -332 -96 -298
rect -62 -332 -50 -298
rect -108 -365 -50 -332
rect 50 -298 108 -265
rect 50 -332 62 -298
rect 96 -332 108 -298
rect 50 -365 108 -332
rect -108 -508 -50 -475
rect -108 -542 -96 -508
rect -62 -542 -50 -508
rect -108 -575 -50 -542
rect 50 -508 108 -475
rect 50 -542 62 -508
rect 96 -542 108 -508
rect 50 -575 108 -542
rect -108 -718 -50 -685
rect -108 -752 -96 -718
rect -62 -752 -50 -718
rect -108 -785 -50 -752
rect 50 -718 108 -685
rect 50 -752 62 -718
rect 96 -752 108 -718
rect 50 -785 108 -752
rect -108 -928 -50 -895
rect -108 -962 -96 -928
rect -62 -962 -50 -928
rect -108 -995 -50 -962
rect 50 -928 108 -895
rect 50 -962 62 -928
rect 96 -962 108 -928
rect 50 -995 108 -962
rect -108 -1138 -50 -1105
rect -108 -1172 -96 -1138
rect -62 -1172 -50 -1138
rect -108 -1205 -50 -1172
rect 50 -1138 108 -1105
rect 50 -1172 62 -1138
rect 96 -1172 108 -1138
rect 50 -1205 108 -1172
<< ndiffc >>
rect -96 1138 -62 1172
rect 62 1138 96 1172
rect -96 928 -62 962
rect 62 928 96 962
rect -96 718 -62 752
rect 62 718 96 752
rect -96 508 -62 542
rect 62 508 96 542
rect -96 298 -62 332
rect 62 298 96 332
rect -96 88 -62 122
rect 62 88 96 122
rect -96 -122 -62 -88
rect 62 -122 96 -88
rect -96 -332 -62 -298
rect 62 -332 96 -298
rect -96 -542 -62 -508
rect 62 -542 96 -508
rect -96 -752 -62 -718
rect 62 -752 96 -718
rect -96 -962 -62 -928
rect 62 -962 96 -928
rect -96 -1172 -62 -1138
rect 62 -1172 96 -1138
<< psubdiff >>
rect -210 1345 -85 1379
rect -51 1345 -17 1379
rect 17 1345 51 1379
rect 85 1345 210 1379
rect -210 1275 -176 1345
rect -210 1207 -176 1241
rect 176 1275 210 1345
rect 176 1207 210 1241
rect -210 1139 -176 1173
rect 176 1139 210 1173
rect -210 1071 -176 1105
rect -210 1003 -176 1037
rect 176 1071 210 1105
rect 176 1003 210 1037
rect -210 935 -176 969
rect -210 867 -176 901
rect 176 935 210 969
rect -210 799 -176 833
rect 176 867 210 901
rect 176 799 210 833
rect -210 731 -176 765
rect -210 663 -176 697
rect 176 731 210 765
rect -210 595 -176 629
rect 176 663 210 697
rect 176 595 210 629
rect -210 527 -176 561
rect -210 459 -176 493
rect 176 527 210 561
rect -210 391 -176 425
rect 176 459 210 493
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect 176 323 210 357
rect -210 187 -176 221
rect 176 255 210 289
rect 176 187 210 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect 176 -85 210 -51
rect 176 -153 210 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect 176 -221 210 -187
rect -210 -357 -176 -323
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect -210 -493 -176 -459
rect 176 -425 210 -391
rect -210 -561 -176 -527
rect 176 -493 210 -459
rect 176 -561 210 -527
rect -210 -629 -176 -595
rect -210 -697 -176 -663
rect 176 -629 210 -595
rect -210 -765 -176 -731
rect 176 -697 210 -663
rect 176 -765 210 -731
rect -210 -833 -176 -799
rect -210 -901 -176 -867
rect 176 -833 210 -799
rect -210 -969 -176 -935
rect 176 -901 210 -867
rect 176 -969 210 -935
rect -210 -1037 -176 -1003
rect -210 -1105 -176 -1071
rect 176 -1037 210 -1003
rect 176 -1105 210 -1071
rect -210 -1173 -176 -1139
rect 176 -1173 210 -1139
rect -210 -1241 -176 -1207
rect -210 -1345 -176 -1275
rect 176 -1241 210 -1207
rect 176 -1345 210 -1275
rect -210 -1379 -85 -1345
rect -51 -1379 -17 -1345
rect 17 -1379 51 -1345
rect 85 -1379 210 -1345
<< psubdiffcont >>
rect -85 1345 -51 1379
rect -17 1345 17 1379
rect 51 1345 85 1379
rect -210 1241 -176 1275
rect -210 1173 -176 1207
rect 176 1241 210 1275
rect -210 1105 -176 1139
rect 176 1173 210 1207
rect 176 1105 210 1139
rect -210 1037 -176 1071
rect -210 969 -176 1003
rect 176 1037 210 1071
rect -210 901 -176 935
rect 176 969 210 1003
rect 176 901 210 935
rect -210 833 -176 867
rect -210 765 -176 799
rect 176 833 210 867
rect -210 697 -176 731
rect 176 765 210 799
rect 176 697 210 731
rect -210 629 -176 663
rect -210 561 -176 595
rect 176 629 210 663
rect -210 493 -176 527
rect 176 561 210 595
rect 176 493 210 527
rect -210 425 -176 459
rect -210 357 -176 391
rect 176 425 210 459
rect -210 289 -176 323
rect 176 357 210 391
rect 176 289 210 323
rect -210 221 -176 255
rect -210 153 -176 187
rect 176 221 210 255
rect -210 85 -176 119
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect 176 -119 210 -85
rect -210 -255 -176 -221
rect 176 -187 210 -153
rect 176 -255 210 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect 176 -323 210 -289
rect -210 -459 -176 -425
rect 176 -391 210 -357
rect 176 -459 210 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect 176 -527 210 -493
rect -210 -663 -176 -629
rect 176 -595 210 -561
rect 176 -663 210 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect 176 -731 210 -697
rect -210 -867 -176 -833
rect 176 -799 210 -765
rect 176 -867 210 -833
rect -210 -935 -176 -901
rect -210 -1003 -176 -969
rect 176 -935 210 -901
rect -210 -1071 -176 -1037
rect 176 -1003 210 -969
rect 176 -1071 210 -1037
rect -210 -1139 -176 -1105
rect -210 -1207 -176 -1173
rect 176 -1139 210 -1105
rect -210 -1275 -176 -1241
rect 176 -1207 210 -1173
rect 176 -1275 210 -1241
rect -85 -1379 -51 -1345
rect -17 -1379 17 -1345
rect 51 -1379 85 -1345
<< poly >>
rect -50 1277 50 1293
rect -50 1243 -17 1277
rect 17 1243 50 1277
rect -50 1205 50 1243
rect -50 1067 50 1105
rect -50 1033 -17 1067
rect 17 1033 50 1067
rect -50 995 50 1033
rect -50 857 50 895
rect -50 823 -17 857
rect 17 823 50 857
rect -50 785 50 823
rect -50 647 50 685
rect -50 613 -17 647
rect 17 613 50 647
rect -50 575 50 613
rect -50 437 50 475
rect -50 403 -17 437
rect 17 403 50 437
rect -50 365 50 403
rect -50 227 50 265
rect -50 193 -17 227
rect 17 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect -50 -265 50 -227
rect -50 -403 50 -365
rect -50 -437 -17 -403
rect 17 -437 50 -403
rect -50 -475 50 -437
rect -50 -613 50 -575
rect -50 -647 -17 -613
rect 17 -647 50 -613
rect -50 -685 50 -647
rect -50 -823 50 -785
rect -50 -857 -17 -823
rect 17 -857 50 -823
rect -50 -895 50 -857
rect -50 -1033 50 -995
rect -50 -1067 -17 -1033
rect 17 -1067 50 -1033
rect -50 -1105 50 -1067
rect -50 -1243 50 -1205
rect -50 -1277 -17 -1243
rect 17 -1277 50 -1243
rect -50 -1293 50 -1277
<< polycont >>
rect -17 1243 17 1277
rect -17 1033 17 1067
rect -17 823 17 857
rect -17 613 17 647
rect -17 403 17 437
rect -17 193 17 227
rect -17 -17 17 17
rect -17 -227 17 -193
rect -17 -437 17 -403
rect -17 -647 17 -613
rect -17 -857 17 -823
rect -17 -1067 17 -1033
rect -17 -1277 17 -1243
<< locali >>
rect -210 1345 -85 1379
rect -51 1345 -17 1379
rect 17 1345 51 1379
rect 85 1345 210 1379
rect -210 1275 -176 1345
rect -50 1243 -17 1277
rect 17 1243 50 1277
rect 176 1275 210 1345
rect -210 1207 -176 1241
rect -210 1139 -176 1173
rect -210 1071 -176 1105
rect -96 1172 -62 1209
rect -96 1101 -62 1138
rect 62 1172 96 1209
rect 62 1101 96 1138
rect 176 1207 210 1241
rect 176 1139 210 1173
rect 176 1071 210 1105
rect -210 1003 -176 1037
rect -50 1033 -17 1067
rect 17 1033 50 1067
rect 176 1003 210 1037
rect -210 935 -176 969
rect -210 867 -176 901
rect -96 962 -62 999
rect -96 891 -62 928
rect 62 962 96 999
rect 62 891 96 928
rect 176 935 210 969
rect 176 867 210 901
rect -210 799 -176 833
rect -50 823 -17 857
rect 17 823 50 857
rect 176 799 210 833
rect -210 731 -176 765
rect -210 663 -176 697
rect -96 752 -62 789
rect -96 681 -62 718
rect 62 752 96 789
rect 62 681 96 718
rect 176 731 210 765
rect 176 663 210 697
rect -210 595 -176 629
rect -50 613 -17 647
rect 17 613 50 647
rect 176 595 210 629
rect -210 527 -176 561
rect -210 459 -176 493
rect -96 542 -62 579
rect -96 471 -62 508
rect 62 542 96 579
rect 62 471 96 508
rect 176 527 210 561
rect 176 459 210 493
rect -210 391 -176 425
rect -50 403 -17 437
rect 17 403 50 437
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -96 332 -62 369
rect -96 261 -62 298
rect 62 332 96 369
rect 62 261 96 298
rect 176 323 210 357
rect 176 255 210 289
rect -210 187 -176 221
rect -50 193 -17 227
rect 17 193 50 227
rect 176 187 210 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -96 122 -62 159
rect -96 51 -62 88
rect 62 122 96 159
rect 62 51 96 88
rect 176 119 210 153
rect 176 51 210 85
rect -210 -17 -176 17
rect -50 -17 -17 17
rect 17 -17 50 17
rect 176 -17 210 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -96 -88 -62 -51
rect -96 -159 -62 -122
rect 62 -88 96 -51
rect 62 -159 96 -122
rect 176 -85 210 -51
rect 176 -153 210 -119
rect -210 -221 -176 -187
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect 176 -221 210 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect -96 -298 -62 -261
rect -96 -369 -62 -332
rect 62 -298 96 -261
rect 62 -369 96 -332
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect -50 -437 -17 -403
rect 17 -437 50 -403
rect 176 -425 210 -391
rect -210 -493 -176 -459
rect -210 -561 -176 -527
rect -96 -508 -62 -471
rect -96 -579 -62 -542
rect 62 -508 96 -471
rect 62 -579 96 -542
rect 176 -493 210 -459
rect 176 -561 210 -527
rect -210 -629 -176 -595
rect -50 -647 -17 -613
rect 17 -647 50 -613
rect 176 -629 210 -595
rect -210 -697 -176 -663
rect -210 -765 -176 -731
rect -96 -718 -62 -681
rect -96 -789 -62 -752
rect 62 -718 96 -681
rect 62 -789 96 -752
rect 176 -697 210 -663
rect 176 -765 210 -731
rect -210 -833 -176 -799
rect -50 -857 -17 -823
rect 17 -857 50 -823
rect 176 -833 210 -799
rect -210 -901 -176 -867
rect -210 -969 -176 -935
rect -96 -928 -62 -891
rect -96 -999 -62 -962
rect 62 -928 96 -891
rect 62 -999 96 -962
rect 176 -901 210 -867
rect 176 -969 210 -935
rect -210 -1037 -176 -1003
rect -50 -1067 -17 -1033
rect 17 -1067 50 -1033
rect 176 -1037 210 -1003
rect -210 -1105 -176 -1071
rect -210 -1173 -176 -1139
rect -210 -1241 -176 -1207
rect -96 -1138 -62 -1101
rect -96 -1209 -62 -1172
rect 62 -1138 96 -1101
rect 62 -1209 96 -1172
rect 176 -1105 210 -1071
rect 176 -1173 210 -1139
rect 176 -1241 210 -1207
rect -210 -1345 -176 -1275
rect -50 -1277 -17 -1243
rect 17 -1277 50 -1243
rect 176 -1345 210 -1275
rect -210 -1379 -85 -1345
rect -51 -1379 -17 -1345
rect 17 -1379 51 -1345
rect 85 -1379 210 -1345
<< viali >>
rect -17 1243 17 1277
rect -96 1138 -62 1172
rect 62 1138 96 1172
rect -17 1033 17 1067
rect -96 928 -62 962
rect 62 928 96 962
rect -17 823 17 857
rect -96 718 -62 752
rect 62 718 96 752
rect -17 613 17 647
rect -96 508 -62 542
rect 62 508 96 542
rect -17 403 17 437
rect -96 298 -62 332
rect 62 298 96 332
rect -17 193 17 227
rect -96 88 -62 122
rect 62 88 96 122
rect -17 -17 17 17
rect -96 -122 -62 -88
rect 62 -122 96 -88
rect -17 -227 17 -193
rect -96 -332 -62 -298
rect 62 -332 96 -298
rect -17 -437 17 -403
rect -96 -542 -62 -508
rect 62 -542 96 -508
rect -17 -647 17 -613
rect -96 -752 -62 -718
rect 62 -752 96 -718
rect -17 -857 17 -823
rect -96 -962 -62 -928
rect 62 -962 96 -928
rect -17 -1067 17 -1033
rect -96 -1172 -62 -1138
rect 62 -1172 96 -1138
rect -17 -1277 17 -1243
<< metal1 >>
rect -46 1277 46 1283
rect -46 1243 -17 1277
rect 17 1243 46 1277
rect -46 1237 46 1243
rect -102 1172 -56 1205
rect -102 1138 -96 1172
rect -62 1138 -56 1172
rect -102 1105 -56 1138
rect 56 1172 102 1205
rect 56 1138 62 1172
rect 96 1138 102 1172
rect 56 1105 102 1138
rect -46 1067 46 1073
rect -46 1033 -17 1067
rect 17 1033 46 1067
rect -46 1027 46 1033
rect -102 962 -56 995
rect -102 928 -96 962
rect -62 928 -56 962
rect -102 895 -56 928
rect 56 962 102 995
rect 56 928 62 962
rect 96 928 102 962
rect 56 895 102 928
rect -46 857 46 863
rect -46 823 -17 857
rect 17 823 46 857
rect -46 817 46 823
rect -102 752 -56 785
rect -102 718 -96 752
rect -62 718 -56 752
rect -102 685 -56 718
rect 56 752 102 785
rect 56 718 62 752
rect 96 718 102 752
rect 56 685 102 718
rect -46 647 46 653
rect -46 613 -17 647
rect 17 613 46 647
rect -46 607 46 613
rect -102 542 -56 575
rect -102 508 -96 542
rect -62 508 -56 542
rect -102 475 -56 508
rect 56 542 102 575
rect 56 508 62 542
rect 96 508 102 542
rect 56 475 102 508
rect -46 437 46 443
rect -46 403 -17 437
rect 17 403 46 437
rect -46 397 46 403
rect -102 332 -56 365
rect -102 298 -96 332
rect -62 298 -56 332
rect -102 265 -56 298
rect 56 332 102 365
rect 56 298 62 332
rect 96 298 102 332
rect 56 265 102 298
rect -46 227 46 233
rect -46 193 -17 227
rect 17 193 46 227
rect -46 187 46 193
rect -102 122 -56 155
rect -102 88 -96 122
rect -62 88 -56 122
rect -102 55 -56 88
rect 56 122 102 155
rect 56 88 62 122
rect 96 88 102 122
rect 56 55 102 88
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -88 -56 -55
rect -102 -122 -96 -88
rect -62 -122 -56 -88
rect -102 -155 -56 -122
rect 56 -88 102 -55
rect 56 -122 62 -88
rect 96 -122 102 -88
rect 56 -155 102 -122
rect -46 -193 46 -187
rect -46 -227 -17 -193
rect 17 -227 46 -193
rect -46 -233 46 -227
rect -102 -298 -56 -265
rect -102 -332 -96 -298
rect -62 -332 -56 -298
rect -102 -365 -56 -332
rect 56 -298 102 -265
rect 56 -332 62 -298
rect 96 -332 102 -298
rect 56 -365 102 -332
rect -46 -403 46 -397
rect -46 -437 -17 -403
rect 17 -437 46 -403
rect -46 -443 46 -437
rect -102 -508 -56 -475
rect -102 -542 -96 -508
rect -62 -542 -56 -508
rect -102 -575 -56 -542
rect 56 -508 102 -475
rect 56 -542 62 -508
rect 96 -542 102 -508
rect 56 -575 102 -542
rect -46 -613 46 -607
rect -46 -647 -17 -613
rect 17 -647 46 -613
rect -46 -653 46 -647
rect -102 -718 -56 -685
rect -102 -752 -96 -718
rect -62 -752 -56 -718
rect -102 -785 -56 -752
rect 56 -718 102 -685
rect 56 -752 62 -718
rect 96 -752 102 -718
rect 56 -785 102 -752
rect -46 -823 46 -817
rect -46 -857 -17 -823
rect 17 -857 46 -823
rect -46 -863 46 -857
rect -102 -928 -56 -895
rect -102 -962 -96 -928
rect -62 -962 -56 -928
rect -102 -995 -56 -962
rect 56 -928 102 -895
rect 56 -962 62 -928
rect 96 -962 102 -928
rect 56 -995 102 -962
rect -46 -1033 46 -1027
rect -46 -1067 -17 -1033
rect 17 -1067 46 -1033
rect -46 -1073 46 -1067
rect -102 -1138 -56 -1105
rect -102 -1172 -96 -1138
rect -62 -1172 -56 -1138
rect -102 -1205 -56 -1172
rect 56 -1138 102 -1105
rect 56 -1172 62 -1138
rect 96 -1172 102 -1138
rect 56 -1205 102 -1172
rect -46 -1243 46 -1237
rect -46 -1277 -17 -1243
rect 17 -1277 46 -1243
rect -46 -1283 46 -1277
<< properties >>
string FIXED_BBOX -193 -1362 193 1362
<< end >>
