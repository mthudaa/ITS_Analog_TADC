magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< error_p >>
rect -29 2041 29 2047
rect -29 2007 -17 2041
rect -29 2001 29 2007
<< pwell >>
rect -201 -2169 201 2169
<< nmos >>
rect -15 -2031 15 1969
<< ndiff >>
rect -73 1924 -15 1969
rect -73 1890 -61 1924
rect -27 1890 -15 1924
rect -73 1856 -15 1890
rect -73 1822 -61 1856
rect -27 1822 -15 1856
rect -73 1788 -15 1822
rect -73 1754 -61 1788
rect -27 1754 -15 1788
rect -73 1720 -15 1754
rect -73 1686 -61 1720
rect -27 1686 -15 1720
rect -73 1652 -15 1686
rect -73 1618 -61 1652
rect -27 1618 -15 1652
rect -73 1584 -15 1618
rect -73 1550 -61 1584
rect -27 1550 -15 1584
rect -73 1516 -15 1550
rect -73 1482 -61 1516
rect -27 1482 -15 1516
rect -73 1448 -15 1482
rect -73 1414 -61 1448
rect -27 1414 -15 1448
rect -73 1380 -15 1414
rect -73 1346 -61 1380
rect -27 1346 -15 1380
rect -73 1312 -15 1346
rect -73 1278 -61 1312
rect -27 1278 -15 1312
rect -73 1244 -15 1278
rect -73 1210 -61 1244
rect -27 1210 -15 1244
rect -73 1176 -15 1210
rect -73 1142 -61 1176
rect -27 1142 -15 1176
rect -73 1108 -15 1142
rect -73 1074 -61 1108
rect -27 1074 -15 1108
rect -73 1040 -15 1074
rect -73 1006 -61 1040
rect -27 1006 -15 1040
rect -73 972 -15 1006
rect -73 938 -61 972
rect -27 938 -15 972
rect -73 904 -15 938
rect -73 870 -61 904
rect -27 870 -15 904
rect -73 836 -15 870
rect -73 802 -61 836
rect -27 802 -15 836
rect -73 768 -15 802
rect -73 734 -61 768
rect -27 734 -15 768
rect -73 700 -15 734
rect -73 666 -61 700
rect -27 666 -15 700
rect -73 632 -15 666
rect -73 598 -61 632
rect -27 598 -15 632
rect -73 564 -15 598
rect -73 530 -61 564
rect -27 530 -15 564
rect -73 496 -15 530
rect -73 462 -61 496
rect -27 462 -15 496
rect -73 428 -15 462
rect -73 394 -61 428
rect -27 394 -15 428
rect -73 360 -15 394
rect -73 326 -61 360
rect -27 326 -15 360
rect -73 292 -15 326
rect -73 258 -61 292
rect -27 258 -15 292
rect -73 224 -15 258
rect -73 190 -61 224
rect -27 190 -15 224
rect -73 156 -15 190
rect -73 122 -61 156
rect -27 122 -15 156
rect -73 88 -15 122
rect -73 54 -61 88
rect -27 54 -15 88
rect -73 20 -15 54
rect -73 -14 -61 20
rect -27 -14 -15 20
rect -73 -48 -15 -14
rect -73 -82 -61 -48
rect -27 -82 -15 -48
rect -73 -116 -15 -82
rect -73 -150 -61 -116
rect -27 -150 -15 -116
rect -73 -184 -15 -150
rect -73 -218 -61 -184
rect -27 -218 -15 -184
rect -73 -252 -15 -218
rect -73 -286 -61 -252
rect -27 -286 -15 -252
rect -73 -320 -15 -286
rect -73 -354 -61 -320
rect -27 -354 -15 -320
rect -73 -388 -15 -354
rect -73 -422 -61 -388
rect -27 -422 -15 -388
rect -73 -456 -15 -422
rect -73 -490 -61 -456
rect -27 -490 -15 -456
rect -73 -524 -15 -490
rect -73 -558 -61 -524
rect -27 -558 -15 -524
rect -73 -592 -15 -558
rect -73 -626 -61 -592
rect -27 -626 -15 -592
rect -73 -660 -15 -626
rect -73 -694 -61 -660
rect -27 -694 -15 -660
rect -73 -728 -15 -694
rect -73 -762 -61 -728
rect -27 -762 -15 -728
rect -73 -796 -15 -762
rect -73 -830 -61 -796
rect -27 -830 -15 -796
rect -73 -864 -15 -830
rect -73 -898 -61 -864
rect -27 -898 -15 -864
rect -73 -932 -15 -898
rect -73 -966 -61 -932
rect -27 -966 -15 -932
rect -73 -1000 -15 -966
rect -73 -1034 -61 -1000
rect -27 -1034 -15 -1000
rect -73 -1068 -15 -1034
rect -73 -1102 -61 -1068
rect -27 -1102 -15 -1068
rect -73 -1136 -15 -1102
rect -73 -1170 -61 -1136
rect -27 -1170 -15 -1136
rect -73 -1204 -15 -1170
rect -73 -1238 -61 -1204
rect -27 -1238 -15 -1204
rect -73 -1272 -15 -1238
rect -73 -1306 -61 -1272
rect -27 -1306 -15 -1272
rect -73 -1340 -15 -1306
rect -73 -1374 -61 -1340
rect -27 -1374 -15 -1340
rect -73 -1408 -15 -1374
rect -73 -1442 -61 -1408
rect -27 -1442 -15 -1408
rect -73 -1476 -15 -1442
rect -73 -1510 -61 -1476
rect -27 -1510 -15 -1476
rect -73 -1544 -15 -1510
rect -73 -1578 -61 -1544
rect -27 -1578 -15 -1544
rect -73 -1612 -15 -1578
rect -73 -1646 -61 -1612
rect -27 -1646 -15 -1612
rect -73 -1680 -15 -1646
rect -73 -1714 -61 -1680
rect -27 -1714 -15 -1680
rect -73 -1748 -15 -1714
rect -73 -1782 -61 -1748
rect -27 -1782 -15 -1748
rect -73 -1816 -15 -1782
rect -73 -1850 -61 -1816
rect -27 -1850 -15 -1816
rect -73 -1884 -15 -1850
rect -73 -1918 -61 -1884
rect -27 -1918 -15 -1884
rect -73 -1952 -15 -1918
rect -73 -1986 -61 -1952
rect -27 -1986 -15 -1952
rect -73 -2031 -15 -1986
rect 15 1924 73 1969
rect 15 1890 27 1924
rect 61 1890 73 1924
rect 15 1856 73 1890
rect 15 1822 27 1856
rect 61 1822 73 1856
rect 15 1788 73 1822
rect 15 1754 27 1788
rect 61 1754 73 1788
rect 15 1720 73 1754
rect 15 1686 27 1720
rect 61 1686 73 1720
rect 15 1652 73 1686
rect 15 1618 27 1652
rect 61 1618 73 1652
rect 15 1584 73 1618
rect 15 1550 27 1584
rect 61 1550 73 1584
rect 15 1516 73 1550
rect 15 1482 27 1516
rect 61 1482 73 1516
rect 15 1448 73 1482
rect 15 1414 27 1448
rect 61 1414 73 1448
rect 15 1380 73 1414
rect 15 1346 27 1380
rect 61 1346 73 1380
rect 15 1312 73 1346
rect 15 1278 27 1312
rect 61 1278 73 1312
rect 15 1244 73 1278
rect 15 1210 27 1244
rect 61 1210 73 1244
rect 15 1176 73 1210
rect 15 1142 27 1176
rect 61 1142 73 1176
rect 15 1108 73 1142
rect 15 1074 27 1108
rect 61 1074 73 1108
rect 15 1040 73 1074
rect 15 1006 27 1040
rect 61 1006 73 1040
rect 15 972 73 1006
rect 15 938 27 972
rect 61 938 73 972
rect 15 904 73 938
rect 15 870 27 904
rect 61 870 73 904
rect 15 836 73 870
rect 15 802 27 836
rect 61 802 73 836
rect 15 768 73 802
rect 15 734 27 768
rect 61 734 73 768
rect 15 700 73 734
rect 15 666 27 700
rect 61 666 73 700
rect 15 632 73 666
rect 15 598 27 632
rect 61 598 73 632
rect 15 564 73 598
rect 15 530 27 564
rect 61 530 73 564
rect 15 496 73 530
rect 15 462 27 496
rect 61 462 73 496
rect 15 428 73 462
rect 15 394 27 428
rect 61 394 73 428
rect 15 360 73 394
rect 15 326 27 360
rect 61 326 73 360
rect 15 292 73 326
rect 15 258 27 292
rect 61 258 73 292
rect 15 224 73 258
rect 15 190 27 224
rect 61 190 73 224
rect 15 156 73 190
rect 15 122 27 156
rect 61 122 73 156
rect 15 88 73 122
rect 15 54 27 88
rect 61 54 73 88
rect 15 20 73 54
rect 15 -14 27 20
rect 61 -14 73 20
rect 15 -48 73 -14
rect 15 -82 27 -48
rect 61 -82 73 -48
rect 15 -116 73 -82
rect 15 -150 27 -116
rect 61 -150 73 -116
rect 15 -184 73 -150
rect 15 -218 27 -184
rect 61 -218 73 -184
rect 15 -252 73 -218
rect 15 -286 27 -252
rect 61 -286 73 -252
rect 15 -320 73 -286
rect 15 -354 27 -320
rect 61 -354 73 -320
rect 15 -388 73 -354
rect 15 -422 27 -388
rect 61 -422 73 -388
rect 15 -456 73 -422
rect 15 -490 27 -456
rect 61 -490 73 -456
rect 15 -524 73 -490
rect 15 -558 27 -524
rect 61 -558 73 -524
rect 15 -592 73 -558
rect 15 -626 27 -592
rect 61 -626 73 -592
rect 15 -660 73 -626
rect 15 -694 27 -660
rect 61 -694 73 -660
rect 15 -728 73 -694
rect 15 -762 27 -728
rect 61 -762 73 -728
rect 15 -796 73 -762
rect 15 -830 27 -796
rect 61 -830 73 -796
rect 15 -864 73 -830
rect 15 -898 27 -864
rect 61 -898 73 -864
rect 15 -932 73 -898
rect 15 -966 27 -932
rect 61 -966 73 -932
rect 15 -1000 73 -966
rect 15 -1034 27 -1000
rect 61 -1034 73 -1000
rect 15 -1068 73 -1034
rect 15 -1102 27 -1068
rect 61 -1102 73 -1068
rect 15 -1136 73 -1102
rect 15 -1170 27 -1136
rect 61 -1170 73 -1136
rect 15 -1204 73 -1170
rect 15 -1238 27 -1204
rect 61 -1238 73 -1204
rect 15 -1272 73 -1238
rect 15 -1306 27 -1272
rect 61 -1306 73 -1272
rect 15 -1340 73 -1306
rect 15 -1374 27 -1340
rect 61 -1374 73 -1340
rect 15 -1408 73 -1374
rect 15 -1442 27 -1408
rect 61 -1442 73 -1408
rect 15 -1476 73 -1442
rect 15 -1510 27 -1476
rect 61 -1510 73 -1476
rect 15 -1544 73 -1510
rect 15 -1578 27 -1544
rect 61 -1578 73 -1544
rect 15 -1612 73 -1578
rect 15 -1646 27 -1612
rect 61 -1646 73 -1612
rect 15 -1680 73 -1646
rect 15 -1714 27 -1680
rect 61 -1714 73 -1680
rect 15 -1748 73 -1714
rect 15 -1782 27 -1748
rect 61 -1782 73 -1748
rect 15 -1816 73 -1782
rect 15 -1850 27 -1816
rect 61 -1850 73 -1816
rect 15 -1884 73 -1850
rect 15 -1918 27 -1884
rect 61 -1918 73 -1884
rect 15 -1952 73 -1918
rect 15 -1986 27 -1952
rect 61 -1986 73 -1952
rect 15 -2031 73 -1986
<< ndiffc >>
rect -61 1890 -27 1924
rect -61 1822 -27 1856
rect -61 1754 -27 1788
rect -61 1686 -27 1720
rect -61 1618 -27 1652
rect -61 1550 -27 1584
rect -61 1482 -27 1516
rect -61 1414 -27 1448
rect -61 1346 -27 1380
rect -61 1278 -27 1312
rect -61 1210 -27 1244
rect -61 1142 -27 1176
rect -61 1074 -27 1108
rect -61 1006 -27 1040
rect -61 938 -27 972
rect -61 870 -27 904
rect -61 802 -27 836
rect -61 734 -27 768
rect -61 666 -27 700
rect -61 598 -27 632
rect -61 530 -27 564
rect -61 462 -27 496
rect -61 394 -27 428
rect -61 326 -27 360
rect -61 258 -27 292
rect -61 190 -27 224
rect -61 122 -27 156
rect -61 54 -27 88
rect -61 -14 -27 20
rect -61 -82 -27 -48
rect -61 -150 -27 -116
rect -61 -218 -27 -184
rect -61 -286 -27 -252
rect -61 -354 -27 -320
rect -61 -422 -27 -388
rect -61 -490 -27 -456
rect -61 -558 -27 -524
rect -61 -626 -27 -592
rect -61 -694 -27 -660
rect -61 -762 -27 -728
rect -61 -830 -27 -796
rect -61 -898 -27 -864
rect -61 -966 -27 -932
rect -61 -1034 -27 -1000
rect -61 -1102 -27 -1068
rect -61 -1170 -27 -1136
rect -61 -1238 -27 -1204
rect -61 -1306 -27 -1272
rect -61 -1374 -27 -1340
rect -61 -1442 -27 -1408
rect -61 -1510 -27 -1476
rect -61 -1578 -27 -1544
rect -61 -1646 -27 -1612
rect -61 -1714 -27 -1680
rect -61 -1782 -27 -1748
rect -61 -1850 -27 -1816
rect -61 -1918 -27 -1884
rect -61 -1986 -27 -1952
rect 27 1890 61 1924
rect 27 1822 61 1856
rect 27 1754 61 1788
rect 27 1686 61 1720
rect 27 1618 61 1652
rect 27 1550 61 1584
rect 27 1482 61 1516
rect 27 1414 61 1448
rect 27 1346 61 1380
rect 27 1278 61 1312
rect 27 1210 61 1244
rect 27 1142 61 1176
rect 27 1074 61 1108
rect 27 1006 61 1040
rect 27 938 61 972
rect 27 870 61 904
rect 27 802 61 836
rect 27 734 61 768
rect 27 666 61 700
rect 27 598 61 632
rect 27 530 61 564
rect 27 462 61 496
rect 27 394 61 428
rect 27 326 61 360
rect 27 258 61 292
rect 27 190 61 224
rect 27 122 61 156
rect 27 54 61 88
rect 27 -14 61 20
rect 27 -82 61 -48
rect 27 -150 61 -116
rect 27 -218 61 -184
rect 27 -286 61 -252
rect 27 -354 61 -320
rect 27 -422 61 -388
rect 27 -490 61 -456
rect 27 -558 61 -524
rect 27 -626 61 -592
rect 27 -694 61 -660
rect 27 -762 61 -728
rect 27 -830 61 -796
rect 27 -898 61 -864
rect 27 -966 61 -932
rect 27 -1034 61 -1000
rect 27 -1102 61 -1068
rect 27 -1170 61 -1136
rect 27 -1238 61 -1204
rect 27 -1306 61 -1272
rect 27 -1374 61 -1340
rect 27 -1442 61 -1408
rect 27 -1510 61 -1476
rect 27 -1578 61 -1544
rect 27 -1646 61 -1612
rect 27 -1714 61 -1680
rect 27 -1782 61 -1748
rect 27 -1850 61 -1816
rect 27 -1918 61 -1884
rect 27 -1986 61 -1952
<< psubdiff >>
rect -175 2109 -51 2143
rect -17 2109 17 2143
rect 51 2109 175 2143
rect -175 2023 -141 2109
rect -175 1955 -141 1989
rect -175 1887 -141 1921
rect -175 1819 -141 1853
rect -175 1751 -141 1785
rect -175 1683 -141 1717
rect -175 1615 -141 1649
rect -175 1547 -141 1581
rect -175 1479 -141 1513
rect -175 1411 -141 1445
rect -175 1343 -141 1377
rect -175 1275 -141 1309
rect -175 1207 -141 1241
rect -175 1139 -141 1173
rect -175 1071 -141 1105
rect -175 1003 -141 1037
rect -175 935 -141 969
rect -175 867 -141 901
rect -175 799 -141 833
rect -175 731 -141 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect -175 -833 -141 -799
rect -175 -901 -141 -867
rect -175 -969 -141 -935
rect -175 -1037 -141 -1003
rect -175 -1105 -141 -1071
rect -175 -1173 -141 -1139
rect -175 -1241 -141 -1207
rect -175 -1309 -141 -1275
rect -175 -1377 -141 -1343
rect -175 -1445 -141 -1411
rect -175 -1513 -141 -1479
rect -175 -1581 -141 -1547
rect -175 -1649 -141 -1615
rect -175 -1717 -141 -1683
rect -175 -1785 -141 -1751
rect -175 -1853 -141 -1819
rect -175 -1921 -141 -1887
rect -175 -1989 -141 -1955
rect -175 -2109 -141 -2023
rect 141 -2109 175 2109
rect -175 -2143 -51 -2109
rect -17 -2143 17 -2109
rect 51 -2143 175 -2109
<< psubdiffcont >>
rect -51 2109 -17 2143
rect 17 2109 51 2143
rect -175 1989 -141 2023
rect -175 1921 -141 1955
rect -175 1853 -141 1887
rect -175 1785 -141 1819
rect -175 1717 -141 1751
rect -175 1649 -141 1683
rect -175 1581 -141 1615
rect -175 1513 -141 1547
rect -175 1445 -141 1479
rect -175 1377 -141 1411
rect -175 1309 -141 1343
rect -175 1241 -141 1275
rect -175 1173 -141 1207
rect -175 1105 -141 1139
rect -175 1037 -141 1071
rect -175 969 -141 1003
rect -175 901 -141 935
rect -175 833 -141 867
rect -175 765 -141 799
rect -175 697 -141 731
rect -175 629 -141 663
rect -175 561 -141 595
rect -175 493 -141 527
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -175 -527 -141 -493
rect -175 -595 -141 -561
rect -175 -663 -141 -629
rect -175 -731 -141 -697
rect -175 -799 -141 -765
rect -175 -867 -141 -833
rect -175 -935 -141 -901
rect -175 -1003 -141 -969
rect -175 -1071 -141 -1037
rect -175 -1139 -141 -1105
rect -175 -1207 -141 -1173
rect -175 -1275 -141 -1241
rect -175 -1343 -141 -1309
rect -175 -1411 -141 -1377
rect -175 -1479 -141 -1445
rect -175 -1547 -141 -1513
rect -175 -1615 -141 -1581
rect -175 -1683 -141 -1649
rect -175 -1751 -141 -1717
rect -175 -1819 -141 -1785
rect -175 -1887 -141 -1853
rect -175 -1955 -141 -1921
rect -175 -2023 -141 -1989
rect -51 -2143 -17 -2109
rect 17 -2143 51 -2109
<< poly >>
rect -33 2041 33 2057
rect -33 2007 -17 2041
rect 17 2007 33 2041
rect -33 1991 33 2007
rect -15 1969 15 1991
rect -15 -2057 15 -2031
<< polycont >>
rect -17 2007 17 2041
<< locali >>
rect -175 2109 -51 2143
rect -17 2109 17 2143
rect 51 2109 175 2143
rect -175 2023 -141 2109
rect -33 2007 -17 2041
rect 17 2007 33 2041
rect -175 1955 -141 1989
rect -175 1887 -141 1921
rect -175 1819 -141 1853
rect -175 1751 -141 1785
rect -175 1683 -141 1717
rect -175 1615 -141 1649
rect -175 1547 -141 1581
rect -175 1479 -141 1513
rect -175 1411 -141 1445
rect -175 1343 -141 1377
rect -175 1275 -141 1309
rect -175 1207 -141 1241
rect -175 1139 -141 1173
rect -175 1071 -141 1105
rect -175 1003 -141 1037
rect -175 935 -141 969
rect -175 867 -141 901
rect -175 799 -141 833
rect -175 731 -141 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect -175 -833 -141 -799
rect -175 -901 -141 -867
rect -175 -969 -141 -935
rect -175 -1037 -141 -1003
rect -175 -1105 -141 -1071
rect -175 -1173 -141 -1139
rect -175 -1241 -141 -1207
rect -175 -1309 -141 -1275
rect -175 -1377 -141 -1343
rect -175 -1445 -141 -1411
rect -175 -1513 -141 -1479
rect -175 -1581 -141 -1547
rect -175 -1649 -141 -1615
rect -175 -1717 -141 -1683
rect -175 -1785 -141 -1751
rect -175 -1853 -141 -1819
rect -175 -1921 -141 -1887
rect -175 -1989 -141 -1955
rect -175 -2109 -141 -2023
rect -61 1930 -27 1973
rect -61 1858 -27 1890
rect -61 1788 -27 1822
rect -61 1720 -27 1752
rect -61 1652 -27 1680
rect -61 1584 -27 1608
rect -61 1516 -27 1536
rect -61 1448 -27 1464
rect -61 1380 -27 1392
rect -61 1312 -27 1320
rect -61 1244 -27 1248
rect -61 1138 -27 1142
rect -61 1066 -27 1074
rect -61 994 -27 1006
rect -61 922 -27 938
rect -61 850 -27 870
rect -61 778 -27 802
rect -61 706 -27 734
rect -61 634 -27 666
rect -61 564 -27 598
rect -61 496 -27 528
rect -61 428 -27 456
rect -61 360 -27 384
rect -61 292 -27 312
rect -61 224 -27 240
rect -61 156 -27 168
rect -61 88 -27 96
rect -61 20 -27 24
rect -61 -86 -27 -82
rect -61 -158 -27 -150
rect -61 -230 -27 -218
rect -61 -302 -27 -286
rect -61 -374 -27 -354
rect -61 -446 -27 -422
rect -61 -518 -27 -490
rect -61 -590 -27 -558
rect -61 -660 -27 -626
rect -61 -728 -27 -696
rect -61 -796 -27 -768
rect -61 -864 -27 -840
rect -61 -932 -27 -912
rect -61 -1000 -27 -984
rect -61 -1068 -27 -1056
rect -61 -1136 -27 -1128
rect -61 -1204 -27 -1200
rect -61 -1310 -27 -1306
rect -61 -1382 -27 -1374
rect -61 -1454 -27 -1442
rect -61 -1526 -27 -1510
rect -61 -1598 -27 -1578
rect -61 -1670 -27 -1646
rect -61 -1742 -27 -1714
rect -61 -1814 -27 -1782
rect -61 -1884 -27 -1850
rect -61 -1952 -27 -1920
rect -61 -2035 -27 -1992
rect 27 1930 61 1973
rect 27 1858 61 1890
rect 27 1788 61 1822
rect 27 1720 61 1752
rect 27 1652 61 1680
rect 27 1584 61 1608
rect 27 1516 61 1536
rect 27 1448 61 1464
rect 27 1380 61 1392
rect 27 1312 61 1320
rect 27 1244 61 1248
rect 27 1138 61 1142
rect 27 1066 61 1074
rect 27 994 61 1006
rect 27 922 61 938
rect 27 850 61 870
rect 27 778 61 802
rect 27 706 61 734
rect 27 634 61 666
rect 27 564 61 598
rect 27 496 61 528
rect 27 428 61 456
rect 27 360 61 384
rect 27 292 61 312
rect 27 224 61 240
rect 27 156 61 168
rect 27 88 61 96
rect 27 20 61 24
rect 27 -86 61 -82
rect 27 -158 61 -150
rect 27 -230 61 -218
rect 27 -302 61 -286
rect 27 -374 61 -354
rect 27 -446 61 -422
rect 27 -518 61 -490
rect 27 -590 61 -558
rect 27 -660 61 -626
rect 27 -728 61 -696
rect 27 -796 61 -768
rect 27 -864 61 -840
rect 27 -932 61 -912
rect 27 -1000 61 -984
rect 27 -1068 61 -1056
rect 27 -1136 61 -1128
rect 27 -1204 61 -1200
rect 27 -1310 61 -1306
rect 27 -1382 61 -1374
rect 27 -1454 61 -1442
rect 27 -1526 61 -1510
rect 27 -1598 61 -1578
rect 27 -1670 61 -1646
rect 27 -1742 61 -1714
rect 27 -1814 61 -1782
rect 27 -1884 61 -1850
rect 27 -1952 61 -1920
rect 27 -2035 61 -1992
rect 141 -2109 175 2109
rect -175 -2143 -51 -2109
rect -17 -2143 17 -2109
rect 51 -2143 175 -2109
<< viali >>
rect -17 2007 17 2041
rect -61 1924 -27 1930
rect -61 1896 -27 1924
rect -61 1856 -27 1858
rect -61 1824 -27 1856
rect -61 1754 -27 1786
rect -61 1752 -27 1754
rect -61 1686 -27 1714
rect -61 1680 -27 1686
rect -61 1618 -27 1642
rect -61 1608 -27 1618
rect -61 1550 -27 1570
rect -61 1536 -27 1550
rect -61 1482 -27 1498
rect -61 1464 -27 1482
rect -61 1414 -27 1426
rect -61 1392 -27 1414
rect -61 1346 -27 1354
rect -61 1320 -27 1346
rect -61 1278 -27 1282
rect -61 1248 -27 1278
rect -61 1176 -27 1210
rect -61 1108 -27 1138
rect -61 1104 -27 1108
rect -61 1040 -27 1066
rect -61 1032 -27 1040
rect -61 972 -27 994
rect -61 960 -27 972
rect -61 904 -27 922
rect -61 888 -27 904
rect -61 836 -27 850
rect -61 816 -27 836
rect -61 768 -27 778
rect -61 744 -27 768
rect -61 700 -27 706
rect -61 672 -27 700
rect -61 632 -27 634
rect -61 600 -27 632
rect -61 530 -27 562
rect -61 528 -27 530
rect -61 462 -27 490
rect -61 456 -27 462
rect -61 394 -27 418
rect -61 384 -27 394
rect -61 326 -27 346
rect -61 312 -27 326
rect -61 258 -27 274
rect -61 240 -27 258
rect -61 190 -27 202
rect -61 168 -27 190
rect -61 122 -27 130
rect -61 96 -27 122
rect -61 54 -27 58
rect -61 24 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -86
rect -61 -120 -27 -116
rect -61 -184 -27 -158
rect -61 -192 -27 -184
rect -61 -252 -27 -230
rect -61 -264 -27 -252
rect -61 -320 -27 -302
rect -61 -336 -27 -320
rect -61 -388 -27 -374
rect -61 -408 -27 -388
rect -61 -456 -27 -446
rect -61 -480 -27 -456
rect -61 -524 -27 -518
rect -61 -552 -27 -524
rect -61 -592 -27 -590
rect -61 -624 -27 -592
rect -61 -694 -27 -662
rect -61 -696 -27 -694
rect -61 -762 -27 -734
rect -61 -768 -27 -762
rect -61 -830 -27 -806
rect -61 -840 -27 -830
rect -61 -898 -27 -878
rect -61 -912 -27 -898
rect -61 -966 -27 -950
rect -61 -984 -27 -966
rect -61 -1034 -27 -1022
rect -61 -1056 -27 -1034
rect -61 -1102 -27 -1094
rect -61 -1128 -27 -1102
rect -61 -1170 -27 -1166
rect -61 -1200 -27 -1170
rect -61 -1272 -27 -1238
rect -61 -1340 -27 -1310
rect -61 -1344 -27 -1340
rect -61 -1408 -27 -1382
rect -61 -1416 -27 -1408
rect -61 -1476 -27 -1454
rect -61 -1488 -27 -1476
rect -61 -1544 -27 -1526
rect -61 -1560 -27 -1544
rect -61 -1612 -27 -1598
rect -61 -1632 -27 -1612
rect -61 -1680 -27 -1670
rect -61 -1704 -27 -1680
rect -61 -1748 -27 -1742
rect -61 -1776 -27 -1748
rect -61 -1816 -27 -1814
rect -61 -1848 -27 -1816
rect -61 -1918 -27 -1886
rect -61 -1920 -27 -1918
rect -61 -1986 -27 -1958
rect -61 -1992 -27 -1986
rect 27 1924 61 1930
rect 27 1896 61 1924
rect 27 1856 61 1858
rect 27 1824 61 1856
rect 27 1754 61 1786
rect 27 1752 61 1754
rect 27 1686 61 1714
rect 27 1680 61 1686
rect 27 1618 61 1642
rect 27 1608 61 1618
rect 27 1550 61 1570
rect 27 1536 61 1550
rect 27 1482 61 1498
rect 27 1464 61 1482
rect 27 1414 61 1426
rect 27 1392 61 1414
rect 27 1346 61 1354
rect 27 1320 61 1346
rect 27 1278 61 1282
rect 27 1248 61 1278
rect 27 1176 61 1210
rect 27 1108 61 1138
rect 27 1104 61 1108
rect 27 1040 61 1066
rect 27 1032 61 1040
rect 27 972 61 994
rect 27 960 61 972
rect 27 904 61 922
rect 27 888 61 904
rect 27 836 61 850
rect 27 816 61 836
rect 27 768 61 778
rect 27 744 61 768
rect 27 700 61 706
rect 27 672 61 700
rect 27 632 61 634
rect 27 600 61 632
rect 27 530 61 562
rect 27 528 61 530
rect 27 462 61 490
rect 27 456 61 462
rect 27 394 61 418
rect 27 384 61 394
rect 27 326 61 346
rect 27 312 61 326
rect 27 258 61 274
rect 27 240 61 258
rect 27 190 61 202
rect 27 168 61 190
rect 27 122 61 130
rect 27 96 61 122
rect 27 54 61 58
rect 27 24 61 54
rect 27 -48 61 -14
rect 27 -116 61 -86
rect 27 -120 61 -116
rect 27 -184 61 -158
rect 27 -192 61 -184
rect 27 -252 61 -230
rect 27 -264 61 -252
rect 27 -320 61 -302
rect 27 -336 61 -320
rect 27 -388 61 -374
rect 27 -408 61 -388
rect 27 -456 61 -446
rect 27 -480 61 -456
rect 27 -524 61 -518
rect 27 -552 61 -524
rect 27 -592 61 -590
rect 27 -624 61 -592
rect 27 -694 61 -662
rect 27 -696 61 -694
rect 27 -762 61 -734
rect 27 -768 61 -762
rect 27 -830 61 -806
rect 27 -840 61 -830
rect 27 -898 61 -878
rect 27 -912 61 -898
rect 27 -966 61 -950
rect 27 -984 61 -966
rect 27 -1034 61 -1022
rect 27 -1056 61 -1034
rect 27 -1102 61 -1094
rect 27 -1128 61 -1102
rect 27 -1170 61 -1166
rect 27 -1200 61 -1170
rect 27 -1272 61 -1238
rect 27 -1340 61 -1310
rect 27 -1344 61 -1340
rect 27 -1408 61 -1382
rect 27 -1416 61 -1408
rect 27 -1476 61 -1454
rect 27 -1488 61 -1476
rect 27 -1544 61 -1526
rect 27 -1560 61 -1544
rect 27 -1612 61 -1598
rect 27 -1632 61 -1612
rect 27 -1680 61 -1670
rect 27 -1704 61 -1680
rect 27 -1748 61 -1742
rect 27 -1776 61 -1748
rect 27 -1816 61 -1814
rect 27 -1848 61 -1816
rect 27 -1918 61 -1886
rect 27 -1920 61 -1918
rect 27 -1986 61 -1958
rect 27 -1992 61 -1986
<< metal1 >>
rect -29 2041 29 2047
rect -29 2007 -17 2041
rect 17 2007 29 2041
rect -29 2001 29 2007
rect -67 1930 -21 1969
rect -67 1896 -61 1930
rect -27 1896 -21 1930
rect -67 1858 -21 1896
rect -67 1824 -61 1858
rect -27 1824 -21 1858
rect -67 1786 -21 1824
rect -67 1752 -61 1786
rect -27 1752 -21 1786
rect -67 1714 -21 1752
rect -67 1680 -61 1714
rect -27 1680 -21 1714
rect -67 1642 -21 1680
rect -67 1608 -61 1642
rect -27 1608 -21 1642
rect -67 1570 -21 1608
rect -67 1536 -61 1570
rect -27 1536 -21 1570
rect -67 1498 -21 1536
rect -67 1464 -61 1498
rect -27 1464 -21 1498
rect -67 1426 -21 1464
rect -67 1392 -61 1426
rect -27 1392 -21 1426
rect -67 1354 -21 1392
rect -67 1320 -61 1354
rect -27 1320 -21 1354
rect -67 1282 -21 1320
rect -67 1248 -61 1282
rect -27 1248 -21 1282
rect -67 1210 -21 1248
rect -67 1176 -61 1210
rect -27 1176 -21 1210
rect -67 1138 -21 1176
rect -67 1104 -61 1138
rect -27 1104 -21 1138
rect -67 1066 -21 1104
rect -67 1032 -61 1066
rect -27 1032 -21 1066
rect -67 994 -21 1032
rect -67 960 -61 994
rect -27 960 -21 994
rect -67 922 -21 960
rect -67 888 -61 922
rect -27 888 -21 922
rect -67 850 -21 888
rect -67 816 -61 850
rect -27 816 -21 850
rect -67 778 -21 816
rect -67 744 -61 778
rect -27 744 -21 778
rect -67 706 -21 744
rect -67 672 -61 706
rect -27 672 -21 706
rect -67 634 -21 672
rect -67 600 -61 634
rect -27 600 -21 634
rect -67 562 -21 600
rect -67 528 -61 562
rect -27 528 -21 562
rect -67 490 -21 528
rect -67 456 -61 490
rect -27 456 -21 490
rect -67 418 -21 456
rect -67 384 -61 418
rect -27 384 -21 418
rect -67 346 -21 384
rect -67 312 -61 346
rect -27 312 -21 346
rect -67 274 -21 312
rect -67 240 -61 274
rect -27 240 -21 274
rect -67 202 -21 240
rect -67 168 -61 202
rect -27 168 -21 202
rect -67 130 -21 168
rect -67 96 -61 130
rect -27 96 -21 130
rect -67 58 -21 96
rect -67 24 -61 58
rect -27 24 -21 58
rect -67 -14 -21 24
rect -67 -48 -61 -14
rect -27 -48 -21 -14
rect -67 -86 -21 -48
rect -67 -120 -61 -86
rect -27 -120 -21 -86
rect -67 -158 -21 -120
rect -67 -192 -61 -158
rect -27 -192 -21 -158
rect -67 -230 -21 -192
rect -67 -264 -61 -230
rect -27 -264 -21 -230
rect -67 -302 -21 -264
rect -67 -336 -61 -302
rect -27 -336 -21 -302
rect -67 -374 -21 -336
rect -67 -408 -61 -374
rect -27 -408 -21 -374
rect -67 -446 -21 -408
rect -67 -480 -61 -446
rect -27 -480 -21 -446
rect -67 -518 -21 -480
rect -67 -552 -61 -518
rect -27 -552 -21 -518
rect -67 -590 -21 -552
rect -67 -624 -61 -590
rect -27 -624 -21 -590
rect -67 -662 -21 -624
rect -67 -696 -61 -662
rect -27 -696 -21 -662
rect -67 -734 -21 -696
rect -67 -768 -61 -734
rect -27 -768 -21 -734
rect -67 -806 -21 -768
rect -67 -840 -61 -806
rect -27 -840 -21 -806
rect -67 -878 -21 -840
rect -67 -912 -61 -878
rect -27 -912 -21 -878
rect -67 -950 -21 -912
rect -67 -984 -61 -950
rect -27 -984 -21 -950
rect -67 -1022 -21 -984
rect -67 -1056 -61 -1022
rect -27 -1056 -21 -1022
rect -67 -1094 -21 -1056
rect -67 -1128 -61 -1094
rect -27 -1128 -21 -1094
rect -67 -1166 -21 -1128
rect -67 -1200 -61 -1166
rect -27 -1200 -21 -1166
rect -67 -1238 -21 -1200
rect -67 -1272 -61 -1238
rect -27 -1272 -21 -1238
rect -67 -1310 -21 -1272
rect -67 -1344 -61 -1310
rect -27 -1344 -21 -1310
rect -67 -1382 -21 -1344
rect -67 -1416 -61 -1382
rect -27 -1416 -21 -1382
rect -67 -1454 -21 -1416
rect -67 -1488 -61 -1454
rect -27 -1488 -21 -1454
rect -67 -1526 -21 -1488
rect -67 -1560 -61 -1526
rect -27 -1560 -21 -1526
rect -67 -1598 -21 -1560
rect -67 -1632 -61 -1598
rect -27 -1632 -21 -1598
rect -67 -1670 -21 -1632
rect -67 -1704 -61 -1670
rect -27 -1704 -21 -1670
rect -67 -1742 -21 -1704
rect -67 -1776 -61 -1742
rect -27 -1776 -21 -1742
rect -67 -1814 -21 -1776
rect -67 -1848 -61 -1814
rect -27 -1848 -21 -1814
rect -67 -1886 -21 -1848
rect -67 -1920 -61 -1886
rect -27 -1920 -21 -1886
rect -67 -1958 -21 -1920
rect -67 -1992 -61 -1958
rect -27 -1992 -21 -1958
rect -67 -2031 -21 -1992
rect 21 1930 67 1969
rect 21 1896 27 1930
rect 61 1896 67 1930
rect 21 1858 67 1896
rect 21 1824 27 1858
rect 61 1824 67 1858
rect 21 1786 67 1824
rect 21 1752 27 1786
rect 61 1752 67 1786
rect 21 1714 67 1752
rect 21 1680 27 1714
rect 61 1680 67 1714
rect 21 1642 67 1680
rect 21 1608 27 1642
rect 61 1608 67 1642
rect 21 1570 67 1608
rect 21 1536 27 1570
rect 61 1536 67 1570
rect 21 1498 67 1536
rect 21 1464 27 1498
rect 61 1464 67 1498
rect 21 1426 67 1464
rect 21 1392 27 1426
rect 61 1392 67 1426
rect 21 1354 67 1392
rect 21 1320 27 1354
rect 61 1320 67 1354
rect 21 1282 67 1320
rect 21 1248 27 1282
rect 61 1248 67 1282
rect 21 1210 67 1248
rect 21 1176 27 1210
rect 61 1176 67 1210
rect 21 1138 67 1176
rect 21 1104 27 1138
rect 61 1104 67 1138
rect 21 1066 67 1104
rect 21 1032 27 1066
rect 61 1032 67 1066
rect 21 994 67 1032
rect 21 960 27 994
rect 61 960 67 994
rect 21 922 67 960
rect 21 888 27 922
rect 61 888 67 922
rect 21 850 67 888
rect 21 816 27 850
rect 61 816 67 850
rect 21 778 67 816
rect 21 744 27 778
rect 61 744 67 778
rect 21 706 67 744
rect 21 672 27 706
rect 61 672 67 706
rect 21 634 67 672
rect 21 600 27 634
rect 61 600 67 634
rect 21 562 67 600
rect 21 528 27 562
rect 61 528 67 562
rect 21 490 67 528
rect 21 456 27 490
rect 61 456 67 490
rect 21 418 67 456
rect 21 384 27 418
rect 61 384 67 418
rect 21 346 67 384
rect 21 312 27 346
rect 61 312 67 346
rect 21 274 67 312
rect 21 240 27 274
rect 61 240 67 274
rect 21 202 67 240
rect 21 168 27 202
rect 61 168 67 202
rect 21 130 67 168
rect 21 96 27 130
rect 61 96 67 130
rect 21 58 67 96
rect 21 24 27 58
rect 61 24 67 58
rect 21 -14 67 24
rect 21 -48 27 -14
rect 61 -48 67 -14
rect 21 -86 67 -48
rect 21 -120 27 -86
rect 61 -120 67 -86
rect 21 -158 67 -120
rect 21 -192 27 -158
rect 61 -192 67 -158
rect 21 -230 67 -192
rect 21 -264 27 -230
rect 61 -264 67 -230
rect 21 -302 67 -264
rect 21 -336 27 -302
rect 61 -336 67 -302
rect 21 -374 67 -336
rect 21 -408 27 -374
rect 61 -408 67 -374
rect 21 -446 67 -408
rect 21 -480 27 -446
rect 61 -480 67 -446
rect 21 -518 67 -480
rect 21 -552 27 -518
rect 61 -552 67 -518
rect 21 -590 67 -552
rect 21 -624 27 -590
rect 61 -624 67 -590
rect 21 -662 67 -624
rect 21 -696 27 -662
rect 61 -696 67 -662
rect 21 -734 67 -696
rect 21 -768 27 -734
rect 61 -768 67 -734
rect 21 -806 67 -768
rect 21 -840 27 -806
rect 61 -840 67 -806
rect 21 -878 67 -840
rect 21 -912 27 -878
rect 61 -912 67 -878
rect 21 -950 67 -912
rect 21 -984 27 -950
rect 61 -984 67 -950
rect 21 -1022 67 -984
rect 21 -1056 27 -1022
rect 61 -1056 67 -1022
rect 21 -1094 67 -1056
rect 21 -1128 27 -1094
rect 61 -1128 67 -1094
rect 21 -1166 67 -1128
rect 21 -1200 27 -1166
rect 61 -1200 67 -1166
rect 21 -1238 67 -1200
rect 21 -1272 27 -1238
rect 61 -1272 67 -1238
rect 21 -1310 67 -1272
rect 21 -1344 27 -1310
rect 61 -1344 67 -1310
rect 21 -1382 67 -1344
rect 21 -1416 27 -1382
rect 61 -1416 67 -1382
rect 21 -1454 67 -1416
rect 21 -1488 27 -1454
rect 61 -1488 67 -1454
rect 21 -1526 67 -1488
rect 21 -1560 27 -1526
rect 61 -1560 67 -1526
rect 21 -1598 67 -1560
rect 21 -1632 27 -1598
rect 61 -1632 67 -1598
rect 21 -1670 67 -1632
rect 21 -1704 27 -1670
rect 61 -1704 67 -1670
rect 21 -1742 67 -1704
rect 21 -1776 27 -1742
rect 61 -1776 67 -1742
rect 21 -1814 67 -1776
rect 21 -1848 27 -1814
rect 61 -1848 67 -1814
rect 21 -1886 67 -1848
rect 21 -1920 27 -1886
rect 61 -1920 67 -1886
rect 21 -1958 67 -1920
rect 21 -1992 27 -1958
rect 61 -1992 67 -1958
rect 21 -2031 67 -1992
<< properties >>
string FIXED_BBOX -158 -2126 158 2126
<< end >>
