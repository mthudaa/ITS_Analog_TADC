magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< pwell >>
rect -211 -198 211 198
<< nmos >>
rect -15 -50 15 50
<< ndiff >>
rect -73 38 -15 50
rect -73 -38 -61 38
rect -27 -38 -15 38
rect -73 -50 -15 -38
rect 15 38 73 50
rect 15 -38 27 38
rect 61 -38 73 38
rect 15 -50 73 -38
<< ndiffc >>
rect -61 -38 -27 38
rect 27 -38 61 38
<< psubdiff >>
rect -175 128 -79 162
rect 79 128 175 162
rect -175 66 -141 128
rect 141 66 175 128
rect -175 -128 -141 -66
rect 141 -128 175 -66
rect -175 -162 -79 -128
rect 79 -162 175 -128
<< psubdiffcont >>
rect -79 128 79 162
rect -175 -66 -141 66
rect 141 -66 175 66
rect -79 -162 79 -128
<< poly >>
rect -15 50 15 76
rect -15 -76 15 -50
<< locali >>
rect -175 128 -79 162
rect 79 128 175 162
rect -175 66 -141 128
rect 141 66 175 128
rect -61 38 -27 54
rect -61 -54 -27 -38
rect 27 38 61 54
rect 27 -54 61 -38
rect -175 -128 -141 -66
rect 141 -128 175 -66
rect -175 -162 -79 -128
rect 79 -162 175 -128
<< viali >>
rect -61 -38 -27 38
rect 27 -38 61 38
<< metal1 >>
rect -67 38 -21 50
rect -67 -38 -61 38
rect -27 -38 -21 38
rect -67 -50 -21 -38
rect 21 38 67 50
rect 21 -38 27 38
rect 61 -38 67 38
rect 21 -50 67 -38
<< properties >>
string FIXED_BBOX -158 -145 158 145
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
