magic
tech sky130A
magscale 1 2
timestamp 1757893939
<< metal1 >>
rect -224 2974 5424 2996
rect -224 2922 -192 2974
rect -140 2922 5340 2974
rect 5392 2922 5424 2974
rect -224 2900 5424 2922
rect -32 2782 5232 2804
rect -32 2730 0 2782
rect 52 2730 2329 2782
rect 2381 2730 5148 2782
rect 5200 2730 5232 2782
rect -32 2708 5232 2730
rect 2195 2590 2414 2612
rect 2195 2538 2329 2590
rect 2381 2538 2414 2590
rect 2195 2516 2414 2538
rect 368 2423 378 2475
rect 430 2466 440 2475
rect 430 2432 609 2466
rect 430 2423 440 2432
rect 2296 2376 2414 2399
rect 2296 2324 2329 2376
rect 2381 2324 2414 2376
rect 2296 2301 2414 2324
rect 2095 1888 2410 1940
rect 160 1379 170 1388
rect -214 1345 170 1379
rect 160 1336 170 1345
rect 222 1379 232 1388
rect 222 1345 613 1379
rect 222 1336 232 1345
rect 264 1305 274 1314
rect -214 1271 274 1305
rect 264 1262 274 1271
rect 326 1305 336 1314
rect 326 1271 636 1305
rect 326 1262 336 1271
rect -224 1206 496 1228
rect -224 1154 -192 1206
rect -140 1154 496 1206
rect -224 1132 496 1154
rect 2210 1132 2306 1228
rect 4990 1206 5424 1228
rect 4990 1154 5340 1206
rect 5392 1154 5424 1206
rect 4990 1132 5424 1154
rect 368 1089 378 1098
rect -214 1055 378 1089
rect 368 1046 378 1055
rect 430 1089 440 1098
rect 430 1055 671 1089
rect 430 1046 440 1055
rect 160 972 170 1024
rect 222 1015 232 1024
rect 222 981 624 1015
rect 222 972 232 981
rect 4983 888 5414 928
rect 4984 676 5414 716
rect 4990 597 5414 637
rect 2095 406 2519 458
rect 2296 36 2414 59
rect 2296 -16 2329 36
rect 2381 -16 2414 36
rect 2296 -39 2414 -16
rect 264 -115 274 -63
rect 326 -72 336 -63
rect 326 -106 637 -72
rect 326 -115 336 -106
rect 2204 -178 2414 -156
rect 2204 -230 2329 -178
rect 2381 -230 2414 -178
rect 2204 -252 2414 -230
rect -32 -370 5232 -348
rect -32 -422 0 -370
rect 52 -422 2329 -370
rect 2381 -422 3574 -370
rect 3626 -422 5148 -370
rect 5200 -422 5232 -370
rect -32 -444 5232 -422
rect -224 -562 5424 -540
rect -224 -614 -192 -562
rect -140 -614 5340 -562
rect 5392 -614 5424 -562
rect -224 -636 5424 -614
<< via1 >>
rect -192 2922 -140 2974
rect 5340 2922 5392 2974
rect 0 2730 52 2782
rect 2329 2730 2381 2782
rect 5148 2730 5200 2782
rect 2329 2538 2381 2590
rect 378 2423 430 2475
rect 2329 2324 2381 2376
rect 170 1336 222 1388
rect 274 1262 326 1314
rect -192 1154 -140 1206
rect 5340 1154 5392 1206
rect 378 1046 430 1098
rect 170 972 222 1024
rect 2329 -16 2381 36
rect 274 -115 326 -63
rect 2329 -230 2381 -178
rect 0 -422 52 -370
rect 2329 -422 2381 -370
rect 3574 -422 3626 -370
rect 5148 -422 5200 -370
rect -192 -614 -140 -562
rect 5340 -614 5392 -562
<< metal2 >>
rect -214 2974 -118 3006
rect -214 2922 -192 2974
rect -140 2922 -118 2974
rect -214 1206 -118 2922
rect 5318 2974 5414 3006
rect 5318 2922 5340 2974
rect 5392 2922 5414 2974
rect -214 1154 -192 1206
rect -140 1154 -118 1206
rect -214 -562 -118 1154
rect -22 2782 74 2814
rect -22 2730 0 2782
rect 52 2730 74 2782
rect -22 -370 74 2730
rect 2306 2782 2404 2814
rect 2306 2730 2329 2782
rect 2381 2730 2404 2782
rect 2306 2590 2404 2730
rect 2306 2538 2329 2590
rect 2381 2538 2404 2590
rect 378 2475 430 2485
rect 170 1388 222 1398
rect 170 1024 222 1336
rect 170 962 222 972
rect 274 1314 326 1324
rect 274 -63 326 1262
rect 378 1098 430 2423
rect 2306 2376 2404 2538
rect 2306 2324 2329 2376
rect 2381 2324 2404 2376
rect 2306 2291 2404 2324
rect 5126 2782 5222 2814
rect 5126 2730 5148 2782
rect 5200 2730 5222 2782
rect 378 1036 430 1046
rect 274 -125 326 -115
rect 2306 36 2404 69
rect 2306 -16 2329 36
rect 2381 -16 2404 36
rect -22 -422 0 -370
rect 52 -422 74 -370
rect -22 -454 74 -422
rect 2306 -178 2404 -16
rect 2306 -230 2329 -178
rect 2381 -230 2404 -178
rect 2306 -370 2404 -230
rect 2306 -422 2329 -370
rect 2381 -422 2404 -370
rect 2306 -454 2404 -422
rect 3552 -370 3648 210
rect 3552 -422 3574 -370
rect 3626 -422 3648 -370
rect 3552 -454 3648 -422
rect 5126 -370 5222 2730
rect 5126 -422 5148 -370
rect 5200 -422 5222 -370
rect 5126 -454 5222 -422
rect 5318 1206 5414 2922
rect 5318 1154 5340 1206
rect 5392 1154 5414 1206
rect -214 -614 -192 -562
rect -140 -614 -118 -562
rect -214 -646 -118 -614
rect 5318 -562 5414 1154
rect 5318 -614 5340 -562
rect 5392 -614 5414 -562
rect 5318 -646 5414 -614
use delay_gate_ori  delay_gate_ori_0
timestamp 1757893504
transform 1 0 1371 0 -1 2130
box -875 -482 853 998
use delay_gate_ori  delay_gate_ori_1
timestamp 1757893504
transform 1 0 1371 0 1 230
box -875 -482 853 998
use phase_detector  phase_detector_0
timestamp 1757893939
transform 1 0 2324 0 1 -47
box -28 -2 2706 2456
<< labels >>
flabel metal1 s 412 2934 442 2964 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 392 2748 422 2778 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -93 1271 -59 1305 0 FreeSans 500 0 0 0 VINP
port 3 nsew
flabel metal1 s -92 1055 -58 1089 0 FreeSans 500 0 0 0 VINN
port 4 nsew
flabel metal1 s 5245 888 5285 928 0 FreeSans 500 0 0 0 RDY
port 5 nsew
flabel metal1 s 5253 676 5293 716 0 FreeSans 500 0 0 0 OUTP
port 6 nsew
flabel metal1 s 5249 597 5289 637 0 FreeSans 500 0 0 0 OUTN
port 7 nsew
flabel metal1 s -103 1345 -69 1379 0 FreeSans 500 0 0 0 CLK
port 8 nsew
<< end >>
