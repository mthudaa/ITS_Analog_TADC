magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -246 -1867 246 1867
<< pmos >>
rect -50 1348 50 1648
rect -50 920 50 1220
rect -50 492 50 792
rect -50 64 50 364
rect -50 -364 50 -64
rect -50 -792 50 -492
rect -50 -1220 50 -920
rect -50 -1648 50 -1348
<< pdiff >>
rect -108 1617 -50 1648
rect -108 1583 -96 1617
rect -62 1583 -50 1617
rect -108 1549 -50 1583
rect -108 1515 -96 1549
rect -62 1515 -50 1549
rect -108 1481 -50 1515
rect -108 1447 -96 1481
rect -62 1447 -50 1481
rect -108 1413 -50 1447
rect -108 1379 -96 1413
rect -62 1379 -50 1413
rect -108 1348 -50 1379
rect 50 1617 108 1648
rect 50 1583 62 1617
rect 96 1583 108 1617
rect 50 1549 108 1583
rect 50 1515 62 1549
rect 96 1515 108 1549
rect 50 1481 108 1515
rect 50 1447 62 1481
rect 96 1447 108 1481
rect 50 1413 108 1447
rect 50 1379 62 1413
rect 96 1379 108 1413
rect 50 1348 108 1379
rect -108 1189 -50 1220
rect -108 1155 -96 1189
rect -62 1155 -50 1189
rect -108 1121 -50 1155
rect -108 1087 -96 1121
rect -62 1087 -50 1121
rect -108 1053 -50 1087
rect -108 1019 -96 1053
rect -62 1019 -50 1053
rect -108 985 -50 1019
rect -108 951 -96 985
rect -62 951 -50 985
rect -108 920 -50 951
rect 50 1189 108 1220
rect 50 1155 62 1189
rect 96 1155 108 1189
rect 50 1121 108 1155
rect 50 1087 62 1121
rect 96 1087 108 1121
rect 50 1053 108 1087
rect 50 1019 62 1053
rect 96 1019 108 1053
rect 50 985 108 1019
rect 50 951 62 985
rect 96 951 108 985
rect 50 920 108 951
rect -108 761 -50 792
rect -108 727 -96 761
rect -62 727 -50 761
rect -108 693 -50 727
rect -108 659 -96 693
rect -62 659 -50 693
rect -108 625 -50 659
rect -108 591 -96 625
rect -62 591 -50 625
rect -108 557 -50 591
rect -108 523 -96 557
rect -62 523 -50 557
rect -108 492 -50 523
rect 50 761 108 792
rect 50 727 62 761
rect 96 727 108 761
rect 50 693 108 727
rect 50 659 62 693
rect 96 659 108 693
rect 50 625 108 659
rect 50 591 62 625
rect 96 591 108 625
rect 50 557 108 591
rect 50 523 62 557
rect 96 523 108 557
rect 50 492 108 523
rect -108 333 -50 364
rect -108 299 -96 333
rect -62 299 -50 333
rect -108 265 -50 299
rect -108 231 -96 265
rect -62 231 -50 265
rect -108 197 -50 231
rect -108 163 -96 197
rect -62 163 -50 197
rect -108 129 -50 163
rect -108 95 -96 129
rect -62 95 -50 129
rect -108 64 -50 95
rect 50 333 108 364
rect 50 299 62 333
rect 96 299 108 333
rect 50 265 108 299
rect 50 231 62 265
rect 96 231 108 265
rect 50 197 108 231
rect 50 163 62 197
rect 96 163 108 197
rect 50 129 108 163
rect 50 95 62 129
rect 96 95 108 129
rect 50 64 108 95
rect -108 -95 -50 -64
rect -108 -129 -96 -95
rect -62 -129 -50 -95
rect -108 -163 -50 -129
rect -108 -197 -96 -163
rect -62 -197 -50 -163
rect -108 -231 -50 -197
rect -108 -265 -96 -231
rect -62 -265 -50 -231
rect -108 -299 -50 -265
rect -108 -333 -96 -299
rect -62 -333 -50 -299
rect -108 -364 -50 -333
rect 50 -95 108 -64
rect 50 -129 62 -95
rect 96 -129 108 -95
rect 50 -163 108 -129
rect 50 -197 62 -163
rect 96 -197 108 -163
rect 50 -231 108 -197
rect 50 -265 62 -231
rect 96 -265 108 -231
rect 50 -299 108 -265
rect 50 -333 62 -299
rect 96 -333 108 -299
rect 50 -364 108 -333
rect -108 -523 -50 -492
rect -108 -557 -96 -523
rect -62 -557 -50 -523
rect -108 -591 -50 -557
rect -108 -625 -96 -591
rect -62 -625 -50 -591
rect -108 -659 -50 -625
rect -108 -693 -96 -659
rect -62 -693 -50 -659
rect -108 -727 -50 -693
rect -108 -761 -96 -727
rect -62 -761 -50 -727
rect -108 -792 -50 -761
rect 50 -523 108 -492
rect 50 -557 62 -523
rect 96 -557 108 -523
rect 50 -591 108 -557
rect 50 -625 62 -591
rect 96 -625 108 -591
rect 50 -659 108 -625
rect 50 -693 62 -659
rect 96 -693 108 -659
rect 50 -727 108 -693
rect 50 -761 62 -727
rect 96 -761 108 -727
rect 50 -792 108 -761
rect -108 -951 -50 -920
rect -108 -985 -96 -951
rect -62 -985 -50 -951
rect -108 -1019 -50 -985
rect -108 -1053 -96 -1019
rect -62 -1053 -50 -1019
rect -108 -1087 -50 -1053
rect -108 -1121 -96 -1087
rect -62 -1121 -50 -1087
rect -108 -1155 -50 -1121
rect -108 -1189 -96 -1155
rect -62 -1189 -50 -1155
rect -108 -1220 -50 -1189
rect 50 -951 108 -920
rect 50 -985 62 -951
rect 96 -985 108 -951
rect 50 -1019 108 -985
rect 50 -1053 62 -1019
rect 96 -1053 108 -1019
rect 50 -1087 108 -1053
rect 50 -1121 62 -1087
rect 96 -1121 108 -1087
rect 50 -1155 108 -1121
rect 50 -1189 62 -1155
rect 96 -1189 108 -1155
rect 50 -1220 108 -1189
rect -108 -1379 -50 -1348
rect -108 -1413 -96 -1379
rect -62 -1413 -50 -1379
rect -108 -1447 -50 -1413
rect -108 -1481 -96 -1447
rect -62 -1481 -50 -1447
rect -108 -1515 -50 -1481
rect -108 -1549 -96 -1515
rect -62 -1549 -50 -1515
rect -108 -1583 -50 -1549
rect -108 -1617 -96 -1583
rect -62 -1617 -50 -1583
rect -108 -1648 -50 -1617
rect 50 -1379 108 -1348
rect 50 -1413 62 -1379
rect 96 -1413 108 -1379
rect 50 -1447 108 -1413
rect 50 -1481 62 -1447
rect 96 -1481 108 -1447
rect 50 -1515 108 -1481
rect 50 -1549 62 -1515
rect 96 -1549 108 -1515
rect 50 -1583 108 -1549
rect 50 -1617 62 -1583
rect 96 -1617 108 -1583
rect 50 -1648 108 -1617
<< pdiffc >>
rect -96 1583 -62 1617
rect -96 1515 -62 1549
rect -96 1447 -62 1481
rect -96 1379 -62 1413
rect 62 1583 96 1617
rect 62 1515 96 1549
rect 62 1447 96 1481
rect 62 1379 96 1413
rect -96 1155 -62 1189
rect -96 1087 -62 1121
rect -96 1019 -62 1053
rect -96 951 -62 985
rect 62 1155 96 1189
rect 62 1087 96 1121
rect 62 1019 96 1053
rect 62 951 96 985
rect -96 727 -62 761
rect -96 659 -62 693
rect -96 591 -62 625
rect -96 523 -62 557
rect 62 727 96 761
rect 62 659 96 693
rect 62 591 96 625
rect 62 523 96 557
rect -96 299 -62 333
rect -96 231 -62 265
rect -96 163 -62 197
rect -96 95 -62 129
rect 62 299 96 333
rect 62 231 96 265
rect 62 163 96 197
rect 62 95 96 129
rect -96 -129 -62 -95
rect -96 -197 -62 -163
rect -96 -265 -62 -231
rect -96 -333 -62 -299
rect 62 -129 96 -95
rect 62 -197 96 -163
rect 62 -265 96 -231
rect 62 -333 96 -299
rect -96 -557 -62 -523
rect -96 -625 -62 -591
rect -96 -693 -62 -659
rect -96 -761 -62 -727
rect 62 -557 96 -523
rect 62 -625 96 -591
rect 62 -693 96 -659
rect 62 -761 96 -727
rect -96 -985 -62 -951
rect -96 -1053 -62 -1019
rect -96 -1121 -62 -1087
rect -96 -1189 -62 -1155
rect 62 -985 96 -951
rect 62 -1053 96 -1019
rect 62 -1121 96 -1087
rect 62 -1189 96 -1155
rect -96 -1413 -62 -1379
rect -96 -1481 -62 -1447
rect -96 -1549 -62 -1515
rect -96 -1617 -62 -1583
rect 62 -1413 96 -1379
rect 62 -1481 96 -1447
rect 62 -1549 96 -1515
rect 62 -1617 96 -1583
<< nsubdiff >>
rect -210 1797 -85 1831
rect -51 1797 -17 1831
rect 17 1797 51 1831
rect 85 1797 210 1831
rect -210 1717 -176 1797
rect -210 1649 -176 1683
rect 176 1717 210 1797
rect 176 1649 210 1683
rect -210 1581 -176 1615
rect -210 1513 -176 1547
rect -210 1445 -176 1479
rect -210 1377 -176 1411
rect 176 1581 210 1615
rect 176 1513 210 1547
rect 176 1445 210 1479
rect 176 1377 210 1411
rect -210 1309 -176 1343
rect -210 1241 -176 1275
rect 176 1309 210 1343
rect 176 1241 210 1275
rect -210 1173 -176 1207
rect -210 1105 -176 1139
rect -210 1037 -176 1071
rect -210 969 -176 1003
rect -210 901 -176 935
rect 176 1173 210 1207
rect 176 1105 210 1139
rect 176 1037 210 1071
rect 176 969 210 1003
rect -210 833 -176 867
rect -210 765 -176 799
rect 176 901 210 935
rect 176 833 210 867
rect -210 697 -176 731
rect -210 629 -176 663
rect -210 561 -176 595
rect -210 493 -176 527
rect 176 765 210 799
rect 176 697 210 731
rect 176 629 210 663
rect 176 561 210 595
rect 176 493 210 527
rect -210 425 -176 459
rect -210 357 -176 391
rect 176 425 210 459
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect -210 -459 -176 -425
rect 176 -391 210 -357
rect 176 -459 210 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -210 -663 -176 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect 176 -527 210 -493
rect 176 -595 210 -561
rect 176 -663 210 -629
rect 176 -731 210 -697
rect -210 -867 -176 -833
rect -210 -935 -176 -901
rect 176 -799 210 -765
rect 176 -867 210 -833
rect -210 -1003 -176 -969
rect -210 -1071 -176 -1037
rect -210 -1139 -176 -1105
rect -210 -1207 -176 -1173
rect 176 -935 210 -901
rect 176 -1003 210 -969
rect 176 -1071 210 -1037
rect 176 -1139 210 -1105
rect 176 -1207 210 -1173
rect -210 -1275 -176 -1241
rect -210 -1343 -176 -1309
rect 176 -1275 210 -1241
rect 176 -1343 210 -1309
rect -210 -1411 -176 -1377
rect -210 -1479 -176 -1445
rect -210 -1547 -176 -1513
rect -210 -1615 -176 -1581
rect 176 -1411 210 -1377
rect 176 -1479 210 -1445
rect 176 -1547 210 -1513
rect 176 -1615 210 -1581
rect -210 -1683 -176 -1649
rect -210 -1797 -176 -1717
rect 176 -1683 210 -1649
rect 176 -1797 210 -1717
rect -210 -1831 -85 -1797
rect -51 -1831 -17 -1797
rect 17 -1831 51 -1797
rect 85 -1831 210 -1797
<< nsubdiffcont >>
rect -85 1797 -51 1831
rect -17 1797 17 1831
rect 51 1797 85 1831
rect -210 1683 -176 1717
rect -210 1615 -176 1649
rect 176 1683 210 1717
rect -210 1547 -176 1581
rect -210 1479 -176 1513
rect -210 1411 -176 1445
rect -210 1343 -176 1377
rect 176 1615 210 1649
rect 176 1547 210 1581
rect 176 1479 210 1513
rect 176 1411 210 1445
rect -210 1275 -176 1309
rect -210 1207 -176 1241
rect 176 1343 210 1377
rect 176 1275 210 1309
rect -210 1139 -176 1173
rect -210 1071 -176 1105
rect -210 1003 -176 1037
rect -210 935 -176 969
rect 176 1207 210 1241
rect 176 1139 210 1173
rect 176 1071 210 1105
rect 176 1003 210 1037
rect 176 935 210 969
rect -210 867 -176 901
rect -210 799 -176 833
rect 176 867 210 901
rect 176 799 210 833
rect -210 731 -176 765
rect -210 663 -176 697
rect -210 595 -176 629
rect -210 527 -176 561
rect -210 459 -176 493
rect 176 731 210 765
rect 176 663 210 697
rect 176 595 210 629
rect 176 527 210 561
rect -210 391 -176 425
rect 176 459 210 493
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect -210 -493 -176 -459
rect 176 -425 210 -391
rect -210 -561 -176 -527
rect -210 -629 -176 -595
rect -210 -697 -176 -663
rect -210 -765 -176 -731
rect 176 -493 210 -459
rect 176 -561 210 -527
rect 176 -629 210 -595
rect 176 -697 210 -663
rect 176 -765 210 -731
rect -210 -833 -176 -799
rect -210 -901 -176 -867
rect 176 -833 210 -799
rect 176 -901 210 -867
rect -210 -969 -176 -935
rect -210 -1037 -176 -1003
rect -210 -1105 -176 -1071
rect -210 -1173 -176 -1139
rect -210 -1241 -176 -1207
rect 176 -969 210 -935
rect 176 -1037 210 -1003
rect 176 -1105 210 -1071
rect 176 -1173 210 -1139
rect -210 -1309 -176 -1275
rect -210 -1377 -176 -1343
rect 176 -1241 210 -1207
rect 176 -1309 210 -1275
rect -210 -1445 -176 -1411
rect -210 -1513 -176 -1479
rect -210 -1581 -176 -1547
rect -210 -1649 -176 -1615
rect 176 -1377 210 -1343
rect 176 -1445 210 -1411
rect 176 -1513 210 -1479
rect 176 -1581 210 -1547
rect -210 -1717 -176 -1683
rect 176 -1649 210 -1615
rect 176 -1717 210 -1683
rect -85 -1831 -51 -1797
rect -17 -1831 17 -1797
rect 51 -1831 85 -1797
<< poly >>
rect -50 1729 50 1745
rect -50 1695 -17 1729
rect 17 1695 50 1729
rect -50 1648 50 1695
rect -50 1301 50 1348
rect -50 1267 -17 1301
rect 17 1267 50 1301
rect -50 1220 50 1267
rect -50 873 50 920
rect -50 839 -17 873
rect 17 839 50 873
rect -50 792 50 839
rect -50 445 50 492
rect -50 411 -17 445
rect 17 411 50 445
rect -50 364 50 411
rect -50 17 50 64
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -64 50 -17
rect -50 -411 50 -364
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect -50 -492 50 -445
rect -50 -839 50 -792
rect -50 -873 -17 -839
rect 17 -873 50 -839
rect -50 -920 50 -873
rect -50 -1267 50 -1220
rect -50 -1301 -17 -1267
rect 17 -1301 50 -1267
rect -50 -1348 50 -1301
rect -50 -1695 50 -1648
rect -50 -1729 -17 -1695
rect 17 -1729 50 -1695
rect -50 -1745 50 -1729
<< polycont >>
rect -17 1695 17 1729
rect -17 1267 17 1301
rect -17 839 17 873
rect -17 411 17 445
rect -17 -17 17 17
rect -17 -445 17 -411
rect -17 -873 17 -839
rect -17 -1301 17 -1267
rect -17 -1729 17 -1695
<< locali >>
rect -210 1797 -85 1831
rect -51 1797 -17 1831
rect 17 1797 51 1831
rect 85 1797 210 1831
rect -210 1717 -176 1797
rect -50 1695 -17 1729
rect 17 1695 50 1729
rect 176 1717 210 1797
rect -210 1649 -176 1683
rect -210 1581 -176 1615
rect -210 1513 -176 1547
rect -210 1445 -176 1479
rect -210 1377 -176 1411
rect -96 1623 -62 1652
rect -96 1551 -62 1583
rect -96 1481 -62 1515
rect -96 1413 -62 1445
rect -96 1344 -62 1373
rect 62 1623 96 1652
rect 62 1551 96 1583
rect 62 1481 96 1515
rect 62 1413 96 1445
rect 62 1344 96 1373
rect 176 1649 210 1683
rect 176 1581 210 1615
rect 176 1513 210 1547
rect 176 1445 210 1479
rect 176 1377 210 1411
rect -210 1309 -176 1343
rect 176 1309 210 1343
rect -210 1241 -176 1275
rect -50 1267 -17 1301
rect 17 1267 50 1301
rect 176 1241 210 1275
rect -210 1173 -176 1207
rect -210 1105 -176 1139
rect -210 1037 -176 1071
rect -210 969 -176 1003
rect -210 901 -176 935
rect -96 1195 -62 1224
rect -96 1123 -62 1155
rect -96 1053 -62 1087
rect -96 985 -62 1017
rect -96 916 -62 945
rect 62 1195 96 1224
rect 62 1123 96 1155
rect 62 1053 96 1087
rect 62 985 96 1017
rect 62 916 96 945
rect 176 1173 210 1207
rect 176 1105 210 1139
rect 176 1037 210 1071
rect 176 969 210 1003
rect 176 901 210 935
rect -210 833 -176 867
rect -50 839 -17 873
rect 17 839 50 873
rect -210 765 -176 799
rect 176 833 210 867
rect -210 697 -176 731
rect -210 629 -176 663
rect -210 561 -176 595
rect -210 493 -176 527
rect -96 767 -62 796
rect -96 695 -62 727
rect -96 625 -62 659
rect -96 557 -62 589
rect -96 488 -62 517
rect 62 767 96 796
rect 62 695 96 727
rect 62 625 96 659
rect 62 557 96 589
rect 62 488 96 517
rect 176 765 210 799
rect 176 697 210 731
rect 176 629 210 663
rect 176 561 210 595
rect 176 493 210 527
rect -210 425 -176 459
rect -50 411 -17 445
rect 17 411 50 445
rect 176 425 210 459
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -96 339 -62 368
rect -96 267 -62 299
rect -96 197 -62 231
rect -96 129 -62 161
rect -96 60 -62 89
rect 62 339 96 368
rect 62 267 96 299
rect 62 197 96 231
rect 62 129 96 161
rect 62 60 96 89
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect 176 17 210 51
rect -50 -17 -17 17
rect 17 -17 50 17
rect -210 -51 -176 -17
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -96 -89 -62 -60
rect -96 -161 -62 -129
rect -96 -231 -62 -197
rect -96 -299 -62 -267
rect -96 -368 -62 -339
rect 62 -89 96 -60
rect 62 -161 96 -129
rect 62 -231 96 -197
rect 62 -299 96 -267
rect 62 -368 96 -339
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect -210 -459 -176 -425
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect 176 -459 210 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -210 -663 -176 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect -96 -517 -62 -488
rect -96 -589 -62 -557
rect -96 -659 -62 -625
rect -96 -727 -62 -695
rect -96 -796 -62 -767
rect 62 -517 96 -488
rect 62 -589 96 -557
rect 62 -659 96 -625
rect 62 -727 96 -695
rect 62 -796 96 -767
rect 176 -527 210 -493
rect 176 -595 210 -561
rect 176 -663 210 -629
rect 176 -731 210 -697
rect -210 -867 -176 -833
rect 176 -799 210 -765
rect -50 -873 -17 -839
rect 17 -873 50 -839
rect 176 -867 210 -833
rect -210 -935 -176 -901
rect -210 -1003 -176 -969
rect -210 -1071 -176 -1037
rect -210 -1139 -176 -1105
rect -210 -1207 -176 -1173
rect -96 -945 -62 -916
rect -96 -1017 -62 -985
rect -96 -1087 -62 -1053
rect -96 -1155 -62 -1123
rect -96 -1224 -62 -1195
rect 62 -945 96 -916
rect 62 -1017 96 -985
rect 62 -1087 96 -1053
rect 62 -1155 96 -1123
rect 62 -1224 96 -1195
rect 176 -935 210 -901
rect 176 -1003 210 -969
rect 176 -1071 210 -1037
rect 176 -1139 210 -1105
rect 176 -1207 210 -1173
rect -210 -1275 -176 -1241
rect -50 -1301 -17 -1267
rect 17 -1301 50 -1267
rect 176 -1275 210 -1241
rect -210 -1343 -176 -1309
rect 176 -1343 210 -1309
rect -210 -1411 -176 -1377
rect -210 -1479 -176 -1445
rect -210 -1547 -176 -1513
rect -210 -1615 -176 -1581
rect -210 -1683 -176 -1649
rect -96 -1373 -62 -1344
rect -96 -1445 -62 -1413
rect -96 -1515 -62 -1481
rect -96 -1583 -62 -1551
rect -96 -1652 -62 -1623
rect 62 -1373 96 -1344
rect 62 -1445 96 -1413
rect 62 -1515 96 -1481
rect 62 -1583 96 -1551
rect 62 -1652 96 -1623
rect 176 -1411 210 -1377
rect 176 -1479 210 -1445
rect 176 -1547 210 -1513
rect 176 -1615 210 -1581
rect 176 -1683 210 -1649
rect -210 -1797 -176 -1717
rect -50 -1729 -17 -1695
rect 17 -1729 50 -1695
rect 176 -1797 210 -1717
rect -210 -1831 -85 -1797
rect -51 -1831 -17 -1797
rect 17 -1831 51 -1797
rect 85 -1831 210 -1797
<< viali >>
rect -17 1695 17 1729
rect -96 1617 -62 1623
rect -96 1589 -62 1617
rect -96 1549 -62 1551
rect -96 1517 -62 1549
rect -96 1447 -62 1479
rect -96 1445 -62 1447
rect -96 1379 -62 1407
rect -96 1373 -62 1379
rect 62 1617 96 1623
rect 62 1589 96 1617
rect 62 1549 96 1551
rect 62 1517 96 1549
rect 62 1447 96 1479
rect 62 1445 96 1447
rect 62 1379 96 1407
rect 62 1373 96 1379
rect -17 1267 17 1301
rect -96 1189 -62 1195
rect -96 1161 -62 1189
rect -96 1121 -62 1123
rect -96 1089 -62 1121
rect -96 1019 -62 1051
rect -96 1017 -62 1019
rect -96 951 -62 979
rect -96 945 -62 951
rect 62 1189 96 1195
rect 62 1161 96 1189
rect 62 1121 96 1123
rect 62 1089 96 1121
rect 62 1019 96 1051
rect 62 1017 96 1019
rect 62 951 96 979
rect 62 945 96 951
rect -17 839 17 873
rect -96 761 -62 767
rect -96 733 -62 761
rect -96 693 -62 695
rect -96 661 -62 693
rect -96 591 -62 623
rect -96 589 -62 591
rect -96 523 -62 551
rect -96 517 -62 523
rect 62 761 96 767
rect 62 733 96 761
rect 62 693 96 695
rect 62 661 96 693
rect 62 591 96 623
rect 62 589 96 591
rect 62 523 96 551
rect 62 517 96 523
rect -17 411 17 445
rect -96 333 -62 339
rect -96 305 -62 333
rect -96 265 -62 267
rect -96 233 -62 265
rect -96 163 -62 195
rect -96 161 -62 163
rect -96 95 -62 123
rect -96 89 -62 95
rect 62 333 96 339
rect 62 305 96 333
rect 62 265 96 267
rect 62 233 96 265
rect 62 163 96 195
rect 62 161 96 163
rect 62 95 96 123
rect 62 89 96 95
rect -17 -17 17 17
rect -96 -95 -62 -89
rect -96 -123 -62 -95
rect -96 -163 -62 -161
rect -96 -195 -62 -163
rect -96 -265 -62 -233
rect -96 -267 -62 -265
rect -96 -333 -62 -305
rect -96 -339 -62 -333
rect 62 -95 96 -89
rect 62 -123 96 -95
rect 62 -163 96 -161
rect 62 -195 96 -163
rect 62 -265 96 -233
rect 62 -267 96 -265
rect 62 -333 96 -305
rect 62 -339 96 -333
rect -17 -445 17 -411
rect -96 -523 -62 -517
rect -96 -551 -62 -523
rect -96 -591 -62 -589
rect -96 -623 -62 -591
rect -96 -693 -62 -661
rect -96 -695 -62 -693
rect -96 -761 -62 -733
rect -96 -767 -62 -761
rect 62 -523 96 -517
rect 62 -551 96 -523
rect 62 -591 96 -589
rect 62 -623 96 -591
rect 62 -693 96 -661
rect 62 -695 96 -693
rect 62 -761 96 -733
rect 62 -767 96 -761
rect -17 -873 17 -839
rect -96 -951 -62 -945
rect -96 -979 -62 -951
rect -96 -1019 -62 -1017
rect -96 -1051 -62 -1019
rect -96 -1121 -62 -1089
rect -96 -1123 -62 -1121
rect -96 -1189 -62 -1161
rect -96 -1195 -62 -1189
rect 62 -951 96 -945
rect 62 -979 96 -951
rect 62 -1019 96 -1017
rect 62 -1051 96 -1019
rect 62 -1121 96 -1089
rect 62 -1123 96 -1121
rect 62 -1189 96 -1161
rect 62 -1195 96 -1189
rect -17 -1301 17 -1267
rect -96 -1379 -62 -1373
rect -96 -1407 -62 -1379
rect -96 -1447 -62 -1445
rect -96 -1479 -62 -1447
rect -96 -1549 -62 -1517
rect -96 -1551 -62 -1549
rect -96 -1617 -62 -1589
rect -96 -1623 -62 -1617
rect 62 -1379 96 -1373
rect 62 -1407 96 -1379
rect 62 -1447 96 -1445
rect 62 -1479 96 -1447
rect 62 -1549 96 -1517
rect 62 -1551 96 -1549
rect 62 -1617 96 -1589
rect 62 -1623 96 -1617
rect -17 -1729 17 -1695
<< metal1 >>
rect -46 1729 46 1735
rect -46 1695 -17 1729
rect 17 1695 46 1729
rect -46 1689 46 1695
rect -102 1623 -56 1648
rect -102 1589 -96 1623
rect -62 1589 -56 1623
rect -102 1551 -56 1589
rect -102 1517 -96 1551
rect -62 1517 -56 1551
rect -102 1479 -56 1517
rect -102 1445 -96 1479
rect -62 1445 -56 1479
rect -102 1407 -56 1445
rect -102 1373 -96 1407
rect -62 1373 -56 1407
rect -102 1348 -56 1373
rect 56 1623 102 1648
rect 56 1589 62 1623
rect 96 1589 102 1623
rect 56 1551 102 1589
rect 56 1517 62 1551
rect 96 1517 102 1551
rect 56 1479 102 1517
rect 56 1445 62 1479
rect 96 1445 102 1479
rect 56 1407 102 1445
rect 56 1373 62 1407
rect 96 1373 102 1407
rect 56 1348 102 1373
rect -46 1301 46 1307
rect -46 1267 -17 1301
rect 17 1267 46 1301
rect -46 1261 46 1267
rect -102 1195 -56 1220
rect -102 1161 -96 1195
rect -62 1161 -56 1195
rect -102 1123 -56 1161
rect -102 1089 -96 1123
rect -62 1089 -56 1123
rect -102 1051 -56 1089
rect -102 1017 -96 1051
rect -62 1017 -56 1051
rect -102 979 -56 1017
rect -102 945 -96 979
rect -62 945 -56 979
rect -102 920 -56 945
rect 56 1195 102 1220
rect 56 1161 62 1195
rect 96 1161 102 1195
rect 56 1123 102 1161
rect 56 1089 62 1123
rect 96 1089 102 1123
rect 56 1051 102 1089
rect 56 1017 62 1051
rect 96 1017 102 1051
rect 56 979 102 1017
rect 56 945 62 979
rect 96 945 102 979
rect 56 920 102 945
rect -46 873 46 879
rect -46 839 -17 873
rect 17 839 46 873
rect -46 833 46 839
rect -102 767 -56 792
rect -102 733 -96 767
rect -62 733 -56 767
rect -102 695 -56 733
rect -102 661 -96 695
rect -62 661 -56 695
rect -102 623 -56 661
rect -102 589 -96 623
rect -62 589 -56 623
rect -102 551 -56 589
rect -102 517 -96 551
rect -62 517 -56 551
rect -102 492 -56 517
rect 56 767 102 792
rect 56 733 62 767
rect 96 733 102 767
rect 56 695 102 733
rect 56 661 62 695
rect 96 661 102 695
rect 56 623 102 661
rect 56 589 62 623
rect 96 589 102 623
rect 56 551 102 589
rect 56 517 62 551
rect 96 517 102 551
rect 56 492 102 517
rect -46 445 46 451
rect -46 411 -17 445
rect 17 411 46 445
rect -46 405 46 411
rect -102 339 -56 364
rect -102 305 -96 339
rect -62 305 -56 339
rect -102 267 -56 305
rect -102 233 -96 267
rect -62 233 -56 267
rect -102 195 -56 233
rect -102 161 -96 195
rect -62 161 -56 195
rect -102 123 -56 161
rect -102 89 -96 123
rect -62 89 -56 123
rect -102 64 -56 89
rect 56 339 102 364
rect 56 305 62 339
rect 96 305 102 339
rect 56 267 102 305
rect 56 233 62 267
rect 96 233 102 267
rect 56 195 102 233
rect 56 161 62 195
rect 96 161 102 195
rect 56 123 102 161
rect 56 89 62 123
rect 96 89 102 123
rect 56 64 102 89
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -89 -56 -64
rect -102 -123 -96 -89
rect -62 -123 -56 -89
rect -102 -161 -56 -123
rect -102 -195 -96 -161
rect -62 -195 -56 -161
rect -102 -233 -56 -195
rect -102 -267 -96 -233
rect -62 -267 -56 -233
rect -102 -305 -56 -267
rect -102 -339 -96 -305
rect -62 -339 -56 -305
rect -102 -364 -56 -339
rect 56 -89 102 -64
rect 56 -123 62 -89
rect 96 -123 102 -89
rect 56 -161 102 -123
rect 56 -195 62 -161
rect 96 -195 102 -161
rect 56 -233 102 -195
rect 56 -267 62 -233
rect 96 -267 102 -233
rect 56 -305 102 -267
rect 56 -339 62 -305
rect 96 -339 102 -305
rect 56 -364 102 -339
rect -46 -411 46 -405
rect -46 -445 -17 -411
rect 17 -445 46 -411
rect -46 -451 46 -445
rect -102 -517 -56 -492
rect -102 -551 -96 -517
rect -62 -551 -56 -517
rect -102 -589 -56 -551
rect -102 -623 -96 -589
rect -62 -623 -56 -589
rect -102 -661 -56 -623
rect -102 -695 -96 -661
rect -62 -695 -56 -661
rect -102 -733 -56 -695
rect -102 -767 -96 -733
rect -62 -767 -56 -733
rect -102 -792 -56 -767
rect 56 -517 102 -492
rect 56 -551 62 -517
rect 96 -551 102 -517
rect 56 -589 102 -551
rect 56 -623 62 -589
rect 96 -623 102 -589
rect 56 -661 102 -623
rect 56 -695 62 -661
rect 96 -695 102 -661
rect 56 -733 102 -695
rect 56 -767 62 -733
rect 96 -767 102 -733
rect 56 -792 102 -767
rect -46 -839 46 -833
rect -46 -873 -17 -839
rect 17 -873 46 -839
rect -46 -879 46 -873
rect -102 -945 -56 -920
rect -102 -979 -96 -945
rect -62 -979 -56 -945
rect -102 -1017 -56 -979
rect -102 -1051 -96 -1017
rect -62 -1051 -56 -1017
rect -102 -1089 -56 -1051
rect -102 -1123 -96 -1089
rect -62 -1123 -56 -1089
rect -102 -1161 -56 -1123
rect -102 -1195 -96 -1161
rect -62 -1195 -56 -1161
rect -102 -1220 -56 -1195
rect 56 -945 102 -920
rect 56 -979 62 -945
rect 96 -979 102 -945
rect 56 -1017 102 -979
rect 56 -1051 62 -1017
rect 96 -1051 102 -1017
rect 56 -1089 102 -1051
rect 56 -1123 62 -1089
rect 96 -1123 102 -1089
rect 56 -1161 102 -1123
rect 56 -1195 62 -1161
rect 96 -1195 102 -1161
rect 56 -1220 102 -1195
rect -46 -1267 46 -1261
rect -46 -1301 -17 -1267
rect 17 -1301 46 -1267
rect -46 -1307 46 -1301
rect -102 -1373 -56 -1348
rect -102 -1407 -96 -1373
rect -62 -1407 -56 -1373
rect -102 -1445 -56 -1407
rect -102 -1479 -96 -1445
rect -62 -1479 -56 -1445
rect -102 -1517 -56 -1479
rect -102 -1551 -96 -1517
rect -62 -1551 -56 -1517
rect -102 -1589 -56 -1551
rect -102 -1623 -96 -1589
rect -62 -1623 -56 -1589
rect -102 -1648 -56 -1623
rect 56 -1373 102 -1348
rect 56 -1407 62 -1373
rect 96 -1407 102 -1373
rect 56 -1445 102 -1407
rect 56 -1479 62 -1445
rect 96 -1479 102 -1445
rect 56 -1517 102 -1479
rect 56 -1551 62 -1517
rect 96 -1551 102 -1517
rect 56 -1589 102 -1551
rect 56 -1623 62 -1589
rect 96 -1623 102 -1589
rect 56 -1648 102 -1623
rect -46 -1695 46 -1689
rect -46 -1729 -17 -1695
rect 17 -1729 46 -1695
rect -46 -1735 46 -1729
<< properties >>
string FIXED_BBOX -193 -1814 193 1814
<< end >>
