magic
tech sky130A
magscale 1 2
timestamp 1757832390
<< metal3 >>
rect -1904 2732 -1132 2760
rect -1904 2308 -1216 2732
rect -1152 2308 -1132 2732
rect -1904 2280 -1132 2308
rect -892 2732 -120 2760
rect -892 2308 -204 2732
rect -140 2308 -120 2732
rect -892 2280 -120 2308
rect 120 2732 892 2760
rect 120 2308 808 2732
rect 872 2308 892 2732
rect 120 2280 892 2308
rect 1132 2732 1904 2760
rect 1132 2308 1820 2732
rect 1884 2308 1904 2732
rect 1132 2280 1904 2308
rect -1904 2012 -1132 2040
rect -1904 1588 -1216 2012
rect -1152 1588 -1132 2012
rect -1904 1560 -1132 1588
rect -892 2012 -120 2040
rect -892 1588 -204 2012
rect -140 1588 -120 2012
rect -892 1560 -120 1588
rect 120 2012 892 2040
rect 120 1588 808 2012
rect 872 1588 892 2012
rect 120 1560 892 1588
rect 1132 2012 1904 2040
rect 1132 1588 1820 2012
rect 1884 1588 1904 2012
rect 1132 1560 1904 1588
rect -1904 1292 -1132 1320
rect -1904 868 -1216 1292
rect -1152 868 -1132 1292
rect -1904 840 -1132 868
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect 1132 1292 1904 1320
rect 1132 868 1820 1292
rect 1884 868 1904 1292
rect 1132 840 1904 868
rect -1904 572 -1132 600
rect -1904 148 -1216 572
rect -1152 148 -1132 572
rect -1904 120 -1132 148
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect 1132 572 1904 600
rect 1132 148 1820 572
rect 1884 148 1904 572
rect 1132 120 1904 148
rect -1904 -148 -1132 -120
rect -1904 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -1904 -600 -1132 -572
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect 1132 -148 1904 -120
rect 1132 -572 1820 -148
rect 1884 -572 1904 -148
rect 1132 -600 1904 -572
rect -1904 -868 -1132 -840
rect -1904 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -1904 -1320 -1132 -1292
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect 1132 -868 1904 -840
rect 1132 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 1132 -1320 1904 -1292
rect -1904 -1588 -1132 -1560
rect -1904 -2012 -1216 -1588
rect -1152 -2012 -1132 -1588
rect -1904 -2040 -1132 -2012
rect -892 -1588 -120 -1560
rect -892 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect -892 -2040 -120 -2012
rect 120 -1588 892 -1560
rect 120 -2012 808 -1588
rect 872 -2012 892 -1588
rect 120 -2040 892 -2012
rect 1132 -1588 1904 -1560
rect 1132 -2012 1820 -1588
rect 1884 -2012 1904 -1588
rect 1132 -2040 1904 -2012
rect -1904 -2308 -1132 -2280
rect -1904 -2732 -1216 -2308
rect -1152 -2732 -1132 -2308
rect -1904 -2760 -1132 -2732
rect -892 -2308 -120 -2280
rect -892 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect -892 -2760 -120 -2732
rect 120 -2308 892 -2280
rect 120 -2732 808 -2308
rect 872 -2732 892 -2308
rect 120 -2760 892 -2732
rect 1132 -2308 1904 -2280
rect 1132 -2732 1820 -2308
rect 1884 -2732 1904 -2308
rect 1132 -2760 1904 -2732
<< via3 >>
rect -1216 2308 -1152 2732
rect -204 2308 -140 2732
rect 808 2308 872 2732
rect 1820 2308 1884 2732
rect -1216 1588 -1152 2012
rect -204 1588 -140 2012
rect 808 1588 872 2012
rect 1820 1588 1884 2012
rect -1216 868 -1152 1292
rect -204 868 -140 1292
rect 808 868 872 1292
rect 1820 868 1884 1292
rect -1216 148 -1152 572
rect -204 148 -140 572
rect 808 148 872 572
rect 1820 148 1884 572
rect -1216 -572 -1152 -148
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect 1820 -572 1884 -148
rect -1216 -1292 -1152 -868
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect 1820 -1292 1884 -868
rect -1216 -2012 -1152 -1588
rect -204 -2012 -140 -1588
rect 808 -2012 872 -1588
rect 1820 -2012 1884 -1588
rect -1216 -2732 -1152 -2308
rect -204 -2732 -140 -2308
rect 808 -2732 872 -2308
rect 1820 -2732 1884 -2308
<< mimcap >>
rect -1864 2680 -1464 2720
rect -1864 2360 -1824 2680
rect -1504 2360 -1464 2680
rect -1864 2320 -1464 2360
rect -852 2680 -452 2720
rect -852 2360 -812 2680
rect -492 2360 -452 2680
rect -852 2320 -452 2360
rect 160 2680 560 2720
rect 160 2360 200 2680
rect 520 2360 560 2680
rect 160 2320 560 2360
rect 1172 2680 1572 2720
rect 1172 2360 1212 2680
rect 1532 2360 1572 2680
rect 1172 2320 1572 2360
rect -1864 1960 -1464 2000
rect -1864 1640 -1824 1960
rect -1504 1640 -1464 1960
rect -1864 1600 -1464 1640
rect -852 1960 -452 2000
rect -852 1640 -812 1960
rect -492 1640 -452 1960
rect -852 1600 -452 1640
rect 160 1960 560 2000
rect 160 1640 200 1960
rect 520 1640 560 1960
rect 160 1600 560 1640
rect 1172 1960 1572 2000
rect 1172 1640 1212 1960
rect 1532 1640 1572 1960
rect 1172 1600 1572 1640
rect -1864 1240 -1464 1280
rect -1864 920 -1824 1240
rect -1504 920 -1464 1240
rect -1864 880 -1464 920
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect 1172 1240 1572 1280
rect 1172 920 1212 1240
rect 1532 920 1572 1240
rect 1172 880 1572 920
rect -1864 520 -1464 560
rect -1864 200 -1824 520
rect -1504 200 -1464 520
rect -1864 160 -1464 200
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect 1172 520 1572 560
rect 1172 200 1212 520
rect 1532 200 1572 520
rect 1172 160 1572 200
rect -1864 -200 -1464 -160
rect -1864 -520 -1824 -200
rect -1504 -520 -1464 -200
rect -1864 -560 -1464 -520
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect 1172 -200 1572 -160
rect 1172 -520 1212 -200
rect 1532 -520 1572 -200
rect 1172 -560 1572 -520
rect -1864 -920 -1464 -880
rect -1864 -1240 -1824 -920
rect -1504 -1240 -1464 -920
rect -1864 -1280 -1464 -1240
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect 1172 -920 1572 -880
rect 1172 -1240 1212 -920
rect 1532 -1240 1572 -920
rect 1172 -1280 1572 -1240
rect -1864 -1640 -1464 -1600
rect -1864 -1960 -1824 -1640
rect -1504 -1960 -1464 -1640
rect -1864 -2000 -1464 -1960
rect -852 -1640 -452 -1600
rect -852 -1960 -812 -1640
rect -492 -1960 -452 -1640
rect -852 -2000 -452 -1960
rect 160 -1640 560 -1600
rect 160 -1960 200 -1640
rect 520 -1960 560 -1640
rect 160 -2000 560 -1960
rect 1172 -1640 1572 -1600
rect 1172 -1960 1212 -1640
rect 1532 -1960 1572 -1640
rect 1172 -2000 1572 -1960
rect -1864 -2360 -1464 -2320
rect -1864 -2680 -1824 -2360
rect -1504 -2680 -1464 -2360
rect -1864 -2720 -1464 -2680
rect -852 -2360 -452 -2320
rect -852 -2680 -812 -2360
rect -492 -2680 -452 -2360
rect -852 -2720 -452 -2680
rect 160 -2360 560 -2320
rect 160 -2680 200 -2360
rect 520 -2680 560 -2360
rect 160 -2720 560 -2680
rect 1172 -2360 1572 -2320
rect 1172 -2680 1212 -2360
rect 1532 -2680 1572 -2360
rect 1172 -2720 1572 -2680
<< mimcapcontact >>
rect -1824 2360 -1504 2680
rect -812 2360 -492 2680
rect 200 2360 520 2680
rect 1212 2360 1532 2680
rect -1824 1640 -1504 1960
rect -812 1640 -492 1960
rect 200 1640 520 1960
rect 1212 1640 1532 1960
rect -1824 920 -1504 1240
rect -812 920 -492 1240
rect 200 920 520 1240
rect 1212 920 1532 1240
rect -1824 200 -1504 520
rect -812 200 -492 520
rect 200 200 520 520
rect 1212 200 1532 520
rect -1824 -520 -1504 -200
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect 1212 -520 1532 -200
rect -1824 -1240 -1504 -920
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect 1212 -1240 1532 -920
rect -1824 -1960 -1504 -1640
rect -812 -1960 -492 -1640
rect 200 -1960 520 -1640
rect 1212 -1960 1532 -1640
rect -1824 -2680 -1504 -2360
rect -812 -2680 -492 -2360
rect 200 -2680 520 -2360
rect 1212 -2680 1532 -2360
<< metal4 >>
rect -1716 2681 -1612 2880
rect -1236 2732 -1132 2880
rect -1825 2680 -1503 2681
rect -1825 2360 -1824 2680
rect -1504 2360 -1503 2680
rect -1825 2359 -1503 2360
rect -1716 1961 -1612 2359
rect -1236 2308 -1216 2732
rect -1152 2308 -1132 2732
rect -704 2681 -600 2880
rect -224 2732 -120 2880
rect -813 2680 -491 2681
rect -813 2360 -812 2680
rect -492 2360 -491 2680
rect -813 2359 -491 2360
rect -1236 2012 -1132 2308
rect -1825 1960 -1503 1961
rect -1825 1640 -1824 1960
rect -1504 1640 -1503 1960
rect -1825 1639 -1503 1640
rect -1716 1241 -1612 1639
rect -1236 1588 -1216 2012
rect -1152 1588 -1132 2012
rect -704 1961 -600 2359
rect -224 2308 -204 2732
rect -140 2308 -120 2732
rect 308 2681 412 2880
rect 788 2732 892 2880
rect 199 2680 521 2681
rect 199 2360 200 2680
rect 520 2360 521 2680
rect 199 2359 521 2360
rect -224 2012 -120 2308
rect -813 1960 -491 1961
rect -813 1640 -812 1960
rect -492 1640 -491 1960
rect -813 1639 -491 1640
rect -1236 1292 -1132 1588
rect -1825 1240 -1503 1241
rect -1825 920 -1824 1240
rect -1504 920 -1503 1240
rect -1825 919 -1503 920
rect -1716 521 -1612 919
rect -1236 868 -1216 1292
rect -1152 868 -1132 1292
rect -704 1241 -600 1639
rect -224 1588 -204 2012
rect -140 1588 -120 2012
rect 308 1961 412 2359
rect 788 2308 808 2732
rect 872 2308 892 2732
rect 1320 2681 1424 2880
rect 1800 2732 1904 2880
rect 1211 2680 1533 2681
rect 1211 2360 1212 2680
rect 1532 2360 1533 2680
rect 1211 2359 1533 2360
rect 788 2012 892 2308
rect 199 1960 521 1961
rect 199 1640 200 1960
rect 520 1640 521 1960
rect 199 1639 521 1640
rect -224 1292 -120 1588
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -1236 572 -1132 868
rect -1825 520 -1503 521
rect -1825 200 -1824 520
rect -1504 200 -1503 520
rect -1825 199 -1503 200
rect -1716 -199 -1612 199
rect -1236 148 -1216 572
rect -1152 148 -1132 572
rect -704 521 -600 919
rect -224 868 -204 1292
rect -140 868 -120 1292
rect 308 1241 412 1639
rect 788 1588 808 2012
rect 872 1588 892 2012
rect 1320 1961 1424 2359
rect 1800 2308 1820 2732
rect 1884 2308 1904 2732
rect 1800 2012 1904 2308
rect 1211 1960 1533 1961
rect 1211 1640 1212 1960
rect 1532 1640 1533 1960
rect 1211 1639 1533 1640
rect 788 1292 892 1588
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -224 572 -120 868
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -1236 -148 -1132 148
rect -1825 -200 -1503 -199
rect -1825 -520 -1824 -200
rect -1504 -520 -1503 -200
rect -1825 -521 -1503 -520
rect -1716 -919 -1612 -521
rect -1236 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -704 -199 -600 199
rect -224 148 -204 572
rect -140 148 -120 572
rect 308 521 412 919
rect 788 868 808 1292
rect 872 868 892 1292
rect 1320 1241 1424 1639
rect 1800 1588 1820 2012
rect 1884 1588 1904 2012
rect 1800 1292 1904 1588
rect 1211 1240 1533 1241
rect 1211 920 1212 1240
rect 1532 920 1533 1240
rect 1211 919 1533 920
rect 788 572 892 868
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -1236 -868 -1132 -572
rect -1825 -920 -1503 -919
rect -1825 -1240 -1824 -920
rect -1504 -1240 -1503 -920
rect -1825 -1241 -1503 -1240
rect -1716 -1639 -1612 -1241
rect -1236 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -704 -919 -600 -521
rect -224 -572 -204 -148
rect -140 -572 -120 -148
rect 308 -199 412 199
rect 788 148 808 572
rect 872 148 892 572
rect 1320 521 1424 919
rect 1800 868 1820 1292
rect 1884 868 1904 1292
rect 1800 572 1904 868
rect 1211 520 1533 521
rect 1211 200 1212 520
rect 1532 200 1533 520
rect 1211 199 1533 200
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -224 -868 -120 -572
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -1236 -1588 -1132 -1292
rect -1825 -1640 -1503 -1639
rect -1825 -1960 -1824 -1640
rect -1504 -1960 -1503 -1640
rect -1825 -1961 -1503 -1960
rect -1716 -2359 -1612 -1961
rect -1236 -2012 -1216 -1588
rect -1152 -2012 -1132 -1588
rect -704 -1639 -600 -1241
rect -224 -1292 -204 -868
rect -140 -1292 -120 -868
rect 308 -919 412 -521
rect 788 -572 808 -148
rect 872 -572 892 -148
rect 1320 -199 1424 199
rect 1800 148 1820 572
rect 1884 148 1904 572
rect 1800 -148 1904 148
rect 1211 -200 1533 -199
rect 1211 -520 1212 -200
rect 1532 -520 1533 -200
rect 1211 -521 1533 -520
rect 788 -868 892 -572
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -224 -1588 -120 -1292
rect -813 -1640 -491 -1639
rect -813 -1960 -812 -1640
rect -492 -1960 -491 -1640
rect -813 -1961 -491 -1960
rect -1236 -2308 -1132 -2012
rect -1825 -2360 -1503 -2359
rect -1825 -2680 -1824 -2360
rect -1504 -2680 -1503 -2360
rect -1825 -2681 -1503 -2680
rect -1716 -2880 -1612 -2681
rect -1236 -2732 -1216 -2308
rect -1152 -2732 -1132 -2308
rect -704 -2359 -600 -1961
rect -224 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect 308 -1639 412 -1241
rect 788 -1292 808 -868
rect 872 -1292 892 -868
rect 1320 -919 1424 -521
rect 1800 -572 1820 -148
rect 1884 -572 1904 -148
rect 1800 -868 1904 -572
rect 1211 -920 1533 -919
rect 1211 -1240 1212 -920
rect 1532 -1240 1533 -920
rect 1211 -1241 1533 -1240
rect 788 -1588 892 -1292
rect 199 -1640 521 -1639
rect 199 -1960 200 -1640
rect 520 -1960 521 -1640
rect 199 -1961 521 -1960
rect -224 -2308 -120 -2012
rect -813 -2360 -491 -2359
rect -813 -2680 -812 -2360
rect -492 -2680 -491 -2360
rect -813 -2681 -491 -2680
rect -1236 -2880 -1132 -2732
rect -704 -2880 -600 -2681
rect -224 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect 308 -2359 412 -1961
rect 788 -2012 808 -1588
rect 872 -2012 892 -1588
rect 1320 -1639 1424 -1241
rect 1800 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 1800 -1588 1904 -1292
rect 1211 -1640 1533 -1639
rect 1211 -1960 1212 -1640
rect 1532 -1960 1533 -1640
rect 1211 -1961 1533 -1960
rect 788 -2308 892 -2012
rect 199 -2360 521 -2359
rect 199 -2680 200 -2360
rect 520 -2680 521 -2360
rect 199 -2681 521 -2680
rect -224 -2880 -120 -2732
rect 308 -2880 412 -2681
rect 788 -2732 808 -2308
rect 872 -2732 892 -2308
rect 1320 -2359 1424 -1961
rect 1800 -2012 1820 -1588
rect 1884 -2012 1904 -1588
rect 1800 -2308 1904 -2012
rect 1211 -2360 1533 -2359
rect 1211 -2680 1212 -2360
rect 1532 -2680 1533 -2360
rect 1211 -2681 1533 -2680
rect 788 -2880 892 -2732
rect 1320 -2880 1424 -2681
rect 1800 -2732 1820 -2308
rect 1884 -2732 1904 -2308
rect 1800 -2880 1904 -2732
<< properties >>
string FIXED_BBOX 1132 2280 1612 2760
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 4 ny 8 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
