magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal3 >>
rect -23884 18312 -22712 18360
rect -23884 18248 -22796 18312
rect -22732 18248 -22712 18312
rect -23884 18232 -22712 18248
rect -23884 18168 -22796 18232
rect -22732 18168 -22712 18232
rect -23884 18152 -22712 18168
rect -23884 18088 -22796 18152
rect -22732 18088 -22712 18152
rect -23884 18072 -22712 18088
rect -23884 18008 -22796 18072
rect -22732 18008 -22712 18072
rect -23884 17992 -22712 18008
rect -23884 17928 -22796 17992
rect -22732 17928 -22712 17992
rect -23884 17912 -22712 17928
rect -23884 17848 -22796 17912
rect -22732 17848 -22712 17912
rect -23884 17832 -22712 17848
rect -23884 17768 -22796 17832
rect -22732 17768 -22712 17832
rect -23884 17752 -22712 17768
rect -23884 17688 -22796 17752
rect -22732 17688 -22712 17752
rect -23884 17672 -22712 17688
rect -23884 17608 -22796 17672
rect -22732 17608 -22712 17672
rect -23884 17592 -22712 17608
rect -23884 17528 -22796 17592
rect -22732 17528 -22712 17592
rect -23884 17480 -22712 17528
rect -22472 18312 -21300 18360
rect -22472 18248 -21384 18312
rect -21320 18248 -21300 18312
rect -22472 18232 -21300 18248
rect -22472 18168 -21384 18232
rect -21320 18168 -21300 18232
rect -22472 18152 -21300 18168
rect -22472 18088 -21384 18152
rect -21320 18088 -21300 18152
rect -22472 18072 -21300 18088
rect -22472 18008 -21384 18072
rect -21320 18008 -21300 18072
rect -22472 17992 -21300 18008
rect -22472 17928 -21384 17992
rect -21320 17928 -21300 17992
rect -22472 17912 -21300 17928
rect -22472 17848 -21384 17912
rect -21320 17848 -21300 17912
rect -22472 17832 -21300 17848
rect -22472 17768 -21384 17832
rect -21320 17768 -21300 17832
rect -22472 17752 -21300 17768
rect -22472 17688 -21384 17752
rect -21320 17688 -21300 17752
rect -22472 17672 -21300 17688
rect -22472 17608 -21384 17672
rect -21320 17608 -21300 17672
rect -22472 17592 -21300 17608
rect -22472 17528 -21384 17592
rect -21320 17528 -21300 17592
rect -22472 17480 -21300 17528
rect -21060 18312 -19888 18360
rect -21060 18248 -19972 18312
rect -19908 18248 -19888 18312
rect -21060 18232 -19888 18248
rect -21060 18168 -19972 18232
rect -19908 18168 -19888 18232
rect -21060 18152 -19888 18168
rect -21060 18088 -19972 18152
rect -19908 18088 -19888 18152
rect -21060 18072 -19888 18088
rect -21060 18008 -19972 18072
rect -19908 18008 -19888 18072
rect -21060 17992 -19888 18008
rect -21060 17928 -19972 17992
rect -19908 17928 -19888 17992
rect -21060 17912 -19888 17928
rect -21060 17848 -19972 17912
rect -19908 17848 -19888 17912
rect -21060 17832 -19888 17848
rect -21060 17768 -19972 17832
rect -19908 17768 -19888 17832
rect -21060 17752 -19888 17768
rect -21060 17688 -19972 17752
rect -19908 17688 -19888 17752
rect -21060 17672 -19888 17688
rect -21060 17608 -19972 17672
rect -19908 17608 -19888 17672
rect -21060 17592 -19888 17608
rect -21060 17528 -19972 17592
rect -19908 17528 -19888 17592
rect -21060 17480 -19888 17528
rect -19648 18312 -18476 18360
rect -19648 18248 -18560 18312
rect -18496 18248 -18476 18312
rect -19648 18232 -18476 18248
rect -19648 18168 -18560 18232
rect -18496 18168 -18476 18232
rect -19648 18152 -18476 18168
rect -19648 18088 -18560 18152
rect -18496 18088 -18476 18152
rect -19648 18072 -18476 18088
rect -19648 18008 -18560 18072
rect -18496 18008 -18476 18072
rect -19648 17992 -18476 18008
rect -19648 17928 -18560 17992
rect -18496 17928 -18476 17992
rect -19648 17912 -18476 17928
rect -19648 17848 -18560 17912
rect -18496 17848 -18476 17912
rect -19648 17832 -18476 17848
rect -19648 17768 -18560 17832
rect -18496 17768 -18476 17832
rect -19648 17752 -18476 17768
rect -19648 17688 -18560 17752
rect -18496 17688 -18476 17752
rect -19648 17672 -18476 17688
rect -19648 17608 -18560 17672
rect -18496 17608 -18476 17672
rect -19648 17592 -18476 17608
rect -19648 17528 -18560 17592
rect -18496 17528 -18476 17592
rect -19648 17480 -18476 17528
rect -18236 18312 -17064 18360
rect -18236 18248 -17148 18312
rect -17084 18248 -17064 18312
rect -18236 18232 -17064 18248
rect -18236 18168 -17148 18232
rect -17084 18168 -17064 18232
rect -18236 18152 -17064 18168
rect -18236 18088 -17148 18152
rect -17084 18088 -17064 18152
rect -18236 18072 -17064 18088
rect -18236 18008 -17148 18072
rect -17084 18008 -17064 18072
rect -18236 17992 -17064 18008
rect -18236 17928 -17148 17992
rect -17084 17928 -17064 17992
rect -18236 17912 -17064 17928
rect -18236 17848 -17148 17912
rect -17084 17848 -17064 17912
rect -18236 17832 -17064 17848
rect -18236 17768 -17148 17832
rect -17084 17768 -17064 17832
rect -18236 17752 -17064 17768
rect -18236 17688 -17148 17752
rect -17084 17688 -17064 17752
rect -18236 17672 -17064 17688
rect -18236 17608 -17148 17672
rect -17084 17608 -17064 17672
rect -18236 17592 -17064 17608
rect -18236 17528 -17148 17592
rect -17084 17528 -17064 17592
rect -18236 17480 -17064 17528
rect -16824 18312 -15652 18360
rect -16824 18248 -15736 18312
rect -15672 18248 -15652 18312
rect -16824 18232 -15652 18248
rect -16824 18168 -15736 18232
rect -15672 18168 -15652 18232
rect -16824 18152 -15652 18168
rect -16824 18088 -15736 18152
rect -15672 18088 -15652 18152
rect -16824 18072 -15652 18088
rect -16824 18008 -15736 18072
rect -15672 18008 -15652 18072
rect -16824 17992 -15652 18008
rect -16824 17928 -15736 17992
rect -15672 17928 -15652 17992
rect -16824 17912 -15652 17928
rect -16824 17848 -15736 17912
rect -15672 17848 -15652 17912
rect -16824 17832 -15652 17848
rect -16824 17768 -15736 17832
rect -15672 17768 -15652 17832
rect -16824 17752 -15652 17768
rect -16824 17688 -15736 17752
rect -15672 17688 -15652 17752
rect -16824 17672 -15652 17688
rect -16824 17608 -15736 17672
rect -15672 17608 -15652 17672
rect -16824 17592 -15652 17608
rect -16824 17528 -15736 17592
rect -15672 17528 -15652 17592
rect -16824 17480 -15652 17528
rect -15412 18312 -14240 18360
rect -15412 18248 -14324 18312
rect -14260 18248 -14240 18312
rect -15412 18232 -14240 18248
rect -15412 18168 -14324 18232
rect -14260 18168 -14240 18232
rect -15412 18152 -14240 18168
rect -15412 18088 -14324 18152
rect -14260 18088 -14240 18152
rect -15412 18072 -14240 18088
rect -15412 18008 -14324 18072
rect -14260 18008 -14240 18072
rect -15412 17992 -14240 18008
rect -15412 17928 -14324 17992
rect -14260 17928 -14240 17992
rect -15412 17912 -14240 17928
rect -15412 17848 -14324 17912
rect -14260 17848 -14240 17912
rect -15412 17832 -14240 17848
rect -15412 17768 -14324 17832
rect -14260 17768 -14240 17832
rect -15412 17752 -14240 17768
rect -15412 17688 -14324 17752
rect -14260 17688 -14240 17752
rect -15412 17672 -14240 17688
rect -15412 17608 -14324 17672
rect -14260 17608 -14240 17672
rect -15412 17592 -14240 17608
rect -15412 17528 -14324 17592
rect -14260 17528 -14240 17592
rect -15412 17480 -14240 17528
rect -14000 18312 -12828 18360
rect -14000 18248 -12912 18312
rect -12848 18248 -12828 18312
rect -14000 18232 -12828 18248
rect -14000 18168 -12912 18232
rect -12848 18168 -12828 18232
rect -14000 18152 -12828 18168
rect -14000 18088 -12912 18152
rect -12848 18088 -12828 18152
rect -14000 18072 -12828 18088
rect -14000 18008 -12912 18072
rect -12848 18008 -12828 18072
rect -14000 17992 -12828 18008
rect -14000 17928 -12912 17992
rect -12848 17928 -12828 17992
rect -14000 17912 -12828 17928
rect -14000 17848 -12912 17912
rect -12848 17848 -12828 17912
rect -14000 17832 -12828 17848
rect -14000 17768 -12912 17832
rect -12848 17768 -12828 17832
rect -14000 17752 -12828 17768
rect -14000 17688 -12912 17752
rect -12848 17688 -12828 17752
rect -14000 17672 -12828 17688
rect -14000 17608 -12912 17672
rect -12848 17608 -12828 17672
rect -14000 17592 -12828 17608
rect -14000 17528 -12912 17592
rect -12848 17528 -12828 17592
rect -14000 17480 -12828 17528
rect -12588 18312 -11416 18360
rect -12588 18248 -11500 18312
rect -11436 18248 -11416 18312
rect -12588 18232 -11416 18248
rect -12588 18168 -11500 18232
rect -11436 18168 -11416 18232
rect -12588 18152 -11416 18168
rect -12588 18088 -11500 18152
rect -11436 18088 -11416 18152
rect -12588 18072 -11416 18088
rect -12588 18008 -11500 18072
rect -11436 18008 -11416 18072
rect -12588 17992 -11416 18008
rect -12588 17928 -11500 17992
rect -11436 17928 -11416 17992
rect -12588 17912 -11416 17928
rect -12588 17848 -11500 17912
rect -11436 17848 -11416 17912
rect -12588 17832 -11416 17848
rect -12588 17768 -11500 17832
rect -11436 17768 -11416 17832
rect -12588 17752 -11416 17768
rect -12588 17688 -11500 17752
rect -11436 17688 -11416 17752
rect -12588 17672 -11416 17688
rect -12588 17608 -11500 17672
rect -11436 17608 -11416 17672
rect -12588 17592 -11416 17608
rect -12588 17528 -11500 17592
rect -11436 17528 -11416 17592
rect -12588 17480 -11416 17528
rect -11176 18312 -10004 18360
rect -11176 18248 -10088 18312
rect -10024 18248 -10004 18312
rect -11176 18232 -10004 18248
rect -11176 18168 -10088 18232
rect -10024 18168 -10004 18232
rect -11176 18152 -10004 18168
rect -11176 18088 -10088 18152
rect -10024 18088 -10004 18152
rect -11176 18072 -10004 18088
rect -11176 18008 -10088 18072
rect -10024 18008 -10004 18072
rect -11176 17992 -10004 18008
rect -11176 17928 -10088 17992
rect -10024 17928 -10004 17992
rect -11176 17912 -10004 17928
rect -11176 17848 -10088 17912
rect -10024 17848 -10004 17912
rect -11176 17832 -10004 17848
rect -11176 17768 -10088 17832
rect -10024 17768 -10004 17832
rect -11176 17752 -10004 17768
rect -11176 17688 -10088 17752
rect -10024 17688 -10004 17752
rect -11176 17672 -10004 17688
rect -11176 17608 -10088 17672
rect -10024 17608 -10004 17672
rect -11176 17592 -10004 17608
rect -11176 17528 -10088 17592
rect -10024 17528 -10004 17592
rect -11176 17480 -10004 17528
rect -9764 18312 -8592 18360
rect -9764 18248 -8676 18312
rect -8612 18248 -8592 18312
rect -9764 18232 -8592 18248
rect -9764 18168 -8676 18232
rect -8612 18168 -8592 18232
rect -9764 18152 -8592 18168
rect -9764 18088 -8676 18152
rect -8612 18088 -8592 18152
rect -9764 18072 -8592 18088
rect -9764 18008 -8676 18072
rect -8612 18008 -8592 18072
rect -9764 17992 -8592 18008
rect -9764 17928 -8676 17992
rect -8612 17928 -8592 17992
rect -9764 17912 -8592 17928
rect -9764 17848 -8676 17912
rect -8612 17848 -8592 17912
rect -9764 17832 -8592 17848
rect -9764 17768 -8676 17832
rect -8612 17768 -8592 17832
rect -9764 17752 -8592 17768
rect -9764 17688 -8676 17752
rect -8612 17688 -8592 17752
rect -9764 17672 -8592 17688
rect -9764 17608 -8676 17672
rect -8612 17608 -8592 17672
rect -9764 17592 -8592 17608
rect -9764 17528 -8676 17592
rect -8612 17528 -8592 17592
rect -9764 17480 -8592 17528
rect -8352 18312 -7180 18360
rect -8352 18248 -7264 18312
rect -7200 18248 -7180 18312
rect -8352 18232 -7180 18248
rect -8352 18168 -7264 18232
rect -7200 18168 -7180 18232
rect -8352 18152 -7180 18168
rect -8352 18088 -7264 18152
rect -7200 18088 -7180 18152
rect -8352 18072 -7180 18088
rect -8352 18008 -7264 18072
rect -7200 18008 -7180 18072
rect -8352 17992 -7180 18008
rect -8352 17928 -7264 17992
rect -7200 17928 -7180 17992
rect -8352 17912 -7180 17928
rect -8352 17848 -7264 17912
rect -7200 17848 -7180 17912
rect -8352 17832 -7180 17848
rect -8352 17768 -7264 17832
rect -7200 17768 -7180 17832
rect -8352 17752 -7180 17768
rect -8352 17688 -7264 17752
rect -7200 17688 -7180 17752
rect -8352 17672 -7180 17688
rect -8352 17608 -7264 17672
rect -7200 17608 -7180 17672
rect -8352 17592 -7180 17608
rect -8352 17528 -7264 17592
rect -7200 17528 -7180 17592
rect -8352 17480 -7180 17528
rect -6940 18312 -5768 18360
rect -6940 18248 -5852 18312
rect -5788 18248 -5768 18312
rect -6940 18232 -5768 18248
rect -6940 18168 -5852 18232
rect -5788 18168 -5768 18232
rect -6940 18152 -5768 18168
rect -6940 18088 -5852 18152
rect -5788 18088 -5768 18152
rect -6940 18072 -5768 18088
rect -6940 18008 -5852 18072
rect -5788 18008 -5768 18072
rect -6940 17992 -5768 18008
rect -6940 17928 -5852 17992
rect -5788 17928 -5768 17992
rect -6940 17912 -5768 17928
rect -6940 17848 -5852 17912
rect -5788 17848 -5768 17912
rect -6940 17832 -5768 17848
rect -6940 17768 -5852 17832
rect -5788 17768 -5768 17832
rect -6940 17752 -5768 17768
rect -6940 17688 -5852 17752
rect -5788 17688 -5768 17752
rect -6940 17672 -5768 17688
rect -6940 17608 -5852 17672
rect -5788 17608 -5768 17672
rect -6940 17592 -5768 17608
rect -6940 17528 -5852 17592
rect -5788 17528 -5768 17592
rect -6940 17480 -5768 17528
rect -5528 18312 -4356 18360
rect -5528 18248 -4440 18312
rect -4376 18248 -4356 18312
rect -5528 18232 -4356 18248
rect -5528 18168 -4440 18232
rect -4376 18168 -4356 18232
rect -5528 18152 -4356 18168
rect -5528 18088 -4440 18152
rect -4376 18088 -4356 18152
rect -5528 18072 -4356 18088
rect -5528 18008 -4440 18072
rect -4376 18008 -4356 18072
rect -5528 17992 -4356 18008
rect -5528 17928 -4440 17992
rect -4376 17928 -4356 17992
rect -5528 17912 -4356 17928
rect -5528 17848 -4440 17912
rect -4376 17848 -4356 17912
rect -5528 17832 -4356 17848
rect -5528 17768 -4440 17832
rect -4376 17768 -4356 17832
rect -5528 17752 -4356 17768
rect -5528 17688 -4440 17752
rect -4376 17688 -4356 17752
rect -5528 17672 -4356 17688
rect -5528 17608 -4440 17672
rect -4376 17608 -4356 17672
rect -5528 17592 -4356 17608
rect -5528 17528 -4440 17592
rect -4376 17528 -4356 17592
rect -5528 17480 -4356 17528
rect -4116 18312 -2944 18360
rect -4116 18248 -3028 18312
rect -2964 18248 -2944 18312
rect -4116 18232 -2944 18248
rect -4116 18168 -3028 18232
rect -2964 18168 -2944 18232
rect -4116 18152 -2944 18168
rect -4116 18088 -3028 18152
rect -2964 18088 -2944 18152
rect -4116 18072 -2944 18088
rect -4116 18008 -3028 18072
rect -2964 18008 -2944 18072
rect -4116 17992 -2944 18008
rect -4116 17928 -3028 17992
rect -2964 17928 -2944 17992
rect -4116 17912 -2944 17928
rect -4116 17848 -3028 17912
rect -2964 17848 -2944 17912
rect -4116 17832 -2944 17848
rect -4116 17768 -3028 17832
rect -2964 17768 -2944 17832
rect -4116 17752 -2944 17768
rect -4116 17688 -3028 17752
rect -2964 17688 -2944 17752
rect -4116 17672 -2944 17688
rect -4116 17608 -3028 17672
rect -2964 17608 -2944 17672
rect -4116 17592 -2944 17608
rect -4116 17528 -3028 17592
rect -2964 17528 -2944 17592
rect -4116 17480 -2944 17528
rect -2704 18312 -1532 18360
rect -2704 18248 -1616 18312
rect -1552 18248 -1532 18312
rect -2704 18232 -1532 18248
rect -2704 18168 -1616 18232
rect -1552 18168 -1532 18232
rect -2704 18152 -1532 18168
rect -2704 18088 -1616 18152
rect -1552 18088 -1532 18152
rect -2704 18072 -1532 18088
rect -2704 18008 -1616 18072
rect -1552 18008 -1532 18072
rect -2704 17992 -1532 18008
rect -2704 17928 -1616 17992
rect -1552 17928 -1532 17992
rect -2704 17912 -1532 17928
rect -2704 17848 -1616 17912
rect -1552 17848 -1532 17912
rect -2704 17832 -1532 17848
rect -2704 17768 -1616 17832
rect -1552 17768 -1532 17832
rect -2704 17752 -1532 17768
rect -2704 17688 -1616 17752
rect -1552 17688 -1532 17752
rect -2704 17672 -1532 17688
rect -2704 17608 -1616 17672
rect -1552 17608 -1532 17672
rect -2704 17592 -1532 17608
rect -2704 17528 -1616 17592
rect -1552 17528 -1532 17592
rect -2704 17480 -1532 17528
rect -1292 18312 -120 18360
rect -1292 18248 -204 18312
rect -140 18248 -120 18312
rect -1292 18232 -120 18248
rect -1292 18168 -204 18232
rect -140 18168 -120 18232
rect -1292 18152 -120 18168
rect -1292 18088 -204 18152
rect -140 18088 -120 18152
rect -1292 18072 -120 18088
rect -1292 18008 -204 18072
rect -140 18008 -120 18072
rect -1292 17992 -120 18008
rect -1292 17928 -204 17992
rect -140 17928 -120 17992
rect -1292 17912 -120 17928
rect -1292 17848 -204 17912
rect -140 17848 -120 17912
rect -1292 17832 -120 17848
rect -1292 17768 -204 17832
rect -140 17768 -120 17832
rect -1292 17752 -120 17768
rect -1292 17688 -204 17752
rect -140 17688 -120 17752
rect -1292 17672 -120 17688
rect -1292 17608 -204 17672
rect -140 17608 -120 17672
rect -1292 17592 -120 17608
rect -1292 17528 -204 17592
rect -140 17528 -120 17592
rect -1292 17480 -120 17528
rect 120 18312 1292 18360
rect 120 18248 1208 18312
rect 1272 18248 1292 18312
rect 120 18232 1292 18248
rect 120 18168 1208 18232
rect 1272 18168 1292 18232
rect 120 18152 1292 18168
rect 120 18088 1208 18152
rect 1272 18088 1292 18152
rect 120 18072 1292 18088
rect 120 18008 1208 18072
rect 1272 18008 1292 18072
rect 120 17992 1292 18008
rect 120 17928 1208 17992
rect 1272 17928 1292 17992
rect 120 17912 1292 17928
rect 120 17848 1208 17912
rect 1272 17848 1292 17912
rect 120 17832 1292 17848
rect 120 17768 1208 17832
rect 1272 17768 1292 17832
rect 120 17752 1292 17768
rect 120 17688 1208 17752
rect 1272 17688 1292 17752
rect 120 17672 1292 17688
rect 120 17608 1208 17672
rect 1272 17608 1292 17672
rect 120 17592 1292 17608
rect 120 17528 1208 17592
rect 1272 17528 1292 17592
rect 120 17480 1292 17528
rect 1532 18312 2704 18360
rect 1532 18248 2620 18312
rect 2684 18248 2704 18312
rect 1532 18232 2704 18248
rect 1532 18168 2620 18232
rect 2684 18168 2704 18232
rect 1532 18152 2704 18168
rect 1532 18088 2620 18152
rect 2684 18088 2704 18152
rect 1532 18072 2704 18088
rect 1532 18008 2620 18072
rect 2684 18008 2704 18072
rect 1532 17992 2704 18008
rect 1532 17928 2620 17992
rect 2684 17928 2704 17992
rect 1532 17912 2704 17928
rect 1532 17848 2620 17912
rect 2684 17848 2704 17912
rect 1532 17832 2704 17848
rect 1532 17768 2620 17832
rect 2684 17768 2704 17832
rect 1532 17752 2704 17768
rect 1532 17688 2620 17752
rect 2684 17688 2704 17752
rect 1532 17672 2704 17688
rect 1532 17608 2620 17672
rect 2684 17608 2704 17672
rect 1532 17592 2704 17608
rect 1532 17528 2620 17592
rect 2684 17528 2704 17592
rect 1532 17480 2704 17528
rect 2944 18312 4116 18360
rect 2944 18248 4032 18312
rect 4096 18248 4116 18312
rect 2944 18232 4116 18248
rect 2944 18168 4032 18232
rect 4096 18168 4116 18232
rect 2944 18152 4116 18168
rect 2944 18088 4032 18152
rect 4096 18088 4116 18152
rect 2944 18072 4116 18088
rect 2944 18008 4032 18072
rect 4096 18008 4116 18072
rect 2944 17992 4116 18008
rect 2944 17928 4032 17992
rect 4096 17928 4116 17992
rect 2944 17912 4116 17928
rect 2944 17848 4032 17912
rect 4096 17848 4116 17912
rect 2944 17832 4116 17848
rect 2944 17768 4032 17832
rect 4096 17768 4116 17832
rect 2944 17752 4116 17768
rect 2944 17688 4032 17752
rect 4096 17688 4116 17752
rect 2944 17672 4116 17688
rect 2944 17608 4032 17672
rect 4096 17608 4116 17672
rect 2944 17592 4116 17608
rect 2944 17528 4032 17592
rect 4096 17528 4116 17592
rect 2944 17480 4116 17528
rect 4356 18312 5528 18360
rect 4356 18248 5444 18312
rect 5508 18248 5528 18312
rect 4356 18232 5528 18248
rect 4356 18168 5444 18232
rect 5508 18168 5528 18232
rect 4356 18152 5528 18168
rect 4356 18088 5444 18152
rect 5508 18088 5528 18152
rect 4356 18072 5528 18088
rect 4356 18008 5444 18072
rect 5508 18008 5528 18072
rect 4356 17992 5528 18008
rect 4356 17928 5444 17992
rect 5508 17928 5528 17992
rect 4356 17912 5528 17928
rect 4356 17848 5444 17912
rect 5508 17848 5528 17912
rect 4356 17832 5528 17848
rect 4356 17768 5444 17832
rect 5508 17768 5528 17832
rect 4356 17752 5528 17768
rect 4356 17688 5444 17752
rect 5508 17688 5528 17752
rect 4356 17672 5528 17688
rect 4356 17608 5444 17672
rect 5508 17608 5528 17672
rect 4356 17592 5528 17608
rect 4356 17528 5444 17592
rect 5508 17528 5528 17592
rect 4356 17480 5528 17528
rect 5768 18312 6940 18360
rect 5768 18248 6856 18312
rect 6920 18248 6940 18312
rect 5768 18232 6940 18248
rect 5768 18168 6856 18232
rect 6920 18168 6940 18232
rect 5768 18152 6940 18168
rect 5768 18088 6856 18152
rect 6920 18088 6940 18152
rect 5768 18072 6940 18088
rect 5768 18008 6856 18072
rect 6920 18008 6940 18072
rect 5768 17992 6940 18008
rect 5768 17928 6856 17992
rect 6920 17928 6940 17992
rect 5768 17912 6940 17928
rect 5768 17848 6856 17912
rect 6920 17848 6940 17912
rect 5768 17832 6940 17848
rect 5768 17768 6856 17832
rect 6920 17768 6940 17832
rect 5768 17752 6940 17768
rect 5768 17688 6856 17752
rect 6920 17688 6940 17752
rect 5768 17672 6940 17688
rect 5768 17608 6856 17672
rect 6920 17608 6940 17672
rect 5768 17592 6940 17608
rect 5768 17528 6856 17592
rect 6920 17528 6940 17592
rect 5768 17480 6940 17528
rect 7180 18312 8352 18360
rect 7180 18248 8268 18312
rect 8332 18248 8352 18312
rect 7180 18232 8352 18248
rect 7180 18168 8268 18232
rect 8332 18168 8352 18232
rect 7180 18152 8352 18168
rect 7180 18088 8268 18152
rect 8332 18088 8352 18152
rect 7180 18072 8352 18088
rect 7180 18008 8268 18072
rect 8332 18008 8352 18072
rect 7180 17992 8352 18008
rect 7180 17928 8268 17992
rect 8332 17928 8352 17992
rect 7180 17912 8352 17928
rect 7180 17848 8268 17912
rect 8332 17848 8352 17912
rect 7180 17832 8352 17848
rect 7180 17768 8268 17832
rect 8332 17768 8352 17832
rect 7180 17752 8352 17768
rect 7180 17688 8268 17752
rect 8332 17688 8352 17752
rect 7180 17672 8352 17688
rect 7180 17608 8268 17672
rect 8332 17608 8352 17672
rect 7180 17592 8352 17608
rect 7180 17528 8268 17592
rect 8332 17528 8352 17592
rect 7180 17480 8352 17528
rect 8592 18312 9764 18360
rect 8592 18248 9680 18312
rect 9744 18248 9764 18312
rect 8592 18232 9764 18248
rect 8592 18168 9680 18232
rect 9744 18168 9764 18232
rect 8592 18152 9764 18168
rect 8592 18088 9680 18152
rect 9744 18088 9764 18152
rect 8592 18072 9764 18088
rect 8592 18008 9680 18072
rect 9744 18008 9764 18072
rect 8592 17992 9764 18008
rect 8592 17928 9680 17992
rect 9744 17928 9764 17992
rect 8592 17912 9764 17928
rect 8592 17848 9680 17912
rect 9744 17848 9764 17912
rect 8592 17832 9764 17848
rect 8592 17768 9680 17832
rect 9744 17768 9764 17832
rect 8592 17752 9764 17768
rect 8592 17688 9680 17752
rect 9744 17688 9764 17752
rect 8592 17672 9764 17688
rect 8592 17608 9680 17672
rect 9744 17608 9764 17672
rect 8592 17592 9764 17608
rect 8592 17528 9680 17592
rect 9744 17528 9764 17592
rect 8592 17480 9764 17528
rect 10004 18312 11176 18360
rect 10004 18248 11092 18312
rect 11156 18248 11176 18312
rect 10004 18232 11176 18248
rect 10004 18168 11092 18232
rect 11156 18168 11176 18232
rect 10004 18152 11176 18168
rect 10004 18088 11092 18152
rect 11156 18088 11176 18152
rect 10004 18072 11176 18088
rect 10004 18008 11092 18072
rect 11156 18008 11176 18072
rect 10004 17992 11176 18008
rect 10004 17928 11092 17992
rect 11156 17928 11176 17992
rect 10004 17912 11176 17928
rect 10004 17848 11092 17912
rect 11156 17848 11176 17912
rect 10004 17832 11176 17848
rect 10004 17768 11092 17832
rect 11156 17768 11176 17832
rect 10004 17752 11176 17768
rect 10004 17688 11092 17752
rect 11156 17688 11176 17752
rect 10004 17672 11176 17688
rect 10004 17608 11092 17672
rect 11156 17608 11176 17672
rect 10004 17592 11176 17608
rect 10004 17528 11092 17592
rect 11156 17528 11176 17592
rect 10004 17480 11176 17528
rect 11416 18312 12588 18360
rect 11416 18248 12504 18312
rect 12568 18248 12588 18312
rect 11416 18232 12588 18248
rect 11416 18168 12504 18232
rect 12568 18168 12588 18232
rect 11416 18152 12588 18168
rect 11416 18088 12504 18152
rect 12568 18088 12588 18152
rect 11416 18072 12588 18088
rect 11416 18008 12504 18072
rect 12568 18008 12588 18072
rect 11416 17992 12588 18008
rect 11416 17928 12504 17992
rect 12568 17928 12588 17992
rect 11416 17912 12588 17928
rect 11416 17848 12504 17912
rect 12568 17848 12588 17912
rect 11416 17832 12588 17848
rect 11416 17768 12504 17832
rect 12568 17768 12588 17832
rect 11416 17752 12588 17768
rect 11416 17688 12504 17752
rect 12568 17688 12588 17752
rect 11416 17672 12588 17688
rect 11416 17608 12504 17672
rect 12568 17608 12588 17672
rect 11416 17592 12588 17608
rect 11416 17528 12504 17592
rect 12568 17528 12588 17592
rect 11416 17480 12588 17528
rect 12828 18312 14000 18360
rect 12828 18248 13916 18312
rect 13980 18248 14000 18312
rect 12828 18232 14000 18248
rect 12828 18168 13916 18232
rect 13980 18168 14000 18232
rect 12828 18152 14000 18168
rect 12828 18088 13916 18152
rect 13980 18088 14000 18152
rect 12828 18072 14000 18088
rect 12828 18008 13916 18072
rect 13980 18008 14000 18072
rect 12828 17992 14000 18008
rect 12828 17928 13916 17992
rect 13980 17928 14000 17992
rect 12828 17912 14000 17928
rect 12828 17848 13916 17912
rect 13980 17848 14000 17912
rect 12828 17832 14000 17848
rect 12828 17768 13916 17832
rect 13980 17768 14000 17832
rect 12828 17752 14000 17768
rect 12828 17688 13916 17752
rect 13980 17688 14000 17752
rect 12828 17672 14000 17688
rect 12828 17608 13916 17672
rect 13980 17608 14000 17672
rect 12828 17592 14000 17608
rect 12828 17528 13916 17592
rect 13980 17528 14000 17592
rect 12828 17480 14000 17528
rect 14240 18312 15412 18360
rect 14240 18248 15328 18312
rect 15392 18248 15412 18312
rect 14240 18232 15412 18248
rect 14240 18168 15328 18232
rect 15392 18168 15412 18232
rect 14240 18152 15412 18168
rect 14240 18088 15328 18152
rect 15392 18088 15412 18152
rect 14240 18072 15412 18088
rect 14240 18008 15328 18072
rect 15392 18008 15412 18072
rect 14240 17992 15412 18008
rect 14240 17928 15328 17992
rect 15392 17928 15412 17992
rect 14240 17912 15412 17928
rect 14240 17848 15328 17912
rect 15392 17848 15412 17912
rect 14240 17832 15412 17848
rect 14240 17768 15328 17832
rect 15392 17768 15412 17832
rect 14240 17752 15412 17768
rect 14240 17688 15328 17752
rect 15392 17688 15412 17752
rect 14240 17672 15412 17688
rect 14240 17608 15328 17672
rect 15392 17608 15412 17672
rect 14240 17592 15412 17608
rect 14240 17528 15328 17592
rect 15392 17528 15412 17592
rect 14240 17480 15412 17528
rect 15652 18312 16824 18360
rect 15652 18248 16740 18312
rect 16804 18248 16824 18312
rect 15652 18232 16824 18248
rect 15652 18168 16740 18232
rect 16804 18168 16824 18232
rect 15652 18152 16824 18168
rect 15652 18088 16740 18152
rect 16804 18088 16824 18152
rect 15652 18072 16824 18088
rect 15652 18008 16740 18072
rect 16804 18008 16824 18072
rect 15652 17992 16824 18008
rect 15652 17928 16740 17992
rect 16804 17928 16824 17992
rect 15652 17912 16824 17928
rect 15652 17848 16740 17912
rect 16804 17848 16824 17912
rect 15652 17832 16824 17848
rect 15652 17768 16740 17832
rect 16804 17768 16824 17832
rect 15652 17752 16824 17768
rect 15652 17688 16740 17752
rect 16804 17688 16824 17752
rect 15652 17672 16824 17688
rect 15652 17608 16740 17672
rect 16804 17608 16824 17672
rect 15652 17592 16824 17608
rect 15652 17528 16740 17592
rect 16804 17528 16824 17592
rect 15652 17480 16824 17528
rect 17064 18312 18236 18360
rect 17064 18248 18152 18312
rect 18216 18248 18236 18312
rect 17064 18232 18236 18248
rect 17064 18168 18152 18232
rect 18216 18168 18236 18232
rect 17064 18152 18236 18168
rect 17064 18088 18152 18152
rect 18216 18088 18236 18152
rect 17064 18072 18236 18088
rect 17064 18008 18152 18072
rect 18216 18008 18236 18072
rect 17064 17992 18236 18008
rect 17064 17928 18152 17992
rect 18216 17928 18236 17992
rect 17064 17912 18236 17928
rect 17064 17848 18152 17912
rect 18216 17848 18236 17912
rect 17064 17832 18236 17848
rect 17064 17768 18152 17832
rect 18216 17768 18236 17832
rect 17064 17752 18236 17768
rect 17064 17688 18152 17752
rect 18216 17688 18236 17752
rect 17064 17672 18236 17688
rect 17064 17608 18152 17672
rect 18216 17608 18236 17672
rect 17064 17592 18236 17608
rect 17064 17528 18152 17592
rect 18216 17528 18236 17592
rect 17064 17480 18236 17528
rect 18476 18312 19648 18360
rect 18476 18248 19564 18312
rect 19628 18248 19648 18312
rect 18476 18232 19648 18248
rect 18476 18168 19564 18232
rect 19628 18168 19648 18232
rect 18476 18152 19648 18168
rect 18476 18088 19564 18152
rect 19628 18088 19648 18152
rect 18476 18072 19648 18088
rect 18476 18008 19564 18072
rect 19628 18008 19648 18072
rect 18476 17992 19648 18008
rect 18476 17928 19564 17992
rect 19628 17928 19648 17992
rect 18476 17912 19648 17928
rect 18476 17848 19564 17912
rect 19628 17848 19648 17912
rect 18476 17832 19648 17848
rect 18476 17768 19564 17832
rect 19628 17768 19648 17832
rect 18476 17752 19648 17768
rect 18476 17688 19564 17752
rect 19628 17688 19648 17752
rect 18476 17672 19648 17688
rect 18476 17608 19564 17672
rect 19628 17608 19648 17672
rect 18476 17592 19648 17608
rect 18476 17528 19564 17592
rect 19628 17528 19648 17592
rect 18476 17480 19648 17528
rect 19888 18312 21060 18360
rect 19888 18248 20976 18312
rect 21040 18248 21060 18312
rect 19888 18232 21060 18248
rect 19888 18168 20976 18232
rect 21040 18168 21060 18232
rect 19888 18152 21060 18168
rect 19888 18088 20976 18152
rect 21040 18088 21060 18152
rect 19888 18072 21060 18088
rect 19888 18008 20976 18072
rect 21040 18008 21060 18072
rect 19888 17992 21060 18008
rect 19888 17928 20976 17992
rect 21040 17928 21060 17992
rect 19888 17912 21060 17928
rect 19888 17848 20976 17912
rect 21040 17848 21060 17912
rect 19888 17832 21060 17848
rect 19888 17768 20976 17832
rect 21040 17768 21060 17832
rect 19888 17752 21060 17768
rect 19888 17688 20976 17752
rect 21040 17688 21060 17752
rect 19888 17672 21060 17688
rect 19888 17608 20976 17672
rect 21040 17608 21060 17672
rect 19888 17592 21060 17608
rect 19888 17528 20976 17592
rect 21040 17528 21060 17592
rect 19888 17480 21060 17528
rect 21300 18312 22472 18360
rect 21300 18248 22388 18312
rect 22452 18248 22472 18312
rect 21300 18232 22472 18248
rect 21300 18168 22388 18232
rect 22452 18168 22472 18232
rect 21300 18152 22472 18168
rect 21300 18088 22388 18152
rect 22452 18088 22472 18152
rect 21300 18072 22472 18088
rect 21300 18008 22388 18072
rect 22452 18008 22472 18072
rect 21300 17992 22472 18008
rect 21300 17928 22388 17992
rect 22452 17928 22472 17992
rect 21300 17912 22472 17928
rect 21300 17848 22388 17912
rect 22452 17848 22472 17912
rect 21300 17832 22472 17848
rect 21300 17768 22388 17832
rect 22452 17768 22472 17832
rect 21300 17752 22472 17768
rect 21300 17688 22388 17752
rect 22452 17688 22472 17752
rect 21300 17672 22472 17688
rect 21300 17608 22388 17672
rect 22452 17608 22472 17672
rect 21300 17592 22472 17608
rect 21300 17528 22388 17592
rect 22452 17528 22472 17592
rect 21300 17480 22472 17528
rect 22712 18312 23884 18360
rect 22712 18248 23800 18312
rect 23864 18248 23884 18312
rect 22712 18232 23884 18248
rect 22712 18168 23800 18232
rect 23864 18168 23884 18232
rect 22712 18152 23884 18168
rect 22712 18088 23800 18152
rect 23864 18088 23884 18152
rect 22712 18072 23884 18088
rect 22712 18008 23800 18072
rect 23864 18008 23884 18072
rect 22712 17992 23884 18008
rect 22712 17928 23800 17992
rect 23864 17928 23884 17992
rect 22712 17912 23884 17928
rect 22712 17848 23800 17912
rect 23864 17848 23884 17912
rect 22712 17832 23884 17848
rect 22712 17768 23800 17832
rect 23864 17768 23884 17832
rect 22712 17752 23884 17768
rect 22712 17688 23800 17752
rect 23864 17688 23884 17752
rect 22712 17672 23884 17688
rect 22712 17608 23800 17672
rect 23864 17608 23884 17672
rect 22712 17592 23884 17608
rect 22712 17528 23800 17592
rect 23864 17528 23884 17592
rect 22712 17480 23884 17528
rect -23884 17192 -22712 17240
rect -23884 17128 -22796 17192
rect -22732 17128 -22712 17192
rect -23884 17112 -22712 17128
rect -23884 17048 -22796 17112
rect -22732 17048 -22712 17112
rect -23884 17032 -22712 17048
rect -23884 16968 -22796 17032
rect -22732 16968 -22712 17032
rect -23884 16952 -22712 16968
rect -23884 16888 -22796 16952
rect -22732 16888 -22712 16952
rect -23884 16872 -22712 16888
rect -23884 16808 -22796 16872
rect -22732 16808 -22712 16872
rect -23884 16792 -22712 16808
rect -23884 16728 -22796 16792
rect -22732 16728 -22712 16792
rect -23884 16712 -22712 16728
rect -23884 16648 -22796 16712
rect -22732 16648 -22712 16712
rect -23884 16632 -22712 16648
rect -23884 16568 -22796 16632
rect -22732 16568 -22712 16632
rect -23884 16552 -22712 16568
rect -23884 16488 -22796 16552
rect -22732 16488 -22712 16552
rect -23884 16472 -22712 16488
rect -23884 16408 -22796 16472
rect -22732 16408 -22712 16472
rect -23884 16360 -22712 16408
rect -22472 17192 -21300 17240
rect -22472 17128 -21384 17192
rect -21320 17128 -21300 17192
rect -22472 17112 -21300 17128
rect -22472 17048 -21384 17112
rect -21320 17048 -21300 17112
rect -22472 17032 -21300 17048
rect -22472 16968 -21384 17032
rect -21320 16968 -21300 17032
rect -22472 16952 -21300 16968
rect -22472 16888 -21384 16952
rect -21320 16888 -21300 16952
rect -22472 16872 -21300 16888
rect -22472 16808 -21384 16872
rect -21320 16808 -21300 16872
rect -22472 16792 -21300 16808
rect -22472 16728 -21384 16792
rect -21320 16728 -21300 16792
rect -22472 16712 -21300 16728
rect -22472 16648 -21384 16712
rect -21320 16648 -21300 16712
rect -22472 16632 -21300 16648
rect -22472 16568 -21384 16632
rect -21320 16568 -21300 16632
rect -22472 16552 -21300 16568
rect -22472 16488 -21384 16552
rect -21320 16488 -21300 16552
rect -22472 16472 -21300 16488
rect -22472 16408 -21384 16472
rect -21320 16408 -21300 16472
rect -22472 16360 -21300 16408
rect -21060 17192 -19888 17240
rect -21060 17128 -19972 17192
rect -19908 17128 -19888 17192
rect -21060 17112 -19888 17128
rect -21060 17048 -19972 17112
rect -19908 17048 -19888 17112
rect -21060 17032 -19888 17048
rect -21060 16968 -19972 17032
rect -19908 16968 -19888 17032
rect -21060 16952 -19888 16968
rect -21060 16888 -19972 16952
rect -19908 16888 -19888 16952
rect -21060 16872 -19888 16888
rect -21060 16808 -19972 16872
rect -19908 16808 -19888 16872
rect -21060 16792 -19888 16808
rect -21060 16728 -19972 16792
rect -19908 16728 -19888 16792
rect -21060 16712 -19888 16728
rect -21060 16648 -19972 16712
rect -19908 16648 -19888 16712
rect -21060 16632 -19888 16648
rect -21060 16568 -19972 16632
rect -19908 16568 -19888 16632
rect -21060 16552 -19888 16568
rect -21060 16488 -19972 16552
rect -19908 16488 -19888 16552
rect -21060 16472 -19888 16488
rect -21060 16408 -19972 16472
rect -19908 16408 -19888 16472
rect -21060 16360 -19888 16408
rect -19648 17192 -18476 17240
rect -19648 17128 -18560 17192
rect -18496 17128 -18476 17192
rect -19648 17112 -18476 17128
rect -19648 17048 -18560 17112
rect -18496 17048 -18476 17112
rect -19648 17032 -18476 17048
rect -19648 16968 -18560 17032
rect -18496 16968 -18476 17032
rect -19648 16952 -18476 16968
rect -19648 16888 -18560 16952
rect -18496 16888 -18476 16952
rect -19648 16872 -18476 16888
rect -19648 16808 -18560 16872
rect -18496 16808 -18476 16872
rect -19648 16792 -18476 16808
rect -19648 16728 -18560 16792
rect -18496 16728 -18476 16792
rect -19648 16712 -18476 16728
rect -19648 16648 -18560 16712
rect -18496 16648 -18476 16712
rect -19648 16632 -18476 16648
rect -19648 16568 -18560 16632
rect -18496 16568 -18476 16632
rect -19648 16552 -18476 16568
rect -19648 16488 -18560 16552
rect -18496 16488 -18476 16552
rect -19648 16472 -18476 16488
rect -19648 16408 -18560 16472
rect -18496 16408 -18476 16472
rect -19648 16360 -18476 16408
rect -18236 17192 -17064 17240
rect -18236 17128 -17148 17192
rect -17084 17128 -17064 17192
rect -18236 17112 -17064 17128
rect -18236 17048 -17148 17112
rect -17084 17048 -17064 17112
rect -18236 17032 -17064 17048
rect -18236 16968 -17148 17032
rect -17084 16968 -17064 17032
rect -18236 16952 -17064 16968
rect -18236 16888 -17148 16952
rect -17084 16888 -17064 16952
rect -18236 16872 -17064 16888
rect -18236 16808 -17148 16872
rect -17084 16808 -17064 16872
rect -18236 16792 -17064 16808
rect -18236 16728 -17148 16792
rect -17084 16728 -17064 16792
rect -18236 16712 -17064 16728
rect -18236 16648 -17148 16712
rect -17084 16648 -17064 16712
rect -18236 16632 -17064 16648
rect -18236 16568 -17148 16632
rect -17084 16568 -17064 16632
rect -18236 16552 -17064 16568
rect -18236 16488 -17148 16552
rect -17084 16488 -17064 16552
rect -18236 16472 -17064 16488
rect -18236 16408 -17148 16472
rect -17084 16408 -17064 16472
rect -18236 16360 -17064 16408
rect -16824 17192 -15652 17240
rect -16824 17128 -15736 17192
rect -15672 17128 -15652 17192
rect -16824 17112 -15652 17128
rect -16824 17048 -15736 17112
rect -15672 17048 -15652 17112
rect -16824 17032 -15652 17048
rect -16824 16968 -15736 17032
rect -15672 16968 -15652 17032
rect -16824 16952 -15652 16968
rect -16824 16888 -15736 16952
rect -15672 16888 -15652 16952
rect -16824 16872 -15652 16888
rect -16824 16808 -15736 16872
rect -15672 16808 -15652 16872
rect -16824 16792 -15652 16808
rect -16824 16728 -15736 16792
rect -15672 16728 -15652 16792
rect -16824 16712 -15652 16728
rect -16824 16648 -15736 16712
rect -15672 16648 -15652 16712
rect -16824 16632 -15652 16648
rect -16824 16568 -15736 16632
rect -15672 16568 -15652 16632
rect -16824 16552 -15652 16568
rect -16824 16488 -15736 16552
rect -15672 16488 -15652 16552
rect -16824 16472 -15652 16488
rect -16824 16408 -15736 16472
rect -15672 16408 -15652 16472
rect -16824 16360 -15652 16408
rect -15412 17192 -14240 17240
rect -15412 17128 -14324 17192
rect -14260 17128 -14240 17192
rect -15412 17112 -14240 17128
rect -15412 17048 -14324 17112
rect -14260 17048 -14240 17112
rect -15412 17032 -14240 17048
rect -15412 16968 -14324 17032
rect -14260 16968 -14240 17032
rect -15412 16952 -14240 16968
rect -15412 16888 -14324 16952
rect -14260 16888 -14240 16952
rect -15412 16872 -14240 16888
rect -15412 16808 -14324 16872
rect -14260 16808 -14240 16872
rect -15412 16792 -14240 16808
rect -15412 16728 -14324 16792
rect -14260 16728 -14240 16792
rect -15412 16712 -14240 16728
rect -15412 16648 -14324 16712
rect -14260 16648 -14240 16712
rect -15412 16632 -14240 16648
rect -15412 16568 -14324 16632
rect -14260 16568 -14240 16632
rect -15412 16552 -14240 16568
rect -15412 16488 -14324 16552
rect -14260 16488 -14240 16552
rect -15412 16472 -14240 16488
rect -15412 16408 -14324 16472
rect -14260 16408 -14240 16472
rect -15412 16360 -14240 16408
rect -14000 17192 -12828 17240
rect -14000 17128 -12912 17192
rect -12848 17128 -12828 17192
rect -14000 17112 -12828 17128
rect -14000 17048 -12912 17112
rect -12848 17048 -12828 17112
rect -14000 17032 -12828 17048
rect -14000 16968 -12912 17032
rect -12848 16968 -12828 17032
rect -14000 16952 -12828 16968
rect -14000 16888 -12912 16952
rect -12848 16888 -12828 16952
rect -14000 16872 -12828 16888
rect -14000 16808 -12912 16872
rect -12848 16808 -12828 16872
rect -14000 16792 -12828 16808
rect -14000 16728 -12912 16792
rect -12848 16728 -12828 16792
rect -14000 16712 -12828 16728
rect -14000 16648 -12912 16712
rect -12848 16648 -12828 16712
rect -14000 16632 -12828 16648
rect -14000 16568 -12912 16632
rect -12848 16568 -12828 16632
rect -14000 16552 -12828 16568
rect -14000 16488 -12912 16552
rect -12848 16488 -12828 16552
rect -14000 16472 -12828 16488
rect -14000 16408 -12912 16472
rect -12848 16408 -12828 16472
rect -14000 16360 -12828 16408
rect -12588 17192 -11416 17240
rect -12588 17128 -11500 17192
rect -11436 17128 -11416 17192
rect -12588 17112 -11416 17128
rect -12588 17048 -11500 17112
rect -11436 17048 -11416 17112
rect -12588 17032 -11416 17048
rect -12588 16968 -11500 17032
rect -11436 16968 -11416 17032
rect -12588 16952 -11416 16968
rect -12588 16888 -11500 16952
rect -11436 16888 -11416 16952
rect -12588 16872 -11416 16888
rect -12588 16808 -11500 16872
rect -11436 16808 -11416 16872
rect -12588 16792 -11416 16808
rect -12588 16728 -11500 16792
rect -11436 16728 -11416 16792
rect -12588 16712 -11416 16728
rect -12588 16648 -11500 16712
rect -11436 16648 -11416 16712
rect -12588 16632 -11416 16648
rect -12588 16568 -11500 16632
rect -11436 16568 -11416 16632
rect -12588 16552 -11416 16568
rect -12588 16488 -11500 16552
rect -11436 16488 -11416 16552
rect -12588 16472 -11416 16488
rect -12588 16408 -11500 16472
rect -11436 16408 -11416 16472
rect -12588 16360 -11416 16408
rect -11176 17192 -10004 17240
rect -11176 17128 -10088 17192
rect -10024 17128 -10004 17192
rect -11176 17112 -10004 17128
rect -11176 17048 -10088 17112
rect -10024 17048 -10004 17112
rect -11176 17032 -10004 17048
rect -11176 16968 -10088 17032
rect -10024 16968 -10004 17032
rect -11176 16952 -10004 16968
rect -11176 16888 -10088 16952
rect -10024 16888 -10004 16952
rect -11176 16872 -10004 16888
rect -11176 16808 -10088 16872
rect -10024 16808 -10004 16872
rect -11176 16792 -10004 16808
rect -11176 16728 -10088 16792
rect -10024 16728 -10004 16792
rect -11176 16712 -10004 16728
rect -11176 16648 -10088 16712
rect -10024 16648 -10004 16712
rect -11176 16632 -10004 16648
rect -11176 16568 -10088 16632
rect -10024 16568 -10004 16632
rect -11176 16552 -10004 16568
rect -11176 16488 -10088 16552
rect -10024 16488 -10004 16552
rect -11176 16472 -10004 16488
rect -11176 16408 -10088 16472
rect -10024 16408 -10004 16472
rect -11176 16360 -10004 16408
rect -9764 17192 -8592 17240
rect -9764 17128 -8676 17192
rect -8612 17128 -8592 17192
rect -9764 17112 -8592 17128
rect -9764 17048 -8676 17112
rect -8612 17048 -8592 17112
rect -9764 17032 -8592 17048
rect -9764 16968 -8676 17032
rect -8612 16968 -8592 17032
rect -9764 16952 -8592 16968
rect -9764 16888 -8676 16952
rect -8612 16888 -8592 16952
rect -9764 16872 -8592 16888
rect -9764 16808 -8676 16872
rect -8612 16808 -8592 16872
rect -9764 16792 -8592 16808
rect -9764 16728 -8676 16792
rect -8612 16728 -8592 16792
rect -9764 16712 -8592 16728
rect -9764 16648 -8676 16712
rect -8612 16648 -8592 16712
rect -9764 16632 -8592 16648
rect -9764 16568 -8676 16632
rect -8612 16568 -8592 16632
rect -9764 16552 -8592 16568
rect -9764 16488 -8676 16552
rect -8612 16488 -8592 16552
rect -9764 16472 -8592 16488
rect -9764 16408 -8676 16472
rect -8612 16408 -8592 16472
rect -9764 16360 -8592 16408
rect -8352 17192 -7180 17240
rect -8352 17128 -7264 17192
rect -7200 17128 -7180 17192
rect -8352 17112 -7180 17128
rect -8352 17048 -7264 17112
rect -7200 17048 -7180 17112
rect -8352 17032 -7180 17048
rect -8352 16968 -7264 17032
rect -7200 16968 -7180 17032
rect -8352 16952 -7180 16968
rect -8352 16888 -7264 16952
rect -7200 16888 -7180 16952
rect -8352 16872 -7180 16888
rect -8352 16808 -7264 16872
rect -7200 16808 -7180 16872
rect -8352 16792 -7180 16808
rect -8352 16728 -7264 16792
rect -7200 16728 -7180 16792
rect -8352 16712 -7180 16728
rect -8352 16648 -7264 16712
rect -7200 16648 -7180 16712
rect -8352 16632 -7180 16648
rect -8352 16568 -7264 16632
rect -7200 16568 -7180 16632
rect -8352 16552 -7180 16568
rect -8352 16488 -7264 16552
rect -7200 16488 -7180 16552
rect -8352 16472 -7180 16488
rect -8352 16408 -7264 16472
rect -7200 16408 -7180 16472
rect -8352 16360 -7180 16408
rect -6940 17192 -5768 17240
rect -6940 17128 -5852 17192
rect -5788 17128 -5768 17192
rect -6940 17112 -5768 17128
rect -6940 17048 -5852 17112
rect -5788 17048 -5768 17112
rect -6940 17032 -5768 17048
rect -6940 16968 -5852 17032
rect -5788 16968 -5768 17032
rect -6940 16952 -5768 16968
rect -6940 16888 -5852 16952
rect -5788 16888 -5768 16952
rect -6940 16872 -5768 16888
rect -6940 16808 -5852 16872
rect -5788 16808 -5768 16872
rect -6940 16792 -5768 16808
rect -6940 16728 -5852 16792
rect -5788 16728 -5768 16792
rect -6940 16712 -5768 16728
rect -6940 16648 -5852 16712
rect -5788 16648 -5768 16712
rect -6940 16632 -5768 16648
rect -6940 16568 -5852 16632
rect -5788 16568 -5768 16632
rect -6940 16552 -5768 16568
rect -6940 16488 -5852 16552
rect -5788 16488 -5768 16552
rect -6940 16472 -5768 16488
rect -6940 16408 -5852 16472
rect -5788 16408 -5768 16472
rect -6940 16360 -5768 16408
rect -5528 17192 -4356 17240
rect -5528 17128 -4440 17192
rect -4376 17128 -4356 17192
rect -5528 17112 -4356 17128
rect -5528 17048 -4440 17112
rect -4376 17048 -4356 17112
rect -5528 17032 -4356 17048
rect -5528 16968 -4440 17032
rect -4376 16968 -4356 17032
rect -5528 16952 -4356 16968
rect -5528 16888 -4440 16952
rect -4376 16888 -4356 16952
rect -5528 16872 -4356 16888
rect -5528 16808 -4440 16872
rect -4376 16808 -4356 16872
rect -5528 16792 -4356 16808
rect -5528 16728 -4440 16792
rect -4376 16728 -4356 16792
rect -5528 16712 -4356 16728
rect -5528 16648 -4440 16712
rect -4376 16648 -4356 16712
rect -5528 16632 -4356 16648
rect -5528 16568 -4440 16632
rect -4376 16568 -4356 16632
rect -5528 16552 -4356 16568
rect -5528 16488 -4440 16552
rect -4376 16488 -4356 16552
rect -5528 16472 -4356 16488
rect -5528 16408 -4440 16472
rect -4376 16408 -4356 16472
rect -5528 16360 -4356 16408
rect -4116 17192 -2944 17240
rect -4116 17128 -3028 17192
rect -2964 17128 -2944 17192
rect -4116 17112 -2944 17128
rect -4116 17048 -3028 17112
rect -2964 17048 -2944 17112
rect -4116 17032 -2944 17048
rect -4116 16968 -3028 17032
rect -2964 16968 -2944 17032
rect -4116 16952 -2944 16968
rect -4116 16888 -3028 16952
rect -2964 16888 -2944 16952
rect -4116 16872 -2944 16888
rect -4116 16808 -3028 16872
rect -2964 16808 -2944 16872
rect -4116 16792 -2944 16808
rect -4116 16728 -3028 16792
rect -2964 16728 -2944 16792
rect -4116 16712 -2944 16728
rect -4116 16648 -3028 16712
rect -2964 16648 -2944 16712
rect -4116 16632 -2944 16648
rect -4116 16568 -3028 16632
rect -2964 16568 -2944 16632
rect -4116 16552 -2944 16568
rect -4116 16488 -3028 16552
rect -2964 16488 -2944 16552
rect -4116 16472 -2944 16488
rect -4116 16408 -3028 16472
rect -2964 16408 -2944 16472
rect -4116 16360 -2944 16408
rect -2704 17192 -1532 17240
rect -2704 17128 -1616 17192
rect -1552 17128 -1532 17192
rect -2704 17112 -1532 17128
rect -2704 17048 -1616 17112
rect -1552 17048 -1532 17112
rect -2704 17032 -1532 17048
rect -2704 16968 -1616 17032
rect -1552 16968 -1532 17032
rect -2704 16952 -1532 16968
rect -2704 16888 -1616 16952
rect -1552 16888 -1532 16952
rect -2704 16872 -1532 16888
rect -2704 16808 -1616 16872
rect -1552 16808 -1532 16872
rect -2704 16792 -1532 16808
rect -2704 16728 -1616 16792
rect -1552 16728 -1532 16792
rect -2704 16712 -1532 16728
rect -2704 16648 -1616 16712
rect -1552 16648 -1532 16712
rect -2704 16632 -1532 16648
rect -2704 16568 -1616 16632
rect -1552 16568 -1532 16632
rect -2704 16552 -1532 16568
rect -2704 16488 -1616 16552
rect -1552 16488 -1532 16552
rect -2704 16472 -1532 16488
rect -2704 16408 -1616 16472
rect -1552 16408 -1532 16472
rect -2704 16360 -1532 16408
rect -1292 17192 -120 17240
rect -1292 17128 -204 17192
rect -140 17128 -120 17192
rect -1292 17112 -120 17128
rect -1292 17048 -204 17112
rect -140 17048 -120 17112
rect -1292 17032 -120 17048
rect -1292 16968 -204 17032
rect -140 16968 -120 17032
rect -1292 16952 -120 16968
rect -1292 16888 -204 16952
rect -140 16888 -120 16952
rect -1292 16872 -120 16888
rect -1292 16808 -204 16872
rect -140 16808 -120 16872
rect -1292 16792 -120 16808
rect -1292 16728 -204 16792
rect -140 16728 -120 16792
rect -1292 16712 -120 16728
rect -1292 16648 -204 16712
rect -140 16648 -120 16712
rect -1292 16632 -120 16648
rect -1292 16568 -204 16632
rect -140 16568 -120 16632
rect -1292 16552 -120 16568
rect -1292 16488 -204 16552
rect -140 16488 -120 16552
rect -1292 16472 -120 16488
rect -1292 16408 -204 16472
rect -140 16408 -120 16472
rect -1292 16360 -120 16408
rect 120 17192 1292 17240
rect 120 17128 1208 17192
rect 1272 17128 1292 17192
rect 120 17112 1292 17128
rect 120 17048 1208 17112
rect 1272 17048 1292 17112
rect 120 17032 1292 17048
rect 120 16968 1208 17032
rect 1272 16968 1292 17032
rect 120 16952 1292 16968
rect 120 16888 1208 16952
rect 1272 16888 1292 16952
rect 120 16872 1292 16888
rect 120 16808 1208 16872
rect 1272 16808 1292 16872
rect 120 16792 1292 16808
rect 120 16728 1208 16792
rect 1272 16728 1292 16792
rect 120 16712 1292 16728
rect 120 16648 1208 16712
rect 1272 16648 1292 16712
rect 120 16632 1292 16648
rect 120 16568 1208 16632
rect 1272 16568 1292 16632
rect 120 16552 1292 16568
rect 120 16488 1208 16552
rect 1272 16488 1292 16552
rect 120 16472 1292 16488
rect 120 16408 1208 16472
rect 1272 16408 1292 16472
rect 120 16360 1292 16408
rect 1532 17192 2704 17240
rect 1532 17128 2620 17192
rect 2684 17128 2704 17192
rect 1532 17112 2704 17128
rect 1532 17048 2620 17112
rect 2684 17048 2704 17112
rect 1532 17032 2704 17048
rect 1532 16968 2620 17032
rect 2684 16968 2704 17032
rect 1532 16952 2704 16968
rect 1532 16888 2620 16952
rect 2684 16888 2704 16952
rect 1532 16872 2704 16888
rect 1532 16808 2620 16872
rect 2684 16808 2704 16872
rect 1532 16792 2704 16808
rect 1532 16728 2620 16792
rect 2684 16728 2704 16792
rect 1532 16712 2704 16728
rect 1532 16648 2620 16712
rect 2684 16648 2704 16712
rect 1532 16632 2704 16648
rect 1532 16568 2620 16632
rect 2684 16568 2704 16632
rect 1532 16552 2704 16568
rect 1532 16488 2620 16552
rect 2684 16488 2704 16552
rect 1532 16472 2704 16488
rect 1532 16408 2620 16472
rect 2684 16408 2704 16472
rect 1532 16360 2704 16408
rect 2944 17192 4116 17240
rect 2944 17128 4032 17192
rect 4096 17128 4116 17192
rect 2944 17112 4116 17128
rect 2944 17048 4032 17112
rect 4096 17048 4116 17112
rect 2944 17032 4116 17048
rect 2944 16968 4032 17032
rect 4096 16968 4116 17032
rect 2944 16952 4116 16968
rect 2944 16888 4032 16952
rect 4096 16888 4116 16952
rect 2944 16872 4116 16888
rect 2944 16808 4032 16872
rect 4096 16808 4116 16872
rect 2944 16792 4116 16808
rect 2944 16728 4032 16792
rect 4096 16728 4116 16792
rect 2944 16712 4116 16728
rect 2944 16648 4032 16712
rect 4096 16648 4116 16712
rect 2944 16632 4116 16648
rect 2944 16568 4032 16632
rect 4096 16568 4116 16632
rect 2944 16552 4116 16568
rect 2944 16488 4032 16552
rect 4096 16488 4116 16552
rect 2944 16472 4116 16488
rect 2944 16408 4032 16472
rect 4096 16408 4116 16472
rect 2944 16360 4116 16408
rect 4356 17192 5528 17240
rect 4356 17128 5444 17192
rect 5508 17128 5528 17192
rect 4356 17112 5528 17128
rect 4356 17048 5444 17112
rect 5508 17048 5528 17112
rect 4356 17032 5528 17048
rect 4356 16968 5444 17032
rect 5508 16968 5528 17032
rect 4356 16952 5528 16968
rect 4356 16888 5444 16952
rect 5508 16888 5528 16952
rect 4356 16872 5528 16888
rect 4356 16808 5444 16872
rect 5508 16808 5528 16872
rect 4356 16792 5528 16808
rect 4356 16728 5444 16792
rect 5508 16728 5528 16792
rect 4356 16712 5528 16728
rect 4356 16648 5444 16712
rect 5508 16648 5528 16712
rect 4356 16632 5528 16648
rect 4356 16568 5444 16632
rect 5508 16568 5528 16632
rect 4356 16552 5528 16568
rect 4356 16488 5444 16552
rect 5508 16488 5528 16552
rect 4356 16472 5528 16488
rect 4356 16408 5444 16472
rect 5508 16408 5528 16472
rect 4356 16360 5528 16408
rect 5768 17192 6940 17240
rect 5768 17128 6856 17192
rect 6920 17128 6940 17192
rect 5768 17112 6940 17128
rect 5768 17048 6856 17112
rect 6920 17048 6940 17112
rect 5768 17032 6940 17048
rect 5768 16968 6856 17032
rect 6920 16968 6940 17032
rect 5768 16952 6940 16968
rect 5768 16888 6856 16952
rect 6920 16888 6940 16952
rect 5768 16872 6940 16888
rect 5768 16808 6856 16872
rect 6920 16808 6940 16872
rect 5768 16792 6940 16808
rect 5768 16728 6856 16792
rect 6920 16728 6940 16792
rect 5768 16712 6940 16728
rect 5768 16648 6856 16712
rect 6920 16648 6940 16712
rect 5768 16632 6940 16648
rect 5768 16568 6856 16632
rect 6920 16568 6940 16632
rect 5768 16552 6940 16568
rect 5768 16488 6856 16552
rect 6920 16488 6940 16552
rect 5768 16472 6940 16488
rect 5768 16408 6856 16472
rect 6920 16408 6940 16472
rect 5768 16360 6940 16408
rect 7180 17192 8352 17240
rect 7180 17128 8268 17192
rect 8332 17128 8352 17192
rect 7180 17112 8352 17128
rect 7180 17048 8268 17112
rect 8332 17048 8352 17112
rect 7180 17032 8352 17048
rect 7180 16968 8268 17032
rect 8332 16968 8352 17032
rect 7180 16952 8352 16968
rect 7180 16888 8268 16952
rect 8332 16888 8352 16952
rect 7180 16872 8352 16888
rect 7180 16808 8268 16872
rect 8332 16808 8352 16872
rect 7180 16792 8352 16808
rect 7180 16728 8268 16792
rect 8332 16728 8352 16792
rect 7180 16712 8352 16728
rect 7180 16648 8268 16712
rect 8332 16648 8352 16712
rect 7180 16632 8352 16648
rect 7180 16568 8268 16632
rect 8332 16568 8352 16632
rect 7180 16552 8352 16568
rect 7180 16488 8268 16552
rect 8332 16488 8352 16552
rect 7180 16472 8352 16488
rect 7180 16408 8268 16472
rect 8332 16408 8352 16472
rect 7180 16360 8352 16408
rect 8592 17192 9764 17240
rect 8592 17128 9680 17192
rect 9744 17128 9764 17192
rect 8592 17112 9764 17128
rect 8592 17048 9680 17112
rect 9744 17048 9764 17112
rect 8592 17032 9764 17048
rect 8592 16968 9680 17032
rect 9744 16968 9764 17032
rect 8592 16952 9764 16968
rect 8592 16888 9680 16952
rect 9744 16888 9764 16952
rect 8592 16872 9764 16888
rect 8592 16808 9680 16872
rect 9744 16808 9764 16872
rect 8592 16792 9764 16808
rect 8592 16728 9680 16792
rect 9744 16728 9764 16792
rect 8592 16712 9764 16728
rect 8592 16648 9680 16712
rect 9744 16648 9764 16712
rect 8592 16632 9764 16648
rect 8592 16568 9680 16632
rect 9744 16568 9764 16632
rect 8592 16552 9764 16568
rect 8592 16488 9680 16552
rect 9744 16488 9764 16552
rect 8592 16472 9764 16488
rect 8592 16408 9680 16472
rect 9744 16408 9764 16472
rect 8592 16360 9764 16408
rect 10004 17192 11176 17240
rect 10004 17128 11092 17192
rect 11156 17128 11176 17192
rect 10004 17112 11176 17128
rect 10004 17048 11092 17112
rect 11156 17048 11176 17112
rect 10004 17032 11176 17048
rect 10004 16968 11092 17032
rect 11156 16968 11176 17032
rect 10004 16952 11176 16968
rect 10004 16888 11092 16952
rect 11156 16888 11176 16952
rect 10004 16872 11176 16888
rect 10004 16808 11092 16872
rect 11156 16808 11176 16872
rect 10004 16792 11176 16808
rect 10004 16728 11092 16792
rect 11156 16728 11176 16792
rect 10004 16712 11176 16728
rect 10004 16648 11092 16712
rect 11156 16648 11176 16712
rect 10004 16632 11176 16648
rect 10004 16568 11092 16632
rect 11156 16568 11176 16632
rect 10004 16552 11176 16568
rect 10004 16488 11092 16552
rect 11156 16488 11176 16552
rect 10004 16472 11176 16488
rect 10004 16408 11092 16472
rect 11156 16408 11176 16472
rect 10004 16360 11176 16408
rect 11416 17192 12588 17240
rect 11416 17128 12504 17192
rect 12568 17128 12588 17192
rect 11416 17112 12588 17128
rect 11416 17048 12504 17112
rect 12568 17048 12588 17112
rect 11416 17032 12588 17048
rect 11416 16968 12504 17032
rect 12568 16968 12588 17032
rect 11416 16952 12588 16968
rect 11416 16888 12504 16952
rect 12568 16888 12588 16952
rect 11416 16872 12588 16888
rect 11416 16808 12504 16872
rect 12568 16808 12588 16872
rect 11416 16792 12588 16808
rect 11416 16728 12504 16792
rect 12568 16728 12588 16792
rect 11416 16712 12588 16728
rect 11416 16648 12504 16712
rect 12568 16648 12588 16712
rect 11416 16632 12588 16648
rect 11416 16568 12504 16632
rect 12568 16568 12588 16632
rect 11416 16552 12588 16568
rect 11416 16488 12504 16552
rect 12568 16488 12588 16552
rect 11416 16472 12588 16488
rect 11416 16408 12504 16472
rect 12568 16408 12588 16472
rect 11416 16360 12588 16408
rect 12828 17192 14000 17240
rect 12828 17128 13916 17192
rect 13980 17128 14000 17192
rect 12828 17112 14000 17128
rect 12828 17048 13916 17112
rect 13980 17048 14000 17112
rect 12828 17032 14000 17048
rect 12828 16968 13916 17032
rect 13980 16968 14000 17032
rect 12828 16952 14000 16968
rect 12828 16888 13916 16952
rect 13980 16888 14000 16952
rect 12828 16872 14000 16888
rect 12828 16808 13916 16872
rect 13980 16808 14000 16872
rect 12828 16792 14000 16808
rect 12828 16728 13916 16792
rect 13980 16728 14000 16792
rect 12828 16712 14000 16728
rect 12828 16648 13916 16712
rect 13980 16648 14000 16712
rect 12828 16632 14000 16648
rect 12828 16568 13916 16632
rect 13980 16568 14000 16632
rect 12828 16552 14000 16568
rect 12828 16488 13916 16552
rect 13980 16488 14000 16552
rect 12828 16472 14000 16488
rect 12828 16408 13916 16472
rect 13980 16408 14000 16472
rect 12828 16360 14000 16408
rect 14240 17192 15412 17240
rect 14240 17128 15328 17192
rect 15392 17128 15412 17192
rect 14240 17112 15412 17128
rect 14240 17048 15328 17112
rect 15392 17048 15412 17112
rect 14240 17032 15412 17048
rect 14240 16968 15328 17032
rect 15392 16968 15412 17032
rect 14240 16952 15412 16968
rect 14240 16888 15328 16952
rect 15392 16888 15412 16952
rect 14240 16872 15412 16888
rect 14240 16808 15328 16872
rect 15392 16808 15412 16872
rect 14240 16792 15412 16808
rect 14240 16728 15328 16792
rect 15392 16728 15412 16792
rect 14240 16712 15412 16728
rect 14240 16648 15328 16712
rect 15392 16648 15412 16712
rect 14240 16632 15412 16648
rect 14240 16568 15328 16632
rect 15392 16568 15412 16632
rect 14240 16552 15412 16568
rect 14240 16488 15328 16552
rect 15392 16488 15412 16552
rect 14240 16472 15412 16488
rect 14240 16408 15328 16472
rect 15392 16408 15412 16472
rect 14240 16360 15412 16408
rect 15652 17192 16824 17240
rect 15652 17128 16740 17192
rect 16804 17128 16824 17192
rect 15652 17112 16824 17128
rect 15652 17048 16740 17112
rect 16804 17048 16824 17112
rect 15652 17032 16824 17048
rect 15652 16968 16740 17032
rect 16804 16968 16824 17032
rect 15652 16952 16824 16968
rect 15652 16888 16740 16952
rect 16804 16888 16824 16952
rect 15652 16872 16824 16888
rect 15652 16808 16740 16872
rect 16804 16808 16824 16872
rect 15652 16792 16824 16808
rect 15652 16728 16740 16792
rect 16804 16728 16824 16792
rect 15652 16712 16824 16728
rect 15652 16648 16740 16712
rect 16804 16648 16824 16712
rect 15652 16632 16824 16648
rect 15652 16568 16740 16632
rect 16804 16568 16824 16632
rect 15652 16552 16824 16568
rect 15652 16488 16740 16552
rect 16804 16488 16824 16552
rect 15652 16472 16824 16488
rect 15652 16408 16740 16472
rect 16804 16408 16824 16472
rect 15652 16360 16824 16408
rect 17064 17192 18236 17240
rect 17064 17128 18152 17192
rect 18216 17128 18236 17192
rect 17064 17112 18236 17128
rect 17064 17048 18152 17112
rect 18216 17048 18236 17112
rect 17064 17032 18236 17048
rect 17064 16968 18152 17032
rect 18216 16968 18236 17032
rect 17064 16952 18236 16968
rect 17064 16888 18152 16952
rect 18216 16888 18236 16952
rect 17064 16872 18236 16888
rect 17064 16808 18152 16872
rect 18216 16808 18236 16872
rect 17064 16792 18236 16808
rect 17064 16728 18152 16792
rect 18216 16728 18236 16792
rect 17064 16712 18236 16728
rect 17064 16648 18152 16712
rect 18216 16648 18236 16712
rect 17064 16632 18236 16648
rect 17064 16568 18152 16632
rect 18216 16568 18236 16632
rect 17064 16552 18236 16568
rect 17064 16488 18152 16552
rect 18216 16488 18236 16552
rect 17064 16472 18236 16488
rect 17064 16408 18152 16472
rect 18216 16408 18236 16472
rect 17064 16360 18236 16408
rect 18476 17192 19648 17240
rect 18476 17128 19564 17192
rect 19628 17128 19648 17192
rect 18476 17112 19648 17128
rect 18476 17048 19564 17112
rect 19628 17048 19648 17112
rect 18476 17032 19648 17048
rect 18476 16968 19564 17032
rect 19628 16968 19648 17032
rect 18476 16952 19648 16968
rect 18476 16888 19564 16952
rect 19628 16888 19648 16952
rect 18476 16872 19648 16888
rect 18476 16808 19564 16872
rect 19628 16808 19648 16872
rect 18476 16792 19648 16808
rect 18476 16728 19564 16792
rect 19628 16728 19648 16792
rect 18476 16712 19648 16728
rect 18476 16648 19564 16712
rect 19628 16648 19648 16712
rect 18476 16632 19648 16648
rect 18476 16568 19564 16632
rect 19628 16568 19648 16632
rect 18476 16552 19648 16568
rect 18476 16488 19564 16552
rect 19628 16488 19648 16552
rect 18476 16472 19648 16488
rect 18476 16408 19564 16472
rect 19628 16408 19648 16472
rect 18476 16360 19648 16408
rect 19888 17192 21060 17240
rect 19888 17128 20976 17192
rect 21040 17128 21060 17192
rect 19888 17112 21060 17128
rect 19888 17048 20976 17112
rect 21040 17048 21060 17112
rect 19888 17032 21060 17048
rect 19888 16968 20976 17032
rect 21040 16968 21060 17032
rect 19888 16952 21060 16968
rect 19888 16888 20976 16952
rect 21040 16888 21060 16952
rect 19888 16872 21060 16888
rect 19888 16808 20976 16872
rect 21040 16808 21060 16872
rect 19888 16792 21060 16808
rect 19888 16728 20976 16792
rect 21040 16728 21060 16792
rect 19888 16712 21060 16728
rect 19888 16648 20976 16712
rect 21040 16648 21060 16712
rect 19888 16632 21060 16648
rect 19888 16568 20976 16632
rect 21040 16568 21060 16632
rect 19888 16552 21060 16568
rect 19888 16488 20976 16552
rect 21040 16488 21060 16552
rect 19888 16472 21060 16488
rect 19888 16408 20976 16472
rect 21040 16408 21060 16472
rect 19888 16360 21060 16408
rect 21300 17192 22472 17240
rect 21300 17128 22388 17192
rect 22452 17128 22472 17192
rect 21300 17112 22472 17128
rect 21300 17048 22388 17112
rect 22452 17048 22472 17112
rect 21300 17032 22472 17048
rect 21300 16968 22388 17032
rect 22452 16968 22472 17032
rect 21300 16952 22472 16968
rect 21300 16888 22388 16952
rect 22452 16888 22472 16952
rect 21300 16872 22472 16888
rect 21300 16808 22388 16872
rect 22452 16808 22472 16872
rect 21300 16792 22472 16808
rect 21300 16728 22388 16792
rect 22452 16728 22472 16792
rect 21300 16712 22472 16728
rect 21300 16648 22388 16712
rect 22452 16648 22472 16712
rect 21300 16632 22472 16648
rect 21300 16568 22388 16632
rect 22452 16568 22472 16632
rect 21300 16552 22472 16568
rect 21300 16488 22388 16552
rect 22452 16488 22472 16552
rect 21300 16472 22472 16488
rect 21300 16408 22388 16472
rect 22452 16408 22472 16472
rect 21300 16360 22472 16408
rect 22712 17192 23884 17240
rect 22712 17128 23800 17192
rect 23864 17128 23884 17192
rect 22712 17112 23884 17128
rect 22712 17048 23800 17112
rect 23864 17048 23884 17112
rect 22712 17032 23884 17048
rect 22712 16968 23800 17032
rect 23864 16968 23884 17032
rect 22712 16952 23884 16968
rect 22712 16888 23800 16952
rect 23864 16888 23884 16952
rect 22712 16872 23884 16888
rect 22712 16808 23800 16872
rect 23864 16808 23884 16872
rect 22712 16792 23884 16808
rect 22712 16728 23800 16792
rect 23864 16728 23884 16792
rect 22712 16712 23884 16728
rect 22712 16648 23800 16712
rect 23864 16648 23884 16712
rect 22712 16632 23884 16648
rect 22712 16568 23800 16632
rect 23864 16568 23884 16632
rect 22712 16552 23884 16568
rect 22712 16488 23800 16552
rect 23864 16488 23884 16552
rect 22712 16472 23884 16488
rect 22712 16408 23800 16472
rect 23864 16408 23884 16472
rect 22712 16360 23884 16408
rect -23884 16072 -22712 16120
rect -23884 16008 -22796 16072
rect -22732 16008 -22712 16072
rect -23884 15992 -22712 16008
rect -23884 15928 -22796 15992
rect -22732 15928 -22712 15992
rect -23884 15912 -22712 15928
rect -23884 15848 -22796 15912
rect -22732 15848 -22712 15912
rect -23884 15832 -22712 15848
rect -23884 15768 -22796 15832
rect -22732 15768 -22712 15832
rect -23884 15752 -22712 15768
rect -23884 15688 -22796 15752
rect -22732 15688 -22712 15752
rect -23884 15672 -22712 15688
rect -23884 15608 -22796 15672
rect -22732 15608 -22712 15672
rect -23884 15592 -22712 15608
rect -23884 15528 -22796 15592
rect -22732 15528 -22712 15592
rect -23884 15512 -22712 15528
rect -23884 15448 -22796 15512
rect -22732 15448 -22712 15512
rect -23884 15432 -22712 15448
rect -23884 15368 -22796 15432
rect -22732 15368 -22712 15432
rect -23884 15352 -22712 15368
rect -23884 15288 -22796 15352
rect -22732 15288 -22712 15352
rect -23884 15240 -22712 15288
rect -22472 16072 -21300 16120
rect -22472 16008 -21384 16072
rect -21320 16008 -21300 16072
rect -22472 15992 -21300 16008
rect -22472 15928 -21384 15992
rect -21320 15928 -21300 15992
rect -22472 15912 -21300 15928
rect -22472 15848 -21384 15912
rect -21320 15848 -21300 15912
rect -22472 15832 -21300 15848
rect -22472 15768 -21384 15832
rect -21320 15768 -21300 15832
rect -22472 15752 -21300 15768
rect -22472 15688 -21384 15752
rect -21320 15688 -21300 15752
rect -22472 15672 -21300 15688
rect -22472 15608 -21384 15672
rect -21320 15608 -21300 15672
rect -22472 15592 -21300 15608
rect -22472 15528 -21384 15592
rect -21320 15528 -21300 15592
rect -22472 15512 -21300 15528
rect -22472 15448 -21384 15512
rect -21320 15448 -21300 15512
rect -22472 15432 -21300 15448
rect -22472 15368 -21384 15432
rect -21320 15368 -21300 15432
rect -22472 15352 -21300 15368
rect -22472 15288 -21384 15352
rect -21320 15288 -21300 15352
rect -22472 15240 -21300 15288
rect -21060 16072 -19888 16120
rect -21060 16008 -19972 16072
rect -19908 16008 -19888 16072
rect -21060 15992 -19888 16008
rect -21060 15928 -19972 15992
rect -19908 15928 -19888 15992
rect -21060 15912 -19888 15928
rect -21060 15848 -19972 15912
rect -19908 15848 -19888 15912
rect -21060 15832 -19888 15848
rect -21060 15768 -19972 15832
rect -19908 15768 -19888 15832
rect -21060 15752 -19888 15768
rect -21060 15688 -19972 15752
rect -19908 15688 -19888 15752
rect -21060 15672 -19888 15688
rect -21060 15608 -19972 15672
rect -19908 15608 -19888 15672
rect -21060 15592 -19888 15608
rect -21060 15528 -19972 15592
rect -19908 15528 -19888 15592
rect -21060 15512 -19888 15528
rect -21060 15448 -19972 15512
rect -19908 15448 -19888 15512
rect -21060 15432 -19888 15448
rect -21060 15368 -19972 15432
rect -19908 15368 -19888 15432
rect -21060 15352 -19888 15368
rect -21060 15288 -19972 15352
rect -19908 15288 -19888 15352
rect -21060 15240 -19888 15288
rect -19648 16072 -18476 16120
rect -19648 16008 -18560 16072
rect -18496 16008 -18476 16072
rect -19648 15992 -18476 16008
rect -19648 15928 -18560 15992
rect -18496 15928 -18476 15992
rect -19648 15912 -18476 15928
rect -19648 15848 -18560 15912
rect -18496 15848 -18476 15912
rect -19648 15832 -18476 15848
rect -19648 15768 -18560 15832
rect -18496 15768 -18476 15832
rect -19648 15752 -18476 15768
rect -19648 15688 -18560 15752
rect -18496 15688 -18476 15752
rect -19648 15672 -18476 15688
rect -19648 15608 -18560 15672
rect -18496 15608 -18476 15672
rect -19648 15592 -18476 15608
rect -19648 15528 -18560 15592
rect -18496 15528 -18476 15592
rect -19648 15512 -18476 15528
rect -19648 15448 -18560 15512
rect -18496 15448 -18476 15512
rect -19648 15432 -18476 15448
rect -19648 15368 -18560 15432
rect -18496 15368 -18476 15432
rect -19648 15352 -18476 15368
rect -19648 15288 -18560 15352
rect -18496 15288 -18476 15352
rect -19648 15240 -18476 15288
rect -18236 16072 -17064 16120
rect -18236 16008 -17148 16072
rect -17084 16008 -17064 16072
rect -18236 15992 -17064 16008
rect -18236 15928 -17148 15992
rect -17084 15928 -17064 15992
rect -18236 15912 -17064 15928
rect -18236 15848 -17148 15912
rect -17084 15848 -17064 15912
rect -18236 15832 -17064 15848
rect -18236 15768 -17148 15832
rect -17084 15768 -17064 15832
rect -18236 15752 -17064 15768
rect -18236 15688 -17148 15752
rect -17084 15688 -17064 15752
rect -18236 15672 -17064 15688
rect -18236 15608 -17148 15672
rect -17084 15608 -17064 15672
rect -18236 15592 -17064 15608
rect -18236 15528 -17148 15592
rect -17084 15528 -17064 15592
rect -18236 15512 -17064 15528
rect -18236 15448 -17148 15512
rect -17084 15448 -17064 15512
rect -18236 15432 -17064 15448
rect -18236 15368 -17148 15432
rect -17084 15368 -17064 15432
rect -18236 15352 -17064 15368
rect -18236 15288 -17148 15352
rect -17084 15288 -17064 15352
rect -18236 15240 -17064 15288
rect -16824 16072 -15652 16120
rect -16824 16008 -15736 16072
rect -15672 16008 -15652 16072
rect -16824 15992 -15652 16008
rect -16824 15928 -15736 15992
rect -15672 15928 -15652 15992
rect -16824 15912 -15652 15928
rect -16824 15848 -15736 15912
rect -15672 15848 -15652 15912
rect -16824 15832 -15652 15848
rect -16824 15768 -15736 15832
rect -15672 15768 -15652 15832
rect -16824 15752 -15652 15768
rect -16824 15688 -15736 15752
rect -15672 15688 -15652 15752
rect -16824 15672 -15652 15688
rect -16824 15608 -15736 15672
rect -15672 15608 -15652 15672
rect -16824 15592 -15652 15608
rect -16824 15528 -15736 15592
rect -15672 15528 -15652 15592
rect -16824 15512 -15652 15528
rect -16824 15448 -15736 15512
rect -15672 15448 -15652 15512
rect -16824 15432 -15652 15448
rect -16824 15368 -15736 15432
rect -15672 15368 -15652 15432
rect -16824 15352 -15652 15368
rect -16824 15288 -15736 15352
rect -15672 15288 -15652 15352
rect -16824 15240 -15652 15288
rect -15412 16072 -14240 16120
rect -15412 16008 -14324 16072
rect -14260 16008 -14240 16072
rect -15412 15992 -14240 16008
rect -15412 15928 -14324 15992
rect -14260 15928 -14240 15992
rect -15412 15912 -14240 15928
rect -15412 15848 -14324 15912
rect -14260 15848 -14240 15912
rect -15412 15832 -14240 15848
rect -15412 15768 -14324 15832
rect -14260 15768 -14240 15832
rect -15412 15752 -14240 15768
rect -15412 15688 -14324 15752
rect -14260 15688 -14240 15752
rect -15412 15672 -14240 15688
rect -15412 15608 -14324 15672
rect -14260 15608 -14240 15672
rect -15412 15592 -14240 15608
rect -15412 15528 -14324 15592
rect -14260 15528 -14240 15592
rect -15412 15512 -14240 15528
rect -15412 15448 -14324 15512
rect -14260 15448 -14240 15512
rect -15412 15432 -14240 15448
rect -15412 15368 -14324 15432
rect -14260 15368 -14240 15432
rect -15412 15352 -14240 15368
rect -15412 15288 -14324 15352
rect -14260 15288 -14240 15352
rect -15412 15240 -14240 15288
rect -14000 16072 -12828 16120
rect -14000 16008 -12912 16072
rect -12848 16008 -12828 16072
rect -14000 15992 -12828 16008
rect -14000 15928 -12912 15992
rect -12848 15928 -12828 15992
rect -14000 15912 -12828 15928
rect -14000 15848 -12912 15912
rect -12848 15848 -12828 15912
rect -14000 15832 -12828 15848
rect -14000 15768 -12912 15832
rect -12848 15768 -12828 15832
rect -14000 15752 -12828 15768
rect -14000 15688 -12912 15752
rect -12848 15688 -12828 15752
rect -14000 15672 -12828 15688
rect -14000 15608 -12912 15672
rect -12848 15608 -12828 15672
rect -14000 15592 -12828 15608
rect -14000 15528 -12912 15592
rect -12848 15528 -12828 15592
rect -14000 15512 -12828 15528
rect -14000 15448 -12912 15512
rect -12848 15448 -12828 15512
rect -14000 15432 -12828 15448
rect -14000 15368 -12912 15432
rect -12848 15368 -12828 15432
rect -14000 15352 -12828 15368
rect -14000 15288 -12912 15352
rect -12848 15288 -12828 15352
rect -14000 15240 -12828 15288
rect -12588 16072 -11416 16120
rect -12588 16008 -11500 16072
rect -11436 16008 -11416 16072
rect -12588 15992 -11416 16008
rect -12588 15928 -11500 15992
rect -11436 15928 -11416 15992
rect -12588 15912 -11416 15928
rect -12588 15848 -11500 15912
rect -11436 15848 -11416 15912
rect -12588 15832 -11416 15848
rect -12588 15768 -11500 15832
rect -11436 15768 -11416 15832
rect -12588 15752 -11416 15768
rect -12588 15688 -11500 15752
rect -11436 15688 -11416 15752
rect -12588 15672 -11416 15688
rect -12588 15608 -11500 15672
rect -11436 15608 -11416 15672
rect -12588 15592 -11416 15608
rect -12588 15528 -11500 15592
rect -11436 15528 -11416 15592
rect -12588 15512 -11416 15528
rect -12588 15448 -11500 15512
rect -11436 15448 -11416 15512
rect -12588 15432 -11416 15448
rect -12588 15368 -11500 15432
rect -11436 15368 -11416 15432
rect -12588 15352 -11416 15368
rect -12588 15288 -11500 15352
rect -11436 15288 -11416 15352
rect -12588 15240 -11416 15288
rect -11176 16072 -10004 16120
rect -11176 16008 -10088 16072
rect -10024 16008 -10004 16072
rect -11176 15992 -10004 16008
rect -11176 15928 -10088 15992
rect -10024 15928 -10004 15992
rect -11176 15912 -10004 15928
rect -11176 15848 -10088 15912
rect -10024 15848 -10004 15912
rect -11176 15832 -10004 15848
rect -11176 15768 -10088 15832
rect -10024 15768 -10004 15832
rect -11176 15752 -10004 15768
rect -11176 15688 -10088 15752
rect -10024 15688 -10004 15752
rect -11176 15672 -10004 15688
rect -11176 15608 -10088 15672
rect -10024 15608 -10004 15672
rect -11176 15592 -10004 15608
rect -11176 15528 -10088 15592
rect -10024 15528 -10004 15592
rect -11176 15512 -10004 15528
rect -11176 15448 -10088 15512
rect -10024 15448 -10004 15512
rect -11176 15432 -10004 15448
rect -11176 15368 -10088 15432
rect -10024 15368 -10004 15432
rect -11176 15352 -10004 15368
rect -11176 15288 -10088 15352
rect -10024 15288 -10004 15352
rect -11176 15240 -10004 15288
rect -9764 16072 -8592 16120
rect -9764 16008 -8676 16072
rect -8612 16008 -8592 16072
rect -9764 15992 -8592 16008
rect -9764 15928 -8676 15992
rect -8612 15928 -8592 15992
rect -9764 15912 -8592 15928
rect -9764 15848 -8676 15912
rect -8612 15848 -8592 15912
rect -9764 15832 -8592 15848
rect -9764 15768 -8676 15832
rect -8612 15768 -8592 15832
rect -9764 15752 -8592 15768
rect -9764 15688 -8676 15752
rect -8612 15688 -8592 15752
rect -9764 15672 -8592 15688
rect -9764 15608 -8676 15672
rect -8612 15608 -8592 15672
rect -9764 15592 -8592 15608
rect -9764 15528 -8676 15592
rect -8612 15528 -8592 15592
rect -9764 15512 -8592 15528
rect -9764 15448 -8676 15512
rect -8612 15448 -8592 15512
rect -9764 15432 -8592 15448
rect -9764 15368 -8676 15432
rect -8612 15368 -8592 15432
rect -9764 15352 -8592 15368
rect -9764 15288 -8676 15352
rect -8612 15288 -8592 15352
rect -9764 15240 -8592 15288
rect -8352 16072 -7180 16120
rect -8352 16008 -7264 16072
rect -7200 16008 -7180 16072
rect -8352 15992 -7180 16008
rect -8352 15928 -7264 15992
rect -7200 15928 -7180 15992
rect -8352 15912 -7180 15928
rect -8352 15848 -7264 15912
rect -7200 15848 -7180 15912
rect -8352 15832 -7180 15848
rect -8352 15768 -7264 15832
rect -7200 15768 -7180 15832
rect -8352 15752 -7180 15768
rect -8352 15688 -7264 15752
rect -7200 15688 -7180 15752
rect -8352 15672 -7180 15688
rect -8352 15608 -7264 15672
rect -7200 15608 -7180 15672
rect -8352 15592 -7180 15608
rect -8352 15528 -7264 15592
rect -7200 15528 -7180 15592
rect -8352 15512 -7180 15528
rect -8352 15448 -7264 15512
rect -7200 15448 -7180 15512
rect -8352 15432 -7180 15448
rect -8352 15368 -7264 15432
rect -7200 15368 -7180 15432
rect -8352 15352 -7180 15368
rect -8352 15288 -7264 15352
rect -7200 15288 -7180 15352
rect -8352 15240 -7180 15288
rect -6940 16072 -5768 16120
rect -6940 16008 -5852 16072
rect -5788 16008 -5768 16072
rect -6940 15992 -5768 16008
rect -6940 15928 -5852 15992
rect -5788 15928 -5768 15992
rect -6940 15912 -5768 15928
rect -6940 15848 -5852 15912
rect -5788 15848 -5768 15912
rect -6940 15832 -5768 15848
rect -6940 15768 -5852 15832
rect -5788 15768 -5768 15832
rect -6940 15752 -5768 15768
rect -6940 15688 -5852 15752
rect -5788 15688 -5768 15752
rect -6940 15672 -5768 15688
rect -6940 15608 -5852 15672
rect -5788 15608 -5768 15672
rect -6940 15592 -5768 15608
rect -6940 15528 -5852 15592
rect -5788 15528 -5768 15592
rect -6940 15512 -5768 15528
rect -6940 15448 -5852 15512
rect -5788 15448 -5768 15512
rect -6940 15432 -5768 15448
rect -6940 15368 -5852 15432
rect -5788 15368 -5768 15432
rect -6940 15352 -5768 15368
rect -6940 15288 -5852 15352
rect -5788 15288 -5768 15352
rect -6940 15240 -5768 15288
rect -5528 16072 -4356 16120
rect -5528 16008 -4440 16072
rect -4376 16008 -4356 16072
rect -5528 15992 -4356 16008
rect -5528 15928 -4440 15992
rect -4376 15928 -4356 15992
rect -5528 15912 -4356 15928
rect -5528 15848 -4440 15912
rect -4376 15848 -4356 15912
rect -5528 15832 -4356 15848
rect -5528 15768 -4440 15832
rect -4376 15768 -4356 15832
rect -5528 15752 -4356 15768
rect -5528 15688 -4440 15752
rect -4376 15688 -4356 15752
rect -5528 15672 -4356 15688
rect -5528 15608 -4440 15672
rect -4376 15608 -4356 15672
rect -5528 15592 -4356 15608
rect -5528 15528 -4440 15592
rect -4376 15528 -4356 15592
rect -5528 15512 -4356 15528
rect -5528 15448 -4440 15512
rect -4376 15448 -4356 15512
rect -5528 15432 -4356 15448
rect -5528 15368 -4440 15432
rect -4376 15368 -4356 15432
rect -5528 15352 -4356 15368
rect -5528 15288 -4440 15352
rect -4376 15288 -4356 15352
rect -5528 15240 -4356 15288
rect -4116 16072 -2944 16120
rect -4116 16008 -3028 16072
rect -2964 16008 -2944 16072
rect -4116 15992 -2944 16008
rect -4116 15928 -3028 15992
rect -2964 15928 -2944 15992
rect -4116 15912 -2944 15928
rect -4116 15848 -3028 15912
rect -2964 15848 -2944 15912
rect -4116 15832 -2944 15848
rect -4116 15768 -3028 15832
rect -2964 15768 -2944 15832
rect -4116 15752 -2944 15768
rect -4116 15688 -3028 15752
rect -2964 15688 -2944 15752
rect -4116 15672 -2944 15688
rect -4116 15608 -3028 15672
rect -2964 15608 -2944 15672
rect -4116 15592 -2944 15608
rect -4116 15528 -3028 15592
rect -2964 15528 -2944 15592
rect -4116 15512 -2944 15528
rect -4116 15448 -3028 15512
rect -2964 15448 -2944 15512
rect -4116 15432 -2944 15448
rect -4116 15368 -3028 15432
rect -2964 15368 -2944 15432
rect -4116 15352 -2944 15368
rect -4116 15288 -3028 15352
rect -2964 15288 -2944 15352
rect -4116 15240 -2944 15288
rect -2704 16072 -1532 16120
rect -2704 16008 -1616 16072
rect -1552 16008 -1532 16072
rect -2704 15992 -1532 16008
rect -2704 15928 -1616 15992
rect -1552 15928 -1532 15992
rect -2704 15912 -1532 15928
rect -2704 15848 -1616 15912
rect -1552 15848 -1532 15912
rect -2704 15832 -1532 15848
rect -2704 15768 -1616 15832
rect -1552 15768 -1532 15832
rect -2704 15752 -1532 15768
rect -2704 15688 -1616 15752
rect -1552 15688 -1532 15752
rect -2704 15672 -1532 15688
rect -2704 15608 -1616 15672
rect -1552 15608 -1532 15672
rect -2704 15592 -1532 15608
rect -2704 15528 -1616 15592
rect -1552 15528 -1532 15592
rect -2704 15512 -1532 15528
rect -2704 15448 -1616 15512
rect -1552 15448 -1532 15512
rect -2704 15432 -1532 15448
rect -2704 15368 -1616 15432
rect -1552 15368 -1532 15432
rect -2704 15352 -1532 15368
rect -2704 15288 -1616 15352
rect -1552 15288 -1532 15352
rect -2704 15240 -1532 15288
rect -1292 16072 -120 16120
rect -1292 16008 -204 16072
rect -140 16008 -120 16072
rect -1292 15992 -120 16008
rect -1292 15928 -204 15992
rect -140 15928 -120 15992
rect -1292 15912 -120 15928
rect -1292 15848 -204 15912
rect -140 15848 -120 15912
rect -1292 15832 -120 15848
rect -1292 15768 -204 15832
rect -140 15768 -120 15832
rect -1292 15752 -120 15768
rect -1292 15688 -204 15752
rect -140 15688 -120 15752
rect -1292 15672 -120 15688
rect -1292 15608 -204 15672
rect -140 15608 -120 15672
rect -1292 15592 -120 15608
rect -1292 15528 -204 15592
rect -140 15528 -120 15592
rect -1292 15512 -120 15528
rect -1292 15448 -204 15512
rect -140 15448 -120 15512
rect -1292 15432 -120 15448
rect -1292 15368 -204 15432
rect -140 15368 -120 15432
rect -1292 15352 -120 15368
rect -1292 15288 -204 15352
rect -140 15288 -120 15352
rect -1292 15240 -120 15288
rect 120 16072 1292 16120
rect 120 16008 1208 16072
rect 1272 16008 1292 16072
rect 120 15992 1292 16008
rect 120 15928 1208 15992
rect 1272 15928 1292 15992
rect 120 15912 1292 15928
rect 120 15848 1208 15912
rect 1272 15848 1292 15912
rect 120 15832 1292 15848
rect 120 15768 1208 15832
rect 1272 15768 1292 15832
rect 120 15752 1292 15768
rect 120 15688 1208 15752
rect 1272 15688 1292 15752
rect 120 15672 1292 15688
rect 120 15608 1208 15672
rect 1272 15608 1292 15672
rect 120 15592 1292 15608
rect 120 15528 1208 15592
rect 1272 15528 1292 15592
rect 120 15512 1292 15528
rect 120 15448 1208 15512
rect 1272 15448 1292 15512
rect 120 15432 1292 15448
rect 120 15368 1208 15432
rect 1272 15368 1292 15432
rect 120 15352 1292 15368
rect 120 15288 1208 15352
rect 1272 15288 1292 15352
rect 120 15240 1292 15288
rect 1532 16072 2704 16120
rect 1532 16008 2620 16072
rect 2684 16008 2704 16072
rect 1532 15992 2704 16008
rect 1532 15928 2620 15992
rect 2684 15928 2704 15992
rect 1532 15912 2704 15928
rect 1532 15848 2620 15912
rect 2684 15848 2704 15912
rect 1532 15832 2704 15848
rect 1532 15768 2620 15832
rect 2684 15768 2704 15832
rect 1532 15752 2704 15768
rect 1532 15688 2620 15752
rect 2684 15688 2704 15752
rect 1532 15672 2704 15688
rect 1532 15608 2620 15672
rect 2684 15608 2704 15672
rect 1532 15592 2704 15608
rect 1532 15528 2620 15592
rect 2684 15528 2704 15592
rect 1532 15512 2704 15528
rect 1532 15448 2620 15512
rect 2684 15448 2704 15512
rect 1532 15432 2704 15448
rect 1532 15368 2620 15432
rect 2684 15368 2704 15432
rect 1532 15352 2704 15368
rect 1532 15288 2620 15352
rect 2684 15288 2704 15352
rect 1532 15240 2704 15288
rect 2944 16072 4116 16120
rect 2944 16008 4032 16072
rect 4096 16008 4116 16072
rect 2944 15992 4116 16008
rect 2944 15928 4032 15992
rect 4096 15928 4116 15992
rect 2944 15912 4116 15928
rect 2944 15848 4032 15912
rect 4096 15848 4116 15912
rect 2944 15832 4116 15848
rect 2944 15768 4032 15832
rect 4096 15768 4116 15832
rect 2944 15752 4116 15768
rect 2944 15688 4032 15752
rect 4096 15688 4116 15752
rect 2944 15672 4116 15688
rect 2944 15608 4032 15672
rect 4096 15608 4116 15672
rect 2944 15592 4116 15608
rect 2944 15528 4032 15592
rect 4096 15528 4116 15592
rect 2944 15512 4116 15528
rect 2944 15448 4032 15512
rect 4096 15448 4116 15512
rect 2944 15432 4116 15448
rect 2944 15368 4032 15432
rect 4096 15368 4116 15432
rect 2944 15352 4116 15368
rect 2944 15288 4032 15352
rect 4096 15288 4116 15352
rect 2944 15240 4116 15288
rect 4356 16072 5528 16120
rect 4356 16008 5444 16072
rect 5508 16008 5528 16072
rect 4356 15992 5528 16008
rect 4356 15928 5444 15992
rect 5508 15928 5528 15992
rect 4356 15912 5528 15928
rect 4356 15848 5444 15912
rect 5508 15848 5528 15912
rect 4356 15832 5528 15848
rect 4356 15768 5444 15832
rect 5508 15768 5528 15832
rect 4356 15752 5528 15768
rect 4356 15688 5444 15752
rect 5508 15688 5528 15752
rect 4356 15672 5528 15688
rect 4356 15608 5444 15672
rect 5508 15608 5528 15672
rect 4356 15592 5528 15608
rect 4356 15528 5444 15592
rect 5508 15528 5528 15592
rect 4356 15512 5528 15528
rect 4356 15448 5444 15512
rect 5508 15448 5528 15512
rect 4356 15432 5528 15448
rect 4356 15368 5444 15432
rect 5508 15368 5528 15432
rect 4356 15352 5528 15368
rect 4356 15288 5444 15352
rect 5508 15288 5528 15352
rect 4356 15240 5528 15288
rect 5768 16072 6940 16120
rect 5768 16008 6856 16072
rect 6920 16008 6940 16072
rect 5768 15992 6940 16008
rect 5768 15928 6856 15992
rect 6920 15928 6940 15992
rect 5768 15912 6940 15928
rect 5768 15848 6856 15912
rect 6920 15848 6940 15912
rect 5768 15832 6940 15848
rect 5768 15768 6856 15832
rect 6920 15768 6940 15832
rect 5768 15752 6940 15768
rect 5768 15688 6856 15752
rect 6920 15688 6940 15752
rect 5768 15672 6940 15688
rect 5768 15608 6856 15672
rect 6920 15608 6940 15672
rect 5768 15592 6940 15608
rect 5768 15528 6856 15592
rect 6920 15528 6940 15592
rect 5768 15512 6940 15528
rect 5768 15448 6856 15512
rect 6920 15448 6940 15512
rect 5768 15432 6940 15448
rect 5768 15368 6856 15432
rect 6920 15368 6940 15432
rect 5768 15352 6940 15368
rect 5768 15288 6856 15352
rect 6920 15288 6940 15352
rect 5768 15240 6940 15288
rect 7180 16072 8352 16120
rect 7180 16008 8268 16072
rect 8332 16008 8352 16072
rect 7180 15992 8352 16008
rect 7180 15928 8268 15992
rect 8332 15928 8352 15992
rect 7180 15912 8352 15928
rect 7180 15848 8268 15912
rect 8332 15848 8352 15912
rect 7180 15832 8352 15848
rect 7180 15768 8268 15832
rect 8332 15768 8352 15832
rect 7180 15752 8352 15768
rect 7180 15688 8268 15752
rect 8332 15688 8352 15752
rect 7180 15672 8352 15688
rect 7180 15608 8268 15672
rect 8332 15608 8352 15672
rect 7180 15592 8352 15608
rect 7180 15528 8268 15592
rect 8332 15528 8352 15592
rect 7180 15512 8352 15528
rect 7180 15448 8268 15512
rect 8332 15448 8352 15512
rect 7180 15432 8352 15448
rect 7180 15368 8268 15432
rect 8332 15368 8352 15432
rect 7180 15352 8352 15368
rect 7180 15288 8268 15352
rect 8332 15288 8352 15352
rect 7180 15240 8352 15288
rect 8592 16072 9764 16120
rect 8592 16008 9680 16072
rect 9744 16008 9764 16072
rect 8592 15992 9764 16008
rect 8592 15928 9680 15992
rect 9744 15928 9764 15992
rect 8592 15912 9764 15928
rect 8592 15848 9680 15912
rect 9744 15848 9764 15912
rect 8592 15832 9764 15848
rect 8592 15768 9680 15832
rect 9744 15768 9764 15832
rect 8592 15752 9764 15768
rect 8592 15688 9680 15752
rect 9744 15688 9764 15752
rect 8592 15672 9764 15688
rect 8592 15608 9680 15672
rect 9744 15608 9764 15672
rect 8592 15592 9764 15608
rect 8592 15528 9680 15592
rect 9744 15528 9764 15592
rect 8592 15512 9764 15528
rect 8592 15448 9680 15512
rect 9744 15448 9764 15512
rect 8592 15432 9764 15448
rect 8592 15368 9680 15432
rect 9744 15368 9764 15432
rect 8592 15352 9764 15368
rect 8592 15288 9680 15352
rect 9744 15288 9764 15352
rect 8592 15240 9764 15288
rect 10004 16072 11176 16120
rect 10004 16008 11092 16072
rect 11156 16008 11176 16072
rect 10004 15992 11176 16008
rect 10004 15928 11092 15992
rect 11156 15928 11176 15992
rect 10004 15912 11176 15928
rect 10004 15848 11092 15912
rect 11156 15848 11176 15912
rect 10004 15832 11176 15848
rect 10004 15768 11092 15832
rect 11156 15768 11176 15832
rect 10004 15752 11176 15768
rect 10004 15688 11092 15752
rect 11156 15688 11176 15752
rect 10004 15672 11176 15688
rect 10004 15608 11092 15672
rect 11156 15608 11176 15672
rect 10004 15592 11176 15608
rect 10004 15528 11092 15592
rect 11156 15528 11176 15592
rect 10004 15512 11176 15528
rect 10004 15448 11092 15512
rect 11156 15448 11176 15512
rect 10004 15432 11176 15448
rect 10004 15368 11092 15432
rect 11156 15368 11176 15432
rect 10004 15352 11176 15368
rect 10004 15288 11092 15352
rect 11156 15288 11176 15352
rect 10004 15240 11176 15288
rect 11416 16072 12588 16120
rect 11416 16008 12504 16072
rect 12568 16008 12588 16072
rect 11416 15992 12588 16008
rect 11416 15928 12504 15992
rect 12568 15928 12588 15992
rect 11416 15912 12588 15928
rect 11416 15848 12504 15912
rect 12568 15848 12588 15912
rect 11416 15832 12588 15848
rect 11416 15768 12504 15832
rect 12568 15768 12588 15832
rect 11416 15752 12588 15768
rect 11416 15688 12504 15752
rect 12568 15688 12588 15752
rect 11416 15672 12588 15688
rect 11416 15608 12504 15672
rect 12568 15608 12588 15672
rect 11416 15592 12588 15608
rect 11416 15528 12504 15592
rect 12568 15528 12588 15592
rect 11416 15512 12588 15528
rect 11416 15448 12504 15512
rect 12568 15448 12588 15512
rect 11416 15432 12588 15448
rect 11416 15368 12504 15432
rect 12568 15368 12588 15432
rect 11416 15352 12588 15368
rect 11416 15288 12504 15352
rect 12568 15288 12588 15352
rect 11416 15240 12588 15288
rect 12828 16072 14000 16120
rect 12828 16008 13916 16072
rect 13980 16008 14000 16072
rect 12828 15992 14000 16008
rect 12828 15928 13916 15992
rect 13980 15928 14000 15992
rect 12828 15912 14000 15928
rect 12828 15848 13916 15912
rect 13980 15848 14000 15912
rect 12828 15832 14000 15848
rect 12828 15768 13916 15832
rect 13980 15768 14000 15832
rect 12828 15752 14000 15768
rect 12828 15688 13916 15752
rect 13980 15688 14000 15752
rect 12828 15672 14000 15688
rect 12828 15608 13916 15672
rect 13980 15608 14000 15672
rect 12828 15592 14000 15608
rect 12828 15528 13916 15592
rect 13980 15528 14000 15592
rect 12828 15512 14000 15528
rect 12828 15448 13916 15512
rect 13980 15448 14000 15512
rect 12828 15432 14000 15448
rect 12828 15368 13916 15432
rect 13980 15368 14000 15432
rect 12828 15352 14000 15368
rect 12828 15288 13916 15352
rect 13980 15288 14000 15352
rect 12828 15240 14000 15288
rect 14240 16072 15412 16120
rect 14240 16008 15328 16072
rect 15392 16008 15412 16072
rect 14240 15992 15412 16008
rect 14240 15928 15328 15992
rect 15392 15928 15412 15992
rect 14240 15912 15412 15928
rect 14240 15848 15328 15912
rect 15392 15848 15412 15912
rect 14240 15832 15412 15848
rect 14240 15768 15328 15832
rect 15392 15768 15412 15832
rect 14240 15752 15412 15768
rect 14240 15688 15328 15752
rect 15392 15688 15412 15752
rect 14240 15672 15412 15688
rect 14240 15608 15328 15672
rect 15392 15608 15412 15672
rect 14240 15592 15412 15608
rect 14240 15528 15328 15592
rect 15392 15528 15412 15592
rect 14240 15512 15412 15528
rect 14240 15448 15328 15512
rect 15392 15448 15412 15512
rect 14240 15432 15412 15448
rect 14240 15368 15328 15432
rect 15392 15368 15412 15432
rect 14240 15352 15412 15368
rect 14240 15288 15328 15352
rect 15392 15288 15412 15352
rect 14240 15240 15412 15288
rect 15652 16072 16824 16120
rect 15652 16008 16740 16072
rect 16804 16008 16824 16072
rect 15652 15992 16824 16008
rect 15652 15928 16740 15992
rect 16804 15928 16824 15992
rect 15652 15912 16824 15928
rect 15652 15848 16740 15912
rect 16804 15848 16824 15912
rect 15652 15832 16824 15848
rect 15652 15768 16740 15832
rect 16804 15768 16824 15832
rect 15652 15752 16824 15768
rect 15652 15688 16740 15752
rect 16804 15688 16824 15752
rect 15652 15672 16824 15688
rect 15652 15608 16740 15672
rect 16804 15608 16824 15672
rect 15652 15592 16824 15608
rect 15652 15528 16740 15592
rect 16804 15528 16824 15592
rect 15652 15512 16824 15528
rect 15652 15448 16740 15512
rect 16804 15448 16824 15512
rect 15652 15432 16824 15448
rect 15652 15368 16740 15432
rect 16804 15368 16824 15432
rect 15652 15352 16824 15368
rect 15652 15288 16740 15352
rect 16804 15288 16824 15352
rect 15652 15240 16824 15288
rect 17064 16072 18236 16120
rect 17064 16008 18152 16072
rect 18216 16008 18236 16072
rect 17064 15992 18236 16008
rect 17064 15928 18152 15992
rect 18216 15928 18236 15992
rect 17064 15912 18236 15928
rect 17064 15848 18152 15912
rect 18216 15848 18236 15912
rect 17064 15832 18236 15848
rect 17064 15768 18152 15832
rect 18216 15768 18236 15832
rect 17064 15752 18236 15768
rect 17064 15688 18152 15752
rect 18216 15688 18236 15752
rect 17064 15672 18236 15688
rect 17064 15608 18152 15672
rect 18216 15608 18236 15672
rect 17064 15592 18236 15608
rect 17064 15528 18152 15592
rect 18216 15528 18236 15592
rect 17064 15512 18236 15528
rect 17064 15448 18152 15512
rect 18216 15448 18236 15512
rect 17064 15432 18236 15448
rect 17064 15368 18152 15432
rect 18216 15368 18236 15432
rect 17064 15352 18236 15368
rect 17064 15288 18152 15352
rect 18216 15288 18236 15352
rect 17064 15240 18236 15288
rect 18476 16072 19648 16120
rect 18476 16008 19564 16072
rect 19628 16008 19648 16072
rect 18476 15992 19648 16008
rect 18476 15928 19564 15992
rect 19628 15928 19648 15992
rect 18476 15912 19648 15928
rect 18476 15848 19564 15912
rect 19628 15848 19648 15912
rect 18476 15832 19648 15848
rect 18476 15768 19564 15832
rect 19628 15768 19648 15832
rect 18476 15752 19648 15768
rect 18476 15688 19564 15752
rect 19628 15688 19648 15752
rect 18476 15672 19648 15688
rect 18476 15608 19564 15672
rect 19628 15608 19648 15672
rect 18476 15592 19648 15608
rect 18476 15528 19564 15592
rect 19628 15528 19648 15592
rect 18476 15512 19648 15528
rect 18476 15448 19564 15512
rect 19628 15448 19648 15512
rect 18476 15432 19648 15448
rect 18476 15368 19564 15432
rect 19628 15368 19648 15432
rect 18476 15352 19648 15368
rect 18476 15288 19564 15352
rect 19628 15288 19648 15352
rect 18476 15240 19648 15288
rect 19888 16072 21060 16120
rect 19888 16008 20976 16072
rect 21040 16008 21060 16072
rect 19888 15992 21060 16008
rect 19888 15928 20976 15992
rect 21040 15928 21060 15992
rect 19888 15912 21060 15928
rect 19888 15848 20976 15912
rect 21040 15848 21060 15912
rect 19888 15832 21060 15848
rect 19888 15768 20976 15832
rect 21040 15768 21060 15832
rect 19888 15752 21060 15768
rect 19888 15688 20976 15752
rect 21040 15688 21060 15752
rect 19888 15672 21060 15688
rect 19888 15608 20976 15672
rect 21040 15608 21060 15672
rect 19888 15592 21060 15608
rect 19888 15528 20976 15592
rect 21040 15528 21060 15592
rect 19888 15512 21060 15528
rect 19888 15448 20976 15512
rect 21040 15448 21060 15512
rect 19888 15432 21060 15448
rect 19888 15368 20976 15432
rect 21040 15368 21060 15432
rect 19888 15352 21060 15368
rect 19888 15288 20976 15352
rect 21040 15288 21060 15352
rect 19888 15240 21060 15288
rect 21300 16072 22472 16120
rect 21300 16008 22388 16072
rect 22452 16008 22472 16072
rect 21300 15992 22472 16008
rect 21300 15928 22388 15992
rect 22452 15928 22472 15992
rect 21300 15912 22472 15928
rect 21300 15848 22388 15912
rect 22452 15848 22472 15912
rect 21300 15832 22472 15848
rect 21300 15768 22388 15832
rect 22452 15768 22472 15832
rect 21300 15752 22472 15768
rect 21300 15688 22388 15752
rect 22452 15688 22472 15752
rect 21300 15672 22472 15688
rect 21300 15608 22388 15672
rect 22452 15608 22472 15672
rect 21300 15592 22472 15608
rect 21300 15528 22388 15592
rect 22452 15528 22472 15592
rect 21300 15512 22472 15528
rect 21300 15448 22388 15512
rect 22452 15448 22472 15512
rect 21300 15432 22472 15448
rect 21300 15368 22388 15432
rect 22452 15368 22472 15432
rect 21300 15352 22472 15368
rect 21300 15288 22388 15352
rect 22452 15288 22472 15352
rect 21300 15240 22472 15288
rect 22712 16072 23884 16120
rect 22712 16008 23800 16072
rect 23864 16008 23884 16072
rect 22712 15992 23884 16008
rect 22712 15928 23800 15992
rect 23864 15928 23884 15992
rect 22712 15912 23884 15928
rect 22712 15848 23800 15912
rect 23864 15848 23884 15912
rect 22712 15832 23884 15848
rect 22712 15768 23800 15832
rect 23864 15768 23884 15832
rect 22712 15752 23884 15768
rect 22712 15688 23800 15752
rect 23864 15688 23884 15752
rect 22712 15672 23884 15688
rect 22712 15608 23800 15672
rect 23864 15608 23884 15672
rect 22712 15592 23884 15608
rect 22712 15528 23800 15592
rect 23864 15528 23884 15592
rect 22712 15512 23884 15528
rect 22712 15448 23800 15512
rect 23864 15448 23884 15512
rect 22712 15432 23884 15448
rect 22712 15368 23800 15432
rect 23864 15368 23884 15432
rect 22712 15352 23884 15368
rect 22712 15288 23800 15352
rect 23864 15288 23884 15352
rect 22712 15240 23884 15288
rect -23884 14952 -22712 15000
rect -23884 14888 -22796 14952
rect -22732 14888 -22712 14952
rect -23884 14872 -22712 14888
rect -23884 14808 -22796 14872
rect -22732 14808 -22712 14872
rect -23884 14792 -22712 14808
rect -23884 14728 -22796 14792
rect -22732 14728 -22712 14792
rect -23884 14712 -22712 14728
rect -23884 14648 -22796 14712
rect -22732 14648 -22712 14712
rect -23884 14632 -22712 14648
rect -23884 14568 -22796 14632
rect -22732 14568 -22712 14632
rect -23884 14552 -22712 14568
rect -23884 14488 -22796 14552
rect -22732 14488 -22712 14552
rect -23884 14472 -22712 14488
rect -23884 14408 -22796 14472
rect -22732 14408 -22712 14472
rect -23884 14392 -22712 14408
rect -23884 14328 -22796 14392
rect -22732 14328 -22712 14392
rect -23884 14312 -22712 14328
rect -23884 14248 -22796 14312
rect -22732 14248 -22712 14312
rect -23884 14232 -22712 14248
rect -23884 14168 -22796 14232
rect -22732 14168 -22712 14232
rect -23884 14120 -22712 14168
rect -22472 14952 -21300 15000
rect -22472 14888 -21384 14952
rect -21320 14888 -21300 14952
rect -22472 14872 -21300 14888
rect -22472 14808 -21384 14872
rect -21320 14808 -21300 14872
rect -22472 14792 -21300 14808
rect -22472 14728 -21384 14792
rect -21320 14728 -21300 14792
rect -22472 14712 -21300 14728
rect -22472 14648 -21384 14712
rect -21320 14648 -21300 14712
rect -22472 14632 -21300 14648
rect -22472 14568 -21384 14632
rect -21320 14568 -21300 14632
rect -22472 14552 -21300 14568
rect -22472 14488 -21384 14552
rect -21320 14488 -21300 14552
rect -22472 14472 -21300 14488
rect -22472 14408 -21384 14472
rect -21320 14408 -21300 14472
rect -22472 14392 -21300 14408
rect -22472 14328 -21384 14392
rect -21320 14328 -21300 14392
rect -22472 14312 -21300 14328
rect -22472 14248 -21384 14312
rect -21320 14248 -21300 14312
rect -22472 14232 -21300 14248
rect -22472 14168 -21384 14232
rect -21320 14168 -21300 14232
rect -22472 14120 -21300 14168
rect -21060 14952 -19888 15000
rect -21060 14888 -19972 14952
rect -19908 14888 -19888 14952
rect -21060 14872 -19888 14888
rect -21060 14808 -19972 14872
rect -19908 14808 -19888 14872
rect -21060 14792 -19888 14808
rect -21060 14728 -19972 14792
rect -19908 14728 -19888 14792
rect -21060 14712 -19888 14728
rect -21060 14648 -19972 14712
rect -19908 14648 -19888 14712
rect -21060 14632 -19888 14648
rect -21060 14568 -19972 14632
rect -19908 14568 -19888 14632
rect -21060 14552 -19888 14568
rect -21060 14488 -19972 14552
rect -19908 14488 -19888 14552
rect -21060 14472 -19888 14488
rect -21060 14408 -19972 14472
rect -19908 14408 -19888 14472
rect -21060 14392 -19888 14408
rect -21060 14328 -19972 14392
rect -19908 14328 -19888 14392
rect -21060 14312 -19888 14328
rect -21060 14248 -19972 14312
rect -19908 14248 -19888 14312
rect -21060 14232 -19888 14248
rect -21060 14168 -19972 14232
rect -19908 14168 -19888 14232
rect -21060 14120 -19888 14168
rect -19648 14952 -18476 15000
rect -19648 14888 -18560 14952
rect -18496 14888 -18476 14952
rect -19648 14872 -18476 14888
rect -19648 14808 -18560 14872
rect -18496 14808 -18476 14872
rect -19648 14792 -18476 14808
rect -19648 14728 -18560 14792
rect -18496 14728 -18476 14792
rect -19648 14712 -18476 14728
rect -19648 14648 -18560 14712
rect -18496 14648 -18476 14712
rect -19648 14632 -18476 14648
rect -19648 14568 -18560 14632
rect -18496 14568 -18476 14632
rect -19648 14552 -18476 14568
rect -19648 14488 -18560 14552
rect -18496 14488 -18476 14552
rect -19648 14472 -18476 14488
rect -19648 14408 -18560 14472
rect -18496 14408 -18476 14472
rect -19648 14392 -18476 14408
rect -19648 14328 -18560 14392
rect -18496 14328 -18476 14392
rect -19648 14312 -18476 14328
rect -19648 14248 -18560 14312
rect -18496 14248 -18476 14312
rect -19648 14232 -18476 14248
rect -19648 14168 -18560 14232
rect -18496 14168 -18476 14232
rect -19648 14120 -18476 14168
rect -18236 14952 -17064 15000
rect -18236 14888 -17148 14952
rect -17084 14888 -17064 14952
rect -18236 14872 -17064 14888
rect -18236 14808 -17148 14872
rect -17084 14808 -17064 14872
rect -18236 14792 -17064 14808
rect -18236 14728 -17148 14792
rect -17084 14728 -17064 14792
rect -18236 14712 -17064 14728
rect -18236 14648 -17148 14712
rect -17084 14648 -17064 14712
rect -18236 14632 -17064 14648
rect -18236 14568 -17148 14632
rect -17084 14568 -17064 14632
rect -18236 14552 -17064 14568
rect -18236 14488 -17148 14552
rect -17084 14488 -17064 14552
rect -18236 14472 -17064 14488
rect -18236 14408 -17148 14472
rect -17084 14408 -17064 14472
rect -18236 14392 -17064 14408
rect -18236 14328 -17148 14392
rect -17084 14328 -17064 14392
rect -18236 14312 -17064 14328
rect -18236 14248 -17148 14312
rect -17084 14248 -17064 14312
rect -18236 14232 -17064 14248
rect -18236 14168 -17148 14232
rect -17084 14168 -17064 14232
rect -18236 14120 -17064 14168
rect -16824 14952 -15652 15000
rect -16824 14888 -15736 14952
rect -15672 14888 -15652 14952
rect -16824 14872 -15652 14888
rect -16824 14808 -15736 14872
rect -15672 14808 -15652 14872
rect -16824 14792 -15652 14808
rect -16824 14728 -15736 14792
rect -15672 14728 -15652 14792
rect -16824 14712 -15652 14728
rect -16824 14648 -15736 14712
rect -15672 14648 -15652 14712
rect -16824 14632 -15652 14648
rect -16824 14568 -15736 14632
rect -15672 14568 -15652 14632
rect -16824 14552 -15652 14568
rect -16824 14488 -15736 14552
rect -15672 14488 -15652 14552
rect -16824 14472 -15652 14488
rect -16824 14408 -15736 14472
rect -15672 14408 -15652 14472
rect -16824 14392 -15652 14408
rect -16824 14328 -15736 14392
rect -15672 14328 -15652 14392
rect -16824 14312 -15652 14328
rect -16824 14248 -15736 14312
rect -15672 14248 -15652 14312
rect -16824 14232 -15652 14248
rect -16824 14168 -15736 14232
rect -15672 14168 -15652 14232
rect -16824 14120 -15652 14168
rect -15412 14952 -14240 15000
rect -15412 14888 -14324 14952
rect -14260 14888 -14240 14952
rect -15412 14872 -14240 14888
rect -15412 14808 -14324 14872
rect -14260 14808 -14240 14872
rect -15412 14792 -14240 14808
rect -15412 14728 -14324 14792
rect -14260 14728 -14240 14792
rect -15412 14712 -14240 14728
rect -15412 14648 -14324 14712
rect -14260 14648 -14240 14712
rect -15412 14632 -14240 14648
rect -15412 14568 -14324 14632
rect -14260 14568 -14240 14632
rect -15412 14552 -14240 14568
rect -15412 14488 -14324 14552
rect -14260 14488 -14240 14552
rect -15412 14472 -14240 14488
rect -15412 14408 -14324 14472
rect -14260 14408 -14240 14472
rect -15412 14392 -14240 14408
rect -15412 14328 -14324 14392
rect -14260 14328 -14240 14392
rect -15412 14312 -14240 14328
rect -15412 14248 -14324 14312
rect -14260 14248 -14240 14312
rect -15412 14232 -14240 14248
rect -15412 14168 -14324 14232
rect -14260 14168 -14240 14232
rect -15412 14120 -14240 14168
rect -14000 14952 -12828 15000
rect -14000 14888 -12912 14952
rect -12848 14888 -12828 14952
rect -14000 14872 -12828 14888
rect -14000 14808 -12912 14872
rect -12848 14808 -12828 14872
rect -14000 14792 -12828 14808
rect -14000 14728 -12912 14792
rect -12848 14728 -12828 14792
rect -14000 14712 -12828 14728
rect -14000 14648 -12912 14712
rect -12848 14648 -12828 14712
rect -14000 14632 -12828 14648
rect -14000 14568 -12912 14632
rect -12848 14568 -12828 14632
rect -14000 14552 -12828 14568
rect -14000 14488 -12912 14552
rect -12848 14488 -12828 14552
rect -14000 14472 -12828 14488
rect -14000 14408 -12912 14472
rect -12848 14408 -12828 14472
rect -14000 14392 -12828 14408
rect -14000 14328 -12912 14392
rect -12848 14328 -12828 14392
rect -14000 14312 -12828 14328
rect -14000 14248 -12912 14312
rect -12848 14248 -12828 14312
rect -14000 14232 -12828 14248
rect -14000 14168 -12912 14232
rect -12848 14168 -12828 14232
rect -14000 14120 -12828 14168
rect -12588 14952 -11416 15000
rect -12588 14888 -11500 14952
rect -11436 14888 -11416 14952
rect -12588 14872 -11416 14888
rect -12588 14808 -11500 14872
rect -11436 14808 -11416 14872
rect -12588 14792 -11416 14808
rect -12588 14728 -11500 14792
rect -11436 14728 -11416 14792
rect -12588 14712 -11416 14728
rect -12588 14648 -11500 14712
rect -11436 14648 -11416 14712
rect -12588 14632 -11416 14648
rect -12588 14568 -11500 14632
rect -11436 14568 -11416 14632
rect -12588 14552 -11416 14568
rect -12588 14488 -11500 14552
rect -11436 14488 -11416 14552
rect -12588 14472 -11416 14488
rect -12588 14408 -11500 14472
rect -11436 14408 -11416 14472
rect -12588 14392 -11416 14408
rect -12588 14328 -11500 14392
rect -11436 14328 -11416 14392
rect -12588 14312 -11416 14328
rect -12588 14248 -11500 14312
rect -11436 14248 -11416 14312
rect -12588 14232 -11416 14248
rect -12588 14168 -11500 14232
rect -11436 14168 -11416 14232
rect -12588 14120 -11416 14168
rect -11176 14952 -10004 15000
rect -11176 14888 -10088 14952
rect -10024 14888 -10004 14952
rect -11176 14872 -10004 14888
rect -11176 14808 -10088 14872
rect -10024 14808 -10004 14872
rect -11176 14792 -10004 14808
rect -11176 14728 -10088 14792
rect -10024 14728 -10004 14792
rect -11176 14712 -10004 14728
rect -11176 14648 -10088 14712
rect -10024 14648 -10004 14712
rect -11176 14632 -10004 14648
rect -11176 14568 -10088 14632
rect -10024 14568 -10004 14632
rect -11176 14552 -10004 14568
rect -11176 14488 -10088 14552
rect -10024 14488 -10004 14552
rect -11176 14472 -10004 14488
rect -11176 14408 -10088 14472
rect -10024 14408 -10004 14472
rect -11176 14392 -10004 14408
rect -11176 14328 -10088 14392
rect -10024 14328 -10004 14392
rect -11176 14312 -10004 14328
rect -11176 14248 -10088 14312
rect -10024 14248 -10004 14312
rect -11176 14232 -10004 14248
rect -11176 14168 -10088 14232
rect -10024 14168 -10004 14232
rect -11176 14120 -10004 14168
rect -9764 14952 -8592 15000
rect -9764 14888 -8676 14952
rect -8612 14888 -8592 14952
rect -9764 14872 -8592 14888
rect -9764 14808 -8676 14872
rect -8612 14808 -8592 14872
rect -9764 14792 -8592 14808
rect -9764 14728 -8676 14792
rect -8612 14728 -8592 14792
rect -9764 14712 -8592 14728
rect -9764 14648 -8676 14712
rect -8612 14648 -8592 14712
rect -9764 14632 -8592 14648
rect -9764 14568 -8676 14632
rect -8612 14568 -8592 14632
rect -9764 14552 -8592 14568
rect -9764 14488 -8676 14552
rect -8612 14488 -8592 14552
rect -9764 14472 -8592 14488
rect -9764 14408 -8676 14472
rect -8612 14408 -8592 14472
rect -9764 14392 -8592 14408
rect -9764 14328 -8676 14392
rect -8612 14328 -8592 14392
rect -9764 14312 -8592 14328
rect -9764 14248 -8676 14312
rect -8612 14248 -8592 14312
rect -9764 14232 -8592 14248
rect -9764 14168 -8676 14232
rect -8612 14168 -8592 14232
rect -9764 14120 -8592 14168
rect -8352 14952 -7180 15000
rect -8352 14888 -7264 14952
rect -7200 14888 -7180 14952
rect -8352 14872 -7180 14888
rect -8352 14808 -7264 14872
rect -7200 14808 -7180 14872
rect -8352 14792 -7180 14808
rect -8352 14728 -7264 14792
rect -7200 14728 -7180 14792
rect -8352 14712 -7180 14728
rect -8352 14648 -7264 14712
rect -7200 14648 -7180 14712
rect -8352 14632 -7180 14648
rect -8352 14568 -7264 14632
rect -7200 14568 -7180 14632
rect -8352 14552 -7180 14568
rect -8352 14488 -7264 14552
rect -7200 14488 -7180 14552
rect -8352 14472 -7180 14488
rect -8352 14408 -7264 14472
rect -7200 14408 -7180 14472
rect -8352 14392 -7180 14408
rect -8352 14328 -7264 14392
rect -7200 14328 -7180 14392
rect -8352 14312 -7180 14328
rect -8352 14248 -7264 14312
rect -7200 14248 -7180 14312
rect -8352 14232 -7180 14248
rect -8352 14168 -7264 14232
rect -7200 14168 -7180 14232
rect -8352 14120 -7180 14168
rect -6940 14952 -5768 15000
rect -6940 14888 -5852 14952
rect -5788 14888 -5768 14952
rect -6940 14872 -5768 14888
rect -6940 14808 -5852 14872
rect -5788 14808 -5768 14872
rect -6940 14792 -5768 14808
rect -6940 14728 -5852 14792
rect -5788 14728 -5768 14792
rect -6940 14712 -5768 14728
rect -6940 14648 -5852 14712
rect -5788 14648 -5768 14712
rect -6940 14632 -5768 14648
rect -6940 14568 -5852 14632
rect -5788 14568 -5768 14632
rect -6940 14552 -5768 14568
rect -6940 14488 -5852 14552
rect -5788 14488 -5768 14552
rect -6940 14472 -5768 14488
rect -6940 14408 -5852 14472
rect -5788 14408 -5768 14472
rect -6940 14392 -5768 14408
rect -6940 14328 -5852 14392
rect -5788 14328 -5768 14392
rect -6940 14312 -5768 14328
rect -6940 14248 -5852 14312
rect -5788 14248 -5768 14312
rect -6940 14232 -5768 14248
rect -6940 14168 -5852 14232
rect -5788 14168 -5768 14232
rect -6940 14120 -5768 14168
rect -5528 14952 -4356 15000
rect -5528 14888 -4440 14952
rect -4376 14888 -4356 14952
rect -5528 14872 -4356 14888
rect -5528 14808 -4440 14872
rect -4376 14808 -4356 14872
rect -5528 14792 -4356 14808
rect -5528 14728 -4440 14792
rect -4376 14728 -4356 14792
rect -5528 14712 -4356 14728
rect -5528 14648 -4440 14712
rect -4376 14648 -4356 14712
rect -5528 14632 -4356 14648
rect -5528 14568 -4440 14632
rect -4376 14568 -4356 14632
rect -5528 14552 -4356 14568
rect -5528 14488 -4440 14552
rect -4376 14488 -4356 14552
rect -5528 14472 -4356 14488
rect -5528 14408 -4440 14472
rect -4376 14408 -4356 14472
rect -5528 14392 -4356 14408
rect -5528 14328 -4440 14392
rect -4376 14328 -4356 14392
rect -5528 14312 -4356 14328
rect -5528 14248 -4440 14312
rect -4376 14248 -4356 14312
rect -5528 14232 -4356 14248
rect -5528 14168 -4440 14232
rect -4376 14168 -4356 14232
rect -5528 14120 -4356 14168
rect -4116 14952 -2944 15000
rect -4116 14888 -3028 14952
rect -2964 14888 -2944 14952
rect -4116 14872 -2944 14888
rect -4116 14808 -3028 14872
rect -2964 14808 -2944 14872
rect -4116 14792 -2944 14808
rect -4116 14728 -3028 14792
rect -2964 14728 -2944 14792
rect -4116 14712 -2944 14728
rect -4116 14648 -3028 14712
rect -2964 14648 -2944 14712
rect -4116 14632 -2944 14648
rect -4116 14568 -3028 14632
rect -2964 14568 -2944 14632
rect -4116 14552 -2944 14568
rect -4116 14488 -3028 14552
rect -2964 14488 -2944 14552
rect -4116 14472 -2944 14488
rect -4116 14408 -3028 14472
rect -2964 14408 -2944 14472
rect -4116 14392 -2944 14408
rect -4116 14328 -3028 14392
rect -2964 14328 -2944 14392
rect -4116 14312 -2944 14328
rect -4116 14248 -3028 14312
rect -2964 14248 -2944 14312
rect -4116 14232 -2944 14248
rect -4116 14168 -3028 14232
rect -2964 14168 -2944 14232
rect -4116 14120 -2944 14168
rect -2704 14952 -1532 15000
rect -2704 14888 -1616 14952
rect -1552 14888 -1532 14952
rect -2704 14872 -1532 14888
rect -2704 14808 -1616 14872
rect -1552 14808 -1532 14872
rect -2704 14792 -1532 14808
rect -2704 14728 -1616 14792
rect -1552 14728 -1532 14792
rect -2704 14712 -1532 14728
rect -2704 14648 -1616 14712
rect -1552 14648 -1532 14712
rect -2704 14632 -1532 14648
rect -2704 14568 -1616 14632
rect -1552 14568 -1532 14632
rect -2704 14552 -1532 14568
rect -2704 14488 -1616 14552
rect -1552 14488 -1532 14552
rect -2704 14472 -1532 14488
rect -2704 14408 -1616 14472
rect -1552 14408 -1532 14472
rect -2704 14392 -1532 14408
rect -2704 14328 -1616 14392
rect -1552 14328 -1532 14392
rect -2704 14312 -1532 14328
rect -2704 14248 -1616 14312
rect -1552 14248 -1532 14312
rect -2704 14232 -1532 14248
rect -2704 14168 -1616 14232
rect -1552 14168 -1532 14232
rect -2704 14120 -1532 14168
rect -1292 14952 -120 15000
rect -1292 14888 -204 14952
rect -140 14888 -120 14952
rect -1292 14872 -120 14888
rect -1292 14808 -204 14872
rect -140 14808 -120 14872
rect -1292 14792 -120 14808
rect -1292 14728 -204 14792
rect -140 14728 -120 14792
rect -1292 14712 -120 14728
rect -1292 14648 -204 14712
rect -140 14648 -120 14712
rect -1292 14632 -120 14648
rect -1292 14568 -204 14632
rect -140 14568 -120 14632
rect -1292 14552 -120 14568
rect -1292 14488 -204 14552
rect -140 14488 -120 14552
rect -1292 14472 -120 14488
rect -1292 14408 -204 14472
rect -140 14408 -120 14472
rect -1292 14392 -120 14408
rect -1292 14328 -204 14392
rect -140 14328 -120 14392
rect -1292 14312 -120 14328
rect -1292 14248 -204 14312
rect -140 14248 -120 14312
rect -1292 14232 -120 14248
rect -1292 14168 -204 14232
rect -140 14168 -120 14232
rect -1292 14120 -120 14168
rect 120 14952 1292 15000
rect 120 14888 1208 14952
rect 1272 14888 1292 14952
rect 120 14872 1292 14888
rect 120 14808 1208 14872
rect 1272 14808 1292 14872
rect 120 14792 1292 14808
rect 120 14728 1208 14792
rect 1272 14728 1292 14792
rect 120 14712 1292 14728
rect 120 14648 1208 14712
rect 1272 14648 1292 14712
rect 120 14632 1292 14648
rect 120 14568 1208 14632
rect 1272 14568 1292 14632
rect 120 14552 1292 14568
rect 120 14488 1208 14552
rect 1272 14488 1292 14552
rect 120 14472 1292 14488
rect 120 14408 1208 14472
rect 1272 14408 1292 14472
rect 120 14392 1292 14408
rect 120 14328 1208 14392
rect 1272 14328 1292 14392
rect 120 14312 1292 14328
rect 120 14248 1208 14312
rect 1272 14248 1292 14312
rect 120 14232 1292 14248
rect 120 14168 1208 14232
rect 1272 14168 1292 14232
rect 120 14120 1292 14168
rect 1532 14952 2704 15000
rect 1532 14888 2620 14952
rect 2684 14888 2704 14952
rect 1532 14872 2704 14888
rect 1532 14808 2620 14872
rect 2684 14808 2704 14872
rect 1532 14792 2704 14808
rect 1532 14728 2620 14792
rect 2684 14728 2704 14792
rect 1532 14712 2704 14728
rect 1532 14648 2620 14712
rect 2684 14648 2704 14712
rect 1532 14632 2704 14648
rect 1532 14568 2620 14632
rect 2684 14568 2704 14632
rect 1532 14552 2704 14568
rect 1532 14488 2620 14552
rect 2684 14488 2704 14552
rect 1532 14472 2704 14488
rect 1532 14408 2620 14472
rect 2684 14408 2704 14472
rect 1532 14392 2704 14408
rect 1532 14328 2620 14392
rect 2684 14328 2704 14392
rect 1532 14312 2704 14328
rect 1532 14248 2620 14312
rect 2684 14248 2704 14312
rect 1532 14232 2704 14248
rect 1532 14168 2620 14232
rect 2684 14168 2704 14232
rect 1532 14120 2704 14168
rect 2944 14952 4116 15000
rect 2944 14888 4032 14952
rect 4096 14888 4116 14952
rect 2944 14872 4116 14888
rect 2944 14808 4032 14872
rect 4096 14808 4116 14872
rect 2944 14792 4116 14808
rect 2944 14728 4032 14792
rect 4096 14728 4116 14792
rect 2944 14712 4116 14728
rect 2944 14648 4032 14712
rect 4096 14648 4116 14712
rect 2944 14632 4116 14648
rect 2944 14568 4032 14632
rect 4096 14568 4116 14632
rect 2944 14552 4116 14568
rect 2944 14488 4032 14552
rect 4096 14488 4116 14552
rect 2944 14472 4116 14488
rect 2944 14408 4032 14472
rect 4096 14408 4116 14472
rect 2944 14392 4116 14408
rect 2944 14328 4032 14392
rect 4096 14328 4116 14392
rect 2944 14312 4116 14328
rect 2944 14248 4032 14312
rect 4096 14248 4116 14312
rect 2944 14232 4116 14248
rect 2944 14168 4032 14232
rect 4096 14168 4116 14232
rect 2944 14120 4116 14168
rect 4356 14952 5528 15000
rect 4356 14888 5444 14952
rect 5508 14888 5528 14952
rect 4356 14872 5528 14888
rect 4356 14808 5444 14872
rect 5508 14808 5528 14872
rect 4356 14792 5528 14808
rect 4356 14728 5444 14792
rect 5508 14728 5528 14792
rect 4356 14712 5528 14728
rect 4356 14648 5444 14712
rect 5508 14648 5528 14712
rect 4356 14632 5528 14648
rect 4356 14568 5444 14632
rect 5508 14568 5528 14632
rect 4356 14552 5528 14568
rect 4356 14488 5444 14552
rect 5508 14488 5528 14552
rect 4356 14472 5528 14488
rect 4356 14408 5444 14472
rect 5508 14408 5528 14472
rect 4356 14392 5528 14408
rect 4356 14328 5444 14392
rect 5508 14328 5528 14392
rect 4356 14312 5528 14328
rect 4356 14248 5444 14312
rect 5508 14248 5528 14312
rect 4356 14232 5528 14248
rect 4356 14168 5444 14232
rect 5508 14168 5528 14232
rect 4356 14120 5528 14168
rect 5768 14952 6940 15000
rect 5768 14888 6856 14952
rect 6920 14888 6940 14952
rect 5768 14872 6940 14888
rect 5768 14808 6856 14872
rect 6920 14808 6940 14872
rect 5768 14792 6940 14808
rect 5768 14728 6856 14792
rect 6920 14728 6940 14792
rect 5768 14712 6940 14728
rect 5768 14648 6856 14712
rect 6920 14648 6940 14712
rect 5768 14632 6940 14648
rect 5768 14568 6856 14632
rect 6920 14568 6940 14632
rect 5768 14552 6940 14568
rect 5768 14488 6856 14552
rect 6920 14488 6940 14552
rect 5768 14472 6940 14488
rect 5768 14408 6856 14472
rect 6920 14408 6940 14472
rect 5768 14392 6940 14408
rect 5768 14328 6856 14392
rect 6920 14328 6940 14392
rect 5768 14312 6940 14328
rect 5768 14248 6856 14312
rect 6920 14248 6940 14312
rect 5768 14232 6940 14248
rect 5768 14168 6856 14232
rect 6920 14168 6940 14232
rect 5768 14120 6940 14168
rect 7180 14952 8352 15000
rect 7180 14888 8268 14952
rect 8332 14888 8352 14952
rect 7180 14872 8352 14888
rect 7180 14808 8268 14872
rect 8332 14808 8352 14872
rect 7180 14792 8352 14808
rect 7180 14728 8268 14792
rect 8332 14728 8352 14792
rect 7180 14712 8352 14728
rect 7180 14648 8268 14712
rect 8332 14648 8352 14712
rect 7180 14632 8352 14648
rect 7180 14568 8268 14632
rect 8332 14568 8352 14632
rect 7180 14552 8352 14568
rect 7180 14488 8268 14552
rect 8332 14488 8352 14552
rect 7180 14472 8352 14488
rect 7180 14408 8268 14472
rect 8332 14408 8352 14472
rect 7180 14392 8352 14408
rect 7180 14328 8268 14392
rect 8332 14328 8352 14392
rect 7180 14312 8352 14328
rect 7180 14248 8268 14312
rect 8332 14248 8352 14312
rect 7180 14232 8352 14248
rect 7180 14168 8268 14232
rect 8332 14168 8352 14232
rect 7180 14120 8352 14168
rect 8592 14952 9764 15000
rect 8592 14888 9680 14952
rect 9744 14888 9764 14952
rect 8592 14872 9764 14888
rect 8592 14808 9680 14872
rect 9744 14808 9764 14872
rect 8592 14792 9764 14808
rect 8592 14728 9680 14792
rect 9744 14728 9764 14792
rect 8592 14712 9764 14728
rect 8592 14648 9680 14712
rect 9744 14648 9764 14712
rect 8592 14632 9764 14648
rect 8592 14568 9680 14632
rect 9744 14568 9764 14632
rect 8592 14552 9764 14568
rect 8592 14488 9680 14552
rect 9744 14488 9764 14552
rect 8592 14472 9764 14488
rect 8592 14408 9680 14472
rect 9744 14408 9764 14472
rect 8592 14392 9764 14408
rect 8592 14328 9680 14392
rect 9744 14328 9764 14392
rect 8592 14312 9764 14328
rect 8592 14248 9680 14312
rect 9744 14248 9764 14312
rect 8592 14232 9764 14248
rect 8592 14168 9680 14232
rect 9744 14168 9764 14232
rect 8592 14120 9764 14168
rect 10004 14952 11176 15000
rect 10004 14888 11092 14952
rect 11156 14888 11176 14952
rect 10004 14872 11176 14888
rect 10004 14808 11092 14872
rect 11156 14808 11176 14872
rect 10004 14792 11176 14808
rect 10004 14728 11092 14792
rect 11156 14728 11176 14792
rect 10004 14712 11176 14728
rect 10004 14648 11092 14712
rect 11156 14648 11176 14712
rect 10004 14632 11176 14648
rect 10004 14568 11092 14632
rect 11156 14568 11176 14632
rect 10004 14552 11176 14568
rect 10004 14488 11092 14552
rect 11156 14488 11176 14552
rect 10004 14472 11176 14488
rect 10004 14408 11092 14472
rect 11156 14408 11176 14472
rect 10004 14392 11176 14408
rect 10004 14328 11092 14392
rect 11156 14328 11176 14392
rect 10004 14312 11176 14328
rect 10004 14248 11092 14312
rect 11156 14248 11176 14312
rect 10004 14232 11176 14248
rect 10004 14168 11092 14232
rect 11156 14168 11176 14232
rect 10004 14120 11176 14168
rect 11416 14952 12588 15000
rect 11416 14888 12504 14952
rect 12568 14888 12588 14952
rect 11416 14872 12588 14888
rect 11416 14808 12504 14872
rect 12568 14808 12588 14872
rect 11416 14792 12588 14808
rect 11416 14728 12504 14792
rect 12568 14728 12588 14792
rect 11416 14712 12588 14728
rect 11416 14648 12504 14712
rect 12568 14648 12588 14712
rect 11416 14632 12588 14648
rect 11416 14568 12504 14632
rect 12568 14568 12588 14632
rect 11416 14552 12588 14568
rect 11416 14488 12504 14552
rect 12568 14488 12588 14552
rect 11416 14472 12588 14488
rect 11416 14408 12504 14472
rect 12568 14408 12588 14472
rect 11416 14392 12588 14408
rect 11416 14328 12504 14392
rect 12568 14328 12588 14392
rect 11416 14312 12588 14328
rect 11416 14248 12504 14312
rect 12568 14248 12588 14312
rect 11416 14232 12588 14248
rect 11416 14168 12504 14232
rect 12568 14168 12588 14232
rect 11416 14120 12588 14168
rect 12828 14952 14000 15000
rect 12828 14888 13916 14952
rect 13980 14888 14000 14952
rect 12828 14872 14000 14888
rect 12828 14808 13916 14872
rect 13980 14808 14000 14872
rect 12828 14792 14000 14808
rect 12828 14728 13916 14792
rect 13980 14728 14000 14792
rect 12828 14712 14000 14728
rect 12828 14648 13916 14712
rect 13980 14648 14000 14712
rect 12828 14632 14000 14648
rect 12828 14568 13916 14632
rect 13980 14568 14000 14632
rect 12828 14552 14000 14568
rect 12828 14488 13916 14552
rect 13980 14488 14000 14552
rect 12828 14472 14000 14488
rect 12828 14408 13916 14472
rect 13980 14408 14000 14472
rect 12828 14392 14000 14408
rect 12828 14328 13916 14392
rect 13980 14328 14000 14392
rect 12828 14312 14000 14328
rect 12828 14248 13916 14312
rect 13980 14248 14000 14312
rect 12828 14232 14000 14248
rect 12828 14168 13916 14232
rect 13980 14168 14000 14232
rect 12828 14120 14000 14168
rect 14240 14952 15412 15000
rect 14240 14888 15328 14952
rect 15392 14888 15412 14952
rect 14240 14872 15412 14888
rect 14240 14808 15328 14872
rect 15392 14808 15412 14872
rect 14240 14792 15412 14808
rect 14240 14728 15328 14792
rect 15392 14728 15412 14792
rect 14240 14712 15412 14728
rect 14240 14648 15328 14712
rect 15392 14648 15412 14712
rect 14240 14632 15412 14648
rect 14240 14568 15328 14632
rect 15392 14568 15412 14632
rect 14240 14552 15412 14568
rect 14240 14488 15328 14552
rect 15392 14488 15412 14552
rect 14240 14472 15412 14488
rect 14240 14408 15328 14472
rect 15392 14408 15412 14472
rect 14240 14392 15412 14408
rect 14240 14328 15328 14392
rect 15392 14328 15412 14392
rect 14240 14312 15412 14328
rect 14240 14248 15328 14312
rect 15392 14248 15412 14312
rect 14240 14232 15412 14248
rect 14240 14168 15328 14232
rect 15392 14168 15412 14232
rect 14240 14120 15412 14168
rect 15652 14952 16824 15000
rect 15652 14888 16740 14952
rect 16804 14888 16824 14952
rect 15652 14872 16824 14888
rect 15652 14808 16740 14872
rect 16804 14808 16824 14872
rect 15652 14792 16824 14808
rect 15652 14728 16740 14792
rect 16804 14728 16824 14792
rect 15652 14712 16824 14728
rect 15652 14648 16740 14712
rect 16804 14648 16824 14712
rect 15652 14632 16824 14648
rect 15652 14568 16740 14632
rect 16804 14568 16824 14632
rect 15652 14552 16824 14568
rect 15652 14488 16740 14552
rect 16804 14488 16824 14552
rect 15652 14472 16824 14488
rect 15652 14408 16740 14472
rect 16804 14408 16824 14472
rect 15652 14392 16824 14408
rect 15652 14328 16740 14392
rect 16804 14328 16824 14392
rect 15652 14312 16824 14328
rect 15652 14248 16740 14312
rect 16804 14248 16824 14312
rect 15652 14232 16824 14248
rect 15652 14168 16740 14232
rect 16804 14168 16824 14232
rect 15652 14120 16824 14168
rect 17064 14952 18236 15000
rect 17064 14888 18152 14952
rect 18216 14888 18236 14952
rect 17064 14872 18236 14888
rect 17064 14808 18152 14872
rect 18216 14808 18236 14872
rect 17064 14792 18236 14808
rect 17064 14728 18152 14792
rect 18216 14728 18236 14792
rect 17064 14712 18236 14728
rect 17064 14648 18152 14712
rect 18216 14648 18236 14712
rect 17064 14632 18236 14648
rect 17064 14568 18152 14632
rect 18216 14568 18236 14632
rect 17064 14552 18236 14568
rect 17064 14488 18152 14552
rect 18216 14488 18236 14552
rect 17064 14472 18236 14488
rect 17064 14408 18152 14472
rect 18216 14408 18236 14472
rect 17064 14392 18236 14408
rect 17064 14328 18152 14392
rect 18216 14328 18236 14392
rect 17064 14312 18236 14328
rect 17064 14248 18152 14312
rect 18216 14248 18236 14312
rect 17064 14232 18236 14248
rect 17064 14168 18152 14232
rect 18216 14168 18236 14232
rect 17064 14120 18236 14168
rect 18476 14952 19648 15000
rect 18476 14888 19564 14952
rect 19628 14888 19648 14952
rect 18476 14872 19648 14888
rect 18476 14808 19564 14872
rect 19628 14808 19648 14872
rect 18476 14792 19648 14808
rect 18476 14728 19564 14792
rect 19628 14728 19648 14792
rect 18476 14712 19648 14728
rect 18476 14648 19564 14712
rect 19628 14648 19648 14712
rect 18476 14632 19648 14648
rect 18476 14568 19564 14632
rect 19628 14568 19648 14632
rect 18476 14552 19648 14568
rect 18476 14488 19564 14552
rect 19628 14488 19648 14552
rect 18476 14472 19648 14488
rect 18476 14408 19564 14472
rect 19628 14408 19648 14472
rect 18476 14392 19648 14408
rect 18476 14328 19564 14392
rect 19628 14328 19648 14392
rect 18476 14312 19648 14328
rect 18476 14248 19564 14312
rect 19628 14248 19648 14312
rect 18476 14232 19648 14248
rect 18476 14168 19564 14232
rect 19628 14168 19648 14232
rect 18476 14120 19648 14168
rect 19888 14952 21060 15000
rect 19888 14888 20976 14952
rect 21040 14888 21060 14952
rect 19888 14872 21060 14888
rect 19888 14808 20976 14872
rect 21040 14808 21060 14872
rect 19888 14792 21060 14808
rect 19888 14728 20976 14792
rect 21040 14728 21060 14792
rect 19888 14712 21060 14728
rect 19888 14648 20976 14712
rect 21040 14648 21060 14712
rect 19888 14632 21060 14648
rect 19888 14568 20976 14632
rect 21040 14568 21060 14632
rect 19888 14552 21060 14568
rect 19888 14488 20976 14552
rect 21040 14488 21060 14552
rect 19888 14472 21060 14488
rect 19888 14408 20976 14472
rect 21040 14408 21060 14472
rect 19888 14392 21060 14408
rect 19888 14328 20976 14392
rect 21040 14328 21060 14392
rect 19888 14312 21060 14328
rect 19888 14248 20976 14312
rect 21040 14248 21060 14312
rect 19888 14232 21060 14248
rect 19888 14168 20976 14232
rect 21040 14168 21060 14232
rect 19888 14120 21060 14168
rect 21300 14952 22472 15000
rect 21300 14888 22388 14952
rect 22452 14888 22472 14952
rect 21300 14872 22472 14888
rect 21300 14808 22388 14872
rect 22452 14808 22472 14872
rect 21300 14792 22472 14808
rect 21300 14728 22388 14792
rect 22452 14728 22472 14792
rect 21300 14712 22472 14728
rect 21300 14648 22388 14712
rect 22452 14648 22472 14712
rect 21300 14632 22472 14648
rect 21300 14568 22388 14632
rect 22452 14568 22472 14632
rect 21300 14552 22472 14568
rect 21300 14488 22388 14552
rect 22452 14488 22472 14552
rect 21300 14472 22472 14488
rect 21300 14408 22388 14472
rect 22452 14408 22472 14472
rect 21300 14392 22472 14408
rect 21300 14328 22388 14392
rect 22452 14328 22472 14392
rect 21300 14312 22472 14328
rect 21300 14248 22388 14312
rect 22452 14248 22472 14312
rect 21300 14232 22472 14248
rect 21300 14168 22388 14232
rect 22452 14168 22472 14232
rect 21300 14120 22472 14168
rect 22712 14952 23884 15000
rect 22712 14888 23800 14952
rect 23864 14888 23884 14952
rect 22712 14872 23884 14888
rect 22712 14808 23800 14872
rect 23864 14808 23884 14872
rect 22712 14792 23884 14808
rect 22712 14728 23800 14792
rect 23864 14728 23884 14792
rect 22712 14712 23884 14728
rect 22712 14648 23800 14712
rect 23864 14648 23884 14712
rect 22712 14632 23884 14648
rect 22712 14568 23800 14632
rect 23864 14568 23884 14632
rect 22712 14552 23884 14568
rect 22712 14488 23800 14552
rect 23864 14488 23884 14552
rect 22712 14472 23884 14488
rect 22712 14408 23800 14472
rect 23864 14408 23884 14472
rect 22712 14392 23884 14408
rect 22712 14328 23800 14392
rect 23864 14328 23884 14392
rect 22712 14312 23884 14328
rect 22712 14248 23800 14312
rect 23864 14248 23884 14312
rect 22712 14232 23884 14248
rect 22712 14168 23800 14232
rect 23864 14168 23884 14232
rect 22712 14120 23884 14168
rect -23884 13832 -22712 13880
rect -23884 13768 -22796 13832
rect -22732 13768 -22712 13832
rect -23884 13752 -22712 13768
rect -23884 13688 -22796 13752
rect -22732 13688 -22712 13752
rect -23884 13672 -22712 13688
rect -23884 13608 -22796 13672
rect -22732 13608 -22712 13672
rect -23884 13592 -22712 13608
rect -23884 13528 -22796 13592
rect -22732 13528 -22712 13592
rect -23884 13512 -22712 13528
rect -23884 13448 -22796 13512
rect -22732 13448 -22712 13512
rect -23884 13432 -22712 13448
rect -23884 13368 -22796 13432
rect -22732 13368 -22712 13432
rect -23884 13352 -22712 13368
rect -23884 13288 -22796 13352
rect -22732 13288 -22712 13352
rect -23884 13272 -22712 13288
rect -23884 13208 -22796 13272
rect -22732 13208 -22712 13272
rect -23884 13192 -22712 13208
rect -23884 13128 -22796 13192
rect -22732 13128 -22712 13192
rect -23884 13112 -22712 13128
rect -23884 13048 -22796 13112
rect -22732 13048 -22712 13112
rect -23884 13000 -22712 13048
rect -22472 13832 -21300 13880
rect -22472 13768 -21384 13832
rect -21320 13768 -21300 13832
rect -22472 13752 -21300 13768
rect -22472 13688 -21384 13752
rect -21320 13688 -21300 13752
rect -22472 13672 -21300 13688
rect -22472 13608 -21384 13672
rect -21320 13608 -21300 13672
rect -22472 13592 -21300 13608
rect -22472 13528 -21384 13592
rect -21320 13528 -21300 13592
rect -22472 13512 -21300 13528
rect -22472 13448 -21384 13512
rect -21320 13448 -21300 13512
rect -22472 13432 -21300 13448
rect -22472 13368 -21384 13432
rect -21320 13368 -21300 13432
rect -22472 13352 -21300 13368
rect -22472 13288 -21384 13352
rect -21320 13288 -21300 13352
rect -22472 13272 -21300 13288
rect -22472 13208 -21384 13272
rect -21320 13208 -21300 13272
rect -22472 13192 -21300 13208
rect -22472 13128 -21384 13192
rect -21320 13128 -21300 13192
rect -22472 13112 -21300 13128
rect -22472 13048 -21384 13112
rect -21320 13048 -21300 13112
rect -22472 13000 -21300 13048
rect -21060 13832 -19888 13880
rect -21060 13768 -19972 13832
rect -19908 13768 -19888 13832
rect -21060 13752 -19888 13768
rect -21060 13688 -19972 13752
rect -19908 13688 -19888 13752
rect -21060 13672 -19888 13688
rect -21060 13608 -19972 13672
rect -19908 13608 -19888 13672
rect -21060 13592 -19888 13608
rect -21060 13528 -19972 13592
rect -19908 13528 -19888 13592
rect -21060 13512 -19888 13528
rect -21060 13448 -19972 13512
rect -19908 13448 -19888 13512
rect -21060 13432 -19888 13448
rect -21060 13368 -19972 13432
rect -19908 13368 -19888 13432
rect -21060 13352 -19888 13368
rect -21060 13288 -19972 13352
rect -19908 13288 -19888 13352
rect -21060 13272 -19888 13288
rect -21060 13208 -19972 13272
rect -19908 13208 -19888 13272
rect -21060 13192 -19888 13208
rect -21060 13128 -19972 13192
rect -19908 13128 -19888 13192
rect -21060 13112 -19888 13128
rect -21060 13048 -19972 13112
rect -19908 13048 -19888 13112
rect -21060 13000 -19888 13048
rect -19648 13832 -18476 13880
rect -19648 13768 -18560 13832
rect -18496 13768 -18476 13832
rect -19648 13752 -18476 13768
rect -19648 13688 -18560 13752
rect -18496 13688 -18476 13752
rect -19648 13672 -18476 13688
rect -19648 13608 -18560 13672
rect -18496 13608 -18476 13672
rect -19648 13592 -18476 13608
rect -19648 13528 -18560 13592
rect -18496 13528 -18476 13592
rect -19648 13512 -18476 13528
rect -19648 13448 -18560 13512
rect -18496 13448 -18476 13512
rect -19648 13432 -18476 13448
rect -19648 13368 -18560 13432
rect -18496 13368 -18476 13432
rect -19648 13352 -18476 13368
rect -19648 13288 -18560 13352
rect -18496 13288 -18476 13352
rect -19648 13272 -18476 13288
rect -19648 13208 -18560 13272
rect -18496 13208 -18476 13272
rect -19648 13192 -18476 13208
rect -19648 13128 -18560 13192
rect -18496 13128 -18476 13192
rect -19648 13112 -18476 13128
rect -19648 13048 -18560 13112
rect -18496 13048 -18476 13112
rect -19648 13000 -18476 13048
rect -18236 13832 -17064 13880
rect -18236 13768 -17148 13832
rect -17084 13768 -17064 13832
rect -18236 13752 -17064 13768
rect -18236 13688 -17148 13752
rect -17084 13688 -17064 13752
rect -18236 13672 -17064 13688
rect -18236 13608 -17148 13672
rect -17084 13608 -17064 13672
rect -18236 13592 -17064 13608
rect -18236 13528 -17148 13592
rect -17084 13528 -17064 13592
rect -18236 13512 -17064 13528
rect -18236 13448 -17148 13512
rect -17084 13448 -17064 13512
rect -18236 13432 -17064 13448
rect -18236 13368 -17148 13432
rect -17084 13368 -17064 13432
rect -18236 13352 -17064 13368
rect -18236 13288 -17148 13352
rect -17084 13288 -17064 13352
rect -18236 13272 -17064 13288
rect -18236 13208 -17148 13272
rect -17084 13208 -17064 13272
rect -18236 13192 -17064 13208
rect -18236 13128 -17148 13192
rect -17084 13128 -17064 13192
rect -18236 13112 -17064 13128
rect -18236 13048 -17148 13112
rect -17084 13048 -17064 13112
rect -18236 13000 -17064 13048
rect -16824 13832 -15652 13880
rect -16824 13768 -15736 13832
rect -15672 13768 -15652 13832
rect -16824 13752 -15652 13768
rect -16824 13688 -15736 13752
rect -15672 13688 -15652 13752
rect -16824 13672 -15652 13688
rect -16824 13608 -15736 13672
rect -15672 13608 -15652 13672
rect -16824 13592 -15652 13608
rect -16824 13528 -15736 13592
rect -15672 13528 -15652 13592
rect -16824 13512 -15652 13528
rect -16824 13448 -15736 13512
rect -15672 13448 -15652 13512
rect -16824 13432 -15652 13448
rect -16824 13368 -15736 13432
rect -15672 13368 -15652 13432
rect -16824 13352 -15652 13368
rect -16824 13288 -15736 13352
rect -15672 13288 -15652 13352
rect -16824 13272 -15652 13288
rect -16824 13208 -15736 13272
rect -15672 13208 -15652 13272
rect -16824 13192 -15652 13208
rect -16824 13128 -15736 13192
rect -15672 13128 -15652 13192
rect -16824 13112 -15652 13128
rect -16824 13048 -15736 13112
rect -15672 13048 -15652 13112
rect -16824 13000 -15652 13048
rect -15412 13832 -14240 13880
rect -15412 13768 -14324 13832
rect -14260 13768 -14240 13832
rect -15412 13752 -14240 13768
rect -15412 13688 -14324 13752
rect -14260 13688 -14240 13752
rect -15412 13672 -14240 13688
rect -15412 13608 -14324 13672
rect -14260 13608 -14240 13672
rect -15412 13592 -14240 13608
rect -15412 13528 -14324 13592
rect -14260 13528 -14240 13592
rect -15412 13512 -14240 13528
rect -15412 13448 -14324 13512
rect -14260 13448 -14240 13512
rect -15412 13432 -14240 13448
rect -15412 13368 -14324 13432
rect -14260 13368 -14240 13432
rect -15412 13352 -14240 13368
rect -15412 13288 -14324 13352
rect -14260 13288 -14240 13352
rect -15412 13272 -14240 13288
rect -15412 13208 -14324 13272
rect -14260 13208 -14240 13272
rect -15412 13192 -14240 13208
rect -15412 13128 -14324 13192
rect -14260 13128 -14240 13192
rect -15412 13112 -14240 13128
rect -15412 13048 -14324 13112
rect -14260 13048 -14240 13112
rect -15412 13000 -14240 13048
rect -14000 13832 -12828 13880
rect -14000 13768 -12912 13832
rect -12848 13768 -12828 13832
rect -14000 13752 -12828 13768
rect -14000 13688 -12912 13752
rect -12848 13688 -12828 13752
rect -14000 13672 -12828 13688
rect -14000 13608 -12912 13672
rect -12848 13608 -12828 13672
rect -14000 13592 -12828 13608
rect -14000 13528 -12912 13592
rect -12848 13528 -12828 13592
rect -14000 13512 -12828 13528
rect -14000 13448 -12912 13512
rect -12848 13448 -12828 13512
rect -14000 13432 -12828 13448
rect -14000 13368 -12912 13432
rect -12848 13368 -12828 13432
rect -14000 13352 -12828 13368
rect -14000 13288 -12912 13352
rect -12848 13288 -12828 13352
rect -14000 13272 -12828 13288
rect -14000 13208 -12912 13272
rect -12848 13208 -12828 13272
rect -14000 13192 -12828 13208
rect -14000 13128 -12912 13192
rect -12848 13128 -12828 13192
rect -14000 13112 -12828 13128
rect -14000 13048 -12912 13112
rect -12848 13048 -12828 13112
rect -14000 13000 -12828 13048
rect -12588 13832 -11416 13880
rect -12588 13768 -11500 13832
rect -11436 13768 -11416 13832
rect -12588 13752 -11416 13768
rect -12588 13688 -11500 13752
rect -11436 13688 -11416 13752
rect -12588 13672 -11416 13688
rect -12588 13608 -11500 13672
rect -11436 13608 -11416 13672
rect -12588 13592 -11416 13608
rect -12588 13528 -11500 13592
rect -11436 13528 -11416 13592
rect -12588 13512 -11416 13528
rect -12588 13448 -11500 13512
rect -11436 13448 -11416 13512
rect -12588 13432 -11416 13448
rect -12588 13368 -11500 13432
rect -11436 13368 -11416 13432
rect -12588 13352 -11416 13368
rect -12588 13288 -11500 13352
rect -11436 13288 -11416 13352
rect -12588 13272 -11416 13288
rect -12588 13208 -11500 13272
rect -11436 13208 -11416 13272
rect -12588 13192 -11416 13208
rect -12588 13128 -11500 13192
rect -11436 13128 -11416 13192
rect -12588 13112 -11416 13128
rect -12588 13048 -11500 13112
rect -11436 13048 -11416 13112
rect -12588 13000 -11416 13048
rect -11176 13832 -10004 13880
rect -11176 13768 -10088 13832
rect -10024 13768 -10004 13832
rect -11176 13752 -10004 13768
rect -11176 13688 -10088 13752
rect -10024 13688 -10004 13752
rect -11176 13672 -10004 13688
rect -11176 13608 -10088 13672
rect -10024 13608 -10004 13672
rect -11176 13592 -10004 13608
rect -11176 13528 -10088 13592
rect -10024 13528 -10004 13592
rect -11176 13512 -10004 13528
rect -11176 13448 -10088 13512
rect -10024 13448 -10004 13512
rect -11176 13432 -10004 13448
rect -11176 13368 -10088 13432
rect -10024 13368 -10004 13432
rect -11176 13352 -10004 13368
rect -11176 13288 -10088 13352
rect -10024 13288 -10004 13352
rect -11176 13272 -10004 13288
rect -11176 13208 -10088 13272
rect -10024 13208 -10004 13272
rect -11176 13192 -10004 13208
rect -11176 13128 -10088 13192
rect -10024 13128 -10004 13192
rect -11176 13112 -10004 13128
rect -11176 13048 -10088 13112
rect -10024 13048 -10004 13112
rect -11176 13000 -10004 13048
rect -9764 13832 -8592 13880
rect -9764 13768 -8676 13832
rect -8612 13768 -8592 13832
rect -9764 13752 -8592 13768
rect -9764 13688 -8676 13752
rect -8612 13688 -8592 13752
rect -9764 13672 -8592 13688
rect -9764 13608 -8676 13672
rect -8612 13608 -8592 13672
rect -9764 13592 -8592 13608
rect -9764 13528 -8676 13592
rect -8612 13528 -8592 13592
rect -9764 13512 -8592 13528
rect -9764 13448 -8676 13512
rect -8612 13448 -8592 13512
rect -9764 13432 -8592 13448
rect -9764 13368 -8676 13432
rect -8612 13368 -8592 13432
rect -9764 13352 -8592 13368
rect -9764 13288 -8676 13352
rect -8612 13288 -8592 13352
rect -9764 13272 -8592 13288
rect -9764 13208 -8676 13272
rect -8612 13208 -8592 13272
rect -9764 13192 -8592 13208
rect -9764 13128 -8676 13192
rect -8612 13128 -8592 13192
rect -9764 13112 -8592 13128
rect -9764 13048 -8676 13112
rect -8612 13048 -8592 13112
rect -9764 13000 -8592 13048
rect -8352 13832 -7180 13880
rect -8352 13768 -7264 13832
rect -7200 13768 -7180 13832
rect -8352 13752 -7180 13768
rect -8352 13688 -7264 13752
rect -7200 13688 -7180 13752
rect -8352 13672 -7180 13688
rect -8352 13608 -7264 13672
rect -7200 13608 -7180 13672
rect -8352 13592 -7180 13608
rect -8352 13528 -7264 13592
rect -7200 13528 -7180 13592
rect -8352 13512 -7180 13528
rect -8352 13448 -7264 13512
rect -7200 13448 -7180 13512
rect -8352 13432 -7180 13448
rect -8352 13368 -7264 13432
rect -7200 13368 -7180 13432
rect -8352 13352 -7180 13368
rect -8352 13288 -7264 13352
rect -7200 13288 -7180 13352
rect -8352 13272 -7180 13288
rect -8352 13208 -7264 13272
rect -7200 13208 -7180 13272
rect -8352 13192 -7180 13208
rect -8352 13128 -7264 13192
rect -7200 13128 -7180 13192
rect -8352 13112 -7180 13128
rect -8352 13048 -7264 13112
rect -7200 13048 -7180 13112
rect -8352 13000 -7180 13048
rect -6940 13832 -5768 13880
rect -6940 13768 -5852 13832
rect -5788 13768 -5768 13832
rect -6940 13752 -5768 13768
rect -6940 13688 -5852 13752
rect -5788 13688 -5768 13752
rect -6940 13672 -5768 13688
rect -6940 13608 -5852 13672
rect -5788 13608 -5768 13672
rect -6940 13592 -5768 13608
rect -6940 13528 -5852 13592
rect -5788 13528 -5768 13592
rect -6940 13512 -5768 13528
rect -6940 13448 -5852 13512
rect -5788 13448 -5768 13512
rect -6940 13432 -5768 13448
rect -6940 13368 -5852 13432
rect -5788 13368 -5768 13432
rect -6940 13352 -5768 13368
rect -6940 13288 -5852 13352
rect -5788 13288 -5768 13352
rect -6940 13272 -5768 13288
rect -6940 13208 -5852 13272
rect -5788 13208 -5768 13272
rect -6940 13192 -5768 13208
rect -6940 13128 -5852 13192
rect -5788 13128 -5768 13192
rect -6940 13112 -5768 13128
rect -6940 13048 -5852 13112
rect -5788 13048 -5768 13112
rect -6940 13000 -5768 13048
rect -5528 13832 -4356 13880
rect -5528 13768 -4440 13832
rect -4376 13768 -4356 13832
rect -5528 13752 -4356 13768
rect -5528 13688 -4440 13752
rect -4376 13688 -4356 13752
rect -5528 13672 -4356 13688
rect -5528 13608 -4440 13672
rect -4376 13608 -4356 13672
rect -5528 13592 -4356 13608
rect -5528 13528 -4440 13592
rect -4376 13528 -4356 13592
rect -5528 13512 -4356 13528
rect -5528 13448 -4440 13512
rect -4376 13448 -4356 13512
rect -5528 13432 -4356 13448
rect -5528 13368 -4440 13432
rect -4376 13368 -4356 13432
rect -5528 13352 -4356 13368
rect -5528 13288 -4440 13352
rect -4376 13288 -4356 13352
rect -5528 13272 -4356 13288
rect -5528 13208 -4440 13272
rect -4376 13208 -4356 13272
rect -5528 13192 -4356 13208
rect -5528 13128 -4440 13192
rect -4376 13128 -4356 13192
rect -5528 13112 -4356 13128
rect -5528 13048 -4440 13112
rect -4376 13048 -4356 13112
rect -5528 13000 -4356 13048
rect -4116 13832 -2944 13880
rect -4116 13768 -3028 13832
rect -2964 13768 -2944 13832
rect -4116 13752 -2944 13768
rect -4116 13688 -3028 13752
rect -2964 13688 -2944 13752
rect -4116 13672 -2944 13688
rect -4116 13608 -3028 13672
rect -2964 13608 -2944 13672
rect -4116 13592 -2944 13608
rect -4116 13528 -3028 13592
rect -2964 13528 -2944 13592
rect -4116 13512 -2944 13528
rect -4116 13448 -3028 13512
rect -2964 13448 -2944 13512
rect -4116 13432 -2944 13448
rect -4116 13368 -3028 13432
rect -2964 13368 -2944 13432
rect -4116 13352 -2944 13368
rect -4116 13288 -3028 13352
rect -2964 13288 -2944 13352
rect -4116 13272 -2944 13288
rect -4116 13208 -3028 13272
rect -2964 13208 -2944 13272
rect -4116 13192 -2944 13208
rect -4116 13128 -3028 13192
rect -2964 13128 -2944 13192
rect -4116 13112 -2944 13128
rect -4116 13048 -3028 13112
rect -2964 13048 -2944 13112
rect -4116 13000 -2944 13048
rect -2704 13832 -1532 13880
rect -2704 13768 -1616 13832
rect -1552 13768 -1532 13832
rect -2704 13752 -1532 13768
rect -2704 13688 -1616 13752
rect -1552 13688 -1532 13752
rect -2704 13672 -1532 13688
rect -2704 13608 -1616 13672
rect -1552 13608 -1532 13672
rect -2704 13592 -1532 13608
rect -2704 13528 -1616 13592
rect -1552 13528 -1532 13592
rect -2704 13512 -1532 13528
rect -2704 13448 -1616 13512
rect -1552 13448 -1532 13512
rect -2704 13432 -1532 13448
rect -2704 13368 -1616 13432
rect -1552 13368 -1532 13432
rect -2704 13352 -1532 13368
rect -2704 13288 -1616 13352
rect -1552 13288 -1532 13352
rect -2704 13272 -1532 13288
rect -2704 13208 -1616 13272
rect -1552 13208 -1532 13272
rect -2704 13192 -1532 13208
rect -2704 13128 -1616 13192
rect -1552 13128 -1532 13192
rect -2704 13112 -1532 13128
rect -2704 13048 -1616 13112
rect -1552 13048 -1532 13112
rect -2704 13000 -1532 13048
rect -1292 13832 -120 13880
rect -1292 13768 -204 13832
rect -140 13768 -120 13832
rect -1292 13752 -120 13768
rect -1292 13688 -204 13752
rect -140 13688 -120 13752
rect -1292 13672 -120 13688
rect -1292 13608 -204 13672
rect -140 13608 -120 13672
rect -1292 13592 -120 13608
rect -1292 13528 -204 13592
rect -140 13528 -120 13592
rect -1292 13512 -120 13528
rect -1292 13448 -204 13512
rect -140 13448 -120 13512
rect -1292 13432 -120 13448
rect -1292 13368 -204 13432
rect -140 13368 -120 13432
rect -1292 13352 -120 13368
rect -1292 13288 -204 13352
rect -140 13288 -120 13352
rect -1292 13272 -120 13288
rect -1292 13208 -204 13272
rect -140 13208 -120 13272
rect -1292 13192 -120 13208
rect -1292 13128 -204 13192
rect -140 13128 -120 13192
rect -1292 13112 -120 13128
rect -1292 13048 -204 13112
rect -140 13048 -120 13112
rect -1292 13000 -120 13048
rect 120 13832 1292 13880
rect 120 13768 1208 13832
rect 1272 13768 1292 13832
rect 120 13752 1292 13768
rect 120 13688 1208 13752
rect 1272 13688 1292 13752
rect 120 13672 1292 13688
rect 120 13608 1208 13672
rect 1272 13608 1292 13672
rect 120 13592 1292 13608
rect 120 13528 1208 13592
rect 1272 13528 1292 13592
rect 120 13512 1292 13528
rect 120 13448 1208 13512
rect 1272 13448 1292 13512
rect 120 13432 1292 13448
rect 120 13368 1208 13432
rect 1272 13368 1292 13432
rect 120 13352 1292 13368
rect 120 13288 1208 13352
rect 1272 13288 1292 13352
rect 120 13272 1292 13288
rect 120 13208 1208 13272
rect 1272 13208 1292 13272
rect 120 13192 1292 13208
rect 120 13128 1208 13192
rect 1272 13128 1292 13192
rect 120 13112 1292 13128
rect 120 13048 1208 13112
rect 1272 13048 1292 13112
rect 120 13000 1292 13048
rect 1532 13832 2704 13880
rect 1532 13768 2620 13832
rect 2684 13768 2704 13832
rect 1532 13752 2704 13768
rect 1532 13688 2620 13752
rect 2684 13688 2704 13752
rect 1532 13672 2704 13688
rect 1532 13608 2620 13672
rect 2684 13608 2704 13672
rect 1532 13592 2704 13608
rect 1532 13528 2620 13592
rect 2684 13528 2704 13592
rect 1532 13512 2704 13528
rect 1532 13448 2620 13512
rect 2684 13448 2704 13512
rect 1532 13432 2704 13448
rect 1532 13368 2620 13432
rect 2684 13368 2704 13432
rect 1532 13352 2704 13368
rect 1532 13288 2620 13352
rect 2684 13288 2704 13352
rect 1532 13272 2704 13288
rect 1532 13208 2620 13272
rect 2684 13208 2704 13272
rect 1532 13192 2704 13208
rect 1532 13128 2620 13192
rect 2684 13128 2704 13192
rect 1532 13112 2704 13128
rect 1532 13048 2620 13112
rect 2684 13048 2704 13112
rect 1532 13000 2704 13048
rect 2944 13832 4116 13880
rect 2944 13768 4032 13832
rect 4096 13768 4116 13832
rect 2944 13752 4116 13768
rect 2944 13688 4032 13752
rect 4096 13688 4116 13752
rect 2944 13672 4116 13688
rect 2944 13608 4032 13672
rect 4096 13608 4116 13672
rect 2944 13592 4116 13608
rect 2944 13528 4032 13592
rect 4096 13528 4116 13592
rect 2944 13512 4116 13528
rect 2944 13448 4032 13512
rect 4096 13448 4116 13512
rect 2944 13432 4116 13448
rect 2944 13368 4032 13432
rect 4096 13368 4116 13432
rect 2944 13352 4116 13368
rect 2944 13288 4032 13352
rect 4096 13288 4116 13352
rect 2944 13272 4116 13288
rect 2944 13208 4032 13272
rect 4096 13208 4116 13272
rect 2944 13192 4116 13208
rect 2944 13128 4032 13192
rect 4096 13128 4116 13192
rect 2944 13112 4116 13128
rect 2944 13048 4032 13112
rect 4096 13048 4116 13112
rect 2944 13000 4116 13048
rect 4356 13832 5528 13880
rect 4356 13768 5444 13832
rect 5508 13768 5528 13832
rect 4356 13752 5528 13768
rect 4356 13688 5444 13752
rect 5508 13688 5528 13752
rect 4356 13672 5528 13688
rect 4356 13608 5444 13672
rect 5508 13608 5528 13672
rect 4356 13592 5528 13608
rect 4356 13528 5444 13592
rect 5508 13528 5528 13592
rect 4356 13512 5528 13528
rect 4356 13448 5444 13512
rect 5508 13448 5528 13512
rect 4356 13432 5528 13448
rect 4356 13368 5444 13432
rect 5508 13368 5528 13432
rect 4356 13352 5528 13368
rect 4356 13288 5444 13352
rect 5508 13288 5528 13352
rect 4356 13272 5528 13288
rect 4356 13208 5444 13272
rect 5508 13208 5528 13272
rect 4356 13192 5528 13208
rect 4356 13128 5444 13192
rect 5508 13128 5528 13192
rect 4356 13112 5528 13128
rect 4356 13048 5444 13112
rect 5508 13048 5528 13112
rect 4356 13000 5528 13048
rect 5768 13832 6940 13880
rect 5768 13768 6856 13832
rect 6920 13768 6940 13832
rect 5768 13752 6940 13768
rect 5768 13688 6856 13752
rect 6920 13688 6940 13752
rect 5768 13672 6940 13688
rect 5768 13608 6856 13672
rect 6920 13608 6940 13672
rect 5768 13592 6940 13608
rect 5768 13528 6856 13592
rect 6920 13528 6940 13592
rect 5768 13512 6940 13528
rect 5768 13448 6856 13512
rect 6920 13448 6940 13512
rect 5768 13432 6940 13448
rect 5768 13368 6856 13432
rect 6920 13368 6940 13432
rect 5768 13352 6940 13368
rect 5768 13288 6856 13352
rect 6920 13288 6940 13352
rect 5768 13272 6940 13288
rect 5768 13208 6856 13272
rect 6920 13208 6940 13272
rect 5768 13192 6940 13208
rect 5768 13128 6856 13192
rect 6920 13128 6940 13192
rect 5768 13112 6940 13128
rect 5768 13048 6856 13112
rect 6920 13048 6940 13112
rect 5768 13000 6940 13048
rect 7180 13832 8352 13880
rect 7180 13768 8268 13832
rect 8332 13768 8352 13832
rect 7180 13752 8352 13768
rect 7180 13688 8268 13752
rect 8332 13688 8352 13752
rect 7180 13672 8352 13688
rect 7180 13608 8268 13672
rect 8332 13608 8352 13672
rect 7180 13592 8352 13608
rect 7180 13528 8268 13592
rect 8332 13528 8352 13592
rect 7180 13512 8352 13528
rect 7180 13448 8268 13512
rect 8332 13448 8352 13512
rect 7180 13432 8352 13448
rect 7180 13368 8268 13432
rect 8332 13368 8352 13432
rect 7180 13352 8352 13368
rect 7180 13288 8268 13352
rect 8332 13288 8352 13352
rect 7180 13272 8352 13288
rect 7180 13208 8268 13272
rect 8332 13208 8352 13272
rect 7180 13192 8352 13208
rect 7180 13128 8268 13192
rect 8332 13128 8352 13192
rect 7180 13112 8352 13128
rect 7180 13048 8268 13112
rect 8332 13048 8352 13112
rect 7180 13000 8352 13048
rect 8592 13832 9764 13880
rect 8592 13768 9680 13832
rect 9744 13768 9764 13832
rect 8592 13752 9764 13768
rect 8592 13688 9680 13752
rect 9744 13688 9764 13752
rect 8592 13672 9764 13688
rect 8592 13608 9680 13672
rect 9744 13608 9764 13672
rect 8592 13592 9764 13608
rect 8592 13528 9680 13592
rect 9744 13528 9764 13592
rect 8592 13512 9764 13528
rect 8592 13448 9680 13512
rect 9744 13448 9764 13512
rect 8592 13432 9764 13448
rect 8592 13368 9680 13432
rect 9744 13368 9764 13432
rect 8592 13352 9764 13368
rect 8592 13288 9680 13352
rect 9744 13288 9764 13352
rect 8592 13272 9764 13288
rect 8592 13208 9680 13272
rect 9744 13208 9764 13272
rect 8592 13192 9764 13208
rect 8592 13128 9680 13192
rect 9744 13128 9764 13192
rect 8592 13112 9764 13128
rect 8592 13048 9680 13112
rect 9744 13048 9764 13112
rect 8592 13000 9764 13048
rect 10004 13832 11176 13880
rect 10004 13768 11092 13832
rect 11156 13768 11176 13832
rect 10004 13752 11176 13768
rect 10004 13688 11092 13752
rect 11156 13688 11176 13752
rect 10004 13672 11176 13688
rect 10004 13608 11092 13672
rect 11156 13608 11176 13672
rect 10004 13592 11176 13608
rect 10004 13528 11092 13592
rect 11156 13528 11176 13592
rect 10004 13512 11176 13528
rect 10004 13448 11092 13512
rect 11156 13448 11176 13512
rect 10004 13432 11176 13448
rect 10004 13368 11092 13432
rect 11156 13368 11176 13432
rect 10004 13352 11176 13368
rect 10004 13288 11092 13352
rect 11156 13288 11176 13352
rect 10004 13272 11176 13288
rect 10004 13208 11092 13272
rect 11156 13208 11176 13272
rect 10004 13192 11176 13208
rect 10004 13128 11092 13192
rect 11156 13128 11176 13192
rect 10004 13112 11176 13128
rect 10004 13048 11092 13112
rect 11156 13048 11176 13112
rect 10004 13000 11176 13048
rect 11416 13832 12588 13880
rect 11416 13768 12504 13832
rect 12568 13768 12588 13832
rect 11416 13752 12588 13768
rect 11416 13688 12504 13752
rect 12568 13688 12588 13752
rect 11416 13672 12588 13688
rect 11416 13608 12504 13672
rect 12568 13608 12588 13672
rect 11416 13592 12588 13608
rect 11416 13528 12504 13592
rect 12568 13528 12588 13592
rect 11416 13512 12588 13528
rect 11416 13448 12504 13512
rect 12568 13448 12588 13512
rect 11416 13432 12588 13448
rect 11416 13368 12504 13432
rect 12568 13368 12588 13432
rect 11416 13352 12588 13368
rect 11416 13288 12504 13352
rect 12568 13288 12588 13352
rect 11416 13272 12588 13288
rect 11416 13208 12504 13272
rect 12568 13208 12588 13272
rect 11416 13192 12588 13208
rect 11416 13128 12504 13192
rect 12568 13128 12588 13192
rect 11416 13112 12588 13128
rect 11416 13048 12504 13112
rect 12568 13048 12588 13112
rect 11416 13000 12588 13048
rect 12828 13832 14000 13880
rect 12828 13768 13916 13832
rect 13980 13768 14000 13832
rect 12828 13752 14000 13768
rect 12828 13688 13916 13752
rect 13980 13688 14000 13752
rect 12828 13672 14000 13688
rect 12828 13608 13916 13672
rect 13980 13608 14000 13672
rect 12828 13592 14000 13608
rect 12828 13528 13916 13592
rect 13980 13528 14000 13592
rect 12828 13512 14000 13528
rect 12828 13448 13916 13512
rect 13980 13448 14000 13512
rect 12828 13432 14000 13448
rect 12828 13368 13916 13432
rect 13980 13368 14000 13432
rect 12828 13352 14000 13368
rect 12828 13288 13916 13352
rect 13980 13288 14000 13352
rect 12828 13272 14000 13288
rect 12828 13208 13916 13272
rect 13980 13208 14000 13272
rect 12828 13192 14000 13208
rect 12828 13128 13916 13192
rect 13980 13128 14000 13192
rect 12828 13112 14000 13128
rect 12828 13048 13916 13112
rect 13980 13048 14000 13112
rect 12828 13000 14000 13048
rect 14240 13832 15412 13880
rect 14240 13768 15328 13832
rect 15392 13768 15412 13832
rect 14240 13752 15412 13768
rect 14240 13688 15328 13752
rect 15392 13688 15412 13752
rect 14240 13672 15412 13688
rect 14240 13608 15328 13672
rect 15392 13608 15412 13672
rect 14240 13592 15412 13608
rect 14240 13528 15328 13592
rect 15392 13528 15412 13592
rect 14240 13512 15412 13528
rect 14240 13448 15328 13512
rect 15392 13448 15412 13512
rect 14240 13432 15412 13448
rect 14240 13368 15328 13432
rect 15392 13368 15412 13432
rect 14240 13352 15412 13368
rect 14240 13288 15328 13352
rect 15392 13288 15412 13352
rect 14240 13272 15412 13288
rect 14240 13208 15328 13272
rect 15392 13208 15412 13272
rect 14240 13192 15412 13208
rect 14240 13128 15328 13192
rect 15392 13128 15412 13192
rect 14240 13112 15412 13128
rect 14240 13048 15328 13112
rect 15392 13048 15412 13112
rect 14240 13000 15412 13048
rect 15652 13832 16824 13880
rect 15652 13768 16740 13832
rect 16804 13768 16824 13832
rect 15652 13752 16824 13768
rect 15652 13688 16740 13752
rect 16804 13688 16824 13752
rect 15652 13672 16824 13688
rect 15652 13608 16740 13672
rect 16804 13608 16824 13672
rect 15652 13592 16824 13608
rect 15652 13528 16740 13592
rect 16804 13528 16824 13592
rect 15652 13512 16824 13528
rect 15652 13448 16740 13512
rect 16804 13448 16824 13512
rect 15652 13432 16824 13448
rect 15652 13368 16740 13432
rect 16804 13368 16824 13432
rect 15652 13352 16824 13368
rect 15652 13288 16740 13352
rect 16804 13288 16824 13352
rect 15652 13272 16824 13288
rect 15652 13208 16740 13272
rect 16804 13208 16824 13272
rect 15652 13192 16824 13208
rect 15652 13128 16740 13192
rect 16804 13128 16824 13192
rect 15652 13112 16824 13128
rect 15652 13048 16740 13112
rect 16804 13048 16824 13112
rect 15652 13000 16824 13048
rect 17064 13832 18236 13880
rect 17064 13768 18152 13832
rect 18216 13768 18236 13832
rect 17064 13752 18236 13768
rect 17064 13688 18152 13752
rect 18216 13688 18236 13752
rect 17064 13672 18236 13688
rect 17064 13608 18152 13672
rect 18216 13608 18236 13672
rect 17064 13592 18236 13608
rect 17064 13528 18152 13592
rect 18216 13528 18236 13592
rect 17064 13512 18236 13528
rect 17064 13448 18152 13512
rect 18216 13448 18236 13512
rect 17064 13432 18236 13448
rect 17064 13368 18152 13432
rect 18216 13368 18236 13432
rect 17064 13352 18236 13368
rect 17064 13288 18152 13352
rect 18216 13288 18236 13352
rect 17064 13272 18236 13288
rect 17064 13208 18152 13272
rect 18216 13208 18236 13272
rect 17064 13192 18236 13208
rect 17064 13128 18152 13192
rect 18216 13128 18236 13192
rect 17064 13112 18236 13128
rect 17064 13048 18152 13112
rect 18216 13048 18236 13112
rect 17064 13000 18236 13048
rect 18476 13832 19648 13880
rect 18476 13768 19564 13832
rect 19628 13768 19648 13832
rect 18476 13752 19648 13768
rect 18476 13688 19564 13752
rect 19628 13688 19648 13752
rect 18476 13672 19648 13688
rect 18476 13608 19564 13672
rect 19628 13608 19648 13672
rect 18476 13592 19648 13608
rect 18476 13528 19564 13592
rect 19628 13528 19648 13592
rect 18476 13512 19648 13528
rect 18476 13448 19564 13512
rect 19628 13448 19648 13512
rect 18476 13432 19648 13448
rect 18476 13368 19564 13432
rect 19628 13368 19648 13432
rect 18476 13352 19648 13368
rect 18476 13288 19564 13352
rect 19628 13288 19648 13352
rect 18476 13272 19648 13288
rect 18476 13208 19564 13272
rect 19628 13208 19648 13272
rect 18476 13192 19648 13208
rect 18476 13128 19564 13192
rect 19628 13128 19648 13192
rect 18476 13112 19648 13128
rect 18476 13048 19564 13112
rect 19628 13048 19648 13112
rect 18476 13000 19648 13048
rect 19888 13832 21060 13880
rect 19888 13768 20976 13832
rect 21040 13768 21060 13832
rect 19888 13752 21060 13768
rect 19888 13688 20976 13752
rect 21040 13688 21060 13752
rect 19888 13672 21060 13688
rect 19888 13608 20976 13672
rect 21040 13608 21060 13672
rect 19888 13592 21060 13608
rect 19888 13528 20976 13592
rect 21040 13528 21060 13592
rect 19888 13512 21060 13528
rect 19888 13448 20976 13512
rect 21040 13448 21060 13512
rect 19888 13432 21060 13448
rect 19888 13368 20976 13432
rect 21040 13368 21060 13432
rect 19888 13352 21060 13368
rect 19888 13288 20976 13352
rect 21040 13288 21060 13352
rect 19888 13272 21060 13288
rect 19888 13208 20976 13272
rect 21040 13208 21060 13272
rect 19888 13192 21060 13208
rect 19888 13128 20976 13192
rect 21040 13128 21060 13192
rect 19888 13112 21060 13128
rect 19888 13048 20976 13112
rect 21040 13048 21060 13112
rect 19888 13000 21060 13048
rect 21300 13832 22472 13880
rect 21300 13768 22388 13832
rect 22452 13768 22472 13832
rect 21300 13752 22472 13768
rect 21300 13688 22388 13752
rect 22452 13688 22472 13752
rect 21300 13672 22472 13688
rect 21300 13608 22388 13672
rect 22452 13608 22472 13672
rect 21300 13592 22472 13608
rect 21300 13528 22388 13592
rect 22452 13528 22472 13592
rect 21300 13512 22472 13528
rect 21300 13448 22388 13512
rect 22452 13448 22472 13512
rect 21300 13432 22472 13448
rect 21300 13368 22388 13432
rect 22452 13368 22472 13432
rect 21300 13352 22472 13368
rect 21300 13288 22388 13352
rect 22452 13288 22472 13352
rect 21300 13272 22472 13288
rect 21300 13208 22388 13272
rect 22452 13208 22472 13272
rect 21300 13192 22472 13208
rect 21300 13128 22388 13192
rect 22452 13128 22472 13192
rect 21300 13112 22472 13128
rect 21300 13048 22388 13112
rect 22452 13048 22472 13112
rect 21300 13000 22472 13048
rect 22712 13832 23884 13880
rect 22712 13768 23800 13832
rect 23864 13768 23884 13832
rect 22712 13752 23884 13768
rect 22712 13688 23800 13752
rect 23864 13688 23884 13752
rect 22712 13672 23884 13688
rect 22712 13608 23800 13672
rect 23864 13608 23884 13672
rect 22712 13592 23884 13608
rect 22712 13528 23800 13592
rect 23864 13528 23884 13592
rect 22712 13512 23884 13528
rect 22712 13448 23800 13512
rect 23864 13448 23884 13512
rect 22712 13432 23884 13448
rect 22712 13368 23800 13432
rect 23864 13368 23884 13432
rect 22712 13352 23884 13368
rect 22712 13288 23800 13352
rect 23864 13288 23884 13352
rect 22712 13272 23884 13288
rect 22712 13208 23800 13272
rect 23864 13208 23884 13272
rect 22712 13192 23884 13208
rect 22712 13128 23800 13192
rect 23864 13128 23884 13192
rect 22712 13112 23884 13128
rect 22712 13048 23800 13112
rect 23864 13048 23884 13112
rect 22712 13000 23884 13048
rect -23884 12712 -22712 12760
rect -23884 12648 -22796 12712
rect -22732 12648 -22712 12712
rect -23884 12632 -22712 12648
rect -23884 12568 -22796 12632
rect -22732 12568 -22712 12632
rect -23884 12552 -22712 12568
rect -23884 12488 -22796 12552
rect -22732 12488 -22712 12552
rect -23884 12472 -22712 12488
rect -23884 12408 -22796 12472
rect -22732 12408 -22712 12472
rect -23884 12392 -22712 12408
rect -23884 12328 -22796 12392
rect -22732 12328 -22712 12392
rect -23884 12312 -22712 12328
rect -23884 12248 -22796 12312
rect -22732 12248 -22712 12312
rect -23884 12232 -22712 12248
rect -23884 12168 -22796 12232
rect -22732 12168 -22712 12232
rect -23884 12152 -22712 12168
rect -23884 12088 -22796 12152
rect -22732 12088 -22712 12152
rect -23884 12072 -22712 12088
rect -23884 12008 -22796 12072
rect -22732 12008 -22712 12072
rect -23884 11992 -22712 12008
rect -23884 11928 -22796 11992
rect -22732 11928 -22712 11992
rect -23884 11880 -22712 11928
rect -22472 12712 -21300 12760
rect -22472 12648 -21384 12712
rect -21320 12648 -21300 12712
rect -22472 12632 -21300 12648
rect -22472 12568 -21384 12632
rect -21320 12568 -21300 12632
rect -22472 12552 -21300 12568
rect -22472 12488 -21384 12552
rect -21320 12488 -21300 12552
rect -22472 12472 -21300 12488
rect -22472 12408 -21384 12472
rect -21320 12408 -21300 12472
rect -22472 12392 -21300 12408
rect -22472 12328 -21384 12392
rect -21320 12328 -21300 12392
rect -22472 12312 -21300 12328
rect -22472 12248 -21384 12312
rect -21320 12248 -21300 12312
rect -22472 12232 -21300 12248
rect -22472 12168 -21384 12232
rect -21320 12168 -21300 12232
rect -22472 12152 -21300 12168
rect -22472 12088 -21384 12152
rect -21320 12088 -21300 12152
rect -22472 12072 -21300 12088
rect -22472 12008 -21384 12072
rect -21320 12008 -21300 12072
rect -22472 11992 -21300 12008
rect -22472 11928 -21384 11992
rect -21320 11928 -21300 11992
rect -22472 11880 -21300 11928
rect -21060 12712 -19888 12760
rect -21060 12648 -19972 12712
rect -19908 12648 -19888 12712
rect -21060 12632 -19888 12648
rect -21060 12568 -19972 12632
rect -19908 12568 -19888 12632
rect -21060 12552 -19888 12568
rect -21060 12488 -19972 12552
rect -19908 12488 -19888 12552
rect -21060 12472 -19888 12488
rect -21060 12408 -19972 12472
rect -19908 12408 -19888 12472
rect -21060 12392 -19888 12408
rect -21060 12328 -19972 12392
rect -19908 12328 -19888 12392
rect -21060 12312 -19888 12328
rect -21060 12248 -19972 12312
rect -19908 12248 -19888 12312
rect -21060 12232 -19888 12248
rect -21060 12168 -19972 12232
rect -19908 12168 -19888 12232
rect -21060 12152 -19888 12168
rect -21060 12088 -19972 12152
rect -19908 12088 -19888 12152
rect -21060 12072 -19888 12088
rect -21060 12008 -19972 12072
rect -19908 12008 -19888 12072
rect -21060 11992 -19888 12008
rect -21060 11928 -19972 11992
rect -19908 11928 -19888 11992
rect -21060 11880 -19888 11928
rect -19648 12712 -18476 12760
rect -19648 12648 -18560 12712
rect -18496 12648 -18476 12712
rect -19648 12632 -18476 12648
rect -19648 12568 -18560 12632
rect -18496 12568 -18476 12632
rect -19648 12552 -18476 12568
rect -19648 12488 -18560 12552
rect -18496 12488 -18476 12552
rect -19648 12472 -18476 12488
rect -19648 12408 -18560 12472
rect -18496 12408 -18476 12472
rect -19648 12392 -18476 12408
rect -19648 12328 -18560 12392
rect -18496 12328 -18476 12392
rect -19648 12312 -18476 12328
rect -19648 12248 -18560 12312
rect -18496 12248 -18476 12312
rect -19648 12232 -18476 12248
rect -19648 12168 -18560 12232
rect -18496 12168 -18476 12232
rect -19648 12152 -18476 12168
rect -19648 12088 -18560 12152
rect -18496 12088 -18476 12152
rect -19648 12072 -18476 12088
rect -19648 12008 -18560 12072
rect -18496 12008 -18476 12072
rect -19648 11992 -18476 12008
rect -19648 11928 -18560 11992
rect -18496 11928 -18476 11992
rect -19648 11880 -18476 11928
rect -18236 12712 -17064 12760
rect -18236 12648 -17148 12712
rect -17084 12648 -17064 12712
rect -18236 12632 -17064 12648
rect -18236 12568 -17148 12632
rect -17084 12568 -17064 12632
rect -18236 12552 -17064 12568
rect -18236 12488 -17148 12552
rect -17084 12488 -17064 12552
rect -18236 12472 -17064 12488
rect -18236 12408 -17148 12472
rect -17084 12408 -17064 12472
rect -18236 12392 -17064 12408
rect -18236 12328 -17148 12392
rect -17084 12328 -17064 12392
rect -18236 12312 -17064 12328
rect -18236 12248 -17148 12312
rect -17084 12248 -17064 12312
rect -18236 12232 -17064 12248
rect -18236 12168 -17148 12232
rect -17084 12168 -17064 12232
rect -18236 12152 -17064 12168
rect -18236 12088 -17148 12152
rect -17084 12088 -17064 12152
rect -18236 12072 -17064 12088
rect -18236 12008 -17148 12072
rect -17084 12008 -17064 12072
rect -18236 11992 -17064 12008
rect -18236 11928 -17148 11992
rect -17084 11928 -17064 11992
rect -18236 11880 -17064 11928
rect -16824 12712 -15652 12760
rect -16824 12648 -15736 12712
rect -15672 12648 -15652 12712
rect -16824 12632 -15652 12648
rect -16824 12568 -15736 12632
rect -15672 12568 -15652 12632
rect -16824 12552 -15652 12568
rect -16824 12488 -15736 12552
rect -15672 12488 -15652 12552
rect -16824 12472 -15652 12488
rect -16824 12408 -15736 12472
rect -15672 12408 -15652 12472
rect -16824 12392 -15652 12408
rect -16824 12328 -15736 12392
rect -15672 12328 -15652 12392
rect -16824 12312 -15652 12328
rect -16824 12248 -15736 12312
rect -15672 12248 -15652 12312
rect -16824 12232 -15652 12248
rect -16824 12168 -15736 12232
rect -15672 12168 -15652 12232
rect -16824 12152 -15652 12168
rect -16824 12088 -15736 12152
rect -15672 12088 -15652 12152
rect -16824 12072 -15652 12088
rect -16824 12008 -15736 12072
rect -15672 12008 -15652 12072
rect -16824 11992 -15652 12008
rect -16824 11928 -15736 11992
rect -15672 11928 -15652 11992
rect -16824 11880 -15652 11928
rect -15412 12712 -14240 12760
rect -15412 12648 -14324 12712
rect -14260 12648 -14240 12712
rect -15412 12632 -14240 12648
rect -15412 12568 -14324 12632
rect -14260 12568 -14240 12632
rect -15412 12552 -14240 12568
rect -15412 12488 -14324 12552
rect -14260 12488 -14240 12552
rect -15412 12472 -14240 12488
rect -15412 12408 -14324 12472
rect -14260 12408 -14240 12472
rect -15412 12392 -14240 12408
rect -15412 12328 -14324 12392
rect -14260 12328 -14240 12392
rect -15412 12312 -14240 12328
rect -15412 12248 -14324 12312
rect -14260 12248 -14240 12312
rect -15412 12232 -14240 12248
rect -15412 12168 -14324 12232
rect -14260 12168 -14240 12232
rect -15412 12152 -14240 12168
rect -15412 12088 -14324 12152
rect -14260 12088 -14240 12152
rect -15412 12072 -14240 12088
rect -15412 12008 -14324 12072
rect -14260 12008 -14240 12072
rect -15412 11992 -14240 12008
rect -15412 11928 -14324 11992
rect -14260 11928 -14240 11992
rect -15412 11880 -14240 11928
rect -14000 12712 -12828 12760
rect -14000 12648 -12912 12712
rect -12848 12648 -12828 12712
rect -14000 12632 -12828 12648
rect -14000 12568 -12912 12632
rect -12848 12568 -12828 12632
rect -14000 12552 -12828 12568
rect -14000 12488 -12912 12552
rect -12848 12488 -12828 12552
rect -14000 12472 -12828 12488
rect -14000 12408 -12912 12472
rect -12848 12408 -12828 12472
rect -14000 12392 -12828 12408
rect -14000 12328 -12912 12392
rect -12848 12328 -12828 12392
rect -14000 12312 -12828 12328
rect -14000 12248 -12912 12312
rect -12848 12248 -12828 12312
rect -14000 12232 -12828 12248
rect -14000 12168 -12912 12232
rect -12848 12168 -12828 12232
rect -14000 12152 -12828 12168
rect -14000 12088 -12912 12152
rect -12848 12088 -12828 12152
rect -14000 12072 -12828 12088
rect -14000 12008 -12912 12072
rect -12848 12008 -12828 12072
rect -14000 11992 -12828 12008
rect -14000 11928 -12912 11992
rect -12848 11928 -12828 11992
rect -14000 11880 -12828 11928
rect -12588 12712 -11416 12760
rect -12588 12648 -11500 12712
rect -11436 12648 -11416 12712
rect -12588 12632 -11416 12648
rect -12588 12568 -11500 12632
rect -11436 12568 -11416 12632
rect -12588 12552 -11416 12568
rect -12588 12488 -11500 12552
rect -11436 12488 -11416 12552
rect -12588 12472 -11416 12488
rect -12588 12408 -11500 12472
rect -11436 12408 -11416 12472
rect -12588 12392 -11416 12408
rect -12588 12328 -11500 12392
rect -11436 12328 -11416 12392
rect -12588 12312 -11416 12328
rect -12588 12248 -11500 12312
rect -11436 12248 -11416 12312
rect -12588 12232 -11416 12248
rect -12588 12168 -11500 12232
rect -11436 12168 -11416 12232
rect -12588 12152 -11416 12168
rect -12588 12088 -11500 12152
rect -11436 12088 -11416 12152
rect -12588 12072 -11416 12088
rect -12588 12008 -11500 12072
rect -11436 12008 -11416 12072
rect -12588 11992 -11416 12008
rect -12588 11928 -11500 11992
rect -11436 11928 -11416 11992
rect -12588 11880 -11416 11928
rect -11176 12712 -10004 12760
rect -11176 12648 -10088 12712
rect -10024 12648 -10004 12712
rect -11176 12632 -10004 12648
rect -11176 12568 -10088 12632
rect -10024 12568 -10004 12632
rect -11176 12552 -10004 12568
rect -11176 12488 -10088 12552
rect -10024 12488 -10004 12552
rect -11176 12472 -10004 12488
rect -11176 12408 -10088 12472
rect -10024 12408 -10004 12472
rect -11176 12392 -10004 12408
rect -11176 12328 -10088 12392
rect -10024 12328 -10004 12392
rect -11176 12312 -10004 12328
rect -11176 12248 -10088 12312
rect -10024 12248 -10004 12312
rect -11176 12232 -10004 12248
rect -11176 12168 -10088 12232
rect -10024 12168 -10004 12232
rect -11176 12152 -10004 12168
rect -11176 12088 -10088 12152
rect -10024 12088 -10004 12152
rect -11176 12072 -10004 12088
rect -11176 12008 -10088 12072
rect -10024 12008 -10004 12072
rect -11176 11992 -10004 12008
rect -11176 11928 -10088 11992
rect -10024 11928 -10004 11992
rect -11176 11880 -10004 11928
rect -9764 12712 -8592 12760
rect -9764 12648 -8676 12712
rect -8612 12648 -8592 12712
rect -9764 12632 -8592 12648
rect -9764 12568 -8676 12632
rect -8612 12568 -8592 12632
rect -9764 12552 -8592 12568
rect -9764 12488 -8676 12552
rect -8612 12488 -8592 12552
rect -9764 12472 -8592 12488
rect -9764 12408 -8676 12472
rect -8612 12408 -8592 12472
rect -9764 12392 -8592 12408
rect -9764 12328 -8676 12392
rect -8612 12328 -8592 12392
rect -9764 12312 -8592 12328
rect -9764 12248 -8676 12312
rect -8612 12248 -8592 12312
rect -9764 12232 -8592 12248
rect -9764 12168 -8676 12232
rect -8612 12168 -8592 12232
rect -9764 12152 -8592 12168
rect -9764 12088 -8676 12152
rect -8612 12088 -8592 12152
rect -9764 12072 -8592 12088
rect -9764 12008 -8676 12072
rect -8612 12008 -8592 12072
rect -9764 11992 -8592 12008
rect -9764 11928 -8676 11992
rect -8612 11928 -8592 11992
rect -9764 11880 -8592 11928
rect -8352 12712 -7180 12760
rect -8352 12648 -7264 12712
rect -7200 12648 -7180 12712
rect -8352 12632 -7180 12648
rect -8352 12568 -7264 12632
rect -7200 12568 -7180 12632
rect -8352 12552 -7180 12568
rect -8352 12488 -7264 12552
rect -7200 12488 -7180 12552
rect -8352 12472 -7180 12488
rect -8352 12408 -7264 12472
rect -7200 12408 -7180 12472
rect -8352 12392 -7180 12408
rect -8352 12328 -7264 12392
rect -7200 12328 -7180 12392
rect -8352 12312 -7180 12328
rect -8352 12248 -7264 12312
rect -7200 12248 -7180 12312
rect -8352 12232 -7180 12248
rect -8352 12168 -7264 12232
rect -7200 12168 -7180 12232
rect -8352 12152 -7180 12168
rect -8352 12088 -7264 12152
rect -7200 12088 -7180 12152
rect -8352 12072 -7180 12088
rect -8352 12008 -7264 12072
rect -7200 12008 -7180 12072
rect -8352 11992 -7180 12008
rect -8352 11928 -7264 11992
rect -7200 11928 -7180 11992
rect -8352 11880 -7180 11928
rect -6940 12712 -5768 12760
rect -6940 12648 -5852 12712
rect -5788 12648 -5768 12712
rect -6940 12632 -5768 12648
rect -6940 12568 -5852 12632
rect -5788 12568 -5768 12632
rect -6940 12552 -5768 12568
rect -6940 12488 -5852 12552
rect -5788 12488 -5768 12552
rect -6940 12472 -5768 12488
rect -6940 12408 -5852 12472
rect -5788 12408 -5768 12472
rect -6940 12392 -5768 12408
rect -6940 12328 -5852 12392
rect -5788 12328 -5768 12392
rect -6940 12312 -5768 12328
rect -6940 12248 -5852 12312
rect -5788 12248 -5768 12312
rect -6940 12232 -5768 12248
rect -6940 12168 -5852 12232
rect -5788 12168 -5768 12232
rect -6940 12152 -5768 12168
rect -6940 12088 -5852 12152
rect -5788 12088 -5768 12152
rect -6940 12072 -5768 12088
rect -6940 12008 -5852 12072
rect -5788 12008 -5768 12072
rect -6940 11992 -5768 12008
rect -6940 11928 -5852 11992
rect -5788 11928 -5768 11992
rect -6940 11880 -5768 11928
rect -5528 12712 -4356 12760
rect -5528 12648 -4440 12712
rect -4376 12648 -4356 12712
rect -5528 12632 -4356 12648
rect -5528 12568 -4440 12632
rect -4376 12568 -4356 12632
rect -5528 12552 -4356 12568
rect -5528 12488 -4440 12552
rect -4376 12488 -4356 12552
rect -5528 12472 -4356 12488
rect -5528 12408 -4440 12472
rect -4376 12408 -4356 12472
rect -5528 12392 -4356 12408
rect -5528 12328 -4440 12392
rect -4376 12328 -4356 12392
rect -5528 12312 -4356 12328
rect -5528 12248 -4440 12312
rect -4376 12248 -4356 12312
rect -5528 12232 -4356 12248
rect -5528 12168 -4440 12232
rect -4376 12168 -4356 12232
rect -5528 12152 -4356 12168
rect -5528 12088 -4440 12152
rect -4376 12088 -4356 12152
rect -5528 12072 -4356 12088
rect -5528 12008 -4440 12072
rect -4376 12008 -4356 12072
rect -5528 11992 -4356 12008
rect -5528 11928 -4440 11992
rect -4376 11928 -4356 11992
rect -5528 11880 -4356 11928
rect -4116 12712 -2944 12760
rect -4116 12648 -3028 12712
rect -2964 12648 -2944 12712
rect -4116 12632 -2944 12648
rect -4116 12568 -3028 12632
rect -2964 12568 -2944 12632
rect -4116 12552 -2944 12568
rect -4116 12488 -3028 12552
rect -2964 12488 -2944 12552
rect -4116 12472 -2944 12488
rect -4116 12408 -3028 12472
rect -2964 12408 -2944 12472
rect -4116 12392 -2944 12408
rect -4116 12328 -3028 12392
rect -2964 12328 -2944 12392
rect -4116 12312 -2944 12328
rect -4116 12248 -3028 12312
rect -2964 12248 -2944 12312
rect -4116 12232 -2944 12248
rect -4116 12168 -3028 12232
rect -2964 12168 -2944 12232
rect -4116 12152 -2944 12168
rect -4116 12088 -3028 12152
rect -2964 12088 -2944 12152
rect -4116 12072 -2944 12088
rect -4116 12008 -3028 12072
rect -2964 12008 -2944 12072
rect -4116 11992 -2944 12008
rect -4116 11928 -3028 11992
rect -2964 11928 -2944 11992
rect -4116 11880 -2944 11928
rect -2704 12712 -1532 12760
rect -2704 12648 -1616 12712
rect -1552 12648 -1532 12712
rect -2704 12632 -1532 12648
rect -2704 12568 -1616 12632
rect -1552 12568 -1532 12632
rect -2704 12552 -1532 12568
rect -2704 12488 -1616 12552
rect -1552 12488 -1532 12552
rect -2704 12472 -1532 12488
rect -2704 12408 -1616 12472
rect -1552 12408 -1532 12472
rect -2704 12392 -1532 12408
rect -2704 12328 -1616 12392
rect -1552 12328 -1532 12392
rect -2704 12312 -1532 12328
rect -2704 12248 -1616 12312
rect -1552 12248 -1532 12312
rect -2704 12232 -1532 12248
rect -2704 12168 -1616 12232
rect -1552 12168 -1532 12232
rect -2704 12152 -1532 12168
rect -2704 12088 -1616 12152
rect -1552 12088 -1532 12152
rect -2704 12072 -1532 12088
rect -2704 12008 -1616 12072
rect -1552 12008 -1532 12072
rect -2704 11992 -1532 12008
rect -2704 11928 -1616 11992
rect -1552 11928 -1532 11992
rect -2704 11880 -1532 11928
rect -1292 12712 -120 12760
rect -1292 12648 -204 12712
rect -140 12648 -120 12712
rect -1292 12632 -120 12648
rect -1292 12568 -204 12632
rect -140 12568 -120 12632
rect -1292 12552 -120 12568
rect -1292 12488 -204 12552
rect -140 12488 -120 12552
rect -1292 12472 -120 12488
rect -1292 12408 -204 12472
rect -140 12408 -120 12472
rect -1292 12392 -120 12408
rect -1292 12328 -204 12392
rect -140 12328 -120 12392
rect -1292 12312 -120 12328
rect -1292 12248 -204 12312
rect -140 12248 -120 12312
rect -1292 12232 -120 12248
rect -1292 12168 -204 12232
rect -140 12168 -120 12232
rect -1292 12152 -120 12168
rect -1292 12088 -204 12152
rect -140 12088 -120 12152
rect -1292 12072 -120 12088
rect -1292 12008 -204 12072
rect -140 12008 -120 12072
rect -1292 11992 -120 12008
rect -1292 11928 -204 11992
rect -140 11928 -120 11992
rect -1292 11880 -120 11928
rect 120 12712 1292 12760
rect 120 12648 1208 12712
rect 1272 12648 1292 12712
rect 120 12632 1292 12648
rect 120 12568 1208 12632
rect 1272 12568 1292 12632
rect 120 12552 1292 12568
rect 120 12488 1208 12552
rect 1272 12488 1292 12552
rect 120 12472 1292 12488
rect 120 12408 1208 12472
rect 1272 12408 1292 12472
rect 120 12392 1292 12408
rect 120 12328 1208 12392
rect 1272 12328 1292 12392
rect 120 12312 1292 12328
rect 120 12248 1208 12312
rect 1272 12248 1292 12312
rect 120 12232 1292 12248
rect 120 12168 1208 12232
rect 1272 12168 1292 12232
rect 120 12152 1292 12168
rect 120 12088 1208 12152
rect 1272 12088 1292 12152
rect 120 12072 1292 12088
rect 120 12008 1208 12072
rect 1272 12008 1292 12072
rect 120 11992 1292 12008
rect 120 11928 1208 11992
rect 1272 11928 1292 11992
rect 120 11880 1292 11928
rect 1532 12712 2704 12760
rect 1532 12648 2620 12712
rect 2684 12648 2704 12712
rect 1532 12632 2704 12648
rect 1532 12568 2620 12632
rect 2684 12568 2704 12632
rect 1532 12552 2704 12568
rect 1532 12488 2620 12552
rect 2684 12488 2704 12552
rect 1532 12472 2704 12488
rect 1532 12408 2620 12472
rect 2684 12408 2704 12472
rect 1532 12392 2704 12408
rect 1532 12328 2620 12392
rect 2684 12328 2704 12392
rect 1532 12312 2704 12328
rect 1532 12248 2620 12312
rect 2684 12248 2704 12312
rect 1532 12232 2704 12248
rect 1532 12168 2620 12232
rect 2684 12168 2704 12232
rect 1532 12152 2704 12168
rect 1532 12088 2620 12152
rect 2684 12088 2704 12152
rect 1532 12072 2704 12088
rect 1532 12008 2620 12072
rect 2684 12008 2704 12072
rect 1532 11992 2704 12008
rect 1532 11928 2620 11992
rect 2684 11928 2704 11992
rect 1532 11880 2704 11928
rect 2944 12712 4116 12760
rect 2944 12648 4032 12712
rect 4096 12648 4116 12712
rect 2944 12632 4116 12648
rect 2944 12568 4032 12632
rect 4096 12568 4116 12632
rect 2944 12552 4116 12568
rect 2944 12488 4032 12552
rect 4096 12488 4116 12552
rect 2944 12472 4116 12488
rect 2944 12408 4032 12472
rect 4096 12408 4116 12472
rect 2944 12392 4116 12408
rect 2944 12328 4032 12392
rect 4096 12328 4116 12392
rect 2944 12312 4116 12328
rect 2944 12248 4032 12312
rect 4096 12248 4116 12312
rect 2944 12232 4116 12248
rect 2944 12168 4032 12232
rect 4096 12168 4116 12232
rect 2944 12152 4116 12168
rect 2944 12088 4032 12152
rect 4096 12088 4116 12152
rect 2944 12072 4116 12088
rect 2944 12008 4032 12072
rect 4096 12008 4116 12072
rect 2944 11992 4116 12008
rect 2944 11928 4032 11992
rect 4096 11928 4116 11992
rect 2944 11880 4116 11928
rect 4356 12712 5528 12760
rect 4356 12648 5444 12712
rect 5508 12648 5528 12712
rect 4356 12632 5528 12648
rect 4356 12568 5444 12632
rect 5508 12568 5528 12632
rect 4356 12552 5528 12568
rect 4356 12488 5444 12552
rect 5508 12488 5528 12552
rect 4356 12472 5528 12488
rect 4356 12408 5444 12472
rect 5508 12408 5528 12472
rect 4356 12392 5528 12408
rect 4356 12328 5444 12392
rect 5508 12328 5528 12392
rect 4356 12312 5528 12328
rect 4356 12248 5444 12312
rect 5508 12248 5528 12312
rect 4356 12232 5528 12248
rect 4356 12168 5444 12232
rect 5508 12168 5528 12232
rect 4356 12152 5528 12168
rect 4356 12088 5444 12152
rect 5508 12088 5528 12152
rect 4356 12072 5528 12088
rect 4356 12008 5444 12072
rect 5508 12008 5528 12072
rect 4356 11992 5528 12008
rect 4356 11928 5444 11992
rect 5508 11928 5528 11992
rect 4356 11880 5528 11928
rect 5768 12712 6940 12760
rect 5768 12648 6856 12712
rect 6920 12648 6940 12712
rect 5768 12632 6940 12648
rect 5768 12568 6856 12632
rect 6920 12568 6940 12632
rect 5768 12552 6940 12568
rect 5768 12488 6856 12552
rect 6920 12488 6940 12552
rect 5768 12472 6940 12488
rect 5768 12408 6856 12472
rect 6920 12408 6940 12472
rect 5768 12392 6940 12408
rect 5768 12328 6856 12392
rect 6920 12328 6940 12392
rect 5768 12312 6940 12328
rect 5768 12248 6856 12312
rect 6920 12248 6940 12312
rect 5768 12232 6940 12248
rect 5768 12168 6856 12232
rect 6920 12168 6940 12232
rect 5768 12152 6940 12168
rect 5768 12088 6856 12152
rect 6920 12088 6940 12152
rect 5768 12072 6940 12088
rect 5768 12008 6856 12072
rect 6920 12008 6940 12072
rect 5768 11992 6940 12008
rect 5768 11928 6856 11992
rect 6920 11928 6940 11992
rect 5768 11880 6940 11928
rect 7180 12712 8352 12760
rect 7180 12648 8268 12712
rect 8332 12648 8352 12712
rect 7180 12632 8352 12648
rect 7180 12568 8268 12632
rect 8332 12568 8352 12632
rect 7180 12552 8352 12568
rect 7180 12488 8268 12552
rect 8332 12488 8352 12552
rect 7180 12472 8352 12488
rect 7180 12408 8268 12472
rect 8332 12408 8352 12472
rect 7180 12392 8352 12408
rect 7180 12328 8268 12392
rect 8332 12328 8352 12392
rect 7180 12312 8352 12328
rect 7180 12248 8268 12312
rect 8332 12248 8352 12312
rect 7180 12232 8352 12248
rect 7180 12168 8268 12232
rect 8332 12168 8352 12232
rect 7180 12152 8352 12168
rect 7180 12088 8268 12152
rect 8332 12088 8352 12152
rect 7180 12072 8352 12088
rect 7180 12008 8268 12072
rect 8332 12008 8352 12072
rect 7180 11992 8352 12008
rect 7180 11928 8268 11992
rect 8332 11928 8352 11992
rect 7180 11880 8352 11928
rect 8592 12712 9764 12760
rect 8592 12648 9680 12712
rect 9744 12648 9764 12712
rect 8592 12632 9764 12648
rect 8592 12568 9680 12632
rect 9744 12568 9764 12632
rect 8592 12552 9764 12568
rect 8592 12488 9680 12552
rect 9744 12488 9764 12552
rect 8592 12472 9764 12488
rect 8592 12408 9680 12472
rect 9744 12408 9764 12472
rect 8592 12392 9764 12408
rect 8592 12328 9680 12392
rect 9744 12328 9764 12392
rect 8592 12312 9764 12328
rect 8592 12248 9680 12312
rect 9744 12248 9764 12312
rect 8592 12232 9764 12248
rect 8592 12168 9680 12232
rect 9744 12168 9764 12232
rect 8592 12152 9764 12168
rect 8592 12088 9680 12152
rect 9744 12088 9764 12152
rect 8592 12072 9764 12088
rect 8592 12008 9680 12072
rect 9744 12008 9764 12072
rect 8592 11992 9764 12008
rect 8592 11928 9680 11992
rect 9744 11928 9764 11992
rect 8592 11880 9764 11928
rect 10004 12712 11176 12760
rect 10004 12648 11092 12712
rect 11156 12648 11176 12712
rect 10004 12632 11176 12648
rect 10004 12568 11092 12632
rect 11156 12568 11176 12632
rect 10004 12552 11176 12568
rect 10004 12488 11092 12552
rect 11156 12488 11176 12552
rect 10004 12472 11176 12488
rect 10004 12408 11092 12472
rect 11156 12408 11176 12472
rect 10004 12392 11176 12408
rect 10004 12328 11092 12392
rect 11156 12328 11176 12392
rect 10004 12312 11176 12328
rect 10004 12248 11092 12312
rect 11156 12248 11176 12312
rect 10004 12232 11176 12248
rect 10004 12168 11092 12232
rect 11156 12168 11176 12232
rect 10004 12152 11176 12168
rect 10004 12088 11092 12152
rect 11156 12088 11176 12152
rect 10004 12072 11176 12088
rect 10004 12008 11092 12072
rect 11156 12008 11176 12072
rect 10004 11992 11176 12008
rect 10004 11928 11092 11992
rect 11156 11928 11176 11992
rect 10004 11880 11176 11928
rect 11416 12712 12588 12760
rect 11416 12648 12504 12712
rect 12568 12648 12588 12712
rect 11416 12632 12588 12648
rect 11416 12568 12504 12632
rect 12568 12568 12588 12632
rect 11416 12552 12588 12568
rect 11416 12488 12504 12552
rect 12568 12488 12588 12552
rect 11416 12472 12588 12488
rect 11416 12408 12504 12472
rect 12568 12408 12588 12472
rect 11416 12392 12588 12408
rect 11416 12328 12504 12392
rect 12568 12328 12588 12392
rect 11416 12312 12588 12328
rect 11416 12248 12504 12312
rect 12568 12248 12588 12312
rect 11416 12232 12588 12248
rect 11416 12168 12504 12232
rect 12568 12168 12588 12232
rect 11416 12152 12588 12168
rect 11416 12088 12504 12152
rect 12568 12088 12588 12152
rect 11416 12072 12588 12088
rect 11416 12008 12504 12072
rect 12568 12008 12588 12072
rect 11416 11992 12588 12008
rect 11416 11928 12504 11992
rect 12568 11928 12588 11992
rect 11416 11880 12588 11928
rect 12828 12712 14000 12760
rect 12828 12648 13916 12712
rect 13980 12648 14000 12712
rect 12828 12632 14000 12648
rect 12828 12568 13916 12632
rect 13980 12568 14000 12632
rect 12828 12552 14000 12568
rect 12828 12488 13916 12552
rect 13980 12488 14000 12552
rect 12828 12472 14000 12488
rect 12828 12408 13916 12472
rect 13980 12408 14000 12472
rect 12828 12392 14000 12408
rect 12828 12328 13916 12392
rect 13980 12328 14000 12392
rect 12828 12312 14000 12328
rect 12828 12248 13916 12312
rect 13980 12248 14000 12312
rect 12828 12232 14000 12248
rect 12828 12168 13916 12232
rect 13980 12168 14000 12232
rect 12828 12152 14000 12168
rect 12828 12088 13916 12152
rect 13980 12088 14000 12152
rect 12828 12072 14000 12088
rect 12828 12008 13916 12072
rect 13980 12008 14000 12072
rect 12828 11992 14000 12008
rect 12828 11928 13916 11992
rect 13980 11928 14000 11992
rect 12828 11880 14000 11928
rect 14240 12712 15412 12760
rect 14240 12648 15328 12712
rect 15392 12648 15412 12712
rect 14240 12632 15412 12648
rect 14240 12568 15328 12632
rect 15392 12568 15412 12632
rect 14240 12552 15412 12568
rect 14240 12488 15328 12552
rect 15392 12488 15412 12552
rect 14240 12472 15412 12488
rect 14240 12408 15328 12472
rect 15392 12408 15412 12472
rect 14240 12392 15412 12408
rect 14240 12328 15328 12392
rect 15392 12328 15412 12392
rect 14240 12312 15412 12328
rect 14240 12248 15328 12312
rect 15392 12248 15412 12312
rect 14240 12232 15412 12248
rect 14240 12168 15328 12232
rect 15392 12168 15412 12232
rect 14240 12152 15412 12168
rect 14240 12088 15328 12152
rect 15392 12088 15412 12152
rect 14240 12072 15412 12088
rect 14240 12008 15328 12072
rect 15392 12008 15412 12072
rect 14240 11992 15412 12008
rect 14240 11928 15328 11992
rect 15392 11928 15412 11992
rect 14240 11880 15412 11928
rect 15652 12712 16824 12760
rect 15652 12648 16740 12712
rect 16804 12648 16824 12712
rect 15652 12632 16824 12648
rect 15652 12568 16740 12632
rect 16804 12568 16824 12632
rect 15652 12552 16824 12568
rect 15652 12488 16740 12552
rect 16804 12488 16824 12552
rect 15652 12472 16824 12488
rect 15652 12408 16740 12472
rect 16804 12408 16824 12472
rect 15652 12392 16824 12408
rect 15652 12328 16740 12392
rect 16804 12328 16824 12392
rect 15652 12312 16824 12328
rect 15652 12248 16740 12312
rect 16804 12248 16824 12312
rect 15652 12232 16824 12248
rect 15652 12168 16740 12232
rect 16804 12168 16824 12232
rect 15652 12152 16824 12168
rect 15652 12088 16740 12152
rect 16804 12088 16824 12152
rect 15652 12072 16824 12088
rect 15652 12008 16740 12072
rect 16804 12008 16824 12072
rect 15652 11992 16824 12008
rect 15652 11928 16740 11992
rect 16804 11928 16824 11992
rect 15652 11880 16824 11928
rect 17064 12712 18236 12760
rect 17064 12648 18152 12712
rect 18216 12648 18236 12712
rect 17064 12632 18236 12648
rect 17064 12568 18152 12632
rect 18216 12568 18236 12632
rect 17064 12552 18236 12568
rect 17064 12488 18152 12552
rect 18216 12488 18236 12552
rect 17064 12472 18236 12488
rect 17064 12408 18152 12472
rect 18216 12408 18236 12472
rect 17064 12392 18236 12408
rect 17064 12328 18152 12392
rect 18216 12328 18236 12392
rect 17064 12312 18236 12328
rect 17064 12248 18152 12312
rect 18216 12248 18236 12312
rect 17064 12232 18236 12248
rect 17064 12168 18152 12232
rect 18216 12168 18236 12232
rect 17064 12152 18236 12168
rect 17064 12088 18152 12152
rect 18216 12088 18236 12152
rect 17064 12072 18236 12088
rect 17064 12008 18152 12072
rect 18216 12008 18236 12072
rect 17064 11992 18236 12008
rect 17064 11928 18152 11992
rect 18216 11928 18236 11992
rect 17064 11880 18236 11928
rect 18476 12712 19648 12760
rect 18476 12648 19564 12712
rect 19628 12648 19648 12712
rect 18476 12632 19648 12648
rect 18476 12568 19564 12632
rect 19628 12568 19648 12632
rect 18476 12552 19648 12568
rect 18476 12488 19564 12552
rect 19628 12488 19648 12552
rect 18476 12472 19648 12488
rect 18476 12408 19564 12472
rect 19628 12408 19648 12472
rect 18476 12392 19648 12408
rect 18476 12328 19564 12392
rect 19628 12328 19648 12392
rect 18476 12312 19648 12328
rect 18476 12248 19564 12312
rect 19628 12248 19648 12312
rect 18476 12232 19648 12248
rect 18476 12168 19564 12232
rect 19628 12168 19648 12232
rect 18476 12152 19648 12168
rect 18476 12088 19564 12152
rect 19628 12088 19648 12152
rect 18476 12072 19648 12088
rect 18476 12008 19564 12072
rect 19628 12008 19648 12072
rect 18476 11992 19648 12008
rect 18476 11928 19564 11992
rect 19628 11928 19648 11992
rect 18476 11880 19648 11928
rect 19888 12712 21060 12760
rect 19888 12648 20976 12712
rect 21040 12648 21060 12712
rect 19888 12632 21060 12648
rect 19888 12568 20976 12632
rect 21040 12568 21060 12632
rect 19888 12552 21060 12568
rect 19888 12488 20976 12552
rect 21040 12488 21060 12552
rect 19888 12472 21060 12488
rect 19888 12408 20976 12472
rect 21040 12408 21060 12472
rect 19888 12392 21060 12408
rect 19888 12328 20976 12392
rect 21040 12328 21060 12392
rect 19888 12312 21060 12328
rect 19888 12248 20976 12312
rect 21040 12248 21060 12312
rect 19888 12232 21060 12248
rect 19888 12168 20976 12232
rect 21040 12168 21060 12232
rect 19888 12152 21060 12168
rect 19888 12088 20976 12152
rect 21040 12088 21060 12152
rect 19888 12072 21060 12088
rect 19888 12008 20976 12072
rect 21040 12008 21060 12072
rect 19888 11992 21060 12008
rect 19888 11928 20976 11992
rect 21040 11928 21060 11992
rect 19888 11880 21060 11928
rect 21300 12712 22472 12760
rect 21300 12648 22388 12712
rect 22452 12648 22472 12712
rect 21300 12632 22472 12648
rect 21300 12568 22388 12632
rect 22452 12568 22472 12632
rect 21300 12552 22472 12568
rect 21300 12488 22388 12552
rect 22452 12488 22472 12552
rect 21300 12472 22472 12488
rect 21300 12408 22388 12472
rect 22452 12408 22472 12472
rect 21300 12392 22472 12408
rect 21300 12328 22388 12392
rect 22452 12328 22472 12392
rect 21300 12312 22472 12328
rect 21300 12248 22388 12312
rect 22452 12248 22472 12312
rect 21300 12232 22472 12248
rect 21300 12168 22388 12232
rect 22452 12168 22472 12232
rect 21300 12152 22472 12168
rect 21300 12088 22388 12152
rect 22452 12088 22472 12152
rect 21300 12072 22472 12088
rect 21300 12008 22388 12072
rect 22452 12008 22472 12072
rect 21300 11992 22472 12008
rect 21300 11928 22388 11992
rect 22452 11928 22472 11992
rect 21300 11880 22472 11928
rect 22712 12712 23884 12760
rect 22712 12648 23800 12712
rect 23864 12648 23884 12712
rect 22712 12632 23884 12648
rect 22712 12568 23800 12632
rect 23864 12568 23884 12632
rect 22712 12552 23884 12568
rect 22712 12488 23800 12552
rect 23864 12488 23884 12552
rect 22712 12472 23884 12488
rect 22712 12408 23800 12472
rect 23864 12408 23884 12472
rect 22712 12392 23884 12408
rect 22712 12328 23800 12392
rect 23864 12328 23884 12392
rect 22712 12312 23884 12328
rect 22712 12248 23800 12312
rect 23864 12248 23884 12312
rect 22712 12232 23884 12248
rect 22712 12168 23800 12232
rect 23864 12168 23884 12232
rect 22712 12152 23884 12168
rect 22712 12088 23800 12152
rect 23864 12088 23884 12152
rect 22712 12072 23884 12088
rect 22712 12008 23800 12072
rect 23864 12008 23884 12072
rect 22712 11992 23884 12008
rect 22712 11928 23800 11992
rect 23864 11928 23884 11992
rect 22712 11880 23884 11928
rect -23884 11592 -22712 11640
rect -23884 11528 -22796 11592
rect -22732 11528 -22712 11592
rect -23884 11512 -22712 11528
rect -23884 11448 -22796 11512
rect -22732 11448 -22712 11512
rect -23884 11432 -22712 11448
rect -23884 11368 -22796 11432
rect -22732 11368 -22712 11432
rect -23884 11352 -22712 11368
rect -23884 11288 -22796 11352
rect -22732 11288 -22712 11352
rect -23884 11272 -22712 11288
rect -23884 11208 -22796 11272
rect -22732 11208 -22712 11272
rect -23884 11192 -22712 11208
rect -23884 11128 -22796 11192
rect -22732 11128 -22712 11192
rect -23884 11112 -22712 11128
rect -23884 11048 -22796 11112
rect -22732 11048 -22712 11112
rect -23884 11032 -22712 11048
rect -23884 10968 -22796 11032
rect -22732 10968 -22712 11032
rect -23884 10952 -22712 10968
rect -23884 10888 -22796 10952
rect -22732 10888 -22712 10952
rect -23884 10872 -22712 10888
rect -23884 10808 -22796 10872
rect -22732 10808 -22712 10872
rect -23884 10760 -22712 10808
rect -22472 11592 -21300 11640
rect -22472 11528 -21384 11592
rect -21320 11528 -21300 11592
rect -22472 11512 -21300 11528
rect -22472 11448 -21384 11512
rect -21320 11448 -21300 11512
rect -22472 11432 -21300 11448
rect -22472 11368 -21384 11432
rect -21320 11368 -21300 11432
rect -22472 11352 -21300 11368
rect -22472 11288 -21384 11352
rect -21320 11288 -21300 11352
rect -22472 11272 -21300 11288
rect -22472 11208 -21384 11272
rect -21320 11208 -21300 11272
rect -22472 11192 -21300 11208
rect -22472 11128 -21384 11192
rect -21320 11128 -21300 11192
rect -22472 11112 -21300 11128
rect -22472 11048 -21384 11112
rect -21320 11048 -21300 11112
rect -22472 11032 -21300 11048
rect -22472 10968 -21384 11032
rect -21320 10968 -21300 11032
rect -22472 10952 -21300 10968
rect -22472 10888 -21384 10952
rect -21320 10888 -21300 10952
rect -22472 10872 -21300 10888
rect -22472 10808 -21384 10872
rect -21320 10808 -21300 10872
rect -22472 10760 -21300 10808
rect -21060 11592 -19888 11640
rect -21060 11528 -19972 11592
rect -19908 11528 -19888 11592
rect -21060 11512 -19888 11528
rect -21060 11448 -19972 11512
rect -19908 11448 -19888 11512
rect -21060 11432 -19888 11448
rect -21060 11368 -19972 11432
rect -19908 11368 -19888 11432
rect -21060 11352 -19888 11368
rect -21060 11288 -19972 11352
rect -19908 11288 -19888 11352
rect -21060 11272 -19888 11288
rect -21060 11208 -19972 11272
rect -19908 11208 -19888 11272
rect -21060 11192 -19888 11208
rect -21060 11128 -19972 11192
rect -19908 11128 -19888 11192
rect -21060 11112 -19888 11128
rect -21060 11048 -19972 11112
rect -19908 11048 -19888 11112
rect -21060 11032 -19888 11048
rect -21060 10968 -19972 11032
rect -19908 10968 -19888 11032
rect -21060 10952 -19888 10968
rect -21060 10888 -19972 10952
rect -19908 10888 -19888 10952
rect -21060 10872 -19888 10888
rect -21060 10808 -19972 10872
rect -19908 10808 -19888 10872
rect -21060 10760 -19888 10808
rect -19648 11592 -18476 11640
rect -19648 11528 -18560 11592
rect -18496 11528 -18476 11592
rect -19648 11512 -18476 11528
rect -19648 11448 -18560 11512
rect -18496 11448 -18476 11512
rect -19648 11432 -18476 11448
rect -19648 11368 -18560 11432
rect -18496 11368 -18476 11432
rect -19648 11352 -18476 11368
rect -19648 11288 -18560 11352
rect -18496 11288 -18476 11352
rect -19648 11272 -18476 11288
rect -19648 11208 -18560 11272
rect -18496 11208 -18476 11272
rect -19648 11192 -18476 11208
rect -19648 11128 -18560 11192
rect -18496 11128 -18476 11192
rect -19648 11112 -18476 11128
rect -19648 11048 -18560 11112
rect -18496 11048 -18476 11112
rect -19648 11032 -18476 11048
rect -19648 10968 -18560 11032
rect -18496 10968 -18476 11032
rect -19648 10952 -18476 10968
rect -19648 10888 -18560 10952
rect -18496 10888 -18476 10952
rect -19648 10872 -18476 10888
rect -19648 10808 -18560 10872
rect -18496 10808 -18476 10872
rect -19648 10760 -18476 10808
rect -18236 11592 -17064 11640
rect -18236 11528 -17148 11592
rect -17084 11528 -17064 11592
rect -18236 11512 -17064 11528
rect -18236 11448 -17148 11512
rect -17084 11448 -17064 11512
rect -18236 11432 -17064 11448
rect -18236 11368 -17148 11432
rect -17084 11368 -17064 11432
rect -18236 11352 -17064 11368
rect -18236 11288 -17148 11352
rect -17084 11288 -17064 11352
rect -18236 11272 -17064 11288
rect -18236 11208 -17148 11272
rect -17084 11208 -17064 11272
rect -18236 11192 -17064 11208
rect -18236 11128 -17148 11192
rect -17084 11128 -17064 11192
rect -18236 11112 -17064 11128
rect -18236 11048 -17148 11112
rect -17084 11048 -17064 11112
rect -18236 11032 -17064 11048
rect -18236 10968 -17148 11032
rect -17084 10968 -17064 11032
rect -18236 10952 -17064 10968
rect -18236 10888 -17148 10952
rect -17084 10888 -17064 10952
rect -18236 10872 -17064 10888
rect -18236 10808 -17148 10872
rect -17084 10808 -17064 10872
rect -18236 10760 -17064 10808
rect -16824 11592 -15652 11640
rect -16824 11528 -15736 11592
rect -15672 11528 -15652 11592
rect -16824 11512 -15652 11528
rect -16824 11448 -15736 11512
rect -15672 11448 -15652 11512
rect -16824 11432 -15652 11448
rect -16824 11368 -15736 11432
rect -15672 11368 -15652 11432
rect -16824 11352 -15652 11368
rect -16824 11288 -15736 11352
rect -15672 11288 -15652 11352
rect -16824 11272 -15652 11288
rect -16824 11208 -15736 11272
rect -15672 11208 -15652 11272
rect -16824 11192 -15652 11208
rect -16824 11128 -15736 11192
rect -15672 11128 -15652 11192
rect -16824 11112 -15652 11128
rect -16824 11048 -15736 11112
rect -15672 11048 -15652 11112
rect -16824 11032 -15652 11048
rect -16824 10968 -15736 11032
rect -15672 10968 -15652 11032
rect -16824 10952 -15652 10968
rect -16824 10888 -15736 10952
rect -15672 10888 -15652 10952
rect -16824 10872 -15652 10888
rect -16824 10808 -15736 10872
rect -15672 10808 -15652 10872
rect -16824 10760 -15652 10808
rect -15412 11592 -14240 11640
rect -15412 11528 -14324 11592
rect -14260 11528 -14240 11592
rect -15412 11512 -14240 11528
rect -15412 11448 -14324 11512
rect -14260 11448 -14240 11512
rect -15412 11432 -14240 11448
rect -15412 11368 -14324 11432
rect -14260 11368 -14240 11432
rect -15412 11352 -14240 11368
rect -15412 11288 -14324 11352
rect -14260 11288 -14240 11352
rect -15412 11272 -14240 11288
rect -15412 11208 -14324 11272
rect -14260 11208 -14240 11272
rect -15412 11192 -14240 11208
rect -15412 11128 -14324 11192
rect -14260 11128 -14240 11192
rect -15412 11112 -14240 11128
rect -15412 11048 -14324 11112
rect -14260 11048 -14240 11112
rect -15412 11032 -14240 11048
rect -15412 10968 -14324 11032
rect -14260 10968 -14240 11032
rect -15412 10952 -14240 10968
rect -15412 10888 -14324 10952
rect -14260 10888 -14240 10952
rect -15412 10872 -14240 10888
rect -15412 10808 -14324 10872
rect -14260 10808 -14240 10872
rect -15412 10760 -14240 10808
rect -14000 11592 -12828 11640
rect -14000 11528 -12912 11592
rect -12848 11528 -12828 11592
rect -14000 11512 -12828 11528
rect -14000 11448 -12912 11512
rect -12848 11448 -12828 11512
rect -14000 11432 -12828 11448
rect -14000 11368 -12912 11432
rect -12848 11368 -12828 11432
rect -14000 11352 -12828 11368
rect -14000 11288 -12912 11352
rect -12848 11288 -12828 11352
rect -14000 11272 -12828 11288
rect -14000 11208 -12912 11272
rect -12848 11208 -12828 11272
rect -14000 11192 -12828 11208
rect -14000 11128 -12912 11192
rect -12848 11128 -12828 11192
rect -14000 11112 -12828 11128
rect -14000 11048 -12912 11112
rect -12848 11048 -12828 11112
rect -14000 11032 -12828 11048
rect -14000 10968 -12912 11032
rect -12848 10968 -12828 11032
rect -14000 10952 -12828 10968
rect -14000 10888 -12912 10952
rect -12848 10888 -12828 10952
rect -14000 10872 -12828 10888
rect -14000 10808 -12912 10872
rect -12848 10808 -12828 10872
rect -14000 10760 -12828 10808
rect -12588 11592 -11416 11640
rect -12588 11528 -11500 11592
rect -11436 11528 -11416 11592
rect -12588 11512 -11416 11528
rect -12588 11448 -11500 11512
rect -11436 11448 -11416 11512
rect -12588 11432 -11416 11448
rect -12588 11368 -11500 11432
rect -11436 11368 -11416 11432
rect -12588 11352 -11416 11368
rect -12588 11288 -11500 11352
rect -11436 11288 -11416 11352
rect -12588 11272 -11416 11288
rect -12588 11208 -11500 11272
rect -11436 11208 -11416 11272
rect -12588 11192 -11416 11208
rect -12588 11128 -11500 11192
rect -11436 11128 -11416 11192
rect -12588 11112 -11416 11128
rect -12588 11048 -11500 11112
rect -11436 11048 -11416 11112
rect -12588 11032 -11416 11048
rect -12588 10968 -11500 11032
rect -11436 10968 -11416 11032
rect -12588 10952 -11416 10968
rect -12588 10888 -11500 10952
rect -11436 10888 -11416 10952
rect -12588 10872 -11416 10888
rect -12588 10808 -11500 10872
rect -11436 10808 -11416 10872
rect -12588 10760 -11416 10808
rect -11176 11592 -10004 11640
rect -11176 11528 -10088 11592
rect -10024 11528 -10004 11592
rect -11176 11512 -10004 11528
rect -11176 11448 -10088 11512
rect -10024 11448 -10004 11512
rect -11176 11432 -10004 11448
rect -11176 11368 -10088 11432
rect -10024 11368 -10004 11432
rect -11176 11352 -10004 11368
rect -11176 11288 -10088 11352
rect -10024 11288 -10004 11352
rect -11176 11272 -10004 11288
rect -11176 11208 -10088 11272
rect -10024 11208 -10004 11272
rect -11176 11192 -10004 11208
rect -11176 11128 -10088 11192
rect -10024 11128 -10004 11192
rect -11176 11112 -10004 11128
rect -11176 11048 -10088 11112
rect -10024 11048 -10004 11112
rect -11176 11032 -10004 11048
rect -11176 10968 -10088 11032
rect -10024 10968 -10004 11032
rect -11176 10952 -10004 10968
rect -11176 10888 -10088 10952
rect -10024 10888 -10004 10952
rect -11176 10872 -10004 10888
rect -11176 10808 -10088 10872
rect -10024 10808 -10004 10872
rect -11176 10760 -10004 10808
rect -9764 11592 -8592 11640
rect -9764 11528 -8676 11592
rect -8612 11528 -8592 11592
rect -9764 11512 -8592 11528
rect -9764 11448 -8676 11512
rect -8612 11448 -8592 11512
rect -9764 11432 -8592 11448
rect -9764 11368 -8676 11432
rect -8612 11368 -8592 11432
rect -9764 11352 -8592 11368
rect -9764 11288 -8676 11352
rect -8612 11288 -8592 11352
rect -9764 11272 -8592 11288
rect -9764 11208 -8676 11272
rect -8612 11208 -8592 11272
rect -9764 11192 -8592 11208
rect -9764 11128 -8676 11192
rect -8612 11128 -8592 11192
rect -9764 11112 -8592 11128
rect -9764 11048 -8676 11112
rect -8612 11048 -8592 11112
rect -9764 11032 -8592 11048
rect -9764 10968 -8676 11032
rect -8612 10968 -8592 11032
rect -9764 10952 -8592 10968
rect -9764 10888 -8676 10952
rect -8612 10888 -8592 10952
rect -9764 10872 -8592 10888
rect -9764 10808 -8676 10872
rect -8612 10808 -8592 10872
rect -9764 10760 -8592 10808
rect -8352 11592 -7180 11640
rect -8352 11528 -7264 11592
rect -7200 11528 -7180 11592
rect -8352 11512 -7180 11528
rect -8352 11448 -7264 11512
rect -7200 11448 -7180 11512
rect -8352 11432 -7180 11448
rect -8352 11368 -7264 11432
rect -7200 11368 -7180 11432
rect -8352 11352 -7180 11368
rect -8352 11288 -7264 11352
rect -7200 11288 -7180 11352
rect -8352 11272 -7180 11288
rect -8352 11208 -7264 11272
rect -7200 11208 -7180 11272
rect -8352 11192 -7180 11208
rect -8352 11128 -7264 11192
rect -7200 11128 -7180 11192
rect -8352 11112 -7180 11128
rect -8352 11048 -7264 11112
rect -7200 11048 -7180 11112
rect -8352 11032 -7180 11048
rect -8352 10968 -7264 11032
rect -7200 10968 -7180 11032
rect -8352 10952 -7180 10968
rect -8352 10888 -7264 10952
rect -7200 10888 -7180 10952
rect -8352 10872 -7180 10888
rect -8352 10808 -7264 10872
rect -7200 10808 -7180 10872
rect -8352 10760 -7180 10808
rect -6940 11592 -5768 11640
rect -6940 11528 -5852 11592
rect -5788 11528 -5768 11592
rect -6940 11512 -5768 11528
rect -6940 11448 -5852 11512
rect -5788 11448 -5768 11512
rect -6940 11432 -5768 11448
rect -6940 11368 -5852 11432
rect -5788 11368 -5768 11432
rect -6940 11352 -5768 11368
rect -6940 11288 -5852 11352
rect -5788 11288 -5768 11352
rect -6940 11272 -5768 11288
rect -6940 11208 -5852 11272
rect -5788 11208 -5768 11272
rect -6940 11192 -5768 11208
rect -6940 11128 -5852 11192
rect -5788 11128 -5768 11192
rect -6940 11112 -5768 11128
rect -6940 11048 -5852 11112
rect -5788 11048 -5768 11112
rect -6940 11032 -5768 11048
rect -6940 10968 -5852 11032
rect -5788 10968 -5768 11032
rect -6940 10952 -5768 10968
rect -6940 10888 -5852 10952
rect -5788 10888 -5768 10952
rect -6940 10872 -5768 10888
rect -6940 10808 -5852 10872
rect -5788 10808 -5768 10872
rect -6940 10760 -5768 10808
rect -5528 11592 -4356 11640
rect -5528 11528 -4440 11592
rect -4376 11528 -4356 11592
rect -5528 11512 -4356 11528
rect -5528 11448 -4440 11512
rect -4376 11448 -4356 11512
rect -5528 11432 -4356 11448
rect -5528 11368 -4440 11432
rect -4376 11368 -4356 11432
rect -5528 11352 -4356 11368
rect -5528 11288 -4440 11352
rect -4376 11288 -4356 11352
rect -5528 11272 -4356 11288
rect -5528 11208 -4440 11272
rect -4376 11208 -4356 11272
rect -5528 11192 -4356 11208
rect -5528 11128 -4440 11192
rect -4376 11128 -4356 11192
rect -5528 11112 -4356 11128
rect -5528 11048 -4440 11112
rect -4376 11048 -4356 11112
rect -5528 11032 -4356 11048
rect -5528 10968 -4440 11032
rect -4376 10968 -4356 11032
rect -5528 10952 -4356 10968
rect -5528 10888 -4440 10952
rect -4376 10888 -4356 10952
rect -5528 10872 -4356 10888
rect -5528 10808 -4440 10872
rect -4376 10808 -4356 10872
rect -5528 10760 -4356 10808
rect -4116 11592 -2944 11640
rect -4116 11528 -3028 11592
rect -2964 11528 -2944 11592
rect -4116 11512 -2944 11528
rect -4116 11448 -3028 11512
rect -2964 11448 -2944 11512
rect -4116 11432 -2944 11448
rect -4116 11368 -3028 11432
rect -2964 11368 -2944 11432
rect -4116 11352 -2944 11368
rect -4116 11288 -3028 11352
rect -2964 11288 -2944 11352
rect -4116 11272 -2944 11288
rect -4116 11208 -3028 11272
rect -2964 11208 -2944 11272
rect -4116 11192 -2944 11208
rect -4116 11128 -3028 11192
rect -2964 11128 -2944 11192
rect -4116 11112 -2944 11128
rect -4116 11048 -3028 11112
rect -2964 11048 -2944 11112
rect -4116 11032 -2944 11048
rect -4116 10968 -3028 11032
rect -2964 10968 -2944 11032
rect -4116 10952 -2944 10968
rect -4116 10888 -3028 10952
rect -2964 10888 -2944 10952
rect -4116 10872 -2944 10888
rect -4116 10808 -3028 10872
rect -2964 10808 -2944 10872
rect -4116 10760 -2944 10808
rect -2704 11592 -1532 11640
rect -2704 11528 -1616 11592
rect -1552 11528 -1532 11592
rect -2704 11512 -1532 11528
rect -2704 11448 -1616 11512
rect -1552 11448 -1532 11512
rect -2704 11432 -1532 11448
rect -2704 11368 -1616 11432
rect -1552 11368 -1532 11432
rect -2704 11352 -1532 11368
rect -2704 11288 -1616 11352
rect -1552 11288 -1532 11352
rect -2704 11272 -1532 11288
rect -2704 11208 -1616 11272
rect -1552 11208 -1532 11272
rect -2704 11192 -1532 11208
rect -2704 11128 -1616 11192
rect -1552 11128 -1532 11192
rect -2704 11112 -1532 11128
rect -2704 11048 -1616 11112
rect -1552 11048 -1532 11112
rect -2704 11032 -1532 11048
rect -2704 10968 -1616 11032
rect -1552 10968 -1532 11032
rect -2704 10952 -1532 10968
rect -2704 10888 -1616 10952
rect -1552 10888 -1532 10952
rect -2704 10872 -1532 10888
rect -2704 10808 -1616 10872
rect -1552 10808 -1532 10872
rect -2704 10760 -1532 10808
rect -1292 11592 -120 11640
rect -1292 11528 -204 11592
rect -140 11528 -120 11592
rect -1292 11512 -120 11528
rect -1292 11448 -204 11512
rect -140 11448 -120 11512
rect -1292 11432 -120 11448
rect -1292 11368 -204 11432
rect -140 11368 -120 11432
rect -1292 11352 -120 11368
rect -1292 11288 -204 11352
rect -140 11288 -120 11352
rect -1292 11272 -120 11288
rect -1292 11208 -204 11272
rect -140 11208 -120 11272
rect -1292 11192 -120 11208
rect -1292 11128 -204 11192
rect -140 11128 -120 11192
rect -1292 11112 -120 11128
rect -1292 11048 -204 11112
rect -140 11048 -120 11112
rect -1292 11032 -120 11048
rect -1292 10968 -204 11032
rect -140 10968 -120 11032
rect -1292 10952 -120 10968
rect -1292 10888 -204 10952
rect -140 10888 -120 10952
rect -1292 10872 -120 10888
rect -1292 10808 -204 10872
rect -140 10808 -120 10872
rect -1292 10760 -120 10808
rect 120 11592 1292 11640
rect 120 11528 1208 11592
rect 1272 11528 1292 11592
rect 120 11512 1292 11528
rect 120 11448 1208 11512
rect 1272 11448 1292 11512
rect 120 11432 1292 11448
rect 120 11368 1208 11432
rect 1272 11368 1292 11432
rect 120 11352 1292 11368
rect 120 11288 1208 11352
rect 1272 11288 1292 11352
rect 120 11272 1292 11288
rect 120 11208 1208 11272
rect 1272 11208 1292 11272
rect 120 11192 1292 11208
rect 120 11128 1208 11192
rect 1272 11128 1292 11192
rect 120 11112 1292 11128
rect 120 11048 1208 11112
rect 1272 11048 1292 11112
rect 120 11032 1292 11048
rect 120 10968 1208 11032
rect 1272 10968 1292 11032
rect 120 10952 1292 10968
rect 120 10888 1208 10952
rect 1272 10888 1292 10952
rect 120 10872 1292 10888
rect 120 10808 1208 10872
rect 1272 10808 1292 10872
rect 120 10760 1292 10808
rect 1532 11592 2704 11640
rect 1532 11528 2620 11592
rect 2684 11528 2704 11592
rect 1532 11512 2704 11528
rect 1532 11448 2620 11512
rect 2684 11448 2704 11512
rect 1532 11432 2704 11448
rect 1532 11368 2620 11432
rect 2684 11368 2704 11432
rect 1532 11352 2704 11368
rect 1532 11288 2620 11352
rect 2684 11288 2704 11352
rect 1532 11272 2704 11288
rect 1532 11208 2620 11272
rect 2684 11208 2704 11272
rect 1532 11192 2704 11208
rect 1532 11128 2620 11192
rect 2684 11128 2704 11192
rect 1532 11112 2704 11128
rect 1532 11048 2620 11112
rect 2684 11048 2704 11112
rect 1532 11032 2704 11048
rect 1532 10968 2620 11032
rect 2684 10968 2704 11032
rect 1532 10952 2704 10968
rect 1532 10888 2620 10952
rect 2684 10888 2704 10952
rect 1532 10872 2704 10888
rect 1532 10808 2620 10872
rect 2684 10808 2704 10872
rect 1532 10760 2704 10808
rect 2944 11592 4116 11640
rect 2944 11528 4032 11592
rect 4096 11528 4116 11592
rect 2944 11512 4116 11528
rect 2944 11448 4032 11512
rect 4096 11448 4116 11512
rect 2944 11432 4116 11448
rect 2944 11368 4032 11432
rect 4096 11368 4116 11432
rect 2944 11352 4116 11368
rect 2944 11288 4032 11352
rect 4096 11288 4116 11352
rect 2944 11272 4116 11288
rect 2944 11208 4032 11272
rect 4096 11208 4116 11272
rect 2944 11192 4116 11208
rect 2944 11128 4032 11192
rect 4096 11128 4116 11192
rect 2944 11112 4116 11128
rect 2944 11048 4032 11112
rect 4096 11048 4116 11112
rect 2944 11032 4116 11048
rect 2944 10968 4032 11032
rect 4096 10968 4116 11032
rect 2944 10952 4116 10968
rect 2944 10888 4032 10952
rect 4096 10888 4116 10952
rect 2944 10872 4116 10888
rect 2944 10808 4032 10872
rect 4096 10808 4116 10872
rect 2944 10760 4116 10808
rect 4356 11592 5528 11640
rect 4356 11528 5444 11592
rect 5508 11528 5528 11592
rect 4356 11512 5528 11528
rect 4356 11448 5444 11512
rect 5508 11448 5528 11512
rect 4356 11432 5528 11448
rect 4356 11368 5444 11432
rect 5508 11368 5528 11432
rect 4356 11352 5528 11368
rect 4356 11288 5444 11352
rect 5508 11288 5528 11352
rect 4356 11272 5528 11288
rect 4356 11208 5444 11272
rect 5508 11208 5528 11272
rect 4356 11192 5528 11208
rect 4356 11128 5444 11192
rect 5508 11128 5528 11192
rect 4356 11112 5528 11128
rect 4356 11048 5444 11112
rect 5508 11048 5528 11112
rect 4356 11032 5528 11048
rect 4356 10968 5444 11032
rect 5508 10968 5528 11032
rect 4356 10952 5528 10968
rect 4356 10888 5444 10952
rect 5508 10888 5528 10952
rect 4356 10872 5528 10888
rect 4356 10808 5444 10872
rect 5508 10808 5528 10872
rect 4356 10760 5528 10808
rect 5768 11592 6940 11640
rect 5768 11528 6856 11592
rect 6920 11528 6940 11592
rect 5768 11512 6940 11528
rect 5768 11448 6856 11512
rect 6920 11448 6940 11512
rect 5768 11432 6940 11448
rect 5768 11368 6856 11432
rect 6920 11368 6940 11432
rect 5768 11352 6940 11368
rect 5768 11288 6856 11352
rect 6920 11288 6940 11352
rect 5768 11272 6940 11288
rect 5768 11208 6856 11272
rect 6920 11208 6940 11272
rect 5768 11192 6940 11208
rect 5768 11128 6856 11192
rect 6920 11128 6940 11192
rect 5768 11112 6940 11128
rect 5768 11048 6856 11112
rect 6920 11048 6940 11112
rect 5768 11032 6940 11048
rect 5768 10968 6856 11032
rect 6920 10968 6940 11032
rect 5768 10952 6940 10968
rect 5768 10888 6856 10952
rect 6920 10888 6940 10952
rect 5768 10872 6940 10888
rect 5768 10808 6856 10872
rect 6920 10808 6940 10872
rect 5768 10760 6940 10808
rect 7180 11592 8352 11640
rect 7180 11528 8268 11592
rect 8332 11528 8352 11592
rect 7180 11512 8352 11528
rect 7180 11448 8268 11512
rect 8332 11448 8352 11512
rect 7180 11432 8352 11448
rect 7180 11368 8268 11432
rect 8332 11368 8352 11432
rect 7180 11352 8352 11368
rect 7180 11288 8268 11352
rect 8332 11288 8352 11352
rect 7180 11272 8352 11288
rect 7180 11208 8268 11272
rect 8332 11208 8352 11272
rect 7180 11192 8352 11208
rect 7180 11128 8268 11192
rect 8332 11128 8352 11192
rect 7180 11112 8352 11128
rect 7180 11048 8268 11112
rect 8332 11048 8352 11112
rect 7180 11032 8352 11048
rect 7180 10968 8268 11032
rect 8332 10968 8352 11032
rect 7180 10952 8352 10968
rect 7180 10888 8268 10952
rect 8332 10888 8352 10952
rect 7180 10872 8352 10888
rect 7180 10808 8268 10872
rect 8332 10808 8352 10872
rect 7180 10760 8352 10808
rect 8592 11592 9764 11640
rect 8592 11528 9680 11592
rect 9744 11528 9764 11592
rect 8592 11512 9764 11528
rect 8592 11448 9680 11512
rect 9744 11448 9764 11512
rect 8592 11432 9764 11448
rect 8592 11368 9680 11432
rect 9744 11368 9764 11432
rect 8592 11352 9764 11368
rect 8592 11288 9680 11352
rect 9744 11288 9764 11352
rect 8592 11272 9764 11288
rect 8592 11208 9680 11272
rect 9744 11208 9764 11272
rect 8592 11192 9764 11208
rect 8592 11128 9680 11192
rect 9744 11128 9764 11192
rect 8592 11112 9764 11128
rect 8592 11048 9680 11112
rect 9744 11048 9764 11112
rect 8592 11032 9764 11048
rect 8592 10968 9680 11032
rect 9744 10968 9764 11032
rect 8592 10952 9764 10968
rect 8592 10888 9680 10952
rect 9744 10888 9764 10952
rect 8592 10872 9764 10888
rect 8592 10808 9680 10872
rect 9744 10808 9764 10872
rect 8592 10760 9764 10808
rect 10004 11592 11176 11640
rect 10004 11528 11092 11592
rect 11156 11528 11176 11592
rect 10004 11512 11176 11528
rect 10004 11448 11092 11512
rect 11156 11448 11176 11512
rect 10004 11432 11176 11448
rect 10004 11368 11092 11432
rect 11156 11368 11176 11432
rect 10004 11352 11176 11368
rect 10004 11288 11092 11352
rect 11156 11288 11176 11352
rect 10004 11272 11176 11288
rect 10004 11208 11092 11272
rect 11156 11208 11176 11272
rect 10004 11192 11176 11208
rect 10004 11128 11092 11192
rect 11156 11128 11176 11192
rect 10004 11112 11176 11128
rect 10004 11048 11092 11112
rect 11156 11048 11176 11112
rect 10004 11032 11176 11048
rect 10004 10968 11092 11032
rect 11156 10968 11176 11032
rect 10004 10952 11176 10968
rect 10004 10888 11092 10952
rect 11156 10888 11176 10952
rect 10004 10872 11176 10888
rect 10004 10808 11092 10872
rect 11156 10808 11176 10872
rect 10004 10760 11176 10808
rect 11416 11592 12588 11640
rect 11416 11528 12504 11592
rect 12568 11528 12588 11592
rect 11416 11512 12588 11528
rect 11416 11448 12504 11512
rect 12568 11448 12588 11512
rect 11416 11432 12588 11448
rect 11416 11368 12504 11432
rect 12568 11368 12588 11432
rect 11416 11352 12588 11368
rect 11416 11288 12504 11352
rect 12568 11288 12588 11352
rect 11416 11272 12588 11288
rect 11416 11208 12504 11272
rect 12568 11208 12588 11272
rect 11416 11192 12588 11208
rect 11416 11128 12504 11192
rect 12568 11128 12588 11192
rect 11416 11112 12588 11128
rect 11416 11048 12504 11112
rect 12568 11048 12588 11112
rect 11416 11032 12588 11048
rect 11416 10968 12504 11032
rect 12568 10968 12588 11032
rect 11416 10952 12588 10968
rect 11416 10888 12504 10952
rect 12568 10888 12588 10952
rect 11416 10872 12588 10888
rect 11416 10808 12504 10872
rect 12568 10808 12588 10872
rect 11416 10760 12588 10808
rect 12828 11592 14000 11640
rect 12828 11528 13916 11592
rect 13980 11528 14000 11592
rect 12828 11512 14000 11528
rect 12828 11448 13916 11512
rect 13980 11448 14000 11512
rect 12828 11432 14000 11448
rect 12828 11368 13916 11432
rect 13980 11368 14000 11432
rect 12828 11352 14000 11368
rect 12828 11288 13916 11352
rect 13980 11288 14000 11352
rect 12828 11272 14000 11288
rect 12828 11208 13916 11272
rect 13980 11208 14000 11272
rect 12828 11192 14000 11208
rect 12828 11128 13916 11192
rect 13980 11128 14000 11192
rect 12828 11112 14000 11128
rect 12828 11048 13916 11112
rect 13980 11048 14000 11112
rect 12828 11032 14000 11048
rect 12828 10968 13916 11032
rect 13980 10968 14000 11032
rect 12828 10952 14000 10968
rect 12828 10888 13916 10952
rect 13980 10888 14000 10952
rect 12828 10872 14000 10888
rect 12828 10808 13916 10872
rect 13980 10808 14000 10872
rect 12828 10760 14000 10808
rect 14240 11592 15412 11640
rect 14240 11528 15328 11592
rect 15392 11528 15412 11592
rect 14240 11512 15412 11528
rect 14240 11448 15328 11512
rect 15392 11448 15412 11512
rect 14240 11432 15412 11448
rect 14240 11368 15328 11432
rect 15392 11368 15412 11432
rect 14240 11352 15412 11368
rect 14240 11288 15328 11352
rect 15392 11288 15412 11352
rect 14240 11272 15412 11288
rect 14240 11208 15328 11272
rect 15392 11208 15412 11272
rect 14240 11192 15412 11208
rect 14240 11128 15328 11192
rect 15392 11128 15412 11192
rect 14240 11112 15412 11128
rect 14240 11048 15328 11112
rect 15392 11048 15412 11112
rect 14240 11032 15412 11048
rect 14240 10968 15328 11032
rect 15392 10968 15412 11032
rect 14240 10952 15412 10968
rect 14240 10888 15328 10952
rect 15392 10888 15412 10952
rect 14240 10872 15412 10888
rect 14240 10808 15328 10872
rect 15392 10808 15412 10872
rect 14240 10760 15412 10808
rect 15652 11592 16824 11640
rect 15652 11528 16740 11592
rect 16804 11528 16824 11592
rect 15652 11512 16824 11528
rect 15652 11448 16740 11512
rect 16804 11448 16824 11512
rect 15652 11432 16824 11448
rect 15652 11368 16740 11432
rect 16804 11368 16824 11432
rect 15652 11352 16824 11368
rect 15652 11288 16740 11352
rect 16804 11288 16824 11352
rect 15652 11272 16824 11288
rect 15652 11208 16740 11272
rect 16804 11208 16824 11272
rect 15652 11192 16824 11208
rect 15652 11128 16740 11192
rect 16804 11128 16824 11192
rect 15652 11112 16824 11128
rect 15652 11048 16740 11112
rect 16804 11048 16824 11112
rect 15652 11032 16824 11048
rect 15652 10968 16740 11032
rect 16804 10968 16824 11032
rect 15652 10952 16824 10968
rect 15652 10888 16740 10952
rect 16804 10888 16824 10952
rect 15652 10872 16824 10888
rect 15652 10808 16740 10872
rect 16804 10808 16824 10872
rect 15652 10760 16824 10808
rect 17064 11592 18236 11640
rect 17064 11528 18152 11592
rect 18216 11528 18236 11592
rect 17064 11512 18236 11528
rect 17064 11448 18152 11512
rect 18216 11448 18236 11512
rect 17064 11432 18236 11448
rect 17064 11368 18152 11432
rect 18216 11368 18236 11432
rect 17064 11352 18236 11368
rect 17064 11288 18152 11352
rect 18216 11288 18236 11352
rect 17064 11272 18236 11288
rect 17064 11208 18152 11272
rect 18216 11208 18236 11272
rect 17064 11192 18236 11208
rect 17064 11128 18152 11192
rect 18216 11128 18236 11192
rect 17064 11112 18236 11128
rect 17064 11048 18152 11112
rect 18216 11048 18236 11112
rect 17064 11032 18236 11048
rect 17064 10968 18152 11032
rect 18216 10968 18236 11032
rect 17064 10952 18236 10968
rect 17064 10888 18152 10952
rect 18216 10888 18236 10952
rect 17064 10872 18236 10888
rect 17064 10808 18152 10872
rect 18216 10808 18236 10872
rect 17064 10760 18236 10808
rect 18476 11592 19648 11640
rect 18476 11528 19564 11592
rect 19628 11528 19648 11592
rect 18476 11512 19648 11528
rect 18476 11448 19564 11512
rect 19628 11448 19648 11512
rect 18476 11432 19648 11448
rect 18476 11368 19564 11432
rect 19628 11368 19648 11432
rect 18476 11352 19648 11368
rect 18476 11288 19564 11352
rect 19628 11288 19648 11352
rect 18476 11272 19648 11288
rect 18476 11208 19564 11272
rect 19628 11208 19648 11272
rect 18476 11192 19648 11208
rect 18476 11128 19564 11192
rect 19628 11128 19648 11192
rect 18476 11112 19648 11128
rect 18476 11048 19564 11112
rect 19628 11048 19648 11112
rect 18476 11032 19648 11048
rect 18476 10968 19564 11032
rect 19628 10968 19648 11032
rect 18476 10952 19648 10968
rect 18476 10888 19564 10952
rect 19628 10888 19648 10952
rect 18476 10872 19648 10888
rect 18476 10808 19564 10872
rect 19628 10808 19648 10872
rect 18476 10760 19648 10808
rect 19888 11592 21060 11640
rect 19888 11528 20976 11592
rect 21040 11528 21060 11592
rect 19888 11512 21060 11528
rect 19888 11448 20976 11512
rect 21040 11448 21060 11512
rect 19888 11432 21060 11448
rect 19888 11368 20976 11432
rect 21040 11368 21060 11432
rect 19888 11352 21060 11368
rect 19888 11288 20976 11352
rect 21040 11288 21060 11352
rect 19888 11272 21060 11288
rect 19888 11208 20976 11272
rect 21040 11208 21060 11272
rect 19888 11192 21060 11208
rect 19888 11128 20976 11192
rect 21040 11128 21060 11192
rect 19888 11112 21060 11128
rect 19888 11048 20976 11112
rect 21040 11048 21060 11112
rect 19888 11032 21060 11048
rect 19888 10968 20976 11032
rect 21040 10968 21060 11032
rect 19888 10952 21060 10968
rect 19888 10888 20976 10952
rect 21040 10888 21060 10952
rect 19888 10872 21060 10888
rect 19888 10808 20976 10872
rect 21040 10808 21060 10872
rect 19888 10760 21060 10808
rect 21300 11592 22472 11640
rect 21300 11528 22388 11592
rect 22452 11528 22472 11592
rect 21300 11512 22472 11528
rect 21300 11448 22388 11512
rect 22452 11448 22472 11512
rect 21300 11432 22472 11448
rect 21300 11368 22388 11432
rect 22452 11368 22472 11432
rect 21300 11352 22472 11368
rect 21300 11288 22388 11352
rect 22452 11288 22472 11352
rect 21300 11272 22472 11288
rect 21300 11208 22388 11272
rect 22452 11208 22472 11272
rect 21300 11192 22472 11208
rect 21300 11128 22388 11192
rect 22452 11128 22472 11192
rect 21300 11112 22472 11128
rect 21300 11048 22388 11112
rect 22452 11048 22472 11112
rect 21300 11032 22472 11048
rect 21300 10968 22388 11032
rect 22452 10968 22472 11032
rect 21300 10952 22472 10968
rect 21300 10888 22388 10952
rect 22452 10888 22472 10952
rect 21300 10872 22472 10888
rect 21300 10808 22388 10872
rect 22452 10808 22472 10872
rect 21300 10760 22472 10808
rect 22712 11592 23884 11640
rect 22712 11528 23800 11592
rect 23864 11528 23884 11592
rect 22712 11512 23884 11528
rect 22712 11448 23800 11512
rect 23864 11448 23884 11512
rect 22712 11432 23884 11448
rect 22712 11368 23800 11432
rect 23864 11368 23884 11432
rect 22712 11352 23884 11368
rect 22712 11288 23800 11352
rect 23864 11288 23884 11352
rect 22712 11272 23884 11288
rect 22712 11208 23800 11272
rect 23864 11208 23884 11272
rect 22712 11192 23884 11208
rect 22712 11128 23800 11192
rect 23864 11128 23884 11192
rect 22712 11112 23884 11128
rect 22712 11048 23800 11112
rect 23864 11048 23884 11112
rect 22712 11032 23884 11048
rect 22712 10968 23800 11032
rect 23864 10968 23884 11032
rect 22712 10952 23884 10968
rect 22712 10888 23800 10952
rect 23864 10888 23884 10952
rect 22712 10872 23884 10888
rect 22712 10808 23800 10872
rect 23864 10808 23884 10872
rect 22712 10760 23884 10808
rect -23884 10472 -22712 10520
rect -23884 10408 -22796 10472
rect -22732 10408 -22712 10472
rect -23884 10392 -22712 10408
rect -23884 10328 -22796 10392
rect -22732 10328 -22712 10392
rect -23884 10312 -22712 10328
rect -23884 10248 -22796 10312
rect -22732 10248 -22712 10312
rect -23884 10232 -22712 10248
rect -23884 10168 -22796 10232
rect -22732 10168 -22712 10232
rect -23884 10152 -22712 10168
rect -23884 10088 -22796 10152
rect -22732 10088 -22712 10152
rect -23884 10072 -22712 10088
rect -23884 10008 -22796 10072
rect -22732 10008 -22712 10072
rect -23884 9992 -22712 10008
rect -23884 9928 -22796 9992
rect -22732 9928 -22712 9992
rect -23884 9912 -22712 9928
rect -23884 9848 -22796 9912
rect -22732 9848 -22712 9912
rect -23884 9832 -22712 9848
rect -23884 9768 -22796 9832
rect -22732 9768 -22712 9832
rect -23884 9752 -22712 9768
rect -23884 9688 -22796 9752
rect -22732 9688 -22712 9752
rect -23884 9640 -22712 9688
rect -22472 10472 -21300 10520
rect -22472 10408 -21384 10472
rect -21320 10408 -21300 10472
rect -22472 10392 -21300 10408
rect -22472 10328 -21384 10392
rect -21320 10328 -21300 10392
rect -22472 10312 -21300 10328
rect -22472 10248 -21384 10312
rect -21320 10248 -21300 10312
rect -22472 10232 -21300 10248
rect -22472 10168 -21384 10232
rect -21320 10168 -21300 10232
rect -22472 10152 -21300 10168
rect -22472 10088 -21384 10152
rect -21320 10088 -21300 10152
rect -22472 10072 -21300 10088
rect -22472 10008 -21384 10072
rect -21320 10008 -21300 10072
rect -22472 9992 -21300 10008
rect -22472 9928 -21384 9992
rect -21320 9928 -21300 9992
rect -22472 9912 -21300 9928
rect -22472 9848 -21384 9912
rect -21320 9848 -21300 9912
rect -22472 9832 -21300 9848
rect -22472 9768 -21384 9832
rect -21320 9768 -21300 9832
rect -22472 9752 -21300 9768
rect -22472 9688 -21384 9752
rect -21320 9688 -21300 9752
rect -22472 9640 -21300 9688
rect -21060 10472 -19888 10520
rect -21060 10408 -19972 10472
rect -19908 10408 -19888 10472
rect -21060 10392 -19888 10408
rect -21060 10328 -19972 10392
rect -19908 10328 -19888 10392
rect -21060 10312 -19888 10328
rect -21060 10248 -19972 10312
rect -19908 10248 -19888 10312
rect -21060 10232 -19888 10248
rect -21060 10168 -19972 10232
rect -19908 10168 -19888 10232
rect -21060 10152 -19888 10168
rect -21060 10088 -19972 10152
rect -19908 10088 -19888 10152
rect -21060 10072 -19888 10088
rect -21060 10008 -19972 10072
rect -19908 10008 -19888 10072
rect -21060 9992 -19888 10008
rect -21060 9928 -19972 9992
rect -19908 9928 -19888 9992
rect -21060 9912 -19888 9928
rect -21060 9848 -19972 9912
rect -19908 9848 -19888 9912
rect -21060 9832 -19888 9848
rect -21060 9768 -19972 9832
rect -19908 9768 -19888 9832
rect -21060 9752 -19888 9768
rect -21060 9688 -19972 9752
rect -19908 9688 -19888 9752
rect -21060 9640 -19888 9688
rect -19648 10472 -18476 10520
rect -19648 10408 -18560 10472
rect -18496 10408 -18476 10472
rect -19648 10392 -18476 10408
rect -19648 10328 -18560 10392
rect -18496 10328 -18476 10392
rect -19648 10312 -18476 10328
rect -19648 10248 -18560 10312
rect -18496 10248 -18476 10312
rect -19648 10232 -18476 10248
rect -19648 10168 -18560 10232
rect -18496 10168 -18476 10232
rect -19648 10152 -18476 10168
rect -19648 10088 -18560 10152
rect -18496 10088 -18476 10152
rect -19648 10072 -18476 10088
rect -19648 10008 -18560 10072
rect -18496 10008 -18476 10072
rect -19648 9992 -18476 10008
rect -19648 9928 -18560 9992
rect -18496 9928 -18476 9992
rect -19648 9912 -18476 9928
rect -19648 9848 -18560 9912
rect -18496 9848 -18476 9912
rect -19648 9832 -18476 9848
rect -19648 9768 -18560 9832
rect -18496 9768 -18476 9832
rect -19648 9752 -18476 9768
rect -19648 9688 -18560 9752
rect -18496 9688 -18476 9752
rect -19648 9640 -18476 9688
rect -18236 10472 -17064 10520
rect -18236 10408 -17148 10472
rect -17084 10408 -17064 10472
rect -18236 10392 -17064 10408
rect -18236 10328 -17148 10392
rect -17084 10328 -17064 10392
rect -18236 10312 -17064 10328
rect -18236 10248 -17148 10312
rect -17084 10248 -17064 10312
rect -18236 10232 -17064 10248
rect -18236 10168 -17148 10232
rect -17084 10168 -17064 10232
rect -18236 10152 -17064 10168
rect -18236 10088 -17148 10152
rect -17084 10088 -17064 10152
rect -18236 10072 -17064 10088
rect -18236 10008 -17148 10072
rect -17084 10008 -17064 10072
rect -18236 9992 -17064 10008
rect -18236 9928 -17148 9992
rect -17084 9928 -17064 9992
rect -18236 9912 -17064 9928
rect -18236 9848 -17148 9912
rect -17084 9848 -17064 9912
rect -18236 9832 -17064 9848
rect -18236 9768 -17148 9832
rect -17084 9768 -17064 9832
rect -18236 9752 -17064 9768
rect -18236 9688 -17148 9752
rect -17084 9688 -17064 9752
rect -18236 9640 -17064 9688
rect -16824 10472 -15652 10520
rect -16824 10408 -15736 10472
rect -15672 10408 -15652 10472
rect -16824 10392 -15652 10408
rect -16824 10328 -15736 10392
rect -15672 10328 -15652 10392
rect -16824 10312 -15652 10328
rect -16824 10248 -15736 10312
rect -15672 10248 -15652 10312
rect -16824 10232 -15652 10248
rect -16824 10168 -15736 10232
rect -15672 10168 -15652 10232
rect -16824 10152 -15652 10168
rect -16824 10088 -15736 10152
rect -15672 10088 -15652 10152
rect -16824 10072 -15652 10088
rect -16824 10008 -15736 10072
rect -15672 10008 -15652 10072
rect -16824 9992 -15652 10008
rect -16824 9928 -15736 9992
rect -15672 9928 -15652 9992
rect -16824 9912 -15652 9928
rect -16824 9848 -15736 9912
rect -15672 9848 -15652 9912
rect -16824 9832 -15652 9848
rect -16824 9768 -15736 9832
rect -15672 9768 -15652 9832
rect -16824 9752 -15652 9768
rect -16824 9688 -15736 9752
rect -15672 9688 -15652 9752
rect -16824 9640 -15652 9688
rect -15412 10472 -14240 10520
rect -15412 10408 -14324 10472
rect -14260 10408 -14240 10472
rect -15412 10392 -14240 10408
rect -15412 10328 -14324 10392
rect -14260 10328 -14240 10392
rect -15412 10312 -14240 10328
rect -15412 10248 -14324 10312
rect -14260 10248 -14240 10312
rect -15412 10232 -14240 10248
rect -15412 10168 -14324 10232
rect -14260 10168 -14240 10232
rect -15412 10152 -14240 10168
rect -15412 10088 -14324 10152
rect -14260 10088 -14240 10152
rect -15412 10072 -14240 10088
rect -15412 10008 -14324 10072
rect -14260 10008 -14240 10072
rect -15412 9992 -14240 10008
rect -15412 9928 -14324 9992
rect -14260 9928 -14240 9992
rect -15412 9912 -14240 9928
rect -15412 9848 -14324 9912
rect -14260 9848 -14240 9912
rect -15412 9832 -14240 9848
rect -15412 9768 -14324 9832
rect -14260 9768 -14240 9832
rect -15412 9752 -14240 9768
rect -15412 9688 -14324 9752
rect -14260 9688 -14240 9752
rect -15412 9640 -14240 9688
rect -14000 10472 -12828 10520
rect -14000 10408 -12912 10472
rect -12848 10408 -12828 10472
rect -14000 10392 -12828 10408
rect -14000 10328 -12912 10392
rect -12848 10328 -12828 10392
rect -14000 10312 -12828 10328
rect -14000 10248 -12912 10312
rect -12848 10248 -12828 10312
rect -14000 10232 -12828 10248
rect -14000 10168 -12912 10232
rect -12848 10168 -12828 10232
rect -14000 10152 -12828 10168
rect -14000 10088 -12912 10152
rect -12848 10088 -12828 10152
rect -14000 10072 -12828 10088
rect -14000 10008 -12912 10072
rect -12848 10008 -12828 10072
rect -14000 9992 -12828 10008
rect -14000 9928 -12912 9992
rect -12848 9928 -12828 9992
rect -14000 9912 -12828 9928
rect -14000 9848 -12912 9912
rect -12848 9848 -12828 9912
rect -14000 9832 -12828 9848
rect -14000 9768 -12912 9832
rect -12848 9768 -12828 9832
rect -14000 9752 -12828 9768
rect -14000 9688 -12912 9752
rect -12848 9688 -12828 9752
rect -14000 9640 -12828 9688
rect -12588 10472 -11416 10520
rect -12588 10408 -11500 10472
rect -11436 10408 -11416 10472
rect -12588 10392 -11416 10408
rect -12588 10328 -11500 10392
rect -11436 10328 -11416 10392
rect -12588 10312 -11416 10328
rect -12588 10248 -11500 10312
rect -11436 10248 -11416 10312
rect -12588 10232 -11416 10248
rect -12588 10168 -11500 10232
rect -11436 10168 -11416 10232
rect -12588 10152 -11416 10168
rect -12588 10088 -11500 10152
rect -11436 10088 -11416 10152
rect -12588 10072 -11416 10088
rect -12588 10008 -11500 10072
rect -11436 10008 -11416 10072
rect -12588 9992 -11416 10008
rect -12588 9928 -11500 9992
rect -11436 9928 -11416 9992
rect -12588 9912 -11416 9928
rect -12588 9848 -11500 9912
rect -11436 9848 -11416 9912
rect -12588 9832 -11416 9848
rect -12588 9768 -11500 9832
rect -11436 9768 -11416 9832
rect -12588 9752 -11416 9768
rect -12588 9688 -11500 9752
rect -11436 9688 -11416 9752
rect -12588 9640 -11416 9688
rect -11176 10472 -10004 10520
rect -11176 10408 -10088 10472
rect -10024 10408 -10004 10472
rect -11176 10392 -10004 10408
rect -11176 10328 -10088 10392
rect -10024 10328 -10004 10392
rect -11176 10312 -10004 10328
rect -11176 10248 -10088 10312
rect -10024 10248 -10004 10312
rect -11176 10232 -10004 10248
rect -11176 10168 -10088 10232
rect -10024 10168 -10004 10232
rect -11176 10152 -10004 10168
rect -11176 10088 -10088 10152
rect -10024 10088 -10004 10152
rect -11176 10072 -10004 10088
rect -11176 10008 -10088 10072
rect -10024 10008 -10004 10072
rect -11176 9992 -10004 10008
rect -11176 9928 -10088 9992
rect -10024 9928 -10004 9992
rect -11176 9912 -10004 9928
rect -11176 9848 -10088 9912
rect -10024 9848 -10004 9912
rect -11176 9832 -10004 9848
rect -11176 9768 -10088 9832
rect -10024 9768 -10004 9832
rect -11176 9752 -10004 9768
rect -11176 9688 -10088 9752
rect -10024 9688 -10004 9752
rect -11176 9640 -10004 9688
rect -9764 10472 -8592 10520
rect -9764 10408 -8676 10472
rect -8612 10408 -8592 10472
rect -9764 10392 -8592 10408
rect -9764 10328 -8676 10392
rect -8612 10328 -8592 10392
rect -9764 10312 -8592 10328
rect -9764 10248 -8676 10312
rect -8612 10248 -8592 10312
rect -9764 10232 -8592 10248
rect -9764 10168 -8676 10232
rect -8612 10168 -8592 10232
rect -9764 10152 -8592 10168
rect -9764 10088 -8676 10152
rect -8612 10088 -8592 10152
rect -9764 10072 -8592 10088
rect -9764 10008 -8676 10072
rect -8612 10008 -8592 10072
rect -9764 9992 -8592 10008
rect -9764 9928 -8676 9992
rect -8612 9928 -8592 9992
rect -9764 9912 -8592 9928
rect -9764 9848 -8676 9912
rect -8612 9848 -8592 9912
rect -9764 9832 -8592 9848
rect -9764 9768 -8676 9832
rect -8612 9768 -8592 9832
rect -9764 9752 -8592 9768
rect -9764 9688 -8676 9752
rect -8612 9688 -8592 9752
rect -9764 9640 -8592 9688
rect -8352 10472 -7180 10520
rect -8352 10408 -7264 10472
rect -7200 10408 -7180 10472
rect -8352 10392 -7180 10408
rect -8352 10328 -7264 10392
rect -7200 10328 -7180 10392
rect -8352 10312 -7180 10328
rect -8352 10248 -7264 10312
rect -7200 10248 -7180 10312
rect -8352 10232 -7180 10248
rect -8352 10168 -7264 10232
rect -7200 10168 -7180 10232
rect -8352 10152 -7180 10168
rect -8352 10088 -7264 10152
rect -7200 10088 -7180 10152
rect -8352 10072 -7180 10088
rect -8352 10008 -7264 10072
rect -7200 10008 -7180 10072
rect -8352 9992 -7180 10008
rect -8352 9928 -7264 9992
rect -7200 9928 -7180 9992
rect -8352 9912 -7180 9928
rect -8352 9848 -7264 9912
rect -7200 9848 -7180 9912
rect -8352 9832 -7180 9848
rect -8352 9768 -7264 9832
rect -7200 9768 -7180 9832
rect -8352 9752 -7180 9768
rect -8352 9688 -7264 9752
rect -7200 9688 -7180 9752
rect -8352 9640 -7180 9688
rect -6940 10472 -5768 10520
rect -6940 10408 -5852 10472
rect -5788 10408 -5768 10472
rect -6940 10392 -5768 10408
rect -6940 10328 -5852 10392
rect -5788 10328 -5768 10392
rect -6940 10312 -5768 10328
rect -6940 10248 -5852 10312
rect -5788 10248 -5768 10312
rect -6940 10232 -5768 10248
rect -6940 10168 -5852 10232
rect -5788 10168 -5768 10232
rect -6940 10152 -5768 10168
rect -6940 10088 -5852 10152
rect -5788 10088 -5768 10152
rect -6940 10072 -5768 10088
rect -6940 10008 -5852 10072
rect -5788 10008 -5768 10072
rect -6940 9992 -5768 10008
rect -6940 9928 -5852 9992
rect -5788 9928 -5768 9992
rect -6940 9912 -5768 9928
rect -6940 9848 -5852 9912
rect -5788 9848 -5768 9912
rect -6940 9832 -5768 9848
rect -6940 9768 -5852 9832
rect -5788 9768 -5768 9832
rect -6940 9752 -5768 9768
rect -6940 9688 -5852 9752
rect -5788 9688 -5768 9752
rect -6940 9640 -5768 9688
rect -5528 10472 -4356 10520
rect -5528 10408 -4440 10472
rect -4376 10408 -4356 10472
rect -5528 10392 -4356 10408
rect -5528 10328 -4440 10392
rect -4376 10328 -4356 10392
rect -5528 10312 -4356 10328
rect -5528 10248 -4440 10312
rect -4376 10248 -4356 10312
rect -5528 10232 -4356 10248
rect -5528 10168 -4440 10232
rect -4376 10168 -4356 10232
rect -5528 10152 -4356 10168
rect -5528 10088 -4440 10152
rect -4376 10088 -4356 10152
rect -5528 10072 -4356 10088
rect -5528 10008 -4440 10072
rect -4376 10008 -4356 10072
rect -5528 9992 -4356 10008
rect -5528 9928 -4440 9992
rect -4376 9928 -4356 9992
rect -5528 9912 -4356 9928
rect -5528 9848 -4440 9912
rect -4376 9848 -4356 9912
rect -5528 9832 -4356 9848
rect -5528 9768 -4440 9832
rect -4376 9768 -4356 9832
rect -5528 9752 -4356 9768
rect -5528 9688 -4440 9752
rect -4376 9688 -4356 9752
rect -5528 9640 -4356 9688
rect -4116 10472 -2944 10520
rect -4116 10408 -3028 10472
rect -2964 10408 -2944 10472
rect -4116 10392 -2944 10408
rect -4116 10328 -3028 10392
rect -2964 10328 -2944 10392
rect -4116 10312 -2944 10328
rect -4116 10248 -3028 10312
rect -2964 10248 -2944 10312
rect -4116 10232 -2944 10248
rect -4116 10168 -3028 10232
rect -2964 10168 -2944 10232
rect -4116 10152 -2944 10168
rect -4116 10088 -3028 10152
rect -2964 10088 -2944 10152
rect -4116 10072 -2944 10088
rect -4116 10008 -3028 10072
rect -2964 10008 -2944 10072
rect -4116 9992 -2944 10008
rect -4116 9928 -3028 9992
rect -2964 9928 -2944 9992
rect -4116 9912 -2944 9928
rect -4116 9848 -3028 9912
rect -2964 9848 -2944 9912
rect -4116 9832 -2944 9848
rect -4116 9768 -3028 9832
rect -2964 9768 -2944 9832
rect -4116 9752 -2944 9768
rect -4116 9688 -3028 9752
rect -2964 9688 -2944 9752
rect -4116 9640 -2944 9688
rect -2704 10472 -1532 10520
rect -2704 10408 -1616 10472
rect -1552 10408 -1532 10472
rect -2704 10392 -1532 10408
rect -2704 10328 -1616 10392
rect -1552 10328 -1532 10392
rect -2704 10312 -1532 10328
rect -2704 10248 -1616 10312
rect -1552 10248 -1532 10312
rect -2704 10232 -1532 10248
rect -2704 10168 -1616 10232
rect -1552 10168 -1532 10232
rect -2704 10152 -1532 10168
rect -2704 10088 -1616 10152
rect -1552 10088 -1532 10152
rect -2704 10072 -1532 10088
rect -2704 10008 -1616 10072
rect -1552 10008 -1532 10072
rect -2704 9992 -1532 10008
rect -2704 9928 -1616 9992
rect -1552 9928 -1532 9992
rect -2704 9912 -1532 9928
rect -2704 9848 -1616 9912
rect -1552 9848 -1532 9912
rect -2704 9832 -1532 9848
rect -2704 9768 -1616 9832
rect -1552 9768 -1532 9832
rect -2704 9752 -1532 9768
rect -2704 9688 -1616 9752
rect -1552 9688 -1532 9752
rect -2704 9640 -1532 9688
rect -1292 10472 -120 10520
rect -1292 10408 -204 10472
rect -140 10408 -120 10472
rect -1292 10392 -120 10408
rect -1292 10328 -204 10392
rect -140 10328 -120 10392
rect -1292 10312 -120 10328
rect -1292 10248 -204 10312
rect -140 10248 -120 10312
rect -1292 10232 -120 10248
rect -1292 10168 -204 10232
rect -140 10168 -120 10232
rect -1292 10152 -120 10168
rect -1292 10088 -204 10152
rect -140 10088 -120 10152
rect -1292 10072 -120 10088
rect -1292 10008 -204 10072
rect -140 10008 -120 10072
rect -1292 9992 -120 10008
rect -1292 9928 -204 9992
rect -140 9928 -120 9992
rect -1292 9912 -120 9928
rect -1292 9848 -204 9912
rect -140 9848 -120 9912
rect -1292 9832 -120 9848
rect -1292 9768 -204 9832
rect -140 9768 -120 9832
rect -1292 9752 -120 9768
rect -1292 9688 -204 9752
rect -140 9688 -120 9752
rect -1292 9640 -120 9688
rect 120 10472 1292 10520
rect 120 10408 1208 10472
rect 1272 10408 1292 10472
rect 120 10392 1292 10408
rect 120 10328 1208 10392
rect 1272 10328 1292 10392
rect 120 10312 1292 10328
rect 120 10248 1208 10312
rect 1272 10248 1292 10312
rect 120 10232 1292 10248
rect 120 10168 1208 10232
rect 1272 10168 1292 10232
rect 120 10152 1292 10168
rect 120 10088 1208 10152
rect 1272 10088 1292 10152
rect 120 10072 1292 10088
rect 120 10008 1208 10072
rect 1272 10008 1292 10072
rect 120 9992 1292 10008
rect 120 9928 1208 9992
rect 1272 9928 1292 9992
rect 120 9912 1292 9928
rect 120 9848 1208 9912
rect 1272 9848 1292 9912
rect 120 9832 1292 9848
rect 120 9768 1208 9832
rect 1272 9768 1292 9832
rect 120 9752 1292 9768
rect 120 9688 1208 9752
rect 1272 9688 1292 9752
rect 120 9640 1292 9688
rect 1532 10472 2704 10520
rect 1532 10408 2620 10472
rect 2684 10408 2704 10472
rect 1532 10392 2704 10408
rect 1532 10328 2620 10392
rect 2684 10328 2704 10392
rect 1532 10312 2704 10328
rect 1532 10248 2620 10312
rect 2684 10248 2704 10312
rect 1532 10232 2704 10248
rect 1532 10168 2620 10232
rect 2684 10168 2704 10232
rect 1532 10152 2704 10168
rect 1532 10088 2620 10152
rect 2684 10088 2704 10152
rect 1532 10072 2704 10088
rect 1532 10008 2620 10072
rect 2684 10008 2704 10072
rect 1532 9992 2704 10008
rect 1532 9928 2620 9992
rect 2684 9928 2704 9992
rect 1532 9912 2704 9928
rect 1532 9848 2620 9912
rect 2684 9848 2704 9912
rect 1532 9832 2704 9848
rect 1532 9768 2620 9832
rect 2684 9768 2704 9832
rect 1532 9752 2704 9768
rect 1532 9688 2620 9752
rect 2684 9688 2704 9752
rect 1532 9640 2704 9688
rect 2944 10472 4116 10520
rect 2944 10408 4032 10472
rect 4096 10408 4116 10472
rect 2944 10392 4116 10408
rect 2944 10328 4032 10392
rect 4096 10328 4116 10392
rect 2944 10312 4116 10328
rect 2944 10248 4032 10312
rect 4096 10248 4116 10312
rect 2944 10232 4116 10248
rect 2944 10168 4032 10232
rect 4096 10168 4116 10232
rect 2944 10152 4116 10168
rect 2944 10088 4032 10152
rect 4096 10088 4116 10152
rect 2944 10072 4116 10088
rect 2944 10008 4032 10072
rect 4096 10008 4116 10072
rect 2944 9992 4116 10008
rect 2944 9928 4032 9992
rect 4096 9928 4116 9992
rect 2944 9912 4116 9928
rect 2944 9848 4032 9912
rect 4096 9848 4116 9912
rect 2944 9832 4116 9848
rect 2944 9768 4032 9832
rect 4096 9768 4116 9832
rect 2944 9752 4116 9768
rect 2944 9688 4032 9752
rect 4096 9688 4116 9752
rect 2944 9640 4116 9688
rect 4356 10472 5528 10520
rect 4356 10408 5444 10472
rect 5508 10408 5528 10472
rect 4356 10392 5528 10408
rect 4356 10328 5444 10392
rect 5508 10328 5528 10392
rect 4356 10312 5528 10328
rect 4356 10248 5444 10312
rect 5508 10248 5528 10312
rect 4356 10232 5528 10248
rect 4356 10168 5444 10232
rect 5508 10168 5528 10232
rect 4356 10152 5528 10168
rect 4356 10088 5444 10152
rect 5508 10088 5528 10152
rect 4356 10072 5528 10088
rect 4356 10008 5444 10072
rect 5508 10008 5528 10072
rect 4356 9992 5528 10008
rect 4356 9928 5444 9992
rect 5508 9928 5528 9992
rect 4356 9912 5528 9928
rect 4356 9848 5444 9912
rect 5508 9848 5528 9912
rect 4356 9832 5528 9848
rect 4356 9768 5444 9832
rect 5508 9768 5528 9832
rect 4356 9752 5528 9768
rect 4356 9688 5444 9752
rect 5508 9688 5528 9752
rect 4356 9640 5528 9688
rect 5768 10472 6940 10520
rect 5768 10408 6856 10472
rect 6920 10408 6940 10472
rect 5768 10392 6940 10408
rect 5768 10328 6856 10392
rect 6920 10328 6940 10392
rect 5768 10312 6940 10328
rect 5768 10248 6856 10312
rect 6920 10248 6940 10312
rect 5768 10232 6940 10248
rect 5768 10168 6856 10232
rect 6920 10168 6940 10232
rect 5768 10152 6940 10168
rect 5768 10088 6856 10152
rect 6920 10088 6940 10152
rect 5768 10072 6940 10088
rect 5768 10008 6856 10072
rect 6920 10008 6940 10072
rect 5768 9992 6940 10008
rect 5768 9928 6856 9992
rect 6920 9928 6940 9992
rect 5768 9912 6940 9928
rect 5768 9848 6856 9912
rect 6920 9848 6940 9912
rect 5768 9832 6940 9848
rect 5768 9768 6856 9832
rect 6920 9768 6940 9832
rect 5768 9752 6940 9768
rect 5768 9688 6856 9752
rect 6920 9688 6940 9752
rect 5768 9640 6940 9688
rect 7180 10472 8352 10520
rect 7180 10408 8268 10472
rect 8332 10408 8352 10472
rect 7180 10392 8352 10408
rect 7180 10328 8268 10392
rect 8332 10328 8352 10392
rect 7180 10312 8352 10328
rect 7180 10248 8268 10312
rect 8332 10248 8352 10312
rect 7180 10232 8352 10248
rect 7180 10168 8268 10232
rect 8332 10168 8352 10232
rect 7180 10152 8352 10168
rect 7180 10088 8268 10152
rect 8332 10088 8352 10152
rect 7180 10072 8352 10088
rect 7180 10008 8268 10072
rect 8332 10008 8352 10072
rect 7180 9992 8352 10008
rect 7180 9928 8268 9992
rect 8332 9928 8352 9992
rect 7180 9912 8352 9928
rect 7180 9848 8268 9912
rect 8332 9848 8352 9912
rect 7180 9832 8352 9848
rect 7180 9768 8268 9832
rect 8332 9768 8352 9832
rect 7180 9752 8352 9768
rect 7180 9688 8268 9752
rect 8332 9688 8352 9752
rect 7180 9640 8352 9688
rect 8592 10472 9764 10520
rect 8592 10408 9680 10472
rect 9744 10408 9764 10472
rect 8592 10392 9764 10408
rect 8592 10328 9680 10392
rect 9744 10328 9764 10392
rect 8592 10312 9764 10328
rect 8592 10248 9680 10312
rect 9744 10248 9764 10312
rect 8592 10232 9764 10248
rect 8592 10168 9680 10232
rect 9744 10168 9764 10232
rect 8592 10152 9764 10168
rect 8592 10088 9680 10152
rect 9744 10088 9764 10152
rect 8592 10072 9764 10088
rect 8592 10008 9680 10072
rect 9744 10008 9764 10072
rect 8592 9992 9764 10008
rect 8592 9928 9680 9992
rect 9744 9928 9764 9992
rect 8592 9912 9764 9928
rect 8592 9848 9680 9912
rect 9744 9848 9764 9912
rect 8592 9832 9764 9848
rect 8592 9768 9680 9832
rect 9744 9768 9764 9832
rect 8592 9752 9764 9768
rect 8592 9688 9680 9752
rect 9744 9688 9764 9752
rect 8592 9640 9764 9688
rect 10004 10472 11176 10520
rect 10004 10408 11092 10472
rect 11156 10408 11176 10472
rect 10004 10392 11176 10408
rect 10004 10328 11092 10392
rect 11156 10328 11176 10392
rect 10004 10312 11176 10328
rect 10004 10248 11092 10312
rect 11156 10248 11176 10312
rect 10004 10232 11176 10248
rect 10004 10168 11092 10232
rect 11156 10168 11176 10232
rect 10004 10152 11176 10168
rect 10004 10088 11092 10152
rect 11156 10088 11176 10152
rect 10004 10072 11176 10088
rect 10004 10008 11092 10072
rect 11156 10008 11176 10072
rect 10004 9992 11176 10008
rect 10004 9928 11092 9992
rect 11156 9928 11176 9992
rect 10004 9912 11176 9928
rect 10004 9848 11092 9912
rect 11156 9848 11176 9912
rect 10004 9832 11176 9848
rect 10004 9768 11092 9832
rect 11156 9768 11176 9832
rect 10004 9752 11176 9768
rect 10004 9688 11092 9752
rect 11156 9688 11176 9752
rect 10004 9640 11176 9688
rect 11416 10472 12588 10520
rect 11416 10408 12504 10472
rect 12568 10408 12588 10472
rect 11416 10392 12588 10408
rect 11416 10328 12504 10392
rect 12568 10328 12588 10392
rect 11416 10312 12588 10328
rect 11416 10248 12504 10312
rect 12568 10248 12588 10312
rect 11416 10232 12588 10248
rect 11416 10168 12504 10232
rect 12568 10168 12588 10232
rect 11416 10152 12588 10168
rect 11416 10088 12504 10152
rect 12568 10088 12588 10152
rect 11416 10072 12588 10088
rect 11416 10008 12504 10072
rect 12568 10008 12588 10072
rect 11416 9992 12588 10008
rect 11416 9928 12504 9992
rect 12568 9928 12588 9992
rect 11416 9912 12588 9928
rect 11416 9848 12504 9912
rect 12568 9848 12588 9912
rect 11416 9832 12588 9848
rect 11416 9768 12504 9832
rect 12568 9768 12588 9832
rect 11416 9752 12588 9768
rect 11416 9688 12504 9752
rect 12568 9688 12588 9752
rect 11416 9640 12588 9688
rect 12828 10472 14000 10520
rect 12828 10408 13916 10472
rect 13980 10408 14000 10472
rect 12828 10392 14000 10408
rect 12828 10328 13916 10392
rect 13980 10328 14000 10392
rect 12828 10312 14000 10328
rect 12828 10248 13916 10312
rect 13980 10248 14000 10312
rect 12828 10232 14000 10248
rect 12828 10168 13916 10232
rect 13980 10168 14000 10232
rect 12828 10152 14000 10168
rect 12828 10088 13916 10152
rect 13980 10088 14000 10152
rect 12828 10072 14000 10088
rect 12828 10008 13916 10072
rect 13980 10008 14000 10072
rect 12828 9992 14000 10008
rect 12828 9928 13916 9992
rect 13980 9928 14000 9992
rect 12828 9912 14000 9928
rect 12828 9848 13916 9912
rect 13980 9848 14000 9912
rect 12828 9832 14000 9848
rect 12828 9768 13916 9832
rect 13980 9768 14000 9832
rect 12828 9752 14000 9768
rect 12828 9688 13916 9752
rect 13980 9688 14000 9752
rect 12828 9640 14000 9688
rect 14240 10472 15412 10520
rect 14240 10408 15328 10472
rect 15392 10408 15412 10472
rect 14240 10392 15412 10408
rect 14240 10328 15328 10392
rect 15392 10328 15412 10392
rect 14240 10312 15412 10328
rect 14240 10248 15328 10312
rect 15392 10248 15412 10312
rect 14240 10232 15412 10248
rect 14240 10168 15328 10232
rect 15392 10168 15412 10232
rect 14240 10152 15412 10168
rect 14240 10088 15328 10152
rect 15392 10088 15412 10152
rect 14240 10072 15412 10088
rect 14240 10008 15328 10072
rect 15392 10008 15412 10072
rect 14240 9992 15412 10008
rect 14240 9928 15328 9992
rect 15392 9928 15412 9992
rect 14240 9912 15412 9928
rect 14240 9848 15328 9912
rect 15392 9848 15412 9912
rect 14240 9832 15412 9848
rect 14240 9768 15328 9832
rect 15392 9768 15412 9832
rect 14240 9752 15412 9768
rect 14240 9688 15328 9752
rect 15392 9688 15412 9752
rect 14240 9640 15412 9688
rect 15652 10472 16824 10520
rect 15652 10408 16740 10472
rect 16804 10408 16824 10472
rect 15652 10392 16824 10408
rect 15652 10328 16740 10392
rect 16804 10328 16824 10392
rect 15652 10312 16824 10328
rect 15652 10248 16740 10312
rect 16804 10248 16824 10312
rect 15652 10232 16824 10248
rect 15652 10168 16740 10232
rect 16804 10168 16824 10232
rect 15652 10152 16824 10168
rect 15652 10088 16740 10152
rect 16804 10088 16824 10152
rect 15652 10072 16824 10088
rect 15652 10008 16740 10072
rect 16804 10008 16824 10072
rect 15652 9992 16824 10008
rect 15652 9928 16740 9992
rect 16804 9928 16824 9992
rect 15652 9912 16824 9928
rect 15652 9848 16740 9912
rect 16804 9848 16824 9912
rect 15652 9832 16824 9848
rect 15652 9768 16740 9832
rect 16804 9768 16824 9832
rect 15652 9752 16824 9768
rect 15652 9688 16740 9752
rect 16804 9688 16824 9752
rect 15652 9640 16824 9688
rect 17064 10472 18236 10520
rect 17064 10408 18152 10472
rect 18216 10408 18236 10472
rect 17064 10392 18236 10408
rect 17064 10328 18152 10392
rect 18216 10328 18236 10392
rect 17064 10312 18236 10328
rect 17064 10248 18152 10312
rect 18216 10248 18236 10312
rect 17064 10232 18236 10248
rect 17064 10168 18152 10232
rect 18216 10168 18236 10232
rect 17064 10152 18236 10168
rect 17064 10088 18152 10152
rect 18216 10088 18236 10152
rect 17064 10072 18236 10088
rect 17064 10008 18152 10072
rect 18216 10008 18236 10072
rect 17064 9992 18236 10008
rect 17064 9928 18152 9992
rect 18216 9928 18236 9992
rect 17064 9912 18236 9928
rect 17064 9848 18152 9912
rect 18216 9848 18236 9912
rect 17064 9832 18236 9848
rect 17064 9768 18152 9832
rect 18216 9768 18236 9832
rect 17064 9752 18236 9768
rect 17064 9688 18152 9752
rect 18216 9688 18236 9752
rect 17064 9640 18236 9688
rect 18476 10472 19648 10520
rect 18476 10408 19564 10472
rect 19628 10408 19648 10472
rect 18476 10392 19648 10408
rect 18476 10328 19564 10392
rect 19628 10328 19648 10392
rect 18476 10312 19648 10328
rect 18476 10248 19564 10312
rect 19628 10248 19648 10312
rect 18476 10232 19648 10248
rect 18476 10168 19564 10232
rect 19628 10168 19648 10232
rect 18476 10152 19648 10168
rect 18476 10088 19564 10152
rect 19628 10088 19648 10152
rect 18476 10072 19648 10088
rect 18476 10008 19564 10072
rect 19628 10008 19648 10072
rect 18476 9992 19648 10008
rect 18476 9928 19564 9992
rect 19628 9928 19648 9992
rect 18476 9912 19648 9928
rect 18476 9848 19564 9912
rect 19628 9848 19648 9912
rect 18476 9832 19648 9848
rect 18476 9768 19564 9832
rect 19628 9768 19648 9832
rect 18476 9752 19648 9768
rect 18476 9688 19564 9752
rect 19628 9688 19648 9752
rect 18476 9640 19648 9688
rect 19888 10472 21060 10520
rect 19888 10408 20976 10472
rect 21040 10408 21060 10472
rect 19888 10392 21060 10408
rect 19888 10328 20976 10392
rect 21040 10328 21060 10392
rect 19888 10312 21060 10328
rect 19888 10248 20976 10312
rect 21040 10248 21060 10312
rect 19888 10232 21060 10248
rect 19888 10168 20976 10232
rect 21040 10168 21060 10232
rect 19888 10152 21060 10168
rect 19888 10088 20976 10152
rect 21040 10088 21060 10152
rect 19888 10072 21060 10088
rect 19888 10008 20976 10072
rect 21040 10008 21060 10072
rect 19888 9992 21060 10008
rect 19888 9928 20976 9992
rect 21040 9928 21060 9992
rect 19888 9912 21060 9928
rect 19888 9848 20976 9912
rect 21040 9848 21060 9912
rect 19888 9832 21060 9848
rect 19888 9768 20976 9832
rect 21040 9768 21060 9832
rect 19888 9752 21060 9768
rect 19888 9688 20976 9752
rect 21040 9688 21060 9752
rect 19888 9640 21060 9688
rect 21300 10472 22472 10520
rect 21300 10408 22388 10472
rect 22452 10408 22472 10472
rect 21300 10392 22472 10408
rect 21300 10328 22388 10392
rect 22452 10328 22472 10392
rect 21300 10312 22472 10328
rect 21300 10248 22388 10312
rect 22452 10248 22472 10312
rect 21300 10232 22472 10248
rect 21300 10168 22388 10232
rect 22452 10168 22472 10232
rect 21300 10152 22472 10168
rect 21300 10088 22388 10152
rect 22452 10088 22472 10152
rect 21300 10072 22472 10088
rect 21300 10008 22388 10072
rect 22452 10008 22472 10072
rect 21300 9992 22472 10008
rect 21300 9928 22388 9992
rect 22452 9928 22472 9992
rect 21300 9912 22472 9928
rect 21300 9848 22388 9912
rect 22452 9848 22472 9912
rect 21300 9832 22472 9848
rect 21300 9768 22388 9832
rect 22452 9768 22472 9832
rect 21300 9752 22472 9768
rect 21300 9688 22388 9752
rect 22452 9688 22472 9752
rect 21300 9640 22472 9688
rect 22712 10472 23884 10520
rect 22712 10408 23800 10472
rect 23864 10408 23884 10472
rect 22712 10392 23884 10408
rect 22712 10328 23800 10392
rect 23864 10328 23884 10392
rect 22712 10312 23884 10328
rect 22712 10248 23800 10312
rect 23864 10248 23884 10312
rect 22712 10232 23884 10248
rect 22712 10168 23800 10232
rect 23864 10168 23884 10232
rect 22712 10152 23884 10168
rect 22712 10088 23800 10152
rect 23864 10088 23884 10152
rect 22712 10072 23884 10088
rect 22712 10008 23800 10072
rect 23864 10008 23884 10072
rect 22712 9992 23884 10008
rect 22712 9928 23800 9992
rect 23864 9928 23884 9992
rect 22712 9912 23884 9928
rect 22712 9848 23800 9912
rect 23864 9848 23884 9912
rect 22712 9832 23884 9848
rect 22712 9768 23800 9832
rect 23864 9768 23884 9832
rect 22712 9752 23884 9768
rect 22712 9688 23800 9752
rect 23864 9688 23884 9752
rect 22712 9640 23884 9688
rect -23884 9352 -22712 9400
rect -23884 9288 -22796 9352
rect -22732 9288 -22712 9352
rect -23884 9272 -22712 9288
rect -23884 9208 -22796 9272
rect -22732 9208 -22712 9272
rect -23884 9192 -22712 9208
rect -23884 9128 -22796 9192
rect -22732 9128 -22712 9192
rect -23884 9112 -22712 9128
rect -23884 9048 -22796 9112
rect -22732 9048 -22712 9112
rect -23884 9032 -22712 9048
rect -23884 8968 -22796 9032
rect -22732 8968 -22712 9032
rect -23884 8952 -22712 8968
rect -23884 8888 -22796 8952
rect -22732 8888 -22712 8952
rect -23884 8872 -22712 8888
rect -23884 8808 -22796 8872
rect -22732 8808 -22712 8872
rect -23884 8792 -22712 8808
rect -23884 8728 -22796 8792
rect -22732 8728 -22712 8792
rect -23884 8712 -22712 8728
rect -23884 8648 -22796 8712
rect -22732 8648 -22712 8712
rect -23884 8632 -22712 8648
rect -23884 8568 -22796 8632
rect -22732 8568 -22712 8632
rect -23884 8520 -22712 8568
rect -22472 9352 -21300 9400
rect -22472 9288 -21384 9352
rect -21320 9288 -21300 9352
rect -22472 9272 -21300 9288
rect -22472 9208 -21384 9272
rect -21320 9208 -21300 9272
rect -22472 9192 -21300 9208
rect -22472 9128 -21384 9192
rect -21320 9128 -21300 9192
rect -22472 9112 -21300 9128
rect -22472 9048 -21384 9112
rect -21320 9048 -21300 9112
rect -22472 9032 -21300 9048
rect -22472 8968 -21384 9032
rect -21320 8968 -21300 9032
rect -22472 8952 -21300 8968
rect -22472 8888 -21384 8952
rect -21320 8888 -21300 8952
rect -22472 8872 -21300 8888
rect -22472 8808 -21384 8872
rect -21320 8808 -21300 8872
rect -22472 8792 -21300 8808
rect -22472 8728 -21384 8792
rect -21320 8728 -21300 8792
rect -22472 8712 -21300 8728
rect -22472 8648 -21384 8712
rect -21320 8648 -21300 8712
rect -22472 8632 -21300 8648
rect -22472 8568 -21384 8632
rect -21320 8568 -21300 8632
rect -22472 8520 -21300 8568
rect -21060 9352 -19888 9400
rect -21060 9288 -19972 9352
rect -19908 9288 -19888 9352
rect -21060 9272 -19888 9288
rect -21060 9208 -19972 9272
rect -19908 9208 -19888 9272
rect -21060 9192 -19888 9208
rect -21060 9128 -19972 9192
rect -19908 9128 -19888 9192
rect -21060 9112 -19888 9128
rect -21060 9048 -19972 9112
rect -19908 9048 -19888 9112
rect -21060 9032 -19888 9048
rect -21060 8968 -19972 9032
rect -19908 8968 -19888 9032
rect -21060 8952 -19888 8968
rect -21060 8888 -19972 8952
rect -19908 8888 -19888 8952
rect -21060 8872 -19888 8888
rect -21060 8808 -19972 8872
rect -19908 8808 -19888 8872
rect -21060 8792 -19888 8808
rect -21060 8728 -19972 8792
rect -19908 8728 -19888 8792
rect -21060 8712 -19888 8728
rect -21060 8648 -19972 8712
rect -19908 8648 -19888 8712
rect -21060 8632 -19888 8648
rect -21060 8568 -19972 8632
rect -19908 8568 -19888 8632
rect -21060 8520 -19888 8568
rect -19648 9352 -18476 9400
rect -19648 9288 -18560 9352
rect -18496 9288 -18476 9352
rect -19648 9272 -18476 9288
rect -19648 9208 -18560 9272
rect -18496 9208 -18476 9272
rect -19648 9192 -18476 9208
rect -19648 9128 -18560 9192
rect -18496 9128 -18476 9192
rect -19648 9112 -18476 9128
rect -19648 9048 -18560 9112
rect -18496 9048 -18476 9112
rect -19648 9032 -18476 9048
rect -19648 8968 -18560 9032
rect -18496 8968 -18476 9032
rect -19648 8952 -18476 8968
rect -19648 8888 -18560 8952
rect -18496 8888 -18476 8952
rect -19648 8872 -18476 8888
rect -19648 8808 -18560 8872
rect -18496 8808 -18476 8872
rect -19648 8792 -18476 8808
rect -19648 8728 -18560 8792
rect -18496 8728 -18476 8792
rect -19648 8712 -18476 8728
rect -19648 8648 -18560 8712
rect -18496 8648 -18476 8712
rect -19648 8632 -18476 8648
rect -19648 8568 -18560 8632
rect -18496 8568 -18476 8632
rect -19648 8520 -18476 8568
rect -18236 9352 -17064 9400
rect -18236 9288 -17148 9352
rect -17084 9288 -17064 9352
rect -18236 9272 -17064 9288
rect -18236 9208 -17148 9272
rect -17084 9208 -17064 9272
rect -18236 9192 -17064 9208
rect -18236 9128 -17148 9192
rect -17084 9128 -17064 9192
rect -18236 9112 -17064 9128
rect -18236 9048 -17148 9112
rect -17084 9048 -17064 9112
rect -18236 9032 -17064 9048
rect -18236 8968 -17148 9032
rect -17084 8968 -17064 9032
rect -18236 8952 -17064 8968
rect -18236 8888 -17148 8952
rect -17084 8888 -17064 8952
rect -18236 8872 -17064 8888
rect -18236 8808 -17148 8872
rect -17084 8808 -17064 8872
rect -18236 8792 -17064 8808
rect -18236 8728 -17148 8792
rect -17084 8728 -17064 8792
rect -18236 8712 -17064 8728
rect -18236 8648 -17148 8712
rect -17084 8648 -17064 8712
rect -18236 8632 -17064 8648
rect -18236 8568 -17148 8632
rect -17084 8568 -17064 8632
rect -18236 8520 -17064 8568
rect -16824 9352 -15652 9400
rect -16824 9288 -15736 9352
rect -15672 9288 -15652 9352
rect -16824 9272 -15652 9288
rect -16824 9208 -15736 9272
rect -15672 9208 -15652 9272
rect -16824 9192 -15652 9208
rect -16824 9128 -15736 9192
rect -15672 9128 -15652 9192
rect -16824 9112 -15652 9128
rect -16824 9048 -15736 9112
rect -15672 9048 -15652 9112
rect -16824 9032 -15652 9048
rect -16824 8968 -15736 9032
rect -15672 8968 -15652 9032
rect -16824 8952 -15652 8968
rect -16824 8888 -15736 8952
rect -15672 8888 -15652 8952
rect -16824 8872 -15652 8888
rect -16824 8808 -15736 8872
rect -15672 8808 -15652 8872
rect -16824 8792 -15652 8808
rect -16824 8728 -15736 8792
rect -15672 8728 -15652 8792
rect -16824 8712 -15652 8728
rect -16824 8648 -15736 8712
rect -15672 8648 -15652 8712
rect -16824 8632 -15652 8648
rect -16824 8568 -15736 8632
rect -15672 8568 -15652 8632
rect -16824 8520 -15652 8568
rect -15412 9352 -14240 9400
rect -15412 9288 -14324 9352
rect -14260 9288 -14240 9352
rect -15412 9272 -14240 9288
rect -15412 9208 -14324 9272
rect -14260 9208 -14240 9272
rect -15412 9192 -14240 9208
rect -15412 9128 -14324 9192
rect -14260 9128 -14240 9192
rect -15412 9112 -14240 9128
rect -15412 9048 -14324 9112
rect -14260 9048 -14240 9112
rect -15412 9032 -14240 9048
rect -15412 8968 -14324 9032
rect -14260 8968 -14240 9032
rect -15412 8952 -14240 8968
rect -15412 8888 -14324 8952
rect -14260 8888 -14240 8952
rect -15412 8872 -14240 8888
rect -15412 8808 -14324 8872
rect -14260 8808 -14240 8872
rect -15412 8792 -14240 8808
rect -15412 8728 -14324 8792
rect -14260 8728 -14240 8792
rect -15412 8712 -14240 8728
rect -15412 8648 -14324 8712
rect -14260 8648 -14240 8712
rect -15412 8632 -14240 8648
rect -15412 8568 -14324 8632
rect -14260 8568 -14240 8632
rect -15412 8520 -14240 8568
rect -14000 9352 -12828 9400
rect -14000 9288 -12912 9352
rect -12848 9288 -12828 9352
rect -14000 9272 -12828 9288
rect -14000 9208 -12912 9272
rect -12848 9208 -12828 9272
rect -14000 9192 -12828 9208
rect -14000 9128 -12912 9192
rect -12848 9128 -12828 9192
rect -14000 9112 -12828 9128
rect -14000 9048 -12912 9112
rect -12848 9048 -12828 9112
rect -14000 9032 -12828 9048
rect -14000 8968 -12912 9032
rect -12848 8968 -12828 9032
rect -14000 8952 -12828 8968
rect -14000 8888 -12912 8952
rect -12848 8888 -12828 8952
rect -14000 8872 -12828 8888
rect -14000 8808 -12912 8872
rect -12848 8808 -12828 8872
rect -14000 8792 -12828 8808
rect -14000 8728 -12912 8792
rect -12848 8728 -12828 8792
rect -14000 8712 -12828 8728
rect -14000 8648 -12912 8712
rect -12848 8648 -12828 8712
rect -14000 8632 -12828 8648
rect -14000 8568 -12912 8632
rect -12848 8568 -12828 8632
rect -14000 8520 -12828 8568
rect -12588 9352 -11416 9400
rect -12588 9288 -11500 9352
rect -11436 9288 -11416 9352
rect -12588 9272 -11416 9288
rect -12588 9208 -11500 9272
rect -11436 9208 -11416 9272
rect -12588 9192 -11416 9208
rect -12588 9128 -11500 9192
rect -11436 9128 -11416 9192
rect -12588 9112 -11416 9128
rect -12588 9048 -11500 9112
rect -11436 9048 -11416 9112
rect -12588 9032 -11416 9048
rect -12588 8968 -11500 9032
rect -11436 8968 -11416 9032
rect -12588 8952 -11416 8968
rect -12588 8888 -11500 8952
rect -11436 8888 -11416 8952
rect -12588 8872 -11416 8888
rect -12588 8808 -11500 8872
rect -11436 8808 -11416 8872
rect -12588 8792 -11416 8808
rect -12588 8728 -11500 8792
rect -11436 8728 -11416 8792
rect -12588 8712 -11416 8728
rect -12588 8648 -11500 8712
rect -11436 8648 -11416 8712
rect -12588 8632 -11416 8648
rect -12588 8568 -11500 8632
rect -11436 8568 -11416 8632
rect -12588 8520 -11416 8568
rect -11176 9352 -10004 9400
rect -11176 9288 -10088 9352
rect -10024 9288 -10004 9352
rect -11176 9272 -10004 9288
rect -11176 9208 -10088 9272
rect -10024 9208 -10004 9272
rect -11176 9192 -10004 9208
rect -11176 9128 -10088 9192
rect -10024 9128 -10004 9192
rect -11176 9112 -10004 9128
rect -11176 9048 -10088 9112
rect -10024 9048 -10004 9112
rect -11176 9032 -10004 9048
rect -11176 8968 -10088 9032
rect -10024 8968 -10004 9032
rect -11176 8952 -10004 8968
rect -11176 8888 -10088 8952
rect -10024 8888 -10004 8952
rect -11176 8872 -10004 8888
rect -11176 8808 -10088 8872
rect -10024 8808 -10004 8872
rect -11176 8792 -10004 8808
rect -11176 8728 -10088 8792
rect -10024 8728 -10004 8792
rect -11176 8712 -10004 8728
rect -11176 8648 -10088 8712
rect -10024 8648 -10004 8712
rect -11176 8632 -10004 8648
rect -11176 8568 -10088 8632
rect -10024 8568 -10004 8632
rect -11176 8520 -10004 8568
rect -9764 9352 -8592 9400
rect -9764 9288 -8676 9352
rect -8612 9288 -8592 9352
rect -9764 9272 -8592 9288
rect -9764 9208 -8676 9272
rect -8612 9208 -8592 9272
rect -9764 9192 -8592 9208
rect -9764 9128 -8676 9192
rect -8612 9128 -8592 9192
rect -9764 9112 -8592 9128
rect -9764 9048 -8676 9112
rect -8612 9048 -8592 9112
rect -9764 9032 -8592 9048
rect -9764 8968 -8676 9032
rect -8612 8968 -8592 9032
rect -9764 8952 -8592 8968
rect -9764 8888 -8676 8952
rect -8612 8888 -8592 8952
rect -9764 8872 -8592 8888
rect -9764 8808 -8676 8872
rect -8612 8808 -8592 8872
rect -9764 8792 -8592 8808
rect -9764 8728 -8676 8792
rect -8612 8728 -8592 8792
rect -9764 8712 -8592 8728
rect -9764 8648 -8676 8712
rect -8612 8648 -8592 8712
rect -9764 8632 -8592 8648
rect -9764 8568 -8676 8632
rect -8612 8568 -8592 8632
rect -9764 8520 -8592 8568
rect -8352 9352 -7180 9400
rect -8352 9288 -7264 9352
rect -7200 9288 -7180 9352
rect -8352 9272 -7180 9288
rect -8352 9208 -7264 9272
rect -7200 9208 -7180 9272
rect -8352 9192 -7180 9208
rect -8352 9128 -7264 9192
rect -7200 9128 -7180 9192
rect -8352 9112 -7180 9128
rect -8352 9048 -7264 9112
rect -7200 9048 -7180 9112
rect -8352 9032 -7180 9048
rect -8352 8968 -7264 9032
rect -7200 8968 -7180 9032
rect -8352 8952 -7180 8968
rect -8352 8888 -7264 8952
rect -7200 8888 -7180 8952
rect -8352 8872 -7180 8888
rect -8352 8808 -7264 8872
rect -7200 8808 -7180 8872
rect -8352 8792 -7180 8808
rect -8352 8728 -7264 8792
rect -7200 8728 -7180 8792
rect -8352 8712 -7180 8728
rect -8352 8648 -7264 8712
rect -7200 8648 -7180 8712
rect -8352 8632 -7180 8648
rect -8352 8568 -7264 8632
rect -7200 8568 -7180 8632
rect -8352 8520 -7180 8568
rect -6940 9352 -5768 9400
rect -6940 9288 -5852 9352
rect -5788 9288 -5768 9352
rect -6940 9272 -5768 9288
rect -6940 9208 -5852 9272
rect -5788 9208 -5768 9272
rect -6940 9192 -5768 9208
rect -6940 9128 -5852 9192
rect -5788 9128 -5768 9192
rect -6940 9112 -5768 9128
rect -6940 9048 -5852 9112
rect -5788 9048 -5768 9112
rect -6940 9032 -5768 9048
rect -6940 8968 -5852 9032
rect -5788 8968 -5768 9032
rect -6940 8952 -5768 8968
rect -6940 8888 -5852 8952
rect -5788 8888 -5768 8952
rect -6940 8872 -5768 8888
rect -6940 8808 -5852 8872
rect -5788 8808 -5768 8872
rect -6940 8792 -5768 8808
rect -6940 8728 -5852 8792
rect -5788 8728 -5768 8792
rect -6940 8712 -5768 8728
rect -6940 8648 -5852 8712
rect -5788 8648 -5768 8712
rect -6940 8632 -5768 8648
rect -6940 8568 -5852 8632
rect -5788 8568 -5768 8632
rect -6940 8520 -5768 8568
rect -5528 9352 -4356 9400
rect -5528 9288 -4440 9352
rect -4376 9288 -4356 9352
rect -5528 9272 -4356 9288
rect -5528 9208 -4440 9272
rect -4376 9208 -4356 9272
rect -5528 9192 -4356 9208
rect -5528 9128 -4440 9192
rect -4376 9128 -4356 9192
rect -5528 9112 -4356 9128
rect -5528 9048 -4440 9112
rect -4376 9048 -4356 9112
rect -5528 9032 -4356 9048
rect -5528 8968 -4440 9032
rect -4376 8968 -4356 9032
rect -5528 8952 -4356 8968
rect -5528 8888 -4440 8952
rect -4376 8888 -4356 8952
rect -5528 8872 -4356 8888
rect -5528 8808 -4440 8872
rect -4376 8808 -4356 8872
rect -5528 8792 -4356 8808
rect -5528 8728 -4440 8792
rect -4376 8728 -4356 8792
rect -5528 8712 -4356 8728
rect -5528 8648 -4440 8712
rect -4376 8648 -4356 8712
rect -5528 8632 -4356 8648
rect -5528 8568 -4440 8632
rect -4376 8568 -4356 8632
rect -5528 8520 -4356 8568
rect -4116 9352 -2944 9400
rect -4116 9288 -3028 9352
rect -2964 9288 -2944 9352
rect -4116 9272 -2944 9288
rect -4116 9208 -3028 9272
rect -2964 9208 -2944 9272
rect -4116 9192 -2944 9208
rect -4116 9128 -3028 9192
rect -2964 9128 -2944 9192
rect -4116 9112 -2944 9128
rect -4116 9048 -3028 9112
rect -2964 9048 -2944 9112
rect -4116 9032 -2944 9048
rect -4116 8968 -3028 9032
rect -2964 8968 -2944 9032
rect -4116 8952 -2944 8968
rect -4116 8888 -3028 8952
rect -2964 8888 -2944 8952
rect -4116 8872 -2944 8888
rect -4116 8808 -3028 8872
rect -2964 8808 -2944 8872
rect -4116 8792 -2944 8808
rect -4116 8728 -3028 8792
rect -2964 8728 -2944 8792
rect -4116 8712 -2944 8728
rect -4116 8648 -3028 8712
rect -2964 8648 -2944 8712
rect -4116 8632 -2944 8648
rect -4116 8568 -3028 8632
rect -2964 8568 -2944 8632
rect -4116 8520 -2944 8568
rect -2704 9352 -1532 9400
rect -2704 9288 -1616 9352
rect -1552 9288 -1532 9352
rect -2704 9272 -1532 9288
rect -2704 9208 -1616 9272
rect -1552 9208 -1532 9272
rect -2704 9192 -1532 9208
rect -2704 9128 -1616 9192
rect -1552 9128 -1532 9192
rect -2704 9112 -1532 9128
rect -2704 9048 -1616 9112
rect -1552 9048 -1532 9112
rect -2704 9032 -1532 9048
rect -2704 8968 -1616 9032
rect -1552 8968 -1532 9032
rect -2704 8952 -1532 8968
rect -2704 8888 -1616 8952
rect -1552 8888 -1532 8952
rect -2704 8872 -1532 8888
rect -2704 8808 -1616 8872
rect -1552 8808 -1532 8872
rect -2704 8792 -1532 8808
rect -2704 8728 -1616 8792
rect -1552 8728 -1532 8792
rect -2704 8712 -1532 8728
rect -2704 8648 -1616 8712
rect -1552 8648 -1532 8712
rect -2704 8632 -1532 8648
rect -2704 8568 -1616 8632
rect -1552 8568 -1532 8632
rect -2704 8520 -1532 8568
rect -1292 9352 -120 9400
rect -1292 9288 -204 9352
rect -140 9288 -120 9352
rect -1292 9272 -120 9288
rect -1292 9208 -204 9272
rect -140 9208 -120 9272
rect -1292 9192 -120 9208
rect -1292 9128 -204 9192
rect -140 9128 -120 9192
rect -1292 9112 -120 9128
rect -1292 9048 -204 9112
rect -140 9048 -120 9112
rect -1292 9032 -120 9048
rect -1292 8968 -204 9032
rect -140 8968 -120 9032
rect -1292 8952 -120 8968
rect -1292 8888 -204 8952
rect -140 8888 -120 8952
rect -1292 8872 -120 8888
rect -1292 8808 -204 8872
rect -140 8808 -120 8872
rect -1292 8792 -120 8808
rect -1292 8728 -204 8792
rect -140 8728 -120 8792
rect -1292 8712 -120 8728
rect -1292 8648 -204 8712
rect -140 8648 -120 8712
rect -1292 8632 -120 8648
rect -1292 8568 -204 8632
rect -140 8568 -120 8632
rect -1292 8520 -120 8568
rect 120 9352 1292 9400
rect 120 9288 1208 9352
rect 1272 9288 1292 9352
rect 120 9272 1292 9288
rect 120 9208 1208 9272
rect 1272 9208 1292 9272
rect 120 9192 1292 9208
rect 120 9128 1208 9192
rect 1272 9128 1292 9192
rect 120 9112 1292 9128
rect 120 9048 1208 9112
rect 1272 9048 1292 9112
rect 120 9032 1292 9048
rect 120 8968 1208 9032
rect 1272 8968 1292 9032
rect 120 8952 1292 8968
rect 120 8888 1208 8952
rect 1272 8888 1292 8952
rect 120 8872 1292 8888
rect 120 8808 1208 8872
rect 1272 8808 1292 8872
rect 120 8792 1292 8808
rect 120 8728 1208 8792
rect 1272 8728 1292 8792
rect 120 8712 1292 8728
rect 120 8648 1208 8712
rect 1272 8648 1292 8712
rect 120 8632 1292 8648
rect 120 8568 1208 8632
rect 1272 8568 1292 8632
rect 120 8520 1292 8568
rect 1532 9352 2704 9400
rect 1532 9288 2620 9352
rect 2684 9288 2704 9352
rect 1532 9272 2704 9288
rect 1532 9208 2620 9272
rect 2684 9208 2704 9272
rect 1532 9192 2704 9208
rect 1532 9128 2620 9192
rect 2684 9128 2704 9192
rect 1532 9112 2704 9128
rect 1532 9048 2620 9112
rect 2684 9048 2704 9112
rect 1532 9032 2704 9048
rect 1532 8968 2620 9032
rect 2684 8968 2704 9032
rect 1532 8952 2704 8968
rect 1532 8888 2620 8952
rect 2684 8888 2704 8952
rect 1532 8872 2704 8888
rect 1532 8808 2620 8872
rect 2684 8808 2704 8872
rect 1532 8792 2704 8808
rect 1532 8728 2620 8792
rect 2684 8728 2704 8792
rect 1532 8712 2704 8728
rect 1532 8648 2620 8712
rect 2684 8648 2704 8712
rect 1532 8632 2704 8648
rect 1532 8568 2620 8632
rect 2684 8568 2704 8632
rect 1532 8520 2704 8568
rect 2944 9352 4116 9400
rect 2944 9288 4032 9352
rect 4096 9288 4116 9352
rect 2944 9272 4116 9288
rect 2944 9208 4032 9272
rect 4096 9208 4116 9272
rect 2944 9192 4116 9208
rect 2944 9128 4032 9192
rect 4096 9128 4116 9192
rect 2944 9112 4116 9128
rect 2944 9048 4032 9112
rect 4096 9048 4116 9112
rect 2944 9032 4116 9048
rect 2944 8968 4032 9032
rect 4096 8968 4116 9032
rect 2944 8952 4116 8968
rect 2944 8888 4032 8952
rect 4096 8888 4116 8952
rect 2944 8872 4116 8888
rect 2944 8808 4032 8872
rect 4096 8808 4116 8872
rect 2944 8792 4116 8808
rect 2944 8728 4032 8792
rect 4096 8728 4116 8792
rect 2944 8712 4116 8728
rect 2944 8648 4032 8712
rect 4096 8648 4116 8712
rect 2944 8632 4116 8648
rect 2944 8568 4032 8632
rect 4096 8568 4116 8632
rect 2944 8520 4116 8568
rect 4356 9352 5528 9400
rect 4356 9288 5444 9352
rect 5508 9288 5528 9352
rect 4356 9272 5528 9288
rect 4356 9208 5444 9272
rect 5508 9208 5528 9272
rect 4356 9192 5528 9208
rect 4356 9128 5444 9192
rect 5508 9128 5528 9192
rect 4356 9112 5528 9128
rect 4356 9048 5444 9112
rect 5508 9048 5528 9112
rect 4356 9032 5528 9048
rect 4356 8968 5444 9032
rect 5508 8968 5528 9032
rect 4356 8952 5528 8968
rect 4356 8888 5444 8952
rect 5508 8888 5528 8952
rect 4356 8872 5528 8888
rect 4356 8808 5444 8872
rect 5508 8808 5528 8872
rect 4356 8792 5528 8808
rect 4356 8728 5444 8792
rect 5508 8728 5528 8792
rect 4356 8712 5528 8728
rect 4356 8648 5444 8712
rect 5508 8648 5528 8712
rect 4356 8632 5528 8648
rect 4356 8568 5444 8632
rect 5508 8568 5528 8632
rect 4356 8520 5528 8568
rect 5768 9352 6940 9400
rect 5768 9288 6856 9352
rect 6920 9288 6940 9352
rect 5768 9272 6940 9288
rect 5768 9208 6856 9272
rect 6920 9208 6940 9272
rect 5768 9192 6940 9208
rect 5768 9128 6856 9192
rect 6920 9128 6940 9192
rect 5768 9112 6940 9128
rect 5768 9048 6856 9112
rect 6920 9048 6940 9112
rect 5768 9032 6940 9048
rect 5768 8968 6856 9032
rect 6920 8968 6940 9032
rect 5768 8952 6940 8968
rect 5768 8888 6856 8952
rect 6920 8888 6940 8952
rect 5768 8872 6940 8888
rect 5768 8808 6856 8872
rect 6920 8808 6940 8872
rect 5768 8792 6940 8808
rect 5768 8728 6856 8792
rect 6920 8728 6940 8792
rect 5768 8712 6940 8728
rect 5768 8648 6856 8712
rect 6920 8648 6940 8712
rect 5768 8632 6940 8648
rect 5768 8568 6856 8632
rect 6920 8568 6940 8632
rect 5768 8520 6940 8568
rect 7180 9352 8352 9400
rect 7180 9288 8268 9352
rect 8332 9288 8352 9352
rect 7180 9272 8352 9288
rect 7180 9208 8268 9272
rect 8332 9208 8352 9272
rect 7180 9192 8352 9208
rect 7180 9128 8268 9192
rect 8332 9128 8352 9192
rect 7180 9112 8352 9128
rect 7180 9048 8268 9112
rect 8332 9048 8352 9112
rect 7180 9032 8352 9048
rect 7180 8968 8268 9032
rect 8332 8968 8352 9032
rect 7180 8952 8352 8968
rect 7180 8888 8268 8952
rect 8332 8888 8352 8952
rect 7180 8872 8352 8888
rect 7180 8808 8268 8872
rect 8332 8808 8352 8872
rect 7180 8792 8352 8808
rect 7180 8728 8268 8792
rect 8332 8728 8352 8792
rect 7180 8712 8352 8728
rect 7180 8648 8268 8712
rect 8332 8648 8352 8712
rect 7180 8632 8352 8648
rect 7180 8568 8268 8632
rect 8332 8568 8352 8632
rect 7180 8520 8352 8568
rect 8592 9352 9764 9400
rect 8592 9288 9680 9352
rect 9744 9288 9764 9352
rect 8592 9272 9764 9288
rect 8592 9208 9680 9272
rect 9744 9208 9764 9272
rect 8592 9192 9764 9208
rect 8592 9128 9680 9192
rect 9744 9128 9764 9192
rect 8592 9112 9764 9128
rect 8592 9048 9680 9112
rect 9744 9048 9764 9112
rect 8592 9032 9764 9048
rect 8592 8968 9680 9032
rect 9744 8968 9764 9032
rect 8592 8952 9764 8968
rect 8592 8888 9680 8952
rect 9744 8888 9764 8952
rect 8592 8872 9764 8888
rect 8592 8808 9680 8872
rect 9744 8808 9764 8872
rect 8592 8792 9764 8808
rect 8592 8728 9680 8792
rect 9744 8728 9764 8792
rect 8592 8712 9764 8728
rect 8592 8648 9680 8712
rect 9744 8648 9764 8712
rect 8592 8632 9764 8648
rect 8592 8568 9680 8632
rect 9744 8568 9764 8632
rect 8592 8520 9764 8568
rect 10004 9352 11176 9400
rect 10004 9288 11092 9352
rect 11156 9288 11176 9352
rect 10004 9272 11176 9288
rect 10004 9208 11092 9272
rect 11156 9208 11176 9272
rect 10004 9192 11176 9208
rect 10004 9128 11092 9192
rect 11156 9128 11176 9192
rect 10004 9112 11176 9128
rect 10004 9048 11092 9112
rect 11156 9048 11176 9112
rect 10004 9032 11176 9048
rect 10004 8968 11092 9032
rect 11156 8968 11176 9032
rect 10004 8952 11176 8968
rect 10004 8888 11092 8952
rect 11156 8888 11176 8952
rect 10004 8872 11176 8888
rect 10004 8808 11092 8872
rect 11156 8808 11176 8872
rect 10004 8792 11176 8808
rect 10004 8728 11092 8792
rect 11156 8728 11176 8792
rect 10004 8712 11176 8728
rect 10004 8648 11092 8712
rect 11156 8648 11176 8712
rect 10004 8632 11176 8648
rect 10004 8568 11092 8632
rect 11156 8568 11176 8632
rect 10004 8520 11176 8568
rect 11416 9352 12588 9400
rect 11416 9288 12504 9352
rect 12568 9288 12588 9352
rect 11416 9272 12588 9288
rect 11416 9208 12504 9272
rect 12568 9208 12588 9272
rect 11416 9192 12588 9208
rect 11416 9128 12504 9192
rect 12568 9128 12588 9192
rect 11416 9112 12588 9128
rect 11416 9048 12504 9112
rect 12568 9048 12588 9112
rect 11416 9032 12588 9048
rect 11416 8968 12504 9032
rect 12568 8968 12588 9032
rect 11416 8952 12588 8968
rect 11416 8888 12504 8952
rect 12568 8888 12588 8952
rect 11416 8872 12588 8888
rect 11416 8808 12504 8872
rect 12568 8808 12588 8872
rect 11416 8792 12588 8808
rect 11416 8728 12504 8792
rect 12568 8728 12588 8792
rect 11416 8712 12588 8728
rect 11416 8648 12504 8712
rect 12568 8648 12588 8712
rect 11416 8632 12588 8648
rect 11416 8568 12504 8632
rect 12568 8568 12588 8632
rect 11416 8520 12588 8568
rect 12828 9352 14000 9400
rect 12828 9288 13916 9352
rect 13980 9288 14000 9352
rect 12828 9272 14000 9288
rect 12828 9208 13916 9272
rect 13980 9208 14000 9272
rect 12828 9192 14000 9208
rect 12828 9128 13916 9192
rect 13980 9128 14000 9192
rect 12828 9112 14000 9128
rect 12828 9048 13916 9112
rect 13980 9048 14000 9112
rect 12828 9032 14000 9048
rect 12828 8968 13916 9032
rect 13980 8968 14000 9032
rect 12828 8952 14000 8968
rect 12828 8888 13916 8952
rect 13980 8888 14000 8952
rect 12828 8872 14000 8888
rect 12828 8808 13916 8872
rect 13980 8808 14000 8872
rect 12828 8792 14000 8808
rect 12828 8728 13916 8792
rect 13980 8728 14000 8792
rect 12828 8712 14000 8728
rect 12828 8648 13916 8712
rect 13980 8648 14000 8712
rect 12828 8632 14000 8648
rect 12828 8568 13916 8632
rect 13980 8568 14000 8632
rect 12828 8520 14000 8568
rect 14240 9352 15412 9400
rect 14240 9288 15328 9352
rect 15392 9288 15412 9352
rect 14240 9272 15412 9288
rect 14240 9208 15328 9272
rect 15392 9208 15412 9272
rect 14240 9192 15412 9208
rect 14240 9128 15328 9192
rect 15392 9128 15412 9192
rect 14240 9112 15412 9128
rect 14240 9048 15328 9112
rect 15392 9048 15412 9112
rect 14240 9032 15412 9048
rect 14240 8968 15328 9032
rect 15392 8968 15412 9032
rect 14240 8952 15412 8968
rect 14240 8888 15328 8952
rect 15392 8888 15412 8952
rect 14240 8872 15412 8888
rect 14240 8808 15328 8872
rect 15392 8808 15412 8872
rect 14240 8792 15412 8808
rect 14240 8728 15328 8792
rect 15392 8728 15412 8792
rect 14240 8712 15412 8728
rect 14240 8648 15328 8712
rect 15392 8648 15412 8712
rect 14240 8632 15412 8648
rect 14240 8568 15328 8632
rect 15392 8568 15412 8632
rect 14240 8520 15412 8568
rect 15652 9352 16824 9400
rect 15652 9288 16740 9352
rect 16804 9288 16824 9352
rect 15652 9272 16824 9288
rect 15652 9208 16740 9272
rect 16804 9208 16824 9272
rect 15652 9192 16824 9208
rect 15652 9128 16740 9192
rect 16804 9128 16824 9192
rect 15652 9112 16824 9128
rect 15652 9048 16740 9112
rect 16804 9048 16824 9112
rect 15652 9032 16824 9048
rect 15652 8968 16740 9032
rect 16804 8968 16824 9032
rect 15652 8952 16824 8968
rect 15652 8888 16740 8952
rect 16804 8888 16824 8952
rect 15652 8872 16824 8888
rect 15652 8808 16740 8872
rect 16804 8808 16824 8872
rect 15652 8792 16824 8808
rect 15652 8728 16740 8792
rect 16804 8728 16824 8792
rect 15652 8712 16824 8728
rect 15652 8648 16740 8712
rect 16804 8648 16824 8712
rect 15652 8632 16824 8648
rect 15652 8568 16740 8632
rect 16804 8568 16824 8632
rect 15652 8520 16824 8568
rect 17064 9352 18236 9400
rect 17064 9288 18152 9352
rect 18216 9288 18236 9352
rect 17064 9272 18236 9288
rect 17064 9208 18152 9272
rect 18216 9208 18236 9272
rect 17064 9192 18236 9208
rect 17064 9128 18152 9192
rect 18216 9128 18236 9192
rect 17064 9112 18236 9128
rect 17064 9048 18152 9112
rect 18216 9048 18236 9112
rect 17064 9032 18236 9048
rect 17064 8968 18152 9032
rect 18216 8968 18236 9032
rect 17064 8952 18236 8968
rect 17064 8888 18152 8952
rect 18216 8888 18236 8952
rect 17064 8872 18236 8888
rect 17064 8808 18152 8872
rect 18216 8808 18236 8872
rect 17064 8792 18236 8808
rect 17064 8728 18152 8792
rect 18216 8728 18236 8792
rect 17064 8712 18236 8728
rect 17064 8648 18152 8712
rect 18216 8648 18236 8712
rect 17064 8632 18236 8648
rect 17064 8568 18152 8632
rect 18216 8568 18236 8632
rect 17064 8520 18236 8568
rect 18476 9352 19648 9400
rect 18476 9288 19564 9352
rect 19628 9288 19648 9352
rect 18476 9272 19648 9288
rect 18476 9208 19564 9272
rect 19628 9208 19648 9272
rect 18476 9192 19648 9208
rect 18476 9128 19564 9192
rect 19628 9128 19648 9192
rect 18476 9112 19648 9128
rect 18476 9048 19564 9112
rect 19628 9048 19648 9112
rect 18476 9032 19648 9048
rect 18476 8968 19564 9032
rect 19628 8968 19648 9032
rect 18476 8952 19648 8968
rect 18476 8888 19564 8952
rect 19628 8888 19648 8952
rect 18476 8872 19648 8888
rect 18476 8808 19564 8872
rect 19628 8808 19648 8872
rect 18476 8792 19648 8808
rect 18476 8728 19564 8792
rect 19628 8728 19648 8792
rect 18476 8712 19648 8728
rect 18476 8648 19564 8712
rect 19628 8648 19648 8712
rect 18476 8632 19648 8648
rect 18476 8568 19564 8632
rect 19628 8568 19648 8632
rect 18476 8520 19648 8568
rect 19888 9352 21060 9400
rect 19888 9288 20976 9352
rect 21040 9288 21060 9352
rect 19888 9272 21060 9288
rect 19888 9208 20976 9272
rect 21040 9208 21060 9272
rect 19888 9192 21060 9208
rect 19888 9128 20976 9192
rect 21040 9128 21060 9192
rect 19888 9112 21060 9128
rect 19888 9048 20976 9112
rect 21040 9048 21060 9112
rect 19888 9032 21060 9048
rect 19888 8968 20976 9032
rect 21040 8968 21060 9032
rect 19888 8952 21060 8968
rect 19888 8888 20976 8952
rect 21040 8888 21060 8952
rect 19888 8872 21060 8888
rect 19888 8808 20976 8872
rect 21040 8808 21060 8872
rect 19888 8792 21060 8808
rect 19888 8728 20976 8792
rect 21040 8728 21060 8792
rect 19888 8712 21060 8728
rect 19888 8648 20976 8712
rect 21040 8648 21060 8712
rect 19888 8632 21060 8648
rect 19888 8568 20976 8632
rect 21040 8568 21060 8632
rect 19888 8520 21060 8568
rect 21300 9352 22472 9400
rect 21300 9288 22388 9352
rect 22452 9288 22472 9352
rect 21300 9272 22472 9288
rect 21300 9208 22388 9272
rect 22452 9208 22472 9272
rect 21300 9192 22472 9208
rect 21300 9128 22388 9192
rect 22452 9128 22472 9192
rect 21300 9112 22472 9128
rect 21300 9048 22388 9112
rect 22452 9048 22472 9112
rect 21300 9032 22472 9048
rect 21300 8968 22388 9032
rect 22452 8968 22472 9032
rect 21300 8952 22472 8968
rect 21300 8888 22388 8952
rect 22452 8888 22472 8952
rect 21300 8872 22472 8888
rect 21300 8808 22388 8872
rect 22452 8808 22472 8872
rect 21300 8792 22472 8808
rect 21300 8728 22388 8792
rect 22452 8728 22472 8792
rect 21300 8712 22472 8728
rect 21300 8648 22388 8712
rect 22452 8648 22472 8712
rect 21300 8632 22472 8648
rect 21300 8568 22388 8632
rect 22452 8568 22472 8632
rect 21300 8520 22472 8568
rect 22712 9352 23884 9400
rect 22712 9288 23800 9352
rect 23864 9288 23884 9352
rect 22712 9272 23884 9288
rect 22712 9208 23800 9272
rect 23864 9208 23884 9272
rect 22712 9192 23884 9208
rect 22712 9128 23800 9192
rect 23864 9128 23884 9192
rect 22712 9112 23884 9128
rect 22712 9048 23800 9112
rect 23864 9048 23884 9112
rect 22712 9032 23884 9048
rect 22712 8968 23800 9032
rect 23864 8968 23884 9032
rect 22712 8952 23884 8968
rect 22712 8888 23800 8952
rect 23864 8888 23884 8952
rect 22712 8872 23884 8888
rect 22712 8808 23800 8872
rect 23864 8808 23884 8872
rect 22712 8792 23884 8808
rect 22712 8728 23800 8792
rect 23864 8728 23884 8792
rect 22712 8712 23884 8728
rect 22712 8648 23800 8712
rect 23864 8648 23884 8712
rect 22712 8632 23884 8648
rect 22712 8568 23800 8632
rect 23864 8568 23884 8632
rect 22712 8520 23884 8568
rect -23884 8232 -22712 8280
rect -23884 8168 -22796 8232
rect -22732 8168 -22712 8232
rect -23884 8152 -22712 8168
rect -23884 8088 -22796 8152
rect -22732 8088 -22712 8152
rect -23884 8072 -22712 8088
rect -23884 8008 -22796 8072
rect -22732 8008 -22712 8072
rect -23884 7992 -22712 8008
rect -23884 7928 -22796 7992
rect -22732 7928 -22712 7992
rect -23884 7912 -22712 7928
rect -23884 7848 -22796 7912
rect -22732 7848 -22712 7912
rect -23884 7832 -22712 7848
rect -23884 7768 -22796 7832
rect -22732 7768 -22712 7832
rect -23884 7752 -22712 7768
rect -23884 7688 -22796 7752
rect -22732 7688 -22712 7752
rect -23884 7672 -22712 7688
rect -23884 7608 -22796 7672
rect -22732 7608 -22712 7672
rect -23884 7592 -22712 7608
rect -23884 7528 -22796 7592
rect -22732 7528 -22712 7592
rect -23884 7512 -22712 7528
rect -23884 7448 -22796 7512
rect -22732 7448 -22712 7512
rect -23884 7400 -22712 7448
rect -22472 8232 -21300 8280
rect -22472 8168 -21384 8232
rect -21320 8168 -21300 8232
rect -22472 8152 -21300 8168
rect -22472 8088 -21384 8152
rect -21320 8088 -21300 8152
rect -22472 8072 -21300 8088
rect -22472 8008 -21384 8072
rect -21320 8008 -21300 8072
rect -22472 7992 -21300 8008
rect -22472 7928 -21384 7992
rect -21320 7928 -21300 7992
rect -22472 7912 -21300 7928
rect -22472 7848 -21384 7912
rect -21320 7848 -21300 7912
rect -22472 7832 -21300 7848
rect -22472 7768 -21384 7832
rect -21320 7768 -21300 7832
rect -22472 7752 -21300 7768
rect -22472 7688 -21384 7752
rect -21320 7688 -21300 7752
rect -22472 7672 -21300 7688
rect -22472 7608 -21384 7672
rect -21320 7608 -21300 7672
rect -22472 7592 -21300 7608
rect -22472 7528 -21384 7592
rect -21320 7528 -21300 7592
rect -22472 7512 -21300 7528
rect -22472 7448 -21384 7512
rect -21320 7448 -21300 7512
rect -22472 7400 -21300 7448
rect -21060 8232 -19888 8280
rect -21060 8168 -19972 8232
rect -19908 8168 -19888 8232
rect -21060 8152 -19888 8168
rect -21060 8088 -19972 8152
rect -19908 8088 -19888 8152
rect -21060 8072 -19888 8088
rect -21060 8008 -19972 8072
rect -19908 8008 -19888 8072
rect -21060 7992 -19888 8008
rect -21060 7928 -19972 7992
rect -19908 7928 -19888 7992
rect -21060 7912 -19888 7928
rect -21060 7848 -19972 7912
rect -19908 7848 -19888 7912
rect -21060 7832 -19888 7848
rect -21060 7768 -19972 7832
rect -19908 7768 -19888 7832
rect -21060 7752 -19888 7768
rect -21060 7688 -19972 7752
rect -19908 7688 -19888 7752
rect -21060 7672 -19888 7688
rect -21060 7608 -19972 7672
rect -19908 7608 -19888 7672
rect -21060 7592 -19888 7608
rect -21060 7528 -19972 7592
rect -19908 7528 -19888 7592
rect -21060 7512 -19888 7528
rect -21060 7448 -19972 7512
rect -19908 7448 -19888 7512
rect -21060 7400 -19888 7448
rect -19648 8232 -18476 8280
rect -19648 8168 -18560 8232
rect -18496 8168 -18476 8232
rect -19648 8152 -18476 8168
rect -19648 8088 -18560 8152
rect -18496 8088 -18476 8152
rect -19648 8072 -18476 8088
rect -19648 8008 -18560 8072
rect -18496 8008 -18476 8072
rect -19648 7992 -18476 8008
rect -19648 7928 -18560 7992
rect -18496 7928 -18476 7992
rect -19648 7912 -18476 7928
rect -19648 7848 -18560 7912
rect -18496 7848 -18476 7912
rect -19648 7832 -18476 7848
rect -19648 7768 -18560 7832
rect -18496 7768 -18476 7832
rect -19648 7752 -18476 7768
rect -19648 7688 -18560 7752
rect -18496 7688 -18476 7752
rect -19648 7672 -18476 7688
rect -19648 7608 -18560 7672
rect -18496 7608 -18476 7672
rect -19648 7592 -18476 7608
rect -19648 7528 -18560 7592
rect -18496 7528 -18476 7592
rect -19648 7512 -18476 7528
rect -19648 7448 -18560 7512
rect -18496 7448 -18476 7512
rect -19648 7400 -18476 7448
rect -18236 8232 -17064 8280
rect -18236 8168 -17148 8232
rect -17084 8168 -17064 8232
rect -18236 8152 -17064 8168
rect -18236 8088 -17148 8152
rect -17084 8088 -17064 8152
rect -18236 8072 -17064 8088
rect -18236 8008 -17148 8072
rect -17084 8008 -17064 8072
rect -18236 7992 -17064 8008
rect -18236 7928 -17148 7992
rect -17084 7928 -17064 7992
rect -18236 7912 -17064 7928
rect -18236 7848 -17148 7912
rect -17084 7848 -17064 7912
rect -18236 7832 -17064 7848
rect -18236 7768 -17148 7832
rect -17084 7768 -17064 7832
rect -18236 7752 -17064 7768
rect -18236 7688 -17148 7752
rect -17084 7688 -17064 7752
rect -18236 7672 -17064 7688
rect -18236 7608 -17148 7672
rect -17084 7608 -17064 7672
rect -18236 7592 -17064 7608
rect -18236 7528 -17148 7592
rect -17084 7528 -17064 7592
rect -18236 7512 -17064 7528
rect -18236 7448 -17148 7512
rect -17084 7448 -17064 7512
rect -18236 7400 -17064 7448
rect -16824 8232 -15652 8280
rect -16824 8168 -15736 8232
rect -15672 8168 -15652 8232
rect -16824 8152 -15652 8168
rect -16824 8088 -15736 8152
rect -15672 8088 -15652 8152
rect -16824 8072 -15652 8088
rect -16824 8008 -15736 8072
rect -15672 8008 -15652 8072
rect -16824 7992 -15652 8008
rect -16824 7928 -15736 7992
rect -15672 7928 -15652 7992
rect -16824 7912 -15652 7928
rect -16824 7848 -15736 7912
rect -15672 7848 -15652 7912
rect -16824 7832 -15652 7848
rect -16824 7768 -15736 7832
rect -15672 7768 -15652 7832
rect -16824 7752 -15652 7768
rect -16824 7688 -15736 7752
rect -15672 7688 -15652 7752
rect -16824 7672 -15652 7688
rect -16824 7608 -15736 7672
rect -15672 7608 -15652 7672
rect -16824 7592 -15652 7608
rect -16824 7528 -15736 7592
rect -15672 7528 -15652 7592
rect -16824 7512 -15652 7528
rect -16824 7448 -15736 7512
rect -15672 7448 -15652 7512
rect -16824 7400 -15652 7448
rect -15412 8232 -14240 8280
rect -15412 8168 -14324 8232
rect -14260 8168 -14240 8232
rect -15412 8152 -14240 8168
rect -15412 8088 -14324 8152
rect -14260 8088 -14240 8152
rect -15412 8072 -14240 8088
rect -15412 8008 -14324 8072
rect -14260 8008 -14240 8072
rect -15412 7992 -14240 8008
rect -15412 7928 -14324 7992
rect -14260 7928 -14240 7992
rect -15412 7912 -14240 7928
rect -15412 7848 -14324 7912
rect -14260 7848 -14240 7912
rect -15412 7832 -14240 7848
rect -15412 7768 -14324 7832
rect -14260 7768 -14240 7832
rect -15412 7752 -14240 7768
rect -15412 7688 -14324 7752
rect -14260 7688 -14240 7752
rect -15412 7672 -14240 7688
rect -15412 7608 -14324 7672
rect -14260 7608 -14240 7672
rect -15412 7592 -14240 7608
rect -15412 7528 -14324 7592
rect -14260 7528 -14240 7592
rect -15412 7512 -14240 7528
rect -15412 7448 -14324 7512
rect -14260 7448 -14240 7512
rect -15412 7400 -14240 7448
rect -14000 8232 -12828 8280
rect -14000 8168 -12912 8232
rect -12848 8168 -12828 8232
rect -14000 8152 -12828 8168
rect -14000 8088 -12912 8152
rect -12848 8088 -12828 8152
rect -14000 8072 -12828 8088
rect -14000 8008 -12912 8072
rect -12848 8008 -12828 8072
rect -14000 7992 -12828 8008
rect -14000 7928 -12912 7992
rect -12848 7928 -12828 7992
rect -14000 7912 -12828 7928
rect -14000 7848 -12912 7912
rect -12848 7848 -12828 7912
rect -14000 7832 -12828 7848
rect -14000 7768 -12912 7832
rect -12848 7768 -12828 7832
rect -14000 7752 -12828 7768
rect -14000 7688 -12912 7752
rect -12848 7688 -12828 7752
rect -14000 7672 -12828 7688
rect -14000 7608 -12912 7672
rect -12848 7608 -12828 7672
rect -14000 7592 -12828 7608
rect -14000 7528 -12912 7592
rect -12848 7528 -12828 7592
rect -14000 7512 -12828 7528
rect -14000 7448 -12912 7512
rect -12848 7448 -12828 7512
rect -14000 7400 -12828 7448
rect -12588 8232 -11416 8280
rect -12588 8168 -11500 8232
rect -11436 8168 -11416 8232
rect -12588 8152 -11416 8168
rect -12588 8088 -11500 8152
rect -11436 8088 -11416 8152
rect -12588 8072 -11416 8088
rect -12588 8008 -11500 8072
rect -11436 8008 -11416 8072
rect -12588 7992 -11416 8008
rect -12588 7928 -11500 7992
rect -11436 7928 -11416 7992
rect -12588 7912 -11416 7928
rect -12588 7848 -11500 7912
rect -11436 7848 -11416 7912
rect -12588 7832 -11416 7848
rect -12588 7768 -11500 7832
rect -11436 7768 -11416 7832
rect -12588 7752 -11416 7768
rect -12588 7688 -11500 7752
rect -11436 7688 -11416 7752
rect -12588 7672 -11416 7688
rect -12588 7608 -11500 7672
rect -11436 7608 -11416 7672
rect -12588 7592 -11416 7608
rect -12588 7528 -11500 7592
rect -11436 7528 -11416 7592
rect -12588 7512 -11416 7528
rect -12588 7448 -11500 7512
rect -11436 7448 -11416 7512
rect -12588 7400 -11416 7448
rect -11176 8232 -10004 8280
rect -11176 8168 -10088 8232
rect -10024 8168 -10004 8232
rect -11176 8152 -10004 8168
rect -11176 8088 -10088 8152
rect -10024 8088 -10004 8152
rect -11176 8072 -10004 8088
rect -11176 8008 -10088 8072
rect -10024 8008 -10004 8072
rect -11176 7992 -10004 8008
rect -11176 7928 -10088 7992
rect -10024 7928 -10004 7992
rect -11176 7912 -10004 7928
rect -11176 7848 -10088 7912
rect -10024 7848 -10004 7912
rect -11176 7832 -10004 7848
rect -11176 7768 -10088 7832
rect -10024 7768 -10004 7832
rect -11176 7752 -10004 7768
rect -11176 7688 -10088 7752
rect -10024 7688 -10004 7752
rect -11176 7672 -10004 7688
rect -11176 7608 -10088 7672
rect -10024 7608 -10004 7672
rect -11176 7592 -10004 7608
rect -11176 7528 -10088 7592
rect -10024 7528 -10004 7592
rect -11176 7512 -10004 7528
rect -11176 7448 -10088 7512
rect -10024 7448 -10004 7512
rect -11176 7400 -10004 7448
rect -9764 8232 -8592 8280
rect -9764 8168 -8676 8232
rect -8612 8168 -8592 8232
rect -9764 8152 -8592 8168
rect -9764 8088 -8676 8152
rect -8612 8088 -8592 8152
rect -9764 8072 -8592 8088
rect -9764 8008 -8676 8072
rect -8612 8008 -8592 8072
rect -9764 7992 -8592 8008
rect -9764 7928 -8676 7992
rect -8612 7928 -8592 7992
rect -9764 7912 -8592 7928
rect -9764 7848 -8676 7912
rect -8612 7848 -8592 7912
rect -9764 7832 -8592 7848
rect -9764 7768 -8676 7832
rect -8612 7768 -8592 7832
rect -9764 7752 -8592 7768
rect -9764 7688 -8676 7752
rect -8612 7688 -8592 7752
rect -9764 7672 -8592 7688
rect -9764 7608 -8676 7672
rect -8612 7608 -8592 7672
rect -9764 7592 -8592 7608
rect -9764 7528 -8676 7592
rect -8612 7528 -8592 7592
rect -9764 7512 -8592 7528
rect -9764 7448 -8676 7512
rect -8612 7448 -8592 7512
rect -9764 7400 -8592 7448
rect -8352 8232 -7180 8280
rect -8352 8168 -7264 8232
rect -7200 8168 -7180 8232
rect -8352 8152 -7180 8168
rect -8352 8088 -7264 8152
rect -7200 8088 -7180 8152
rect -8352 8072 -7180 8088
rect -8352 8008 -7264 8072
rect -7200 8008 -7180 8072
rect -8352 7992 -7180 8008
rect -8352 7928 -7264 7992
rect -7200 7928 -7180 7992
rect -8352 7912 -7180 7928
rect -8352 7848 -7264 7912
rect -7200 7848 -7180 7912
rect -8352 7832 -7180 7848
rect -8352 7768 -7264 7832
rect -7200 7768 -7180 7832
rect -8352 7752 -7180 7768
rect -8352 7688 -7264 7752
rect -7200 7688 -7180 7752
rect -8352 7672 -7180 7688
rect -8352 7608 -7264 7672
rect -7200 7608 -7180 7672
rect -8352 7592 -7180 7608
rect -8352 7528 -7264 7592
rect -7200 7528 -7180 7592
rect -8352 7512 -7180 7528
rect -8352 7448 -7264 7512
rect -7200 7448 -7180 7512
rect -8352 7400 -7180 7448
rect -6940 8232 -5768 8280
rect -6940 8168 -5852 8232
rect -5788 8168 -5768 8232
rect -6940 8152 -5768 8168
rect -6940 8088 -5852 8152
rect -5788 8088 -5768 8152
rect -6940 8072 -5768 8088
rect -6940 8008 -5852 8072
rect -5788 8008 -5768 8072
rect -6940 7992 -5768 8008
rect -6940 7928 -5852 7992
rect -5788 7928 -5768 7992
rect -6940 7912 -5768 7928
rect -6940 7848 -5852 7912
rect -5788 7848 -5768 7912
rect -6940 7832 -5768 7848
rect -6940 7768 -5852 7832
rect -5788 7768 -5768 7832
rect -6940 7752 -5768 7768
rect -6940 7688 -5852 7752
rect -5788 7688 -5768 7752
rect -6940 7672 -5768 7688
rect -6940 7608 -5852 7672
rect -5788 7608 -5768 7672
rect -6940 7592 -5768 7608
rect -6940 7528 -5852 7592
rect -5788 7528 -5768 7592
rect -6940 7512 -5768 7528
rect -6940 7448 -5852 7512
rect -5788 7448 -5768 7512
rect -6940 7400 -5768 7448
rect -5528 8232 -4356 8280
rect -5528 8168 -4440 8232
rect -4376 8168 -4356 8232
rect -5528 8152 -4356 8168
rect -5528 8088 -4440 8152
rect -4376 8088 -4356 8152
rect -5528 8072 -4356 8088
rect -5528 8008 -4440 8072
rect -4376 8008 -4356 8072
rect -5528 7992 -4356 8008
rect -5528 7928 -4440 7992
rect -4376 7928 -4356 7992
rect -5528 7912 -4356 7928
rect -5528 7848 -4440 7912
rect -4376 7848 -4356 7912
rect -5528 7832 -4356 7848
rect -5528 7768 -4440 7832
rect -4376 7768 -4356 7832
rect -5528 7752 -4356 7768
rect -5528 7688 -4440 7752
rect -4376 7688 -4356 7752
rect -5528 7672 -4356 7688
rect -5528 7608 -4440 7672
rect -4376 7608 -4356 7672
rect -5528 7592 -4356 7608
rect -5528 7528 -4440 7592
rect -4376 7528 -4356 7592
rect -5528 7512 -4356 7528
rect -5528 7448 -4440 7512
rect -4376 7448 -4356 7512
rect -5528 7400 -4356 7448
rect -4116 8232 -2944 8280
rect -4116 8168 -3028 8232
rect -2964 8168 -2944 8232
rect -4116 8152 -2944 8168
rect -4116 8088 -3028 8152
rect -2964 8088 -2944 8152
rect -4116 8072 -2944 8088
rect -4116 8008 -3028 8072
rect -2964 8008 -2944 8072
rect -4116 7992 -2944 8008
rect -4116 7928 -3028 7992
rect -2964 7928 -2944 7992
rect -4116 7912 -2944 7928
rect -4116 7848 -3028 7912
rect -2964 7848 -2944 7912
rect -4116 7832 -2944 7848
rect -4116 7768 -3028 7832
rect -2964 7768 -2944 7832
rect -4116 7752 -2944 7768
rect -4116 7688 -3028 7752
rect -2964 7688 -2944 7752
rect -4116 7672 -2944 7688
rect -4116 7608 -3028 7672
rect -2964 7608 -2944 7672
rect -4116 7592 -2944 7608
rect -4116 7528 -3028 7592
rect -2964 7528 -2944 7592
rect -4116 7512 -2944 7528
rect -4116 7448 -3028 7512
rect -2964 7448 -2944 7512
rect -4116 7400 -2944 7448
rect -2704 8232 -1532 8280
rect -2704 8168 -1616 8232
rect -1552 8168 -1532 8232
rect -2704 8152 -1532 8168
rect -2704 8088 -1616 8152
rect -1552 8088 -1532 8152
rect -2704 8072 -1532 8088
rect -2704 8008 -1616 8072
rect -1552 8008 -1532 8072
rect -2704 7992 -1532 8008
rect -2704 7928 -1616 7992
rect -1552 7928 -1532 7992
rect -2704 7912 -1532 7928
rect -2704 7848 -1616 7912
rect -1552 7848 -1532 7912
rect -2704 7832 -1532 7848
rect -2704 7768 -1616 7832
rect -1552 7768 -1532 7832
rect -2704 7752 -1532 7768
rect -2704 7688 -1616 7752
rect -1552 7688 -1532 7752
rect -2704 7672 -1532 7688
rect -2704 7608 -1616 7672
rect -1552 7608 -1532 7672
rect -2704 7592 -1532 7608
rect -2704 7528 -1616 7592
rect -1552 7528 -1532 7592
rect -2704 7512 -1532 7528
rect -2704 7448 -1616 7512
rect -1552 7448 -1532 7512
rect -2704 7400 -1532 7448
rect -1292 8232 -120 8280
rect -1292 8168 -204 8232
rect -140 8168 -120 8232
rect -1292 8152 -120 8168
rect -1292 8088 -204 8152
rect -140 8088 -120 8152
rect -1292 8072 -120 8088
rect -1292 8008 -204 8072
rect -140 8008 -120 8072
rect -1292 7992 -120 8008
rect -1292 7928 -204 7992
rect -140 7928 -120 7992
rect -1292 7912 -120 7928
rect -1292 7848 -204 7912
rect -140 7848 -120 7912
rect -1292 7832 -120 7848
rect -1292 7768 -204 7832
rect -140 7768 -120 7832
rect -1292 7752 -120 7768
rect -1292 7688 -204 7752
rect -140 7688 -120 7752
rect -1292 7672 -120 7688
rect -1292 7608 -204 7672
rect -140 7608 -120 7672
rect -1292 7592 -120 7608
rect -1292 7528 -204 7592
rect -140 7528 -120 7592
rect -1292 7512 -120 7528
rect -1292 7448 -204 7512
rect -140 7448 -120 7512
rect -1292 7400 -120 7448
rect 120 8232 1292 8280
rect 120 8168 1208 8232
rect 1272 8168 1292 8232
rect 120 8152 1292 8168
rect 120 8088 1208 8152
rect 1272 8088 1292 8152
rect 120 8072 1292 8088
rect 120 8008 1208 8072
rect 1272 8008 1292 8072
rect 120 7992 1292 8008
rect 120 7928 1208 7992
rect 1272 7928 1292 7992
rect 120 7912 1292 7928
rect 120 7848 1208 7912
rect 1272 7848 1292 7912
rect 120 7832 1292 7848
rect 120 7768 1208 7832
rect 1272 7768 1292 7832
rect 120 7752 1292 7768
rect 120 7688 1208 7752
rect 1272 7688 1292 7752
rect 120 7672 1292 7688
rect 120 7608 1208 7672
rect 1272 7608 1292 7672
rect 120 7592 1292 7608
rect 120 7528 1208 7592
rect 1272 7528 1292 7592
rect 120 7512 1292 7528
rect 120 7448 1208 7512
rect 1272 7448 1292 7512
rect 120 7400 1292 7448
rect 1532 8232 2704 8280
rect 1532 8168 2620 8232
rect 2684 8168 2704 8232
rect 1532 8152 2704 8168
rect 1532 8088 2620 8152
rect 2684 8088 2704 8152
rect 1532 8072 2704 8088
rect 1532 8008 2620 8072
rect 2684 8008 2704 8072
rect 1532 7992 2704 8008
rect 1532 7928 2620 7992
rect 2684 7928 2704 7992
rect 1532 7912 2704 7928
rect 1532 7848 2620 7912
rect 2684 7848 2704 7912
rect 1532 7832 2704 7848
rect 1532 7768 2620 7832
rect 2684 7768 2704 7832
rect 1532 7752 2704 7768
rect 1532 7688 2620 7752
rect 2684 7688 2704 7752
rect 1532 7672 2704 7688
rect 1532 7608 2620 7672
rect 2684 7608 2704 7672
rect 1532 7592 2704 7608
rect 1532 7528 2620 7592
rect 2684 7528 2704 7592
rect 1532 7512 2704 7528
rect 1532 7448 2620 7512
rect 2684 7448 2704 7512
rect 1532 7400 2704 7448
rect 2944 8232 4116 8280
rect 2944 8168 4032 8232
rect 4096 8168 4116 8232
rect 2944 8152 4116 8168
rect 2944 8088 4032 8152
rect 4096 8088 4116 8152
rect 2944 8072 4116 8088
rect 2944 8008 4032 8072
rect 4096 8008 4116 8072
rect 2944 7992 4116 8008
rect 2944 7928 4032 7992
rect 4096 7928 4116 7992
rect 2944 7912 4116 7928
rect 2944 7848 4032 7912
rect 4096 7848 4116 7912
rect 2944 7832 4116 7848
rect 2944 7768 4032 7832
rect 4096 7768 4116 7832
rect 2944 7752 4116 7768
rect 2944 7688 4032 7752
rect 4096 7688 4116 7752
rect 2944 7672 4116 7688
rect 2944 7608 4032 7672
rect 4096 7608 4116 7672
rect 2944 7592 4116 7608
rect 2944 7528 4032 7592
rect 4096 7528 4116 7592
rect 2944 7512 4116 7528
rect 2944 7448 4032 7512
rect 4096 7448 4116 7512
rect 2944 7400 4116 7448
rect 4356 8232 5528 8280
rect 4356 8168 5444 8232
rect 5508 8168 5528 8232
rect 4356 8152 5528 8168
rect 4356 8088 5444 8152
rect 5508 8088 5528 8152
rect 4356 8072 5528 8088
rect 4356 8008 5444 8072
rect 5508 8008 5528 8072
rect 4356 7992 5528 8008
rect 4356 7928 5444 7992
rect 5508 7928 5528 7992
rect 4356 7912 5528 7928
rect 4356 7848 5444 7912
rect 5508 7848 5528 7912
rect 4356 7832 5528 7848
rect 4356 7768 5444 7832
rect 5508 7768 5528 7832
rect 4356 7752 5528 7768
rect 4356 7688 5444 7752
rect 5508 7688 5528 7752
rect 4356 7672 5528 7688
rect 4356 7608 5444 7672
rect 5508 7608 5528 7672
rect 4356 7592 5528 7608
rect 4356 7528 5444 7592
rect 5508 7528 5528 7592
rect 4356 7512 5528 7528
rect 4356 7448 5444 7512
rect 5508 7448 5528 7512
rect 4356 7400 5528 7448
rect 5768 8232 6940 8280
rect 5768 8168 6856 8232
rect 6920 8168 6940 8232
rect 5768 8152 6940 8168
rect 5768 8088 6856 8152
rect 6920 8088 6940 8152
rect 5768 8072 6940 8088
rect 5768 8008 6856 8072
rect 6920 8008 6940 8072
rect 5768 7992 6940 8008
rect 5768 7928 6856 7992
rect 6920 7928 6940 7992
rect 5768 7912 6940 7928
rect 5768 7848 6856 7912
rect 6920 7848 6940 7912
rect 5768 7832 6940 7848
rect 5768 7768 6856 7832
rect 6920 7768 6940 7832
rect 5768 7752 6940 7768
rect 5768 7688 6856 7752
rect 6920 7688 6940 7752
rect 5768 7672 6940 7688
rect 5768 7608 6856 7672
rect 6920 7608 6940 7672
rect 5768 7592 6940 7608
rect 5768 7528 6856 7592
rect 6920 7528 6940 7592
rect 5768 7512 6940 7528
rect 5768 7448 6856 7512
rect 6920 7448 6940 7512
rect 5768 7400 6940 7448
rect 7180 8232 8352 8280
rect 7180 8168 8268 8232
rect 8332 8168 8352 8232
rect 7180 8152 8352 8168
rect 7180 8088 8268 8152
rect 8332 8088 8352 8152
rect 7180 8072 8352 8088
rect 7180 8008 8268 8072
rect 8332 8008 8352 8072
rect 7180 7992 8352 8008
rect 7180 7928 8268 7992
rect 8332 7928 8352 7992
rect 7180 7912 8352 7928
rect 7180 7848 8268 7912
rect 8332 7848 8352 7912
rect 7180 7832 8352 7848
rect 7180 7768 8268 7832
rect 8332 7768 8352 7832
rect 7180 7752 8352 7768
rect 7180 7688 8268 7752
rect 8332 7688 8352 7752
rect 7180 7672 8352 7688
rect 7180 7608 8268 7672
rect 8332 7608 8352 7672
rect 7180 7592 8352 7608
rect 7180 7528 8268 7592
rect 8332 7528 8352 7592
rect 7180 7512 8352 7528
rect 7180 7448 8268 7512
rect 8332 7448 8352 7512
rect 7180 7400 8352 7448
rect 8592 8232 9764 8280
rect 8592 8168 9680 8232
rect 9744 8168 9764 8232
rect 8592 8152 9764 8168
rect 8592 8088 9680 8152
rect 9744 8088 9764 8152
rect 8592 8072 9764 8088
rect 8592 8008 9680 8072
rect 9744 8008 9764 8072
rect 8592 7992 9764 8008
rect 8592 7928 9680 7992
rect 9744 7928 9764 7992
rect 8592 7912 9764 7928
rect 8592 7848 9680 7912
rect 9744 7848 9764 7912
rect 8592 7832 9764 7848
rect 8592 7768 9680 7832
rect 9744 7768 9764 7832
rect 8592 7752 9764 7768
rect 8592 7688 9680 7752
rect 9744 7688 9764 7752
rect 8592 7672 9764 7688
rect 8592 7608 9680 7672
rect 9744 7608 9764 7672
rect 8592 7592 9764 7608
rect 8592 7528 9680 7592
rect 9744 7528 9764 7592
rect 8592 7512 9764 7528
rect 8592 7448 9680 7512
rect 9744 7448 9764 7512
rect 8592 7400 9764 7448
rect 10004 8232 11176 8280
rect 10004 8168 11092 8232
rect 11156 8168 11176 8232
rect 10004 8152 11176 8168
rect 10004 8088 11092 8152
rect 11156 8088 11176 8152
rect 10004 8072 11176 8088
rect 10004 8008 11092 8072
rect 11156 8008 11176 8072
rect 10004 7992 11176 8008
rect 10004 7928 11092 7992
rect 11156 7928 11176 7992
rect 10004 7912 11176 7928
rect 10004 7848 11092 7912
rect 11156 7848 11176 7912
rect 10004 7832 11176 7848
rect 10004 7768 11092 7832
rect 11156 7768 11176 7832
rect 10004 7752 11176 7768
rect 10004 7688 11092 7752
rect 11156 7688 11176 7752
rect 10004 7672 11176 7688
rect 10004 7608 11092 7672
rect 11156 7608 11176 7672
rect 10004 7592 11176 7608
rect 10004 7528 11092 7592
rect 11156 7528 11176 7592
rect 10004 7512 11176 7528
rect 10004 7448 11092 7512
rect 11156 7448 11176 7512
rect 10004 7400 11176 7448
rect 11416 8232 12588 8280
rect 11416 8168 12504 8232
rect 12568 8168 12588 8232
rect 11416 8152 12588 8168
rect 11416 8088 12504 8152
rect 12568 8088 12588 8152
rect 11416 8072 12588 8088
rect 11416 8008 12504 8072
rect 12568 8008 12588 8072
rect 11416 7992 12588 8008
rect 11416 7928 12504 7992
rect 12568 7928 12588 7992
rect 11416 7912 12588 7928
rect 11416 7848 12504 7912
rect 12568 7848 12588 7912
rect 11416 7832 12588 7848
rect 11416 7768 12504 7832
rect 12568 7768 12588 7832
rect 11416 7752 12588 7768
rect 11416 7688 12504 7752
rect 12568 7688 12588 7752
rect 11416 7672 12588 7688
rect 11416 7608 12504 7672
rect 12568 7608 12588 7672
rect 11416 7592 12588 7608
rect 11416 7528 12504 7592
rect 12568 7528 12588 7592
rect 11416 7512 12588 7528
rect 11416 7448 12504 7512
rect 12568 7448 12588 7512
rect 11416 7400 12588 7448
rect 12828 8232 14000 8280
rect 12828 8168 13916 8232
rect 13980 8168 14000 8232
rect 12828 8152 14000 8168
rect 12828 8088 13916 8152
rect 13980 8088 14000 8152
rect 12828 8072 14000 8088
rect 12828 8008 13916 8072
rect 13980 8008 14000 8072
rect 12828 7992 14000 8008
rect 12828 7928 13916 7992
rect 13980 7928 14000 7992
rect 12828 7912 14000 7928
rect 12828 7848 13916 7912
rect 13980 7848 14000 7912
rect 12828 7832 14000 7848
rect 12828 7768 13916 7832
rect 13980 7768 14000 7832
rect 12828 7752 14000 7768
rect 12828 7688 13916 7752
rect 13980 7688 14000 7752
rect 12828 7672 14000 7688
rect 12828 7608 13916 7672
rect 13980 7608 14000 7672
rect 12828 7592 14000 7608
rect 12828 7528 13916 7592
rect 13980 7528 14000 7592
rect 12828 7512 14000 7528
rect 12828 7448 13916 7512
rect 13980 7448 14000 7512
rect 12828 7400 14000 7448
rect 14240 8232 15412 8280
rect 14240 8168 15328 8232
rect 15392 8168 15412 8232
rect 14240 8152 15412 8168
rect 14240 8088 15328 8152
rect 15392 8088 15412 8152
rect 14240 8072 15412 8088
rect 14240 8008 15328 8072
rect 15392 8008 15412 8072
rect 14240 7992 15412 8008
rect 14240 7928 15328 7992
rect 15392 7928 15412 7992
rect 14240 7912 15412 7928
rect 14240 7848 15328 7912
rect 15392 7848 15412 7912
rect 14240 7832 15412 7848
rect 14240 7768 15328 7832
rect 15392 7768 15412 7832
rect 14240 7752 15412 7768
rect 14240 7688 15328 7752
rect 15392 7688 15412 7752
rect 14240 7672 15412 7688
rect 14240 7608 15328 7672
rect 15392 7608 15412 7672
rect 14240 7592 15412 7608
rect 14240 7528 15328 7592
rect 15392 7528 15412 7592
rect 14240 7512 15412 7528
rect 14240 7448 15328 7512
rect 15392 7448 15412 7512
rect 14240 7400 15412 7448
rect 15652 8232 16824 8280
rect 15652 8168 16740 8232
rect 16804 8168 16824 8232
rect 15652 8152 16824 8168
rect 15652 8088 16740 8152
rect 16804 8088 16824 8152
rect 15652 8072 16824 8088
rect 15652 8008 16740 8072
rect 16804 8008 16824 8072
rect 15652 7992 16824 8008
rect 15652 7928 16740 7992
rect 16804 7928 16824 7992
rect 15652 7912 16824 7928
rect 15652 7848 16740 7912
rect 16804 7848 16824 7912
rect 15652 7832 16824 7848
rect 15652 7768 16740 7832
rect 16804 7768 16824 7832
rect 15652 7752 16824 7768
rect 15652 7688 16740 7752
rect 16804 7688 16824 7752
rect 15652 7672 16824 7688
rect 15652 7608 16740 7672
rect 16804 7608 16824 7672
rect 15652 7592 16824 7608
rect 15652 7528 16740 7592
rect 16804 7528 16824 7592
rect 15652 7512 16824 7528
rect 15652 7448 16740 7512
rect 16804 7448 16824 7512
rect 15652 7400 16824 7448
rect 17064 8232 18236 8280
rect 17064 8168 18152 8232
rect 18216 8168 18236 8232
rect 17064 8152 18236 8168
rect 17064 8088 18152 8152
rect 18216 8088 18236 8152
rect 17064 8072 18236 8088
rect 17064 8008 18152 8072
rect 18216 8008 18236 8072
rect 17064 7992 18236 8008
rect 17064 7928 18152 7992
rect 18216 7928 18236 7992
rect 17064 7912 18236 7928
rect 17064 7848 18152 7912
rect 18216 7848 18236 7912
rect 17064 7832 18236 7848
rect 17064 7768 18152 7832
rect 18216 7768 18236 7832
rect 17064 7752 18236 7768
rect 17064 7688 18152 7752
rect 18216 7688 18236 7752
rect 17064 7672 18236 7688
rect 17064 7608 18152 7672
rect 18216 7608 18236 7672
rect 17064 7592 18236 7608
rect 17064 7528 18152 7592
rect 18216 7528 18236 7592
rect 17064 7512 18236 7528
rect 17064 7448 18152 7512
rect 18216 7448 18236 7512
rect 17064 7400 18236 7448
rect 18476 8232 19648 8280
rect 18476 8168 19564 8232
rect 19628 8168 19648 8232
rect 18476 8152 19648 8168
rect 18476 8088 19564 8152
rect 19628 8088 19648 8152
rect 18476 8072 19648 8088
rect 18476 8008 19564 8072
rect 19628 8008 19648 8072
rect 18476 7992 19648 8008
rect 18476 7928 19564 7992
rect 19628 7928 19648 7992
rect 18476 7912 19648 7928
rect 18476 7848 19564 7912
rect 19628 7848 19648 7912
rect 18476 7832 19648 7848
rect 18476 7768 19564 7832
rect 19628 7768 19648 7832
rect 18476 7752 19648 7768
rect 18476 7688 19564 7752
rect 19628 7688 19648 7752
rect 18476 7672 19648 7688
rect 18476 7608 19564 7672
rect 19628 7608 19648 7672
rect 18476 7592 19648 7608
rect 18476 7528 19564 7592
rect 19628 7528 19648 7592
rect 18476 7512 19648 7528
rect 18476 7448 19564 7512
rect 19628 7448 19648 7512
rect 18476 7400 19648 7448
rect 19888 8232 21060 8280
rect 19888 8168 20976 8232
rect 21040 8168 21060 8232
rect 19888 8152 21060 8168
rect 19888 8088 20976 8152
rect 21040 8088 21060 8152
rect 19888 8072 21060 8088
rect 19888 8008 20976 8072
rect 21040 8008 21060 8072
rect 19888 7992 21060 8008
rect 19888 7928 20976 7992
rect 21040 7928 21060 7992
rect 19888 7912 21060 7928
rect 19888 7848 20976 7912
rect 21040 7848 21060 7912
rect 19888 7832 21060 7848
rect 19888 7768 20976 7832
rect 21040 7768 21060 7832
rect 19888 7752 21060 7768
rect 19888 7688 20976 7752
rect 21040 7688 21060 7752
rect 19888 7672 21060 7688
rect 19888 7608 20976 7672
rect 21040 7608 21060 7672
rect 19888 7592 21060 7608
rect 19888 7528 20976 7592
rect 21040 7528 21060 7592
rect 19888 7512 21060 7528
rect 19888 7448 20976 7512
rect 21040 7448 21060 7512
rect 19888 7400 21060 7448
rect 21300 8232 22472 8280
rect 21300 8168 22388 8232
rect 22452 8168 22472 8232
rect 21300 8152 22472 8168
rect 21300 8088 22388 8152
rect 22452 8088 22472 8152
rect 21300 8072 22472 8088
rect 21300 8008 22388 8072
rect 22452 8008 22472 8072
rect 21300 7992 22472 8008
rect 21300 7928 22388 7992
rect 22452 7928 22472 7992
rect 21300 7912 22472 7928
rect 21300 7848 22388 7912
rect 22452 7848 22472 7912
rect 21300 7832 22472 7848
rect 21300 7768 22388 7832
rect 22452 7768 22472 7832
rect 21300 7752 22472 7768
rect 21300 7688 22388 7752
rect 22452 7688 22472 7752
rect 21300 7672 22472 7688
rect 21300 7608 22388 7672
rect 22452 7608 22472 7672
rect 21300 7592 22472 7608
rect 21300 7528 22388 7592
rect 22452 7528 22472 7592
rect 21300 7512 22472 7528
rect 21300 7448 22388 7512
rect 22452 7448 22472 7512
rect 21300 7400 22472 7448
rect 22712 8232 23884 8280
rect 22712 8168 23800 8232
rect 23864 8168 23884 8232
rect 22712 8152 23884 8168
rect 22712 8088 23800 8152
rect 23864 8088 23884 8152
rect 22712 8072 23884 8088
rect 22712 8008 23800 8072
rect 23864 8008 23884 8072
rect 22712 7992 23884 8008
rect 22712 7928 23800 7992
rect 23864 7928 23884 7992
rect 22712 7912 23884 7928
rect 22712 7848 23800 7912
rect 23864 7848 23884 7912
rect 22712 7832 23884 7848
rect 22712 7768 23800 7832
rect 23864 7768 23884 7832
rect 22712 7752 23884 7768
rect 22712 7688 23800 7752
rect 23864 7688 23884 7752
rect 22712 7672 23884 7688
rect 22712 7608 23800 7672
rect 23864 7608 23884 7672
rect 22712 7592 23884 7608
rect 22712 7528 23800 7592
rect 23864 7528 23884 7592
rect 22712 7512 23884 7528
rect 22712 7448 23800 7512
rect 23864 7448 23884 7512
rect 22712 7400 23884 7448
rect -23884 7112 -22712 7160
rect -23884 7048 -22796 7112
rect -22732 7048 -22712 7112
rect -23884 7032 -22712 7048
rect -23884 6968 -22796 7032
rect -22732 6968 -22712 7032
rect -23884 6952 -22712 6968
rect -23884 6888 -22796 6952
rect -22732 6888 -22712 6952
rect -23884 6872 -22712 6888
rect -23884 6808 -22796 6872
rect -22732 6808 -22712 6872
rect -23884 6792 -22712 6808
rect -23884 6728 -22796 6792
rect -22732 6728 -22712 6792
rect -23884 6712 -22712 6728
rect -23884 6648 -22796 6712
rect -22732 6648 -22712 6712
rect -23884 6632 -22712 6648
rect -23884 6568 -22796 6632
rect -22732 6568 -22712 6632
rect -23884 6552 -22712 6568
rect -23884 6488 -22796 6552
rect -22732 6488 -22712 6552
rect -23884 6472 -22712 6488
rect -23884 6408 -22796 6472
rect -22732 6408 -22712 6472
rect -23884 6392 -22712 6408
rect -23884 6328 -22796 6392
rect -22732 6328 -22712 6392
rect -23884 6280 -22712 6328
rect -22472 7112 -21300 7160
rect -22472 7048 -21384 7112
rect -21320 7048 -21300 7112
rect -22472 7032 -21300 7048
rect -22472 6968 -21384 7032
rect -21320 6968 -21300 7032
rect -22472 6952 -21300 6968
rect -22472 6888 -21384 6952
rect -21320 6888 -21300 6952
rect -22472 6872 -21300 6888
rect -22472 6808 -21384 6872
rect -21320 6808 -21300 6872
rect -22472 6792 -21300 6808
rect -22472 6728 -21384 6792
rect -21320 6728 -21300 6792
rect -22472 6712 -21300 6728
rect -22472 6648 -21384 6712
rect -21320 6648 -21300 6712
rect -22472 6632 -21300 6648
rect -22472 6568 -21384 6632
rect -21320 6568 -21300 6632
rect -22472 6552 -21300 6568
rect -22472 6488 -21384 6552
rect -21320 6488 -21300 6552
rect -22472 6472 -21300 6488
rect -22472 6408 -21384 6472
rect -21320 6408 -21300 6472
rect -22472 6392 -21300 6408
rect -22472 6328 -21384 6392
rect -21320 6328 -21300 6392
rect -22472 6280 -21300 6328
rect -21060 7112 -19888 7160
rect -21060 7048 -19972 7112
rect -19908 7048 -19888 7112
rect -21060 7032 -19888 7048
rect -21060 6968 -19972 7032
rect -19908 6968 -19888 7032
rect -21060 6952 -19888 6968
rect -21060 6888 -19972 6952
rect -19908 6888 -19888 6952
rect -21060 6872 -19888 6888
rect -21060 6808 -19972 6872
rect -19908 6808 -19888 6872
rect -21060 6792 -19888 6808
rect -21060 6728 -19972 6792
rect -19908 6728 -19888 6792
rect -21060 6712 -19888 6728
rect -21060 6648 -19972 6712
rect -19908 6648 -19888 6712
rect -21060 6632 -19888 6648
rect -21060 6568 -19972 6632
rect -19908 6568 -19888 6632
rect -21060 6552 -19888 6568
rect -21060 6488 -19972 6552
rect -19908 6488 -19888 6552
rect -21060 6472 -19888 6488
rect -21060 6408 -19972 6472
rect -19908 6408 -19888 6472
rect -21060 6392 -19888 6408
rect -21060 6328 -19972 6392
rect -19908 6328 -19888 6392
rect -21060 6280 -19888 6328
rect -19648 7112 -18476 7160
rect -19648 7048 -18560 7112
rect -18496 7048 -18476 7112
rect -19648 7032 -18476 7048
rect -19648 6968 -18560 7032
rect -18496 6968 -18476 7032
rect -19648 6952 -18476 6968
rect -19648 6888 -18560 6952
rect -18496 6888 -18476 6952
rect -19648 6872 -18476 6888
rect -19648 6808 -18560 6872
rect -18496 6808 -18476 6872
rect -19648 6792 -18476 6808
rect -19648 6728 -18560 6792
rect -18496 6728 -18476 6792
rect -19648 6712 -18476 6728
rect -19648 6648 -18560 6712
rect -18496 6648 -18476 6712
rect -19648 6632 -18476 6648
rect -19648 6568 -18560 6632
rect -18496 6568 -18476 6632
rect -19648 6552 -18476 6568
rect -19648 6488 -18560 6552
rect -18496 6488 -18476 6552
rect -19648 6472 -18476 6488
rect -19648 6408 -18560 6472
rect -18496 6408 -18476 6472
rect -19648 6392 -18476 6408
rect -19648 6328 -18560 6392
rect -18496 6328 -18476 6392
rect -19648 6280 -18476 6328
rect -18236 7112 -17064 7160
rect -18236 7048 -17148 7112
rect -17084 7048 -17064 7112
rect -18236 7032 -17064 7048
rect -18236 6968 -17148 7032
rect -17084 6968 -17064 7032
rect -18236 6952 -17064 6968
rect -18236 6888 -17148 6952
rect -17084 6888 -17064 6952
rect -18236 6872 -17064 6888
rect -18236 6808 -17148 6872
rect -17084 6808 -17064 6872
rect -18236 6792 -17064 6808
rect -18236 6728 -17148 6792
rect -17084 6728 -17064 6792
rect -18236 6712 -17064 6728
rect -18236 6648 -17148 6712
rect -17084 6648 -17064 6712
rect -18236 6632 -17064 6648
rect -18236 6568 -17148 6632
rect -17084 6568 -17064 6632
rect -18236 6552 -17064 6568
rect -18236 6488 -17148 6552
rect -17084 6488 -17064 6552
rect -18236 6472 -17064 6488
rect -18236 6408 -17148 6472
rect -17084 6408 -17064 6472
rect -18236 6392 -17064 6408
rect -18236 6328 -17148 6392
rect -17084 6328 -17064 6392
rect -18236 6280 -17064 6328
rect -16824 7112 -15652 7160
rect -16824 7048 -15736 7112
rect -15672 7048 -15652 7112
rect -16824 7032 -15652 7048
rect -16824 6968 -15736 7032
rect -15672 6968 -15652 7032
rect -16824 6952 -15652 6968
rect -16824 6888 -15736 6952
rect -15672 6888 -15652 6952
rect -16824 6872 -15652 6888
rect -16824 6808 -15736 6872
rect -15672 6808 -15652 6872
rect -16824 6792 -15652 6808
rect -16824 6728 -15736 6792
rect -15672 6728 -15652 6792
rect -16824 6712 -15652 6728
rect -16824 6648 -15736 6712
rect -15672 6648 -15652 6712
rect -16824 6632 -15652 6648
rect -16824 6568 -15736 6632
rect -15672 6568 -15652 6632
rect -16824 6552 -15652 6568
rect -16824 6488 -15736 6552
rect -15672 6488 -15652 6552
rect -16824 6472 -15652 6488
rect -16824 6408 -15736 6472
rect -15672 6408 -15652 6472
rect -16824 6392 -15652 6408
rect -16824 6328 -15736 6392
rect -15672 6328 -15652 6392
rect -16824 6280 -15652 6328
rect -15412 7112 -14240 7160
rect -15412 7048 -14324 7112
rect -14260 7048 -14240 7112
rect -15412 7032 -14240 7048
rect -15412 6968 -14324 7032
rect -14260 6968 -14240 7032
rect -15412 6952 -14240 6968
rect -15412 6888 -14324 6952
rect -14260 6888 -14240 6952
rect -15412 6872 -14240 6888
rect -15412 6808 -14324 6872
rect -14260 6808 -14240 6872
rect -15412 6792 -14240 6808
rect -15412 6728 -14324 6792
rect -14260 6728 -14240 6792
rect -15412 6712 -14240 6728
rect -15412 6648 -14324 6712
rect -14260 6648 -14240 6712
rect -15412 6632 -14240 6648
rect -15412 6568 -14324 6632
rect -14260 6568 -14240 6632
rect -15412 6552 -14240 6568
rect -15412 6488 -14324 6552
rect -14260 6488 -14240 6552
rect -15412 6472 -14240 6488
rect -15412 6408 -14324 6472
rect -14260 6408 -14240 6472
rect -15412 6392 -14240 6408
rect -15412 6328 -14324 6392
rect -14260 6328 -14240 6392
rect -15412 6280 -14240 6328
rect -14000 7112 -12828 7160
rect -14000 7048 -12912 7112
rect -12848 7048 -12828 7112
rect -14000 7032 -12828 7048
rect -14000 6968 -12912 7032
rect -12848 6968 -12828 7032
rect -14000 6952 -12828 6968
rect -14000 6888 -12912 6952
rect -12848 6888 -12828 6952
rect -14000 6872 -12828 6888
rect -14000 6808 -12912 6872
rect -12848 6808 -12828 6872
rect -14000 6792 -12828 6808
rect -14000 6728 -12912 6792
rect -12848 6728 -12828 6792
rect -14000 6712 -12828 6728
rect -14000 6648 -12912 6712
rect -12848 6648 -12828 6712
rect -14000 6632 -12828 6648
rect -14000 6568 -12912 6632
rect -12848 6568 -12828 6632
rect -14000 6552 -12828 6568
rect -14000 6488 -12912 6552
rect -12848 6488 -12828 6552
rect -14000 6472 -12828 6488
rect -14000 6408 -12912 6472
rect -12848 6408 -12828 6472
rect -14000 6392 -12828 6408
rect -14000 6328 -12912 6392
rect -12848 6328 -12828 6392
rect -14000 6280 -12828 6328
rect -12588 7112 -11416 7160
rect -12588 7048 -11500 7112
rect -11436 7048 -11416 7112
rect -12588 7032 -11416 7048
rect -12588 6968 -11500 7032
rect -11436 6968 -11416 7032
rect -12588 6952 -11416 6968
rect -12588 6888 -11500 6952
rect -11436 6888 -11416 6952
rect -12588 6872 -11416 6888
rect -12588 6808 -11500 6872
rect -11436 6808 -11416 6872
rect -12588 6792 -11416 6808
rect -12588 6728 -11500 6792
rect -11436 6728 -11416 6792
rect -12588 6712 -11416 6728
rect -12588 6648 -11500 6712
rect -11436 6648 -11416 6712
rect -12588 6632 -11416 6648
rect -12588 6568 -11500 6632
rect -11436 6568 -11416 6632
rect -12588 6552 -11416 6568
rect -12588 6488 -11500 6552
rect -11436 6488 -11416 6552
rect -12588 6472 -11416 6488
rect -12588 6408 -11500 6472
rect -11436 6408 -11416 6472
rect -12588 6392 -11416 6408
rect -12588 6328 -11500 6392
rect -11436 6328 -11416 6392
rect -12588 6280 -11416 6328
rect -11176 7112 -10004 7160
rect -11176 7048 -10088 7112
rect -10024 7048 -10004 7112
rect -11176 7032 -10004 7048
rect -11176 6968 -10088 7032
rect -10024 6968 -10004 7032
rect -11176 6952 -10004 6968
rect -11176 6888 -10088 6952
rect -10024 6888 -10004 6952
rect -11176 6872 -10004 6888
rect -11176 6808 -10088 6872
rect -10024 6808 -10004 6872
rect -11176 6792 -10004 6808
rect -11176 6728 -10088 6792
rect -10024 6728 -10004 6792
rect -11176 6712 -10004 6728
rect -11176 6648 -10088 6712
rect -10024 6648 -10004 6712
rect -11176 6632 -10004 6648
rect -11176 6568 -10088 6632
rect -10024 6568 -10004 6632
rect -11176 6552 -10004 6568
rect -11176 6488 -10088 6552
rect -10024 6488 -10004 6552
rect -11176 6472 -10004 6488
rect -11176 6408 -10088 6472
rect -10024 6408 -10004 6472
rect -11176 6392 -10004 6408
rect -11176 6328 -10088 6392
rect -10024 6328 -10004 6392
rect -11176 6280 -10004 6328
rect -9764 7112 -8592 7160
rect -9764 7048 -8676 7112
rect -8612 7048 -8592 7112
rect -9764 7032 -8592 7048
rect -9764 6968 -8676 7032
rect -8612 6968 -8592 7032
rect -9764 6952 -8592 6968
rect -9764 6888 -8676 6952
rect -8612 6888 -8592 6952
rect -9764 6872 -8592 6888
rect -9764 6808 -8676 6872
rect -8612 6808 -8592 6872
rect -9764 6792 -8592 6808
rect -9764 6728 -8676 6792
rect -8612 6728 -8592 6792
rect -9764 6712 -8592 6728
rect -9764 6648 -8676 6712
rect -8612 6648 -8592 6712
rect -9764 6632 -8592 6648
rect -9764 6568 -8676 6632
rect -8612 6568 -8592 6632
rect -9764 6552 -8592 6568
rect -9764 6488 -8676 6552
rect -8612 6488 -8592 6552
rect -9764 6472 -8592 6488
rect -9764 6408 -8676 6472
rect -8612 6408 -8592 6472
rect -9764 6392 -8592 6408
rect -9764 6328 -8676 6392
rect -8612 6328 -8592 6392
rect -9764 6280 -8592 6328
rect -8352 7112 -7180 7160
rect -8352 7048 -7264 7112
rect -7200 7048 -7180 7112
rect -8352 7032 -7180 7048
rect -8352 6968 -7264 7032
rect -7200 6968 -7180 7032
rect -8352 6952 -7180 6968
rect -8352 6888 -7264 6952
rect -7200 6888 -7180 6952
rect -8352 6872 -7180 6888
rect -8352 6808 -7264 6872
rect -7200 6808 -7180 6872
rect -8352 6792 -7180 6808
rect -8352 6728 -7264 6792
rect -7200 6728 -7180 6792
rect -8352 6712 -7180 6728
rect -8352 6648 -7264 6712
rect -7200 6648 -7180 6712
rect -8352 6632 -7180 6648
rect -8352 6568 -7264 6632
rect -7200 6568 -7180 6632
rect -8352 6552 -7180 6568
rect -8352 6488 -7264 6552
rect -7200 6488 -7180 6552
rect -8352 6472 -7180 6488
rect -8352 6408 -7264 6472
rect -7200 6408 -7180 6472
rect -8352 6392 -7180 6408
rect -8352 6328 -7264 6392
rect -7200 6328 -7180 6392
rect -8352 6280 -7180 6328
rect -6940 7112 -5768 7160
rect -6940 7048 -5852 7112
rect -5788 7048 -5768 7112
rect -6940 7032 -5768 7048
rect -6940 6968 -5852 7032
rect -5788 6968 -5768 7032
rect -6940 6952 -5768 6968
rect -6940 6888 -5852 6952
rect -5788 6888 -5768 6952
rect -6940 6872 -5768 6888
rect -6940 6808 -5852 6872
rect -5788 6808 -5768 6872
rect -6940 6792 -5768 6808
rect -6940 6728 -5852 6792
rect -5788 6728 -5768 6792
rect -6940 6712 -5768 6728
rect -6940 6648 -5852 6712
rect -5788 6648 -5768 6712
rect -6940 6632 -5768 6648
rect -6940 6568 -5852 6632
rect -5788 6568 -5768 6632
rect -6940 6552 -5768 6568
rect -6940 6488 -5852 6552
rect -5788 6488 -5768 6552
rect -6940 6472 -5768 6488
rect -6940 6408 -5852 6472
rect -5788 6408 -5768 6472
rect -6940 6392 -5768 6408
rect -6940 6328 -5852 6392
rect -5788 6328 -5768 6392
rect -6940 6280 -5768 6328
rect -5528 7112 -4356 7160
rect -5528 7048 -4440 7112
rect -4376 7048 -4356 7112
rect -5528 7032 -4356 7048
rect -5528 6968 -4440 7032
rect -4376 6968 -4356 7032
rect -5528 6952 -4356 6968
rect -5528 6888 -4440 6952
rect -4376 6888 -4356 6952
rect -5528 6872 -4356 6888
rect -5528 6808 -4440 6872
rect -4376 6808 -4356 6872
rect -5528 6792 -4356 6808
rect -5528 6728 -4440 6792
rect -4376 6728 -4356 6792
rect -5528 6712 -4356 6728
rect -5528 6648 -4440 6712
rect -4376 6648 -4356 6712
rect -5528 6632 -4356 6648
rect -5528 6568 -4440 6632
rect -4376 6568 -4356 6632
rect -5528 6552 -4356 6568
rect -5528 6488 -4440 6552
rect -4376 6488 -4356 6552
rect -5528 6472 -4356 6488
rect -5528 6408 -4440 6472
rect -4376 6408 -4356 6472
rect -5528 6392 -4356 6408
rect -5528 6328 -4440 6392
rect -4376 6328 -4356 6392
rect -5528 6280 -4356 6328
rect -4116 7112 -2944 7160
rect -4116 7048 -3028 7112
rect -2964 7048 -2944 7112
rect -4116 7032 -2944 7048
rect -4116 6968 -3028 7032
rect -2964 6968 -2944 7032
rect -4116 6952 -2944 6968
rect -4116 6888 -3028 6952
rect -2964 6888 -2944 6952
rect -4116 6872 -2944 6888
rect -4116 6808 -3028 6872
rect -2964 6808 -2944 6872
rect -4116 6792 -2944 6808
rect -4116 6728 -3028 6792
rect -2964 6728 -2944 6792
rect -4116 6712 -2944 6728
rect -4116 6648 -3028 6712
rect -2964 6648 -2944 6712
rect -4116 6632 -2944 6648
rect -4116 6568 -3028 6632
rect -2964 6568 -2944 6632
rect -4116 6552 -2944 6568
rect -4116 6488 -3028 6552
rect -2964 6488 -2944 6552
rect -4116 6472 -2944 6488
rect -4116 6408 -3028 6472
rect -2964 6408 -2944 6472
rect -4116 6392 -2944 6408
rect -4116 6328 -3028 6392
rect -2964 6328 -2944 6392
rect -4116 6280 -2944 6328
rect -2704 7112 -1532 7160
rect -2704 7048 -1616 7112
rect -1552 7048 -1532 7112
rect -2704 7032 -1532 7048
rect -2704 6968 -1616 7032
rect -1552 6968 -1532 7032
rect -2704 6952 -1532 6968
rect -2704 6888 -1616 6952
rect -1552 6888 -1532 6952
rect -2704 6872 -1532 6888
rect -2704 6808 -1616 6872
rect -1552 6808 -1532 6872
rect -2704 6792 -1532 6808
rect -2704 6728 -1616 6792
rect -1552 6728 -1532 6792
rect -2704 6712 -1532 6728
rect -2704 6648 -1616 6712
rect -1552 6648 -1532 6712
rect -2704 6632 -1532 6648
rect -2704 6568 -1616 6632
rect -1552 6568 -1532 6632
rect -2704 6552 -1532 6568
rect -2704 6488 -1616 6552
rect -1552 6488 -1532 6552
rect -2704 6472 -1532 6488
rect -2704 6408 -1616 6472
rect -1552 6408 -1532 6472
rect -2704 6392 -1532 6408
rect -2704 6328 -1616 6392
rect -1552 6328 -1532 6392
rect -2704 6280 -1532 6328
rect -1292 7112 -120 7160
rect -1292 7048 -204 7112
rect -140 7048 -120 7112
rect -1292 7032 -120 7048
rect -1292 6968 -204 7032
rect -140 6968 -120 7032
rect -1292 6952 -120 6968
rect -1292 6888 -204 6952
rect -140 6888 -120 6952
rect -1292 6872 -120 6888
rect -1292 6808 -204 6872
rect -140 6808 -120 6872
rect -1292 6792 -120 6808
rect -1292 6728 -204 6792
rect -140 6728 -120 6792
rect -1292 6712 -120 6728
rect -1292 6648 -204 6712
rect -140 6648 -120 6712
rect -1292 6632 -120 6648
rect -1292 6568 -204 6632
rect -140 6568 -120 6632
rect -1292 6552 -120 6568
rect -1292 6488 -204 6552
rect -140 6488 -120 6552
rect -1292 6472 -120 6488
rect -1292 6408 -204 6472
rect -140 6408 -120 6472
rect -1292 6392 -120 6408
rect -1292 6328 -204 6392
rect -140 6328 -120 6392
rect -1292 6280 -120 6328
rect 120 7112 1292 7160
rect 120 7048 1208 7112
rect 1272 7048 1292 7112
rect 120 7032 1292 7048
rect 120 6968 1208 7032
rect 1272 6968 1292 7032
rect 120 6952 1292 6968
rect 120 6888 1208 6952
rect 1272 6888 1292 6952
rect 120 6872 1292 6888
rect 120 6808 1208 6872
rect 1272 6808 1292 6872
rect 120 6792 1292 6808
rect 120 6728 1208 6792
rect 1272 6728 1292 6792
rect 120 6712 1292 6728
rect 120 6648 1208 6712
rect 1272 6648 1292 6712
rect 120 6632 1292 6648
rect 120 6568 1208 6632
rect 1272 6568 1292 6632
rect 120 6552 1292 6568
rect 120 6488 1208 6552
rect 1272 6488 1292 6552
rect 120 6472 1292 6488
rect 120 6408 1208 6472
rect 1272 6408 1292 6472
rect 120 6392 1292 6408
rect 120 6328 1208 6392
rect 1272 6328 1292 6392
rect 120 6280 1292 6328
rect 1532 7112 2704 7160
rect 1532 7048 2620 7112
rect 2684 7048 2704 7112
rect 1532 7032 2704 7048
rect 1532 6968 2620 7032
rect 2684 6968 2704 7032
rect 1532 6952 2704 6968
rect 1532 6888 2620 6952
rect 2684 6888 2704 6952
rect 1532 6872 2704 6888
rect 1532 6808 2620 6872
rect 2684 6808 2704 6872
rect 1532 6792 2704 6808
rect 1532 6728 2620 6792
rect 2684 6728 2704 6792
rect 1532 6712 2704 6728
rect 1532 6648 2620 6712
rect 2684 6648 2704 6712
rect 1532 6632 2704 6648
rect 1532 6568 2620 6632
rect 2684 6568 2704 6632
rect 1532 6552 2704 6568
rect 1532 6488 2620 6552
rect 2684 6488 2704 6552
rect 1532 6472 2704 6488
rect 1532 6408 2620 6472
rect 2684 6408 2704 6472
rect 1532 6392 2704 6408
rect 1532 6328 2620 6392
rect 2684 6328 2704 6392
rect 1532 6280 2704 6328
rect 2944 7112 4116 7160
rect 2944 7048 4032 7112
rect 4096 7048 4116 7112
rect 2944 7032 4116 7048
rect 2944 6968 4032 7032
rect 4096 6968 4116 7032
rect 2944 6952 4116 6968
rect 2944 6888 4032 6952
rect 4096 6888 4116 6952
rect 2944 6872 4116 6888
rect 2944 6808 4032 6872
rect 4096 6808 4116 6872
rect 2944 6792 4116 6808
rect 2944 6728 4032 6792
rect 4096 6728 4116 6792
rect 2944 6712 4116 6728
rect 2944 6648 4032 6712
rect 4096 6648 4116 6712
rect 2944 6632 4116 6648
rect 2944 6568 4032 6632
rect 4096 6568 4116 6632
rect 2944 6552 4116 6568
rect 2944 6488 4032 6552
rect 4096 6488 4116 6552
rect 2944 6472 4116 6488
rect 2944 6408 4032 6472
rect 4096 6408 4116 6472
rect 2944 6392 4116 6408
rect 2944 6328 4032 6392
rect 4096 6328 4116 6392
rect 2944 6280 4116 6328
rect 4356 7112 5528 7160
rect 4356 7048 5444 7112
rect 5508 7048 5528 7112
rect 4356 7032 5528 7048
rect 4356 6968 5444 7032
rect 5508 6968 5528 7032
rect 4356 6952 5528 6968
rect 4356 6888 5444 6952
rect 5508 6888 5528 6952
rect 4356 6872 5528 6888
rect 4356 6808 5444 6872
rect 5508 6808 5528 6872
rect 4356 6792 5528 6808
rect 4356 6728 5444 6792
rect 5508 6728 5528 6792
rect 4356 6712 5528 6728
rect 4356 6648 5444 6712
rect 5508 6648 5528 6712
rect 4356 6632 5528 6648
rect 4356 6568 5444 6632
rect 5508 6568 5528 6632
rect 4356 6552 5528 6568
rect 4356 6488 5444 6552
rect 5508 6488 5528 6552
rect 4356 6472 5528 6488
rect 4356 6408 5444 6472
rect 5508 6408 5528 6472
rect 4356 6392 5528 6408
rect 4356 6328 5444 6392
rect 5508 6328 5528 6392
rect 4356 6280 5528 6328
rect 5768 7112 6940 7160
rect 5768 7048 6856 7112
rect 6920 7048 6940 7112
rect 5768 7032 6940 7048
rect 5768 6968 6856 7032
rect 6920 6968 6940 7032
rect 5768 6952 6940 6968
rect 5768 6888 6856 6952
rect 6920 6888 6940 6952
rect 5768 6872 6940 6888
rect 5768 6808 6856 6872
rect 6920 6808 6940 6872
rect 5768 6792 6940 6808
rect 5768 6728 6856 6792
rect 6920 6728 6940 6792
rect 5768 6712 6940 6728
rect 5768 6648 6856 6712
rect 6920 6648 6940 6712
rect 5768 6632 6940 6648
rect 5768 6568 6856 6632
rect 6920 6568 6940 6632
rect 5768 6552 6940 6568
rect 5768 6488 6856 6552
rect 6920 6488 6940 6552
rect 5768 6472 6940 6488
rect 5768 6408 6856 6472
rect 6920 6408 6940 6472
rect 5768 6392 6940 6408
rect 5768 6328 6856 6392
rect 6920 6328 6940 6392
rect 5768 6280 6940 6328
rect 7180 7112 8352 7160
rect 7180 7048 8268 7112
rect 8332 7048 8352 7112
rect 7180 7032 8352 7048
rect 7180 6968 8268 7032
rect 8332 6968 8352 7032
rect 7180 6952 8352 6968
rect 7180 6888 8268 6952
rect 8332 6888 8352 6952
rect 7180 6872 8352 6888
rect 7180 6808 8268 6872
rect 8332 6808 8352 6872
rect 7180 6792 8352 6808
rect 7180 6728 8268 6792
rect 8332 6728 8352 6792
rect 7180 6712 8352 6728
rect 7180 6648 8268 6712
rect 8332 6648 8352 6712
rect 7180 6632 8352 6648
rect 7180 6568 8268 6632
rect 8332 6568 8352 6632
rect 7180 6552 8352 6568
rect 7180 6488 8268 6552
rect 8332 6488 8352 6552
rect 7180 6472 8352 6488
rect 7180 6408 8268 6472
rect 8332 6408 8352 6472
rect 7180 6392 8352 6408
rect 7180 6328 8268 6392
rect 8332 6328 8352 6392
rect 7180 6280 8352 6328
rect 8592 7112 9764 7160
rect 8592 7048 9680 7112
rect 9744 7048 9764 7112
rect 8592 7032 9764 7048
rect 8592 6968 9680 7032
rect 9744 6968 9764 7032
rect 8592 6952 9764 6968
rect 8592 6888 9680 6952
rect 9744 6888 9764 6952
rect 8592 6872 9764 6888
rect 8592 6808 9680 6872
rect 9744 6808 9764 6872
rect 8592 6792 9764 6808
rect 8592 6728 9680 6792
rect 9744 6728 9764 6792
rect 8592 6712 9764 6728
rect 8592 6648 9680 6712
rect 9744 6648 9764 6712
rect 8592 6632 9764 6648
rect 8592 6568 9680 6632
rect 9744 6568 9764 6632
rect 8592 6552 9764 6568
rect 8592 6488 9680 6552
rect 9744 6488 9764 6552
rect 8592 6472 9764 6488
rect 8592 6408 9680 6472
rect 9744 6408 9764 6472
rect 8592 6392 9764 6408
rect 8592 6328 9680 6392
rect 9744 6328 9764 6392
rect 8592 6280 9764 6328
rect 10004 7112 11176 7160
rect 10004 7048 11092 7112
rect 11156 7048 11176 7112
rect 10004 7032 11176 7048
rect 10004 6968 11092 7032
rect 11156 6968 11176 7032
rect 10004 6952 11176 6968
rect 10004 6888 11092 6952
rect 11156 6888 11176 6952
rect 10004 6872 11176 6888
rect 10004 6808 11092 6872
rect 11156 6808 11176 6872
rect 10004 6792 11176 6808
rect 10004 6728 11092 6792
rect 11156 6728 11176 6792
rect 10004 6712 11176 6728
rect 10004 6648 11092 6712
rect 11156 6648 11176 6712
rect 10004 6632 11176 6648
rect 10004 6568 11092 6632
rect 11156 6568 11176 6632
rect 10004 6552 11176 6568
rect 10004 6488 11092 6552
rect 11156 6488 11176 6552
rect 10004 6472 11176 6488
rect 10004 6408 11092 6472
rect 11156 6408 11176 6472
rect 10004 6392 11176 6408
rect 10004 6328 11092 6392
rect 11156 6328 11176 6392
rect 10004 6280 11176 6328
rect 11416 7112 12588 7160
rect 11416 7048 12504 7112
rect 12568 7048 12588 7112
rect 11416 7032 12588 7048
rect 11416 6968 12504 7032
rect 12568 6968 12588 7032
rect 11416 6952 12588 6968
rect 11416 6888 12504 6952
rect 12568 6888 12588 6952
rect 11416 6872 12588 6888
rect 11416 6808 12504 6872
rect 12568 6808 12588 6872
rect 11416 6792 12588 6808
rect 11416 6728 12504 6792
rect 12568 6728 12588 6792
rect 11416 6712 12588 6728
rect 11416 6648 12504 6712
rect 12568 6648 12588 6712
rect 11416 6632 12588 6648
rect 11416 6568 12504 6632
rect 12568 6568 12588 6632
rect 11416 6552 12588 6568
rect 11416 6488 12504 6552
rect 12568 6488 12588 6552
rect 11416 6472 12588 6488
rect 11416 6408 12504 6472
rect 12568 6408 12588 6472
rect 11416 6392 12588 6408
rect 11416 6328 12504 6392
rect 12568 6328 12588 6392
rect 11416 6280 12588 6328
rect 12828 7112 14000 7160
rect 12828 7048 13916 7112
rect 13980 7048 14000 7112
rect 12828 7032 14000 7048
rect 12828 6968 13916 7032
rect 13980 6968 14000 7032
rect 12828 6952 14000 6968
rect 12828 6888 13916 6952
rect 13980 6888 14000 6952
rect 12828 6872 14000 6888
rect 12828 6808 13916 6872
rect 13980 6808 14000 6872
rect 12828 6792 14000 6808
rect 12828 6728 13916 6792
rect 13980 6728 14000 6792
rect 12828 6712 14000 6728
rect 12828 6648 13916 6712
rect 13980 6648 14000 6712
rect 12828 6632 14000 6648
rect 12828 6568 13916 6632
rect 13980 6568 14000 6632
rect 12828 6552 14000 6568
rect 12828 6488 13916 6552
rect 13980 6488 14000 6552
rect 12828 6472 14000 6488
rect 12828 6408 13916 6472
rect 13980 6408 14000 6472
rect 12828 6392 14000 6408
rect 12828 6328 13916 6392
rect 13980 6328 14000 6392
rect 12828 6280 14000 6328
rect 14240 7112 15412 7160
rect 14240 7048 15328 7112
rect 15392 7048 15412 7112
rect 14240 7032 15412 7048
rect 14240 6968 15328 7032
rect 15392 6968 15412 7032
rect 14240 6952 15412 6968
rect 14240 6888 15328 6952
rect 15392 6888 15412 6952
rect 14240 6872 15412 6888
rect 14240 6808 15328 6872
rect 15392 6808 15412 6872
rect 14240 6792 15412 6808
rect 14240 6728 15328 6792
rect 15392 6728 15412 6792
rect 14240 6712 15412 6728
rect 14240 6648 15328 6712
rect 15392 6648 15412 6712
rect 14240 6632 15412 6648
rect 14240 6568 15328 6632
rect 15392 6568 15412 6632
rect 14240 6552 15412 6568
rect 14240 6488 15328 6552
rect 15392 6488 15412 6552
rect 14240 6472 15412 6488
rect 14240 6408 15328 6472
rect 15392 6408 15412 6472
rect 14240 6392 15412 6408
rect 14240 6328 15328 6392
rect 15392 6328 15412 6392
rect 14240 6280 15412 6328
rect 15652 7112 16824 7160
rect 15652 7048 16740 7112
rect 16804 7048 16824 7112
rect 15652 7032 16824 7048
rect 15652 6968 16740 7032
rect 16804 6968 16824 7032
rect 15652 6952 16824 6968
rect 15652 6888 16740 6952
rect 16804 6888 16824 6952
rect 15652 6872 16824 6888
rect 15652 6808 16740 6872
rect 16804 6808 16824 6872
rect 15652 6792 16824 6808
rect 15652 6728 16740 6792
rect 16804 6728 16824 6792
rect 15652 6712 16824 6728
rect 15652 6648 16740 6712
rect 16804 6648 16824 6712
rect 15652 6632 16824 6648
rect 15652 6568 16740 6632
rect 16804 6568 16824 6632
rect 15652 6552 16824 6568
rect 15652 6488 16740 6552
rect 16804 6488 16824 6552
rect 15652 6472 16824 6488
rect 15652 6408 16740 6472
rect 16804 6408 16824 6472
rect 15652 6392 16824 6408
rect 15652 6328 16740 6392
rect 16804 6328 16824 6392
rect 15652 6280 16824 6328
rect 17064 7112 18236 7160
rect 17064 7048 18152 7112
rect 18216 7048 18236 7112
rect 17064 7032 18236 7048
rect 17064 6968 18152 7032
rect 18216 6968 18236 7032
rect 17064 6952 18236 6968
rect 17064 6888 18152 6952
rect 18216 6888 18236 6952
rect 17064 6872 18236 6888
rect 17064 6808 18152 6872
rect 18216 6808 18236 6872
rect 17064 6792 18236 6808
rect 17064 6728 18152 6792
rect 18216 6728 18236 6792
rect 17064 6712 18236 6728
rect 17064 6648 18152 6712
rect 18216 6648 18236 6712
rect 17064 6632 18236 6648
rect 17064 6568 18152 6632
rect 18216 6568 18236 6632
rect 17064 6552 18236 6568
rect 17064 6488 18152 6552
rect 18216 6488 18236 6552
rect 17064 6472 18236 6488
rect 17064 6408 18152 6472
rect 18216 6408 18236 6472
rect 17064 6392 18236 6408
rect 17064 6328 18152 6392
rect 18216 6328 18236 6392
rect 17064 6280 18236 6328
rect 18476 7112 19648 7160
rect 18476 7048 19564 7112
rect 19628 7048 19648 7112
rect 18476 7032 19648 7048
rect 18476 6968 19564 7032
rect 19628 6968 19648 7032
rect 18476 6952 19648 6968
rect 18476 6888 19564 6952
rect 19628 6888 19648 6952
rect 18476 6872 19648 6888
rect 18476 6808 19564 6872
rect 19628 6808 19648 6872
rect 18476 6792 19648 6808
rect 18476 6728 19564 6792
rect 19628 6728 19648 6792
rect 18476 6712 19648 6728
rect 18476 6648 19564 6712
rect 19628 6648 19648 6712
rect 18476 6632 19648 6648
rect 18476 6568 19564 6632
rect 19628 6568 19648 6632
rect 18476 6552 19648 6568
rect 18476 6488 19564 6552
rect 19628 6488 19648 6552
rect 18476 6472 19648 6488
rect 18476 6408 19564 6472
rect 19628 6408 19648 6472
rect 18476 6392 19648 6408
rect 18476 6328 19564 6392
rect 19628 6328 19648 6392
rect 18476 6280 19648 6328
rect 19888 7112 21060 7160
rect 19888 7048 20976 7112
rect 21040 7048 21060 7112
rect 19888 7032 21060 7048
rect 19888 6968 20976 7032
rect 21040 6968 21060 7032
rect 19888 6952 21060 6968
rect 19888 6888 20976 6952
rect 21040 6888 21060 6952
rect 19888 6872 21060 6888
rect 19888 6808 20976 6872
rect 21040 6808 21060 6872
rect 19888 6792 21060 6808
rect 19888 6728 20976 6792
rect 21040 6728 21060 6792
rect 19888 6712 21060 6728
rect 19888 6648 20976 6712
rect 21040 6648 21060 6712
rect 19888 6632 21060 6648
rect 19888 6568 20976 6632
rect 21040 6568 21060 6632
rect 19888 6552 21060 6568
rect 19888 6488 20976 6552
rect 21040 6488 21060 6552
rect 19888 6472 21060 6488
rect 19888 6408 20976 6472
rect 21040 6408 21060 6472
rect 19888 6392 21060 6408
rect 19888 6328 20976 6392
rect 21040 6328 21060 6392
rect 19888 6280 21060 6328
rect 21300 7112 22472 7160
rect 21300 7048 22388 7112
rect 22452 7048 22472 7112
rect 21300 7032 22472 7048
rect 21300 6968 22388 7032
rect 22452 6968 22472 7032
rect 21300 6952 22472 6968
rect 21300 6888 22388 6952
rect 22452 6888 22472 6952
rect 21300 6872 22472 6888
rect 21300 6808 22388 6872
rect 22452 6808 22472 6872
rect 21300 6792 22472 6808
rect 21300 6728 22388 6792
rect 22452 6728 22472 6792
rect 21300 6712 22472 6728
rect 21300 6648 22388 6712
rect 22452 6648 22472 6712
rect 21300 6632 22472 6648
rect 21300 6568 22388 6632
rect 22452 6568 22472 6632
rect 21300 6552 22472 6568
rect 21300 6488 22388 6552
rect 22452 6488 22472 6552
rect 21300 6472 22472 6488
rect 21300 6408 22388 6472
rect 22452 6408 22472 6472
rect 21300 6392 22472 6408
rect 21300 6328 22388 6392
rect 22452 6328 22472 6392
rect 21300 6280 22472 6328
rect 22712 7112 23884 7160
rect 22712 7048 23800 7112
rect 23864 7048 23884 7112
rect 22712 7032 23884 7048
rect 22712 6968 23800 7032
rect 23864 6968 23884 7032
rect 22712 6952 23884 6968
rect 22712 6888 23800 6952
rect 23864 6888 23884 6952
rect 22712 6872 23884 6888
rect 22712 6808 23800 6872
rect 23864 6808 23884 6872
rect 22712 6792 23884 6808
rect 22712 6728 23800 6792
rect 23864 6728 23884 6792
rect 22712 6712 23884 6728
rect 22712 6648 23800 6712
rect 23864 6648 23884 6712
rect 22712 6632 23884 6648
rect 22712 6568 23800 6632
rect 23864 6568 23884 6632
rect 22712 6552 23884 6568
rect 22712 6488 23800 6552
rect 23864 6488 23884 6552
rect 22712 6472 23884 6488
rect 22712 6408 23800 6472
rect 23864 6408 23884 6472
rect 22712 6392 23884 6408
rect 22712 6328 23800 6392
rect 23864 6328 23884 6392
rect 22712 6280 23884 6328
rect -23884 5992 -22712 6040
rect -23884 5928 -22796 5992
rect -22732 5928 -22712 5992
rect -23884 5912 -22712 5928
rect -23884 5848 -22796 5912
rect -22732 5848 -22712 5912
rect -23884 5832 -22712 5848
rect -23884 5768 -22796 5832
rect -22732 5768 -22712 5832
rect -23884 5752 -22712 5768
rect -23884 5688 -22796 5752
rect -22732 5688 -22712 5752
rect -23884 5672 -22712 5688
rect -23884 5608 -22796 5672
rect -22732 5608 -22712 5672
rect -23884 5592 -22712 5608
rect -23884 5528 -22796 5592
rect -22732 5528 -22712 5592
rect -23884 5512 -22712 5528
rect -23884 5448 -22796 5512
rect -22732 5448 -22712 5512
rect -23884 5432 -22712 5448
rect -23884 5368 -22796 5432
rect -22732 5368 -22712 5432
rect -23884 5352 -22712 5368
rect -23884 5288 -22796 5352
rect -22732 5288 -22712 5352
rect -23884 5272 -22712 5288
rect -23884 5208 -22796 5272
rect -22732 5208 -22712 5272
rect -23884 5160 -22712 5208
rect -22472 5992 -21300 6040
rect -22472 5928 -21384 5992
rect -21320 5928 -21300 5992
rect -22472 5912 -21300 5928
rect -22472 5848 -21384 5912
rect -21320 5848 -21300 5912
rect -22472 5832 -21300 5848
rect -22472 5768 -21384 5832
rect -21320 5768 -21300 5832
rect -22472 5752 -21300 5768
rect -22472 5688 -21384 5752
rect -21320 5688 -21300 5752
rect -22472 5672 -21300 5688
rect -22472 5608 -21384 5672
rect -21320 5608 -21300 5672
rect -22472 5592 -21300 5608
rect -22472 5528 -21384 5592
rect -21320 5528 -21300 5592
rect -22472 5512 -21300 5528
rect -22472 5448 -21384 5512
rect -21320 5448 -21300 5512
rect -22472 5432 -21300 5448
rect -22472 5368 -21384 5432
rect -21320 5368 -21300 5432
rect -22472 5352 -21300 5368
rect -22472 5288 -21384 5352
rect -21320 5288 -21300 5352
rect -22472 5272 -21300 5288
rect -22472 5208 -21384 5272
rect -21320 5208 -21300 5272
rect -22472 5160 -21300 5208
rect -21060 5992 -19888 6040
rect -21060 5928 -19972 5992
rect -19908 5928 -19888 5992
rect -21060 5912 -19888 5928
rect -21060 5848 -19972 5912
rect -19908 5848 -19888 5912
rect -21060 5832 -19888 5848
rect -21060 5768 -19972 5832
rect -19908 5768 -19888 5832
rect -21060 5752 -19888 5768
rect -21060 5688 -19972 5752
rect -19908 5688 -19888 5752
rect -21060 5672 -19888 5688
rect -21060 5608 -19972 5672
rect -19908 5608 -19888 5672
rect -21060 5592 -19888 5608
rect -21060 5528 -19972 5592
rect -19908 5528 -19888 5592
rect -21060 5512 -19888 5528
rect -21060 5448 -19972 5512
rect -19908 5448 -19888 5512
rect -21060 5432 -19888 5448
rect -21060 5368 -19972 5432
rect -19908 5368 -19888 5432
rect -21060 5352 -19888 5368
rect -21060 5288 -19972 5352
rect -19908 5288 -19888 5352
rect -21060 5272 -19888 5288
rect -21060 5208 -19972 5272
rect -19908 5208 -19888 5272
rect -21060 5160 -19888 5208
rect -19648 5992 -18476 6040
rect -19648 5928 -18560 5992
rect -18496 5928 -18476 5992
rect -19648 5912 -18476 5928
rect -19648 5848 -18560 5912
rect -18496 5848 -18476 5912
rect -19648 5832 -18476 5848
rect -19648 5768 -18560 5832
rect -18496 5768 -18476 5832
rect -19648 5752 -18476 5768
rect -19648 5688 -18560 5752
rect -18496 5688 -18476 5752
rect -19648 5672 -18476 5688
rect -19648 5608 -18560 5672
rect -18496 5608 -18476 5672
rect -19648 5592 -18476 5608
rect -19648 5528 -18560 5592
rect -18496 5528 -18476 5592
rect -19648 5512 -18476 5528
rect -19648 5448 -18560 5512
rect -18496 5448 -18476 5512
rect -19648 5432 -18476 5448
rect -19648 5368 -18560 5432
rect -18496 5368 -18476 5432
rect -19648 5352 -18476 5368
rect -19648 5288 -18560 5352
rect -18496 5288 -18476 5352
rect -19648 5272 -18476 5288
rect -19648 5208 -18560 5272
rect -18496 5208 -18476 5272
rect -19648 5160 -18476 5208
rect -18236 5992 -17064 6040
rect -18236 5928 -17148 5992
rect -17084 5928 -17064 5992
rect -18236 5912 -17064 5928
rect -18236 5848 -17148 5912
rect -17084 5848 -17064 5912
rect -18236 5832 -17064 5848
rect -18236 5768 -17148 5832
rect -17084 5768 -17064 5832
rect -18236 5752 -17064 5768
rect -18236 5688 -17148 5752
rect -17084 5688 -17064 5752
rect -18236 5672 -17064 5688
rect -18236 5608 -17148 5672
rect -17084 5608 -17064 5672
rect -18236 5592 -17064 5608
rect -18236 5528 -17148 5592
rect -17084 5528 -17064 5592
rect -18236 5512 -17064 5528
rect -18236 5448 -17148 5512
rect -17084 5448 -17064 5512
rect -18236 5432 -17064 5448
rect -18236 5368 -17148 5432
rect -17084 5368 -17064 5432
rect -18236 5352 -17064 5368
rect -18236 5288 -17148 5352
rect -17084 5288 -17064 5352
rect -18236 5272 -17064 5288
rect -18236 5208 -17148 5272
rect -17084 5208 -17064 5272
rect -18236 5160 -17064 5208
rect -16824 5992 -15652 6040
rect -16824 5928 -15736 5992
rect -15672 5928 -15652 5992
rect -16824 5912 -15652 5928
rect -16824 5848 -15736 5912
rect -15672 5848 -15652 5912
rect -16824 5832 -15652 5848
rect -16824 5768 -15736 5832
rect -15672 5768 -15652 5832
rect -16824 5752 -15652 5768
rect -16824 5688 -15736 5752
rect -15672 5688 -15652 5752
rect -16824 5672 -15652 5688
rect -16824 5608 -15736 5672
rect -15672 5608 -15652 5672
rect -16824 5592 -15652 5608
rect -16824 5528 -15736 5592
rect -15672 5528 -15652 5592
rect -16824 5512 -15652 5528
rect -16824 5448 -15736 5512
rect -15672 5448 -15652 5512
rect -16824 5432 -15652 5448
rect -16824 5368 -15736 5432
rect -15672 5368 -15652 5432
rect -16824 5352 -15652 5368
rect -16824 5288 -15736 5352
rect -15672 5288 -15652 5352
rect -16824 5272 -15652 5288
rect -16824 5208 -15736 5272
rect -15672 5208 -15652 5272
rect -16824 5160 -15652 5208
rect -15412 5992 -14240 6040
rect -15412 5928 -14324 5992
rect -14260 5928 -14240 5992
rect -15412 5912 -14240 5928
rect -15412 5848 -14324 5912
rect -14260 5848 -14240 5912
rect -15412 5832 -14240 5848
rect -15412 5768 -14324 5832
rect -14260 5768 -14240 5832
rect -15412 5752 -14240 5768
rect -15412 5688 -14324 5752
rect -14260 5688 -14240 5752
rect -15412 5672 -14240 5688
rect -15412 5608 -14324 5672
rect -14260 5608 -14240 5672
rect -15412 5592 -14240 5608
rect -15412 5528 -14324 5592
rect -14260 5528 -14240 5592
rect -15412 5512 -14240 5528
rect -15412 5448 -14324 5512
rect -14260 5448 -14240 5512
rect -15412 5432 -14240 5448
rect -15412 5368 -14324 5432
rect -14260 5368 -14240 5432
rect -15412 5352 -14240 5368
rect -15412 5288 -14324 5352
rect -14260 5288 -14240 5352
rect -15412 5272 -14240 5288
rect -15412 5208 -14324 5272
rect -14260 5208 -14240 5272
rect -15412 5160 -14240 5208
rect -14000 5992 -12828 6040
rect -14000 5928 -12912 5992
rect -12848 5928 -12828 5992
rect -14000 5912 -12828 5928
rect -14000 5848 -12912 5912
rect -12848 5848 -12828 5912
rect -14000 5832 -12828 5848
rect -14000 5768 -12912 5832
rect -12848 5768 -12828 5832
rect -14000 5752 -12828 5768
rect -14000 5688 -12912 5752
rect -12848 5688 -12828 5752
rect -14000 5672 -12828 5688
rect -14000 5608 -12912 5672
rect -12848 5608 -12828 5672
rect -14000 5592 -12828 5608
rect -14000 5528 -12912 5592
rect -12848 5528 -12828 5592
rect -14000 5512 -12828 5528
rect -14000 5448 -12912 5512
rect -12848 5448 -12828 5512
rect -14000 5432 -12828 5448
rect -14000 5368 -12912 5432
rect -12848 5368 -12828 5432
rect -14000 5352 -12828 5368
rect -14000 5288 -12912 5352
rect -12848 5288 -12828 5352
rect -14000 5272 -12828 5288
rect -14000 5208 -12912 5272
rect -12848 5208 -12828 5272
rect -14000 5160 -12828 5208
rect -12588 5992 -11416 6040
rect -12588 5928 -11500 5992
rect -11436 5928 -11416 5992
rect -12588 5912 -11416 5928
rect -12588 5848 -11500 5912
rect -11436 5848 -11416 5912
rect -12588 5832 -11416 5848
rect -12588 5768 -11500 5832
rect -11436 5768 -11416 5832
rect -12588 5752 -11416 5768
rect -12588 5688 -11500 5752
rect -11436 5688 -11416 5752
rect -12588 5672 -11416 5688
rect -12588 5608 -11500 5672
rect -11436 5608 -11416 5672
rect -12588 5592 -11416 5608
rect -12588 5528 -11500 5592
rect -11436 5528 -11416 5592
rect -12588 5512 -11416 5528
rect -12588 5448 -11500 5512
rect -11436 5448 -11416 5512
rect -12588 5432 -11416 5448
rect -12588 5368 -11500 5432
rect -11436 5368 -11416 5432
rect -12588 5352 -11416 5368
rect -12588 5288 -11500 5352
rect -11436 5288 -11416 5352
rect -12588 5272 -11416 5288
rect -12588 5208 -11500 5272
rect -11436 5208 -11416 5272
rect -12588 5160 -11416 5208
rect -11176 5992 -10004 6040
rect -11176 5928 -10088 5992
rect -10024 5928 -10004 5992
rect -11176 5912 -10004 5928
rect -11176 5848 -10088 5912
rect -10024 5848 -10004 5912
rect -11176 5832 -10004 5848
rect -11176 5768 -10088 5832
rect -10024 5768 -10004 5832
rect -11176 5752 -10004 5768
rect -11176 5688 -10088 5752
rect -10024 5688 -10004 5752
rect -11176 5672 -10004 5688
rect -11176 5608 -10088 5672
rect -10024 5608 -10004 5672
rect -11176 5592 -10004 5608
rect -11176 5528 -10088 5592
rect -10024 5528 -10004 5592
rect -11176 5512 -10004 5528
rect -11176 5448 -10088 5512
rect -10024 5448 -10004 5512
rect -11176 5432 -10004 5448
rect -11176 5368 -10088 5432
rect -10024 5368 -10004 5432
rect -11176 5352 -10004 5368
rect -11176 5288 -10088 5352
rect -10024 5288 -10004 5352
rect -11176 5272 -10004 5288
rect -11176 5208 -10088 5272
rect -10024 5208 -10004 5272
rect -11176 5160 -10004 5208
rect -9764 5992 -8592 6040
rect -9764 5928 -8676 5992
rect -8612 5928 -8592 5992
rect -9764 5912 -8592 5928
rect -9764 5848 -8676 5912
rect -8612 5848 -8592 5912
rect -9764 5832 -8592 5848
rect -9764 5768 -8676 5832
rect -8612 5768 -8592 5832
rect -9764 5752 -8592 5768
rect -9764 5688 -8676 5752
rect -8612 5688 -8592 5752
rect -9764 5672 -8592 5688
rect -9764 5608 -8676 5672
rect -8612 5608 -8592 5672
rect -9764 5592 -8592 5608
rect -9764 5528 -8676 5592
rect -8612 5528 -8592 5592
rect -9764 5512 -8592 5528
rect -9764 5448 -8676 5512
rect -8612 5448 -8592 5512
rect -9764 5432 -8592 5448
rect -9764 5368 -8676 5432
rect -8612 5368 -8592 5432
rect -9764 5352 -8592 5368
rect -9764 5288 -8676 5352
rect -8612 5288 -8592 5352
rect -9764 5272 -8592 5288
rect -9764 5208 -8676 5272
rect -8612 5208 -8592 5272
rect -9764 5160 -8592 5208
rect -8352 5992 -7180 6040
rect -8352 5928 -7264 5992
rect -7200 5928 -7180 5992
rect -8352 5912 -7180 5928
rect -8352 5848 -7264 5912
rect -7200 5848 -7180 5912
rect -8352 5832 -7180 5848
rect -8352 5768 -7264 5832
rect -7200 5768 -7180 5832
rect -8352 5752 -7180 5768
rect -8352 5688 -7264 5752
rect -7200 5688 -7180 5752
rect -8352 5672 -7180 5688
rect -8352 5608 -7264 5672
rect -7200 5608 -7180 5672
rect -8352 5592 -7180 5608
rect -8352 5528 -7264 5592
rect -7200 5528 -7180 5592
rect -8352 5512 -7180 5528
rect -8352 5448 -7264 5512
rect -7200 5448 -7180 5512
rect -8352 5432 -7180 5448
rect -8352 5368 -7264 5432
rect -7200 5368 -7180 5432
rect -8352 5352 -7180 5368
rect -8352 5288 -7264 5352
rect -7200 5288 -7180 5352
rect -8352 5272 -7180 5288
rect -8352 5208 -7264 5272
rect -7200 5208 -7180 5272
rect -8352 5160 -7180 5208
rect -6940 5992 -5768 6040
rect -6940 5928 -5852 5992
rect -5788 5928 -5768 5992
rect -6940 5912 -5768 5928
rect -6940 5848 -5852 5912
rect -5788 5848 -5768 5912
rect -6940 5832 -5768 5848
rect -6940 5768 -5852 5832
rect -5788 5768 -5768 5832
rect -6940 5752 -5768 5768
rect -6940 5688 -5852 5752
rect -5788 5688 -5768 5752
rect -6940 5672 -5768 5688
rect -6940 5608 -5852 5672
rect -5788 5608 -5768 5672
rect -6940 5592 -5768 5608
rect -6940 5528 -5852 5592
rect -5788 5528 -5768 5592
rect -6940 5512 -5768 5528
rect -6940 5448 -5852 5512
rect -5788 5448 -5768 5512
rect -6940 5432 -5768 5448
rect -6940 5368 -5852 5432
rect -5788 5368 -5768 5432
rect -6940 5352 -5768 5368
rect -6940 5288 -5852 5352
rect -5788 5288 -5768 5352
rect -6940 5272 -5768 5288
rect -6940 5208 -5852 5272
rect -5788 5208 -5768 5272
rect -6940 5160 -5768 5208
rect -5528 5992 -4356 6040
rect -5528 5928 -4440 5992
rect -4376 5928 -4356 5992
rect -5528 5912 -4356 5928
rect -5528 5848 -4440 5912
rect -4376 5848 -4356 5912
rect -5528 5832 -4356 5848
rect -5528 5768 -4440 5832
rect -4376 5768 -4356 5832
rect -5528 5752 -4356 5768
rect -5528 5688 -4440 5752
rect -4376 5688 -4356 5752
rect -5528 5672 -4356 5688
rect -5528 5608 -4440 5672
rect -4376 5608 -4356 5672
rect -5528 5592 -4356 5608
rect -5528 5528 -4440 5592
rect -4376 5528 -4356 5592
rect -5528 5512 -4356 5528
rect -5528 5448 -4440 5512
rect -4376 5448 -4356 5512
rect -5528 5432 -4356 5448
rect -5528 5368 -4440 5432
rect -4376 5368 -4356 5432
rect -5528 5352 -4356 5368
rect -5528 5288 -4440 5352
rect -4376 5288 -4356 5352
rect -5528 5272 -4356 5288
rect -5528 5208 -4440 5272
rect -4376 5208 -4356 5272
rect -5528 5160 -4356 5208
rect -4116 5992 -2944 6040
rect -4116 5928 -3028 5992
rect -2964 5928 -2944 5992
rect -4116 5912 -2944 5928
rect -4116 5848 -3028 5912
rect -2964 5848 -2944 5912
rect -4116 5832 -2944 5848
rect -4116 5768 -3028 5832
rect -2964 5768 -2944 5832
rect -4116 5752 -2944 5768
rect -4116 5688 -3028 5752
rect -2964 5688 -2944 5752
rect -4116 5672 -2944 5688
rect -4116 5608 -3028 5672
rect -2964 5608 -2944 5672
rect -4116 5592 -2944 5608
rect -4116 5528 -3028 5592
rect -2964 5528 -2944 5592
rect -4116 5512 -2944 5528
rect -4116 5448 -3028 5512
rect -2964 5448 -2944 5512
rect -4116 5432 -2944 5448
rect -4116 5368 -3028 5432
rect -2964 5368 -2944 5432
rect -4116 5352 -2944 5368
rect -4116 5288 -3028 5352
rect -2964 5288 -2944 5352
rect -4116 5272 -2944 5288
rect -4116 5208 -3028 5272
rect -2964 5208 -2944 5272
rect -4116 5160 -2944 5208
rect -2704 5992 -1532 6040
rect -2704 5928 -1616 5992
rect -1552 5928 -1532 5992
rect -2704 5912 -1532 5928
rect -2704 5848 -1616 5912
rect -1552 5848 -1532 5912
rect -2704 5832 -1532 5848
rect -2704 5768 -1616 5832
rect -1552 5768 -1532 5832
rect -2704 5752 -1532 5768
rect -2704 5688 -1616 5752
rect -1552 5688 -1532 5752
rect -2704 5672 -1532 5688
rect -2704 5608 -1616 5672
rect -1552 5608 -1532 5672
rect -2704 5592 -1532 5608
rect -2704 5528 -1616 5592
rect -1552 5528 -1532 5592
rect -2704 5512 -1532 5528
rect -2704 5448 -1616 5512
rect -1552 5448 -1532 5512
rect -2704 5432 -1532 5448
rect -2704 5368 -1616 5432
rect -1552 5368 -1532 5432
rect -2704 5352 -1532 5368
rect -2704 5288 -1616 5352
rect -1552 5288 -1532 5352
rect -2704 5272 -1532 5288
rect -2704 5208 -1616 5272
rect -1552 5208 -1532 5272
rect -2704 5160 -1532 5208
rect -1292 5992 -120 6040
rect -1292 5928 -204 5992
rect -140 5928 -120 5992
rect -1292 5912 -120 5928
rect -1292 5848 -204 5912
rect -140 5848 -120 5912
rect -1292 5832 -120 5848
rect -1292 5768 -204 5832
rect -140 5768 -120 5832
rect -1292 5752 -120 5768
rect -1292 5688 -204 5752
rect -140 5688 -120 5752
rect -1292 5672 -120 5688
rect -1292 5608 -204 5672
rect -140 5608 -120 5672
rect -1292 5592 -120 5608
rect -1292 5528 -204 5592
rect -140 5528 -120 5592
rect -1292 5512 -120 5528
rect -1292 5448 -204 5512
rect -140 5448 -120 5512
rect -1292 5432 -120 5448
rect -1292 5368 -204 5432
rect -140 5368 -120 5432
rect -1292 5352 -120 5368
rect -1292 5288 -204 5352
rect -140 5288 -120 5352
rect -1292 5272 -120 5288
rect -1292 5208 -204 5272
rect -140 5208 -120 5272
rect -1292 5160 -120 5208
rect 120 5992 1292 6040
rect 120 5928 1208 5992
rect 1272 5928 1292 5992
rect 120 5912 1292 5928
rect 120 5848 1208 5912
rect 1272 5848 1292 5912
rect 120 5832 1292 5848
rect 120 5768 1208 5832
rect 1272 5768 1292 5832
rect 120 5752 1292 5768
rect 120 5688 1208 5752
rect 1272 5688 1292 5752
rect 120 5672 1292 5688
rect 120 5608 1208 5672
rect 1272 5608 1292 5672
rect 120 5592 1292 5608
rect 120 5528 1208 5592
rect 1272 5528 1292 5592
rect 120 5512 1292 5528
rect 120 5448 1208 5512
rect 1272 5448 1292 5512
rect 120 5432 1292 5448
rect 120 5368 1208 5432
rect 1272 5368 1292 5432
rect 120 5352 1292 5368
rect 120 5288 1208 5352
rect 1272 5288 1292 5352
rect 120 5272 1292 5288
rect 120 5208 1208 5272
rect 1272 5208 1292 5272
rect 120 5160 1292 5208
rect 1532 5992 2704 6040
rect 1532 5928 2620 5992
rect 2684 5928 2704 5992
rect 1532 5912 2704 5928
rect 1532 5848 2620 5912
rect 2684 5848 2704 5912
rect 1532 5832 2704 5848
rect 1532 5768 2620 5832
rect 2684 5768 2704 5832
rect 1532 5752 2704 5768
rect 1532 5688 2620 5752
rect 2684 5688 2704 5752
rect 1532 5672 2704 5688
rect 1532 5608 2620 5672
rect 2684 5608 2704 5672
rect 1532 5592 2704 5608
rect 1532 5528 2620 5592
rect 2684 5528 2704 5592
rect 1532 5512 2704 5528
rect 1532 5448 2620 5512
rect 2684 5448 2704 5512
rect 1532 5432 2704 5448
rect 1532 5368 2620 5432
rect 2684 5368 2704 5432
rect 1532 5352 2704 5368
rect 1532 5288 2620 5352
rect 2684 5288 2704 5352
rect 1532 5272 2704 5288
rect 1532 5208 2620 5272
rect 2684 5208 2704 5272
rect 1532 5160 2704 5208
rect 2944 5992 4116 6040
rect 2944 5928 4032 5992
rect 4096 5928 4116 5992
rect 2944 5912 4116 5928
rect 2944 5848 4032 5912
rect 4096 5848 4116 5912
rect 2944 5832 4116 5848
rect 2944 5768 4032 5832
rect 4096 5768 4116 5832
rect 2944 5752 4116 5768
rect 2944 5688 4032 5752
rect 4096 5688 4116 5752
rect 2944 5672 4116 5688
rect 2944 5608 4032 5672
rect 4096 5608 4116 5672
rect 2944 5592 4116 5608
rect 2944 5528 4032 5592
rect 4096 5528 4116 5592
rect 2944 5512 4116 5528
rect 2944 5448 4032 5512
rect 4096 5448 4116 5512
rect 2944 5432 4116 5448
rect 2944 5368 4032 5432
rect 4096 5368 4116 5432
rect 2944 5352 4116 5368
rect 2944 5288 4032 5352
rect 4096 5288 4116 5352
rect 2944 5272 4116 5288
rect 2944 5208 4032 5272
rect 4096 5208 4116 5272
rect 2944 5160 4116 5208
rect 4356 5992 5528 6040
rect 4356 5928 5444 5992
rect 5508 5928 5528 5992
rect 4356 5912 5528 5928
rect 4356 5848 5444 5912
rect 5508 5848 5528 5912
rect 4356 5832 5528 5848
rect 4356 5768 5444 5832
rect 5508 5768 5528 5832
rect 4356 5752 5528 5768
rect 4356 5688 5444 5752
rect 5508 5688 5528 5752
rect 4356 5672 5528 5688
rect 4356 5608 5444 5672
rect 5508 5608 5528 5672
rect 4356 5592 5528 5608
rect 4356 5528 5444 5592
rect 5508 5528 5528 5592
rect 4356 5512 5528 5528
rect 4356 5448 5444 5512
rect 5508 5448 5528 5512
rect 4356 5432 5528 5448
rect 4356 5368 5444 5432
rect 5508 5368 5528 5432
rect 4356 5352 5528 5368
rect 4356 5288 5444 5352
rect 5508 5288 5528 5352
rect 4356 5272 5528 5288
rect 4356 5208 5444 5272
rect 5508 5208 5528 5272
rect 4356 5160 5528 5208
rect 5768 5992 6940 6040
rect 5768 5928 6856 5992
rect 6920 5928 6940 5992
rect 5768 5912 6940 5928
rect 5768 5848 6856 5912
rect 6920 5848 6940 5912
rect 5768 5832 6940 5848
rect 5768 5768 6856 5832
rect 6920 5768 6940 5832
rect 5768 5752 6940 5768
rect 5768 5688 6856 5752
rect 6920 5688 6940 5752
rect 5768 5672 6940 5688
rect 5768 5608 6856 5672
rect 6920 5608 6940 5672
rect 5768 5592 6940 5608
rect 5768 5528 6856 5592
rect 6920 5528 6940 5592
rect 5768 5512 6940 5528
rect 5768 5448 6856 5512
rect 6920 5448 6940 5512
rect 5768 5432 6940 5448
rect 5768 5368 6856 5432
rect 6920 5368 6940 5432
rect 5768 5352 6940 5368
rect 5768 5288 6856 5352
rect 6920 5288 6940 5352
rect 5768 5272 6940 5288
rect 5768 5208 6856 5272
rect 6920 5208 6940 5272
rect 5768 5160 6940 5208
rect 7180 5992 8352 6040
rect 7180 5928 8268 5992
rect 8332 5928 8352 5992
rect 7180 5912 8352 5928
rect 7180 5848 8268 5912
rect 8332 5848 8352 5912
rect 7180 5832 8352 5848
rect 7180 5768 8268 5832
rect 8332 5768 8352 5832
rect 7180 5752 8352 5768
rect 7180 5688 8268 5752
rect 8332 5688 8352 5752
rect 7180 5672 8352 5688
rect 7180 5608 8268 5672
rect 8332 5608 8352 5672
rect 7180 5592 8352 5608
rect 7180 5528 8268 5592
rect 8332 5528 8352 5592
rect 7180 5512 8352 5528
rect 7180 5448 8268 5512
rect 8332 5448 8352 5512
rect 7180 5432 8352 5448
rect 7180 5368 8268 5432
rect 8332 5368 8352 5432
rect 7180 5352 8352 5368
rect 7180 5288 8268 5352
rect 8332 5288 8352 5352
rect 7180 5272 8352 5288
rect 7180 5208 8268 5272
rect 8332 5208 8352 5272
rect 7180 5160 8352 5208
rect 8592 5992 9764 6040
rect 8592 5928 9680 5992
rect 9744 5928 9764 5992
rect 8592 5912 9764 5928
rect 8592 5848 9680 5912
rect 9744 5848 9764 5912
rect 8592 5832 9764 5848
rect 8592 5768 9680 5832
rect 9744 5768 9764 5832
rect 8592 5752 9764 5768
rect 8592 5688 9680 5752
rect 9744 5688 9764 5752
rect 8592 5672 9764 5688
rect 8592 5608 9680 5672
rect 9744 5608 9764 5672
rect 8592 5592 9764 5608
rect 8592 5528 9680 5592
rect 9744 5528 9764 5592
rect 8592 5512 9764 5528
rect 8592 5448 9680 5512
rect 9744 5448 9764 5512
rect 8592 5432 9764 5448
rect 8592 5368 9680 5432
rect 9744 5368 9764 5432
rect 8592 5352 9764 5368
rect 8592 5288 9680 5352
rect 9744 5288 9764 5352
rect 8592 5272 9764 5288
rect 8592 5208 9680 5272
rect 9744 5208 9764 5272
rect 8592 5160 9764 5208
rect 10004 5992 11176 6040
rect 10004 5928 11092 5992
rect 11156 5928 11176 5992
rect 10004 5912 11176 5928
rect 10004 5848 11092 5912
rect 11156 5848 11176 5912
rect 10004 5832 11176 5848
rect 10004 5768 11092 5832
rect 11156 5768 11176 5832
rect 10004 5752 11176 5768
rect 10004 5688 11092 5752
rect 11156 5688 11176 5752
rect 10004 5672 11176 5688
rect 10004 5608 11092 5672
rect 11156 5608 11176 5672
rect 10004 5592 11176 5608
rect 10004 5528 11092 5592
rect 11156 5528 11176 5592
rect 10004 5512 11176 5528
rect 10004 5448 11092 5512
rect 11156 5448 11176 5512
rect 10004 5432 11176 5448
rect 10004 5368 11092 5432
rect 11156 5368 11176 5432
rect 10004 5352 11176 5368
rect 10004 5288 11092 5352
rect 11156 5288 11176 5352
rect 10004 5272 11176 5288
rect 10004 5208 11092 5272
rect 11156 5208 11176 5272
rect 10004 5160 11176 5208
rect 11416 5992 12588 6040
rect 11416 5928 12504 5992
rect 12568 5928 12588 5992
rect 11416 5912 12588 5928
rect 11416 5848 12504 5912
rect 12568 5848 12588 5912
rect 11416 5832 12588 5848
rect 11416 5768 12504 5832
rect 12568 5768 12588 5832
rect 11416 5752 12588 5768
rect 11416 5688 12504 5752
rect 12568 5688 12588 5752
rect 11416 5672 12588 5688
rect 11416 5608 12504 5672
rect 12568 5608 12588 5672
rect 11416 5592 12588 5608
rect 11416 5528 12504 5592
rect 12568 5528 12588 5592
rect 11416 5512 12588 5528
rect 11416 5448 12504 5512
rect 12568 5448 12588 5512
rect 11416 5432 12588 5448
rect 11416 5368 12504 5432
rect 12568 5368 12588 5432
rect 11416 5352 12588 5368
rect 11416 5288 12504 5352
rect 12568 5288 12588 5352
rect 11416 5272 12588 5288
rect 11416 5208 12504 5272
rect 12568 5208 12588 5272
rect 11416 5160 12588 5208
rect 12828 5992 14000 6040
rect 12828 5928 13916 5992
rect 13980 5928 14000 5992
rect 12828 5912 14000 5928
rect 12828 5848 13916 5912
rect 13980 5848 14000 5912
rect 12828 5832 14000 5848
rect 12828 5768 13916 5832
rect 13980 5768 14000 5832
rect 12828 5752 14000 5768
rect 12828 5688 13916 5752
rect 13980 5688 14000 5752
rect 12828 5672 14000 5688
rect 12828 5608 13916 5672
rect 13980 5608 14000 5672
rect 12828 5592 14000 5608
rect 12828 5528 13916 5592
rect 13980 5528 14000 5592
rect 12828 5512 14000 5528
rect 12828 5448 13916 5512
rect 13980 5448 14000 5512
rect 12828 5432 14000 5448
rect 12828 5368 13916 5432
rect 13980 5368 14000 5432
rect 12828 5352 14000 5368
rect 12828 5288 13916 5352
rect 13980 5288 14000 5352
rect 12828 5272 14000 5288
rect 12828 5208 13916 5272
rect 13980 5208 14000 5272
rect 12828 5160 14000 5208
rect 14240 5992 15412 6040
rect 14240 5928 15328 5992
rect 15392 5928 15412 5992
rect 14240 5912 15412 5928
rect 14240 5848 15328 5912
rect 15392 5848 15412 5912
rect 14240 5832 15412 5848
rect 14240 5768 15328 5832
rect 15392 5768 15412 5832
rect 14240 5752 15412 5768
rect 14240 5688 15328 5752
rect 15392 5688 15412 5752
rect 14240 5672 15412 5688
rect 14240 5608 15328 5672
rect 15392 5608 15412 5672
rect 14240 5592 15412 5608
rect 14240 5528 15328 5592
rect 15392 5528 15412 5592
rect 14240 5512 15412 5528
rect 14240 5448 15328 5512
rect 15392 5448 15412 5512
rect 14240 5432 15412 5448
rect 14240 5368 15328 5432
rect 15392 5368 15412 5432
rect 14240 5352 15412 5368
rect 14240 5288 15328 5352
rect 15392 5288 15412 5352
rect 14240 5272 15412 5288
rect 14240 5208 15328 5272
rect 15392 5208 15412 5272
rect 14240 5160 15412 5208
rect 15652 5992 16824 6040
rect 15652 5928 16740 5992
rect 16804 5928 16824 5992
rect 15652 5912 16824 5928
rect 15652 5848 16740 5912
rect 16804 5848 16824 5912
rect 15652 5832 16824 5848
rect 15652 5768 16740 5832
rect 16804 5768 16824 5832
rect 15652 5752 16824 5768
rect 15652 5688 16740 5752
rect 16804 5688 16824 5752
rect 15652 5672 16824 5688
rect 15652 5608 16740 5672
rect 16804 5608 16824 5672
rect 15652 5592 16824 5608
rect 15652 5528 16740 5592
rect 16804 5528 16824 5592
rect 15652 5512 16824 5528
rect 15652 5448 16740 5512
rect 16804 5448 16824 5512
rect 15652 5432 16824 5448
rect 15652 5368 16740 5432
rect 16804 5368 16824 5432
rect 15652 5352 16824 5368
rect 15652 5288 16740 5352
rect 16804 5288 16824 5352
rect 15652 5272 16824 5288
rect 15652 5208 16740 5272
rect 16804 5208 16824 5272
rect 15652 5160 16824 5208
rect 17064 5992 18236 6040
rect 17064 5928 18152 5992
rect 18216 5928 18236 5992
rect 17064 5912 18236 5928
rect 17064 5848 18152 5912
rect 18216 5848 18236 5912
rect 17064 5832 18236 5848
rect 17064 5768 18152 5832
rect 18216 5768 18236 5832
rect 17064 5752 18236 5768
rect 17064 5688 18152 5752
rect 18216 5688 18236 5752
rect 17064 5672 18236 5688
rect 17064 5608 18152 5672
rect 18216 5608 18236 5672
rect 17064 5592 18236 5608
rect 17064 5528 18152 5592
rect 18216 5528 18236 5592
rect 17064 5512 18236 5528
rect 17064 5448 18152 5512
rect 18216 5448 18236 5512
rect 17064 5432 18236 5448
rect 17064 5368 18152 5432
rect 18216 5368 18236 5432
rect 17064 5352 18236 5368
rect 17064 5288 18152 5352
rect 18216 5288 18236 5352
rect 17064 5272 18236 5288
rect 17064 5208 18152 5272
rect 18216 5208 18236 5272
rect 17064 5160 18236 5208
rect 18476 5992 19648 6040
rect 18476 5928 19564 5992
rect 19628 5928 19648 5992
rect 18476 5912 19648 5928
rect 18476 5848 19564 5912
rect 19628 5848 19648 5912
rect 18476 5832 19648 5848
rect 18476 5768 19564 5832
rect 19628 5768 19648 5832
rect 18476 5752 19648 5768
rect 18476 5688 19564 5752
rect 19628 5688 19648 5752
rect 18476 5672 19648 5688
rect 18476 5608 19564 5672
rect 19628 5608 19648 5672
rect 18476 5592 19648 5608
rect 18476 5528 19564 5592
rect 19628 5528 19648 5592
rect 18476 5512 19648 5528
rect 18476 5448 19564 5512
rect 19628 5448 19648 5512
rect 18476 5432 19648 5448
rect 18476 5368 19564 5432
rect 19628 5368 19648 5432
rect 18476 5352 19648 5368
rect 18476 5288 19564 5352
rect 19628 5288 19648 5352
rect 18476 5272 19648 5288
rect 18476 5208 19564 5272
rect 19628 5208 19648 5272
rect 18476 5160 19648 5208
rect 19888 5992 21060 6040
rect 19888 5928 20976 5992
rect 21040 5928 21060 5992
rect 19888 5912 21060 5928
rect 19888 5848 20976 5912
rect 21040 5848 21060 5912
rect 19888 5832 21060 5848
rect 19888 5768 20976 5832
rect 21040 5768 21060 5832
rect 19888 5752 21060 5768
rect 19888 5688 20976 5752
rect 21040 5688 21060 5752
rect 19888 5672 21060 5688
rect 19888 5608 20976 5672
rect 21040 5608 21060 5672
rect 19888 5592 21060 5608
rect 19888 5528 20976 5592
rect 21040 5528 21060 5592
rect 19888 5512 21060 5528
rect 19888 5448 20976 5512
rect 21040 5448 21060 5512
rect 19888 5432 21060 5448
rect 19888 5368 20976 5432
rect 21040 5368 21060 5432
rect 19888 5352 21060 5368
rect 19888 5288 20976 5352
rect 21040 5288 21060 5352
rect 19888 5272 21060 5288
rect 19888 5208 20976 5272
rect 21040 5208 21060 5272
rect 19888 5160 21060 5208
rect 21300 5992 22472 6040
rect 21300 5928 22388 5992
rect 22452 5928 22472 5992
rect 21300 5912 22472 5928
rect 21300 5848 22388 5912
rect 22452 5848 22472 5912
rect 21300 5832 22472 5848
rect 21300 5768 22388 5832
rect 22452 5768 22472 5832
rect 21300 5752 22472 5768
rect 21300 5688 22388 5752
rect 22452 5688 22472 5752
rect 21300 5672 22472 5688
rect 21300 5608 22388 5672
rect 22452 5608 22472 5672
rect 21300 5592 22472 5608
rect 21300 5528 22388 5592
rect 22452 5528 22472 5592
rect 21300 5512 22472 5528
rect 21300 5448 22388 5512
rect 22452 5448 22472 5512
rect 21300 5432 22472 5448
rect 21300 5368 22388 5432
rect 22452 5368 22472 5432
rect 21300 5352 22472 5368
rect 21300 5288 22388 5352
rect 22452 5288 22472 5352
rect 21300 5272 22472 5288
rect 21300 5208 22388 5272
rect 22452 5208 22472 5272
rect 21300 5160 22472 5208
rect 22712 5992 23884 6040
rect 22712 5928 23800 5992
rect 23864 5928 23884 5992
rect 22712 5912 23884 5928
rect 22712 5848 23800 5912
rect 23864 5848 23884 5912
rect 22712 5832 23884 5848
rect 22712 5768 23800 5832
rect 23864 5768 23884 5832
rect 22712 5752 23884 5768
rect 22712 5688 23800 5752
rect 23864 5688 23884 5752
rect 22712 5672 23884 5688
rect 22712 5608 23800 5672
rect 23864 5608 23884 5672
rect 22712 5592 23884 5608
rect 22712 5528 23800 5592
rect 23864 5528 23884 5592
rect 22712 5512 23884 5528
rect 22712 5448 23800 5512
rect 23864 5448 23884 5512
rect 22712 5432 23884 5448
rect 22712 5368 23800 5432
rect 23864 5368 23884 5432
rect 22712 5352 23884 5368
rect 22712 5288 23800 5352
rect 23864 5288 23884 5352
rect 22712 5272 23884 5288
rect 22712 5208 23800 5272
rect 23864 5208 23884 5272
rect 22712 5160 23884 5208
rect -23884 4872 -22712 4920
rect -23884 4808 -22796 4872
rect -22732 4808 -22712 4872
rect -23884 4792 -22712 4808
rect -23884 4728 -22796 4792
rect -22732 4728 -22712 4792
rect -23884 4712 -22712 4728
rect -23884 4648 -22796 4712
rect -22732 4648 -22712 4712
rect -23884 4632 -22712 4648
rect -23884 4568 -22796 4632
rect -22732 4568 -22712 4632
rect -23884 4552 -22712 4568
rect -23884 4488 -22796 4552
rect -22732 4488 -22712 4552
rect -23884 4472 -22712 4488
rect -23884 4408 -22796 4472
rect -22732 4408 -22712 4472
rect -23884 4392 -22712 4408
rect -23884 4328 -22796 4392
rect -22732 4328 -22712 4392
rect -23884 4312 -22712 4328
rect -23884 4248 -22796 4312
rect -22732 4248 -22712 4312
rect -23884 4232 -22712 4248
rect -23884 4168 -22796 4232
rect -22732 4168 -22712 4232
rect -23884 4152 -22712 4168
rect -23884 4088 -22796 4152
rect -22732 4088 -22712 4152
rect -23884 4040 -22712 4088
rect -22472 4872 -21300 4920
rect -22472 4808 -21384 4872
rect -21320 4808 -21300 4872
rect -22472 4792 -21300 4808
rect -22472 4728 -21384 4792
rect -21320 4728 -21300 4792
rect -22472 4712 -21300 4728
rect -22472 4648 -21384 4712
rect -21320 4648 -21300 4712
rect -22472 4632 -21300 4648
rect -22472 4568 -21384 4632
rect -21320 4568 -21300 4632
rect -22472 4552 -21300 4568
rect -22472 4488 -21384 4552
rect -21320 4488 -21300 4552
rect -22472 4472 -21300 4488
rect -22472 4408 -21384 4472
rect -21320 4408 -21300 4472
rect -22472 4392 -21300 4408
rect -22472 4328 -21384 4392
rect -21320 4328 -21300 4392
rect -22472 4312 -21300 4328
rect -22472 4248 -21384 4312
rect -21320 4248 -21300 4312
rect -22472 4232 -21300 4248
rect -22472 4168 -21384 4232
rect -21320 4168 -21300 4232
rect -22472 4152 -21300 4168
rect -22472 4088 -21384 4152
rect -21320 4088 -21300 4152
rect -22472 4040 -21300 4088
rect -21060 4872 -19888 4920
rect -21060 4808 -19972 4872
rect -19908 4808 -19888 4872
rect -21060 4792 -19888 4808
rect -21060 4728 -19972 4792
rect -19908 4728 -19888 4792
rect -21060 4712 -19888 4728
rect -21060 4648 -19972 4712
rect -19908 4648 -19888 4712
rect -21060 4632 -19888 4648
rect -21060 4568 -19972 4632
rect -19908 4568 -19888 4632
rect -21060 4552 -19888 4568
rect -21060 4488 -19972 4552
rect -19908 4488 -19888 4552
rect -21060 4472 -19888 4488
rect -21060 4408 -19972 4472
rect -19908 4408 -19888 4472
rect -21060 4392 -19888 4408
rect -21060 4328 -19972 4392
rect -19908 4328 -19888 4392
rect -21060 4312 -19888 4328
rect -21060 4248 -19972 4312
rect -19908 4248 -19888 4312
rect -21060 4232 -19888 4248
rect -21060 4168 -19972 4232
rect -19908 4168 -19888 4232
rect -21060 4152 -19888 4168
rect -21060 4088 -19972 4152
rect -19908 4088 -19888 4152
rect -21060 4040 -19888 4088
rect -19648 4872 -18476 4920
rect -19648 4808 -18560 4872
rect -18496 4808 -18476 4872
rect -19648 4792 -18476 4808
rect -19648 4728 -18560 4792
rect -18496 4728 -18476 4792
rect -19648 4712 -18476 4728
rect -19648 4648 -18560 4712
rect -18496 4648 -18476 4712
rect -19648 4632 -18476 4648
rect -19648 4568 -18560 4632
rect -18496 4568 -18476 4632
rect -19648 4552 -18476 4568
rect -19648 4488 -18560 4552
rect -18496 4488 -18476 4552
rect -19648 4472 -18476 4488
rect -19648 4408 -18560 4472
rect -18496 4408 -18476 4472
rect -19648 4392 -18476 4408
rect -19648 4328 -18560 4392
rect -18496 4328 -18476 4392
rect -19648 4312 -18476 4328
rect -19648 4248 -18560 4312
rect -18496 4248 -18476 4312
rect -19648 4232 -18476 4248
rect -19648 4168 -18560 4232
rect -18496 4168 -18476 4232
rect -19648 4152 -18476 4168
rect -19648 4088 -18560 4152
rect -18496 4088 -18476 4152
rect -19648 4040 -18476 4088
rect -18236 4872 -17064 4920
rect -18236 4808 -17148 4872
rect -17084 4808 -17064 4872
rect -18236 4792 -17064 4808
rect -18236 4728 -17148 4792
rect -17084 4728 -17064 4792
rect -18236 4712 -17064 4728
rect -18236 4648 -17148 4712
rect -17084 4648 -17064 4712
rect -18236 4632 -17064 4648
rect -18236 4568 -17148 4632
rect -17084 4568 -17064 4632
rect -18236 4552 -17064 4568
rect -18236 4488 -17148 4552
rect -17084 4488 -17064 4552
rect -18236 4472 -17064 4488
rect -18236 4408 -17148 4472
rect -17084 4408 -17064 4472
rect -18236 4392 -17064 4408
rect -18236 4328 -17148 4392
rect -17084 4328 -17064 4392
rect -18236 4312 -17064 4328
rect -18236 4248 -17148 4312
rect -17084 4248 -17064 4312
rect -18236 4232 -17064 4248
rect -18236 4168 -17148 4232
rect -17084 4168 -17064 4232
rect -18236 4152 -17064 4168
rect -18236 4088 -17148 4152
rect -17084 4088 -17064 4152
rect -18236 4040 -17064 4088
rect -16824 4872 -15652 4920
rect -16824 4808 -15736 4872
rect -15672 4808 -15652 4872
rect -16824 4792 -15652 4808
rect -16824 4728 -15736 4792
rect -15672 4728 -15652 4792
rect -16824 4712 -15652 4728
rect -16824 4648 -15736 4712
rect -15672 4648 -15652 4712
rect -16824 4632 -15652 4648
rect -16824 4568 -15736 4632
rect -15672 4568 -15652 4632
rect -16824 4552 -15652 4568
rect -16824 4488 -15736 4552
rect -15672 4488 -15652 4552
rect -16824 4472 -15652 4488
rect -16824 4408 -15736 4472
rect -15672 4408 -15652 4472
rect -16824 4392 -15652 4408
rect -16824 4328 -15736 4392
rect -15672 4328 -15652 4392
rect -16824 4312 -15652 4328
rect -16824 4248 -15736 4312
rect -15672 4248 -15652 4312
rect -16824 4232 -15652 4248
rect -16824 4168 -15736 4232
rect -15672 4168 -15652 4232
rect -16824 4152 -15652 4168
rect -16824 4088 -15736 4152
rect -15672 4088 -15652 4152
rect -16824 4040 -15652 4088
rect -15412 4872 -14240 4920
rect -15412 4808 -14324 4872
rect -14260 4808 -14240 4872
rect -15412 4792 -14240 4808
rect -15412 4728 -14324 4792
rect -14260 4728 -14240 4792
rect -15412 4712 -14240 4728
rect -15412 4648 -14324 4712
rect -14260 4648 -14240 4712
rect -15412 4632 -14240 4648
rect -15412 4568 -14324 4632
rect -14260 4568 -14240 4632
rect -15412 4552 -14240 4568
rect -15412 4488 -14324 4552
rect -14260 4488 -14240 4552
rect -15412 4472 -14240 4488
rect -15412 4408 -14324 4472
rect -14260 4408 -14240 4472
rect -15412 4392 -14240 4408
rect -15412 4328 -14324 4392
rect -14260 4328 -14240 4392
rect -15412 4312 -14240 4328
rect -15412 4248 -14324 4312
rect -14260 4248 -14240 4312
rect -15412 4232 -14240 4248
rect -15412 4168 -14324 4232
rect -14260 4168 -14240 4232
rect -15412 4152 -14240 4168
rect -15412 4088 -14324 4152
rect -14260 4088 -14240 4152
rect -15412 4040 -14240 4088
rect -14000 4872 -12828 4920
rect -14000 4808 -12912 4872
rect -12848 4808 -12828 4872
rect -14000 4792 -12828 4808
rect -14000 4728 -12912 4792
rect -12848 4728 -12828 4792
rect -14000 4712 -12828 4728
rect -14000 4648 -12912 4712
rect -12848 4648 -12828 4712
rect -14000 4632 -12828 4648
rect -14000 4568 -12912 4632
rect -12848 4568 -12828 4632
rect -14000 4552 -12828 4568
rect -14000 4488 -12912 4552
rect -12848 4488 -12828 4552
rect -14000 4472 -12828 4488
rect -14000 4408 -12912 4472
rect -12848 4408 -12828 4472
rect -14000 4392 -12828 4408
rect -14000 4328 -12912 4392
rect -12848 4328 -12828 4392
rect -14000 4312 -12828 4328
rect -14000 4248 -12912 4312
rect -12848 4248 -12828 4312
rect -14000 4232 -12828 4248
rect -14000 4168 -12912 4232
rect -12848 4168 -12828 4232
rect -14000 4152 -12828 4168
rect -14000 4088 -12912 4152
rect -12848 4088 -12828 4152
rect -14000 4040 -12828 4088
rect -12588 4872 -11416 4920
rect -12588 4808 -11500 4872
rect -11436 4808 -11416 4872
rect -12588 4792 -11416 4808
rect -12588 4728 -11500 4792
rect -11436 4728 -11416 4792
rect -12588 4712 -11416 4728
rect -12588 4648 -11500 4712
rect -11436 4648 -11416 4712
rect -12588 4632 -11416 4648
rect -12588 4568 -11500 4632
rect -11436 4568 -11416 4632
rect -12588 4552 -11416 4568
rect -12588 4488 -11500 4552
rect -11436 4488 -11416 4552
rect -12588 4472 -11416 4488
rect -12588 4408 -11500 4472
rect -11436 4408 -11416 4472
rect -12588 4392 -11416 4408
rect -12588 4328 -11500 4392
rect -11436 4328 -11416 4392
rect -12588 4312 -11416 4328
rect -12588 4248 -11500 4312
rect -11436 4248 -11416 4312
rect -12588 4232 -11416 4248
rect -12588 4168 -11500 4232
rect -11436 4168 -11416 4232
rect -12588 4152 -11416 4168
rect -12588 4088 -11500 4152
rect -11436 4088 -11416 4152
rect -12588 4040 -11416 4088
rect -11176 4872 -10004 4920
rect -11176 4808 -10088 4872
rect -10024 4808 -10004 4872
rect -11176 4792 -10004 4808
rect -11176 4728 -10088 4792
rect -10024 4728 -10004 4792
rect -11176 4712 -10004 4728
rect -11176 4648 -10088 4712
rect -10024 4648 -10004 4712
rect -11176 4632 -10004 4648
rect -11176 4568 -10088 4632
rect -10024 4568 -10004 4632
rect -11176 4552 -10004 4568
rect -11176 4488 -10088 4552
rect -10024 4488 -10004 4552
rect -11176 4472 -10004 4488
rect -11176 4408 -10088 4472
rect -10024 4408 -10004 4472
rect -11176 4392 -10004 4408
rect -11176 4328 -10088 4392
rect -10024 4328 -10004 4392
rect -11176 4312 -10004 4328
rect -11176 4248 -10088 4312
rect -10024 4248 -10004 4312
rect -11176 4232 -10004 4248
rect -11176 4168 -10088 4232
rect -10024 4168 -10004 4232
rect -11176 4152 -10004 4168
rect -11176 4088 -10088 4152
rect -10024 4088 -10004 4152
rect -11176 4040 -10004 4088
rect -9764 4872 -8592 4920
rect -9764 4808 -8676 4872
rect -8612 4808 -8592 4872
rect -9764 4792 -8592 4808
rect -9764 4728 -8676 4792
rect -8612 4728 -8592 4792
rect -9764 4712 -8592 4728
rect -9764 4648 -8676 4712
rect -8612 4648 -8592 4712
rect -9764 4632 -8592 4648
rect -9764 4568 -8676 4632
rect -8612 4568 -8592 4632
rect -9764 4552 -8592 4568
rect -9764 4488 -8676 4552
rect -8612 4488 -8592 4552
rect -9764 4472 -8592 4488
rect -9764 4408 -8676 4472
rect -8612 4408 -8592 4472
rect -9764 4392 -8592 4408
rect -9764 4328 -8676 4392
rect -8612 4328 -8592 4392
rect -9764 4312 -8592 4328
rect -9764 4248 -8676 4312
rect -8612 4248 -8592 4312
rect -9764 4232 -8592 4248
rect -9764 4168 -8676 4232
rect -8612 4168 -8592 4232
rect -9764 4152 -8592 4168
rect -9764 4088 -8676 4152
rect -8612 4088 -8592 4152
rect -9764 4040 -8592 4088
rect -8352 4872 -7180 4920
rect -8352 4808 -7264 4872
rect -7200 4808 -7180 4872
rect -8352 4792 -7180 4808
rect -8352 4728 -7264 4792
rect -7200 4728 -7180 4792
rect -8352 4712 -7180 4728
rect -8352 4648 -7264 4712
rect -7200 4648 -7180 4712
rect -8352 4632 -7180 4648
rect -8352 4568 -7264 4632
rect -7200 4568 -7180 4632
rect -8352 4552 -7180 4568
rect -8352 4488 -7264 4552
rect -7200 4488 -7180 4552
rect -8352 4472 -7180 4488
rect -8352 4408 -7264 4472
rect -7200 4408 -7180 4472
rect -8352 4392 -7180 4408
rect -8352 4328 -7264 4392
rect -7200 4328 -7180 4392
rect -8352 4312 -7180 4328
rect -8352 4248 -7264 4312
rect -7200 4248 -7180 4312
rect -8352 4232 -7180 4248
rect -8352 4168 -7264 4232
rect -7200 4168 -7180 4232
rect -8352 4152 -7180 4168
rect -8352 4088 -7264 4152
rect -7200 4088 -7180 4152
rect -8352 4040 -7180 4088
rect -6940 4872 -5768 4920
rect -6940 4808 -5852 4872
rect -5788 4808 -5768 4872
rect -6940 4792 -5768 4808
rect -6940 4728 -5852 4792
rect -5788 4728 -5768 4792
rect -6940 4712 -5768 4728
rect -6940 4648 -5852 4712
rect -5788 4648 -5768 4712
rect -6940 4632 -5768 4648
rect -6940 4568 -5852 4632
rect -5788 4568 -5768 4632
rect -6940 4552 -5768 4568
rect -6940 4488 -5852 4552
rect -5788 4488 -5768 4552
rect -6940 4472 -5768 4488
rect -6940 4408 -5852 4472
rect -5788 4408 -5768 4472
rect -6940 4392 -5768 4408
rect -6940 4328 -5852 4392
rect -5788 4328 -5768 4392
rect -6940 4312 -5768 4328
rect -6940 4248 -5852 4312
rect -5788 4248 -5768 4312
rect -6940 4232 -5768 4248
rect -6940 4168 -5852 4232
rect -5788 4168 -5768 4232
rect -6940 4152 -5768 4168
rect -6940 4088 -5852 4152
rect -5788 4088 -5768 4152
rect -6940 4040 -5768 4088
rect -5528 4872 -4356 4920
rect -5528 4808 -4440 4872
rect -4376 4808 -4356 4872
rect -5528 4792 -4356 4808
rect -5528 4728 -4440 4792
rect -4376 4728 -4356 4792
rect -5528 4712 -4356 4728
rect -5528 4648 -4440 4712
rect -4376 4648 -4356 4712
rect -5528 4632 -4356 4648
rect -5528 4568 -4440 4632
rect -4376 4568 -4356 4632
rect -5528 4552 -4356 4568
rect -5528 4488 -4440 4552
rect -4376 4488 -4356 4552
rect -5528 4472 -4356 4488
rect -5528 4408 -4440 4472
rect -4376 4408 -4356 4472
rect -5528 4392 -4356 4408
rect -5528 4328 -4440 4392
rect -4376 4328 -4356 4392
rect -5528 4312 -4356 4328
rect -5528 4248 -4440 4312
rect -4376 4248 -4356 4312
rect -5528 4232 -4356 4248
rect -5528 4168 -4440 4232
rect -4376 4168 -4356 4232
rect -5528 4152 -4356 4168
rect -5528 4088 -4440 4152
rect -4376 4088 -4356 4152
rect -5528 4040 -4356 4088
rect -4116 4872 -2944 4920
rect -4116 4808 -3028 4872
rect -2964 4808 -2944 4872
rect -4116 4792 -2944 4808
rect -4116 4728 -3028 4792
rect -2964 4728 -2944 4792
rect -4116 4712 -2944 4728
rect -4116 4648 -3028 4712
rect -2964 4648 -2944 4712
rect -4116 4632 -2944 4648
rect -4116 4568 -3028 4632
rect -2964 4568 -2944 4632
rect -4116 4552 -2944 4568
rect -4116 4488 -3028 4552
rect -2964 4488 -2944 4552
rect -4116 4472 -2944 4488
rect -4116 4408 -3028 4472
rect -2964 4408 -2944 4472
rect -4116 4392 -2944 4408
rect -4116 4328 -3028 4392
rect -2964 4328 -2944 4392
rect -4116 4312 -2944 4328
rect -4116 4248 -3028 4312
rect -2964 4248 -2944 4312
rect -4116 4232 -2944 4248
rect -4116 4168 -3028 4232
rect -2964 4168 -2944 4232
rect -4116 4152 -2944 4168
rect -4116 4088 -3028 4152
rect -2964 4088 -2944 4152
rect -4116 4040 -2944 4088
rect -2704 4872 -1532 4920
rect -2704 4808 -1616 4872
rect -1552 4808 -1532 4872
rect -2704 4792 -1532 4808
rect -2704 4728 -1616 4792
rect -1552 4728 -1532 4792
rect -2704 4712 -1532 4728
rect -2704 4648 -1616 4712
rect -1552 4648 -1532 4712
rect -2704 4632 -1532 4648
rect -2704 4568 -1616 4632
rect -1552 4568 -1532 4632
rect -2704 4552 -1532 4568
rect -2704 4488 -1616 4552
rect -1552 4488 -1532 4552
rect -2704 4472 -1532 4488
rect -2704 4408 -1616 4472
rect -1552 4408 -1532 4472
rect -2704 4392 -1532 4408
rect -2704 4328 -1616 4392
rect -1552 4328 -1532 4392
rect -2704 4312 -1532 4328
rect -2704 4248 -1616 4312
rect -1552 4248 -1532 4312
rect -2704 4232 -1532 4248
rect -2704 4168 -1616 4232
rect -1552 4168 -1532 4232
rect -2704 4152 -1532 4168
rect -2704 4088 -1616 4152
rect -1552 4088 -1532 4152
rect -2704 4040 -1532 4088
rect -1292 4872 -120 4920
rect -1292 4808 -204 4872
rect -140 4808 -120 4872
rect -1292 4792 -120 4808
rect -1292 4728 -204 4792
rect -140 4728 -120 4792
rect -1292 4712 -120 4728
rect -1292 4648 -204 4712
rect -140 4648 -120 4712
rect -1292 4632 -120 4648
rect -1292 4568 -204 4632
rect -140 4568 -120 4632
rect -1292 4552 -120 4568
rect -1292 4488 -204 4552
rect -140 4488 -120 4552
rect -1292 4472 -120 4488
rect -1292 4408 -204 4472
rect -140 4408 -120 4472
rect -1292 4392 -120 4408
rect -1292 4328 -204 4392
rect -140 4328 -120 4392
rect -1292 4312 -120 4328
rect -1292 4248 -204 4312
rect -140 4248 -120 4312
rect -1292 4232 -120 4248
rect -1292 4168 -204 4232
rect -140 4168 -120 4232
rect -1292 4152 -120 4168
rect -1292 4088 -204 4152
rect -140 4088 -120 4152
rect -1292 4040 -120 4088
rect 120 4872 1292 4920
rect 120 4808 1208 4872
rect 1272 4808 1292 4872
rect 120 4792 1292 4808
rect 120 4728 1208 4792
rect 1272 4728 1292 4792
rect 120 4712 1292 4728
rect 120 4648 1208 4712
rect 1272 4648 1292 4712
rect 120 4632 1292 4648
rect 120 4568 1208 4632
rect 1272 4568 1292 4632
rect 120 4552 1292 4568
rect 120 4488 1208 4552
rect 1272 4488 1292 4552
rect 120 4472 1292 4488
rect 120 4408 1208 4472
rect 1272 4408 1292 4472
rect 120 4392 1292 4408
rect 120 4328 1208 4392
rect 1272 4328 1292 4392
rect 120 4312 1292 4328
rect 120 4248 1208 4312
rect 1272 4248 1292 4312
rect 120 4232 1292 4248
rect 120 4168 1208 4232
rect 1272 4168 1292 4232
rect 120 4152 1292 4168
rect 120 4088 1208 4152
rect 1272 4088 1292 4152
rect 120 4040 1292 4088
rect 1532 4872 2704 4920
rect 1532 4808 2620 4872
rect 2684 4808 2704 4872
rect 1532 4792 2704 4808
rect 1532 4728 2620 4792
rect 2684 4728 2704 4792
rect 1532 4712 2704 4728
rect 1532 4648 2620 4712
rect 2684 4648 2704 4712
rect 1532 4632 2704 4648
rect 1532 4568 2620 4632
rect 2684 4568 2704 4632
rect 1532 4552 2704 4568
rect 1532 4488 2620 4552
rect 2684 4488 2704 4552
rect 1532 4472 2704 4488
rect 1532 4408 2620 4472
rect 2684 4408 2704 4472
rect 1532 4392 2704 4408
rect 1532 4328 2620 4392
rect 2684 4328 2704 4392
rect 1532 4312 2704 4328
rect 1532 4248 2620 4312
rect 2684 4248 2704 4312
rect 1532 4232 2704 4248
rect 1532 4168 2620 4232
rect 2684 4168 2704 4232
rect 1532 4152 2704 4168
rect 1532 4088 2620 4152
rect 2684 4088 2704 4152
rect 1532 4040 2704 4088
rect 2944 4872 4116 4920
rect 2944 4808 4032 4872
rect 4096 4808 4116 4872
rect 2944 4792 4116 4808
rect 2944 4728 4032 4792
rect 4096 4728 4116 4792
rect 2944 4712 4116 4728
rect 2944 4648 4032 4712
rect 4096 4648 4116 4712
rect 2944 4632 4116 4648
rect 2944 4568 4032 4632
rect 4096 4568 4116 4632
rect 2944 4552 4116 4568
rect 2944 4488 4032 4552
rect 4096 4488 4116 4552
rect 2944 4472 4116 4488
rect 2944 4408 4032 4472
rect 4096 4408 4116 4472
rect 2944 4392 4116 4408
rect 2944 4328 4032 4392
rect 4096 4328 4116 4392
rect 2944 4312 4116 4328
rect 2944 4248 4032 4312
rect 4096 4248 4116 4312
rect 2944 4232 4116 4248
rect 2944 4168 4032 4232
rect 4096 4168 4116 4232
rect 2944 4152 4116 4168
rect 2944 4088 4032 4152
rect 4096 4088 4116 4152
rect 2944 4040 4116 4088
rect 4356 4872 5528 4920
rect 4356 4808 5444 4872
rect 5508 4808 5528 4872
rect 4356 4792 5528 4808
rect 4356 4728 5444 4792
rect 5508 4728 5528 4792
rect 4356 4712 5528 4728
rect 4356 4648 5444 4712
rect 5508 4648 5528 4712
rect 4356 4632 5528 4648
rect 4356 4568 5444 4632
rect 5508 4568 5528 4632
rect 4356 4552 5528 4568
rect 4356 4488 5444 4552
rect 5508 4488 5528 4552
rect 4356 4472 5528 4488
rect 4356 4408 5444 4472
rect 5508 4408 5528 4472
rect 4356 4392 5528 4408
rect 4356 4328 5444 4392
rect 5508 4328 5528 4392
rect 4356 4312 5528 4328
rect 4356 4248 5444 4312
rect 5508 4248 5528 4312
rect 4356 4232 5528 4248
rect 4356 4168 5444 4232
rect 5508 4168 5528 4232
rect 4356 4152 5528 4168
rect 4356 4088 5444 4152
rect 5508 4088 5528 4152
rect 4356 4040 5528 4088
rect 5768 4872 6940 4920
rect 5768 4808 6856 4872
rect 6920 4808 6940 4872
rect 5768 4792 6940 4808
rect 5768 4728 6856 4792
rect 6920 4728 6940 4792
rect 5768 4712 6940 4728
rect 5768 4648 6856 4712
rect 6920 4648 6940 4712
rect 5768 4632 6940 4648
rect 5768 4568 6856 4632
rect 6920 4568 6940 4632
rect 5768 4552 6940 4568
rect 5768 4488 6856 4552
rect 6920 4488 6940 4552
rect 5768 4472 6940 4488
rect 5768 4408 6856 4472
rect 6920 4408 6940 4472
rect 5768 4392 6940 4408
rect 5768 4328 6856 4392
rect 6920 4328 6940 4392
rect 5768 4312 6940 4328
rect 5768 4248 6856 4312
rect 6920 4248 6940 4312
rect 5768 4232 6940 4248
rect 5768 4168 6856 4232
rect 6920 4168 6940 4232
rect 5768 4152 6940 4168
rect 5768 4088 6856 4152
rect 6920 4088 6940 4152
rect 5768 4040 6940 4088
rect 7180 4872 8352 4920
rect 7180 4808 8268 4872
rect 8332 4808 8352 4872
rect 7180 4792 8352 4808
rect 7180 4728 8268 4792
rect 8332 4728 8352 4792
rect 7180 4712 8352 4728
rect 7180 4648 8268 4712
rect 8332 4648 8352 4712
rect 7180 4632 8352 4648
rect 7180 4568 8268 4632
rect 8332 4568 8352 4632
rect 7180 4552 8352 4568
rect 7180 4488 8268 4552
rect 8332 4488 8352 4552
rect 7180 4472 8352 4488
rect 7180 4408 8268 4472
rect 8332 4408 8352 4472
rect 7180 4392 8352 4408
rect 7180 4328 8268 4392
rect 8332 4328 8352 4392
rect 7180 4312 8352 4328
rect 7180 4248 8268 4312
rect 8332 4248 8352 4312
rect 7180 4232 8352 4248
rect 7180 4168 8268 4232
rect 8332 4168 8352 4232
rect 7180 4152 8352 4168
rect 7180 4088 8268 4152
rect 8332 4088 8352 4152
rect 7180 4040 8352 4088
rect 8592 4872 9764 4920
rect 8592 4808 9680 4872
rect 9744 4808 9764 4872
rect 8592 4792 9764 4808
rect 8592 4728 9680 4792
rect 9744 4728 9764 4792
rect 8592 4712 9764 4728
rect 8592 4648 9680 4712
rect 9744 4648 9764 4712
rect 8592 4632 9764 4648
rect 8592 4568 9680 4632
rect 9744 4568 9764 4632
rect 8592 4552 9764 4568
rect 8592 4488 9680 4552
rect 9744 4488 9764 4552
rect 8592 4472 9764 4488
rect 8592 4408 9680 4472
rect 9744 4408 9764 4472
rect 8592 4392 9764 4408
rect 8592 4328 9680 4392
rect 9744 4328 9764 4392
rect 8592 4312 9764 4328
rect 8592 4248 9680 4312
rect 9744 4248 9764 4312
rect 8592 4232 9764 4248
rect 8592 4168 9680 4232
rect 9744 4168 9764 4232
rect 8592 4152 9764 4168
rect 8592 4088 9680 4152
rect 9744 4088 9764 4152
rect 8592 4040 9764 4088
rect 10004 4872 11176 4920
rect 10004 4808 11092 4872
rect 11156 4808 11176 4872
rect 10004 4792 11176 4808
rect 10004 4728 11092 4792
rect 11156 4728 11176 4792
rect 10004 4712 11176 4728
rect 10004 4648 11092 4712
rect 11156 4648 11176 4712
rect 10004 4632 11176 4648
rect 10004 4568 11092 4632
rect 11156 4568 11176 4632
rect 10004 4552 11176 4568
rect 10004 4488 11092 4552
rect 11156 4488 11176 4552
rect 10004 4472 11176 4488
rect 10004 4408 11092 4472
rect 11156 4408 11176 4472
rect 10004 4392 11176 4408
rect 10004 4328 11092 4392
rect 11156 4328 11176 4392
rect 10004 4312 11176 4328
rect 10004 4248 11092 4312
rect 11156 4248 11176 4312
rect 10004 4232 11176 4248
rect 10004 4168 11092 4232
rect 11156 4168 11176 4232
rect 10004 4152 11176 4168
rect 10004 4088 11092 4152
rect 11156 4088 11176 4152
rect 10004 4040 11176 4088
rect 11416 4872 12588 4920
rect 11416 4808 12504 4872
rect 12568 4808 12588 4872
rect 11416 4792 12588 4808
rect 11416 4728 12504 4792
rect 12568 4728 12588 4792
rect 11416 4712 12588 4728
rect 11416 4648 12504 4712
rect 12568 4648 12588 4712
rect 11416 4632 12588 4648
rect 11416 4568 12504 4632
rect 12568 4568 12588 4632
rect 11416 4552 12588 4568
rect 11416 4488 12504 4552
rect 12568 4488 12588 4552
rect 11416 4472 12588 4488
rect 11416 4408 12504 4472
rect 12568 4408 12588 4472
rect 11416 4392 12588 4408
rect 11416 4328 12504 4392
rect 12568 4328 12588 4392
rect 11416 4312 12588 4328
rect 11416 4248 12504 4312
rect 12568 4248 12588 4312
rect 11416 4232 12588 4248
rect 11416 4168 12504 4232
rect 12568 4168 12588 4232
rect 11416 4152 12588 4168
rect 11416 4088 12504 4152
rect 12568 4088 12588 4152
rect 11416 4040 12588 4088
rect 12828 4872 14000 4920
rect 12828 4808 13916 4872
rect 13980 4808 14000 4872
rect 12828 4792 14000 4808
rect 12828 4728 13916 4792
rect 13980 4728 14000 4792
rect 12828 4712 14000 4728
rect 12828 4648 13916 4712
rect 13980 4648 14000 4712
rect 12828 4632 14000 4648
rect 12828 4568 13916 4632
rect 13980 4568 14000 4632
rect 12828 4552 14000 4568
rect 12828 4488 13916 4552
rect 13980 4488 14000 4552
rect 12828 4472 14000 4488
rect 12828 4408 13916 4472
rect 13980 4408 14000 4472
rect 12828 4392 14000 4408
rect 12828 4328 13916 4392
rect 13980 4328 14000 4392
rect 12828 4312 14000 4328
rect 12828 4248 13916 4312
rect 13980 4248 14000 4312
rect 12828 4232 14000 4248
rect 12828 4168 13916 4232
rect 13980 4168 14000 4232
rect 12828 4152 14000 4168
rect 12828 4088 13916 4152
rect 13980 4088 14000 4152
rect 12828 4040 14000 4088
rect 14240 4872 15412 4920
rect 14240 4808 15328 4872
rect 15392 4808 15412 4872
rect 14240 4792 15412 4808
rect 14240 4728 15328 4792
rect 15392 4728 15412 4792
rect 14240 4712 15412 4728
rect 14240 4648 15328 4712
rect 15392 4648 15412 4712
rect 14240 4632 15412 4648
rect 14240 4568 15328 4632
rect 15392 4568 15412 4632
rect 14240 4552 15412 4568
rect 14240 4488 15328 4552
rect 15392 4488 15412 4552
rect 14240 4472 15412 4488
rect 14240 4408 15328 4472
rect 15392 4408 15412 4472
rect 14240 4392 15412 4408
rect 14240 4328 15328 4392
rect 15392 4328 15412 4392
rect 14240 4312 15412 4328
rect 14240 4248 15328 4312
rect 15392 4248 15412 4312
rect 14240 4232 15412 4248
rect 14240 4168 15328 4232
rect 15392 4168 15412 4232
rect 14240 4152 15412 4168
rect 14240 4088 15328 4152
rect 15392 4088 15412 4152
rect 14240 4040 15412 4088
rect 15652 4872 16824 4920
rect 15652 4808 16740 4872
rect 16804 4808 16824 4872
rect 15652 4792 16824 4808
rect 15652 4728 16740 4792
rect 16804 4728 16824 4792
rect 15652 4712 16824 4728
rect 15652 4648 16740 4712
rect 16804 4648 16824 4712
rect 15652 4632 16824 4648
rect 15652 4568 16740 4632
rect 16804 4568 16824 4632
rect 15652 4552 16824 4568
rect 15652 4488 16740 4552
rect 16804 4488 16824 4552
rect 15652 4472 16824 4488
rect 15652 4408 16740 4472
rect 16804 4408 16824 4472
rect 15652 4392 16824 4408
rect 15652 4328 16740 4392
rect 16804 4328 16824 4392
rect 15652 4312 16824 4328
rect 15652 4248 16740 4312
rect 16804 4248 16824 4312
rect 15652 4232 16824 4248
rect 15652 4168 16740 4232
rect 16804 4168 16824 4232
rect 15652 4152 16824 4168
rect 15652 4088 16740 4152
rect 16804 4088 16824 4152
rect 15652 4040 16824 4088
rect 17064 4872 18236 4920
rect 17064 4808 18152 4872
rect 18216 4808 18236 4872
rect 17064 4792 18236 4808
rect 17064 4728 18152 4792
rect 18216 4728 18236 4792
rect 17064 4712 18236 4728
rect 17064 4648 18152 4712
rect 18216 4648 18236 4712
rect 17064 4632 18236 4648
rect 17064 4568 18152 4632
rect 18216 4568 18236 4632
rect 17064 4552 18236 4568
rect 17064 4488 18152 4552
rect 18216 4488 18236 4552
rect 17064 4472 18236 4488
rect 17064 4408 18152 4472
rect 18216 4408 18236 4472
rect 17064 4392 18236 4408
rect 17064 4328 18152 4392
rect 18216 4328 18236 4392
rect 17064 4312 18236 4328
rect 17064 4248 18152 4312
rect 18216 4248 18236 4312
rect 17064 4232 18236 4248
rect 17064 4168 18152 4232
rect 18216 4168 18236 4232
rect 17064 4152 18236 4168
rect 17064 4088 18152 4152
rect 18216 4088 18236 4152
rect 17064 4040 18236 4088
rect 18476 4872 19648 4920
rect 18476 4808 19564 4872
rect 19628 4808 19648 4872
rect 18476 4792 19648 4808
rect 18476 4728 19564 4792
rect 19628 4728 19648 4792
rect 18476 4712 19648 4728
rect 18476 4648 19564 4712
rect 19628 4648 19648 4712
rect 18476 4632 19648 4648
rect 18476 4568 19564 4632
rect 19628 4568 19648 4632
rect 18476 4552 19648 4568
rect 18476 4488 19564 4552
rect 19628 4488 19648 4552
rect 18476 4472 19648 4488
rect 18476 4408 19564 4472
rect 19628 4408 19648 4472
rect 18476 4392 19648 4408
rect 18476 4328 19564 4392
rect 19628 4328 19648 4392
rect 18476 4312 19648 4328
rect 18476 4248 19564 4312
rect 19628 4248 19648 4312
rect 18476 4232 19648 4248
rect 18476 4168 19564 4232
rect 19628 4168 19648 4232
rect 18476 4152 19648 4168
rect 18476 4088 19564 4152
rect 19628 4088 19648 4152
rect 18476 4040 19648 4088
rect 19888 4872 21060 4920
rect 19888 4808 20976 4872
rect 21040 4808 21060 4872
rect 19888 4792 21060 4808
rect 19888 4728 20976 4792
rect 21040 4728 21060 4792
rect 19888 4712 21060 4728
rect 19888 4648 20976 4712
rect 21040 4648 21060 4712
rect 19888 4632 21060 4648
rect 19888 4568 20976 4632
rect 21040 4568 21060 4632
rect 19888 4552 21060 4568
rect 19888 4488 20976 4552
rect 21040 4488 21060 4552
rect 19888 4472 21060 4488
rect 19888 4408 20976 4472
rect 21040 4408 21060 4472
rect 19888 4392 21060 4408
rect 19888 4328 20976 4392
rect 21040 4328 21060 4392
rect 19888 4312 21060 4328
rect 19888 4248 20976 4312
rect 21040 4248 21060 4312
rect 19888 4232 21060 4248
rect 19888 4168 20976 4232
rect 21040 4168 21060 4232
rect 19888 4152 21060 4168
rect 19888 4088 20976 4152
rect 21040 4088 21060 4152
rect 19888 4040 21060 4088
rect 21300 4872 22472 4920
rect 21300 4808 22388 4872
rect 22452 4808 22472 4872
rect 21300 4792 22472 4808
rect 21300 4728 22388 4792
rect 22452 4728 22472 4792
rect 21300 4712 22472 4728
rect 21300 4648 22388 4712
rect 22452 4648 22472 4712
rect 21300 4632 22472 4648
rect 21300 4568 22388 4632
rect 22452 4568 22472 4632
rect 21300 4552 22472 4568
rect 21300 4488 22388 4552
rect 22452 4488 22472 4552
rect 21300 4472 22472 4488
rect 21300 4408 22388 4472
rect 22452 4408 22472 4472
rect 21300 4392 22472 4408
rect 21300 4328 22388 4392
rect 22452 4328 22472 4392
rect 21300 4312 22472 4328
rect 21300 4248 22388 4312
rect 22452 4248 22472 4312
rect 21300 4232 22472 4248
rect 21300 4168 22388 4232
rect 22452 4168 22472 4232
rect 21300 4152 22472 4168
rect 21300 4088 22388 4152
rect 22452 4088 22472 4152
rect 21300 4040 22472 4088
rect 22712 4872 23884 4920
rect 22712 4808 23800 4872
rect 23864 4808 23884 4872
rect 22712 4792 23884 4808
rect 22712 4728 23800 4792
rect 23864 4728 23884 4792
rect 22712 4712 23884 4728
rect 22712 4648 23800 4712
rect 23864 4648 23884 4712
rect 22712 4632 23884 4648
rect 22712 4568 23800 4632
rect 23864 4568 23884 4632
rect 22712 4552 23884 4568
rect 22712 4488 23800 4552
rect 23864 4488 23884 4552
rect 22712 4472 23884 4488
rect 22712 4408 23800 4472
rect 23864 4408 23884 4472
rect 22712 4392 23884 4408
rect 22712 4328 23800 4392
rect 23864 4328 23884 4392
rect 22712 4312 23884 4328
rect 22712 4248 23800 4312
rect 23864 4248 23884 4312
rect 22712 4232 23884 4248
rect 22712 4168 23800 4232
rect 23864 4168 23884 4232
rect 22712 4152 23884 4168
rect 22712 4088 23800 4152
rect 23864 4088 23884 4152
rect 22712 4040 23884 4088
rect -23884 3752 -22712 3800
rect -23884 3688 -22796 3752
rect -22732 3688 -22712 3752
rect -23884 3672 -22712 3688
rect -23884 3608 -22796 3672
rect -22732 3608 -22712 3672
rect -23884 3592 -22712 3608
rect -23884 3528 -22796 3592
rect -22732 3528 -22712 3592
rect -23884 3512 -22712 3528
rect -23884 3448 -22796 3512
rect -22732 3448 -22712 3512
rect -23884 3432 -22712 3448
rect -23884 3368 -22796 3432
rect -22732 3368 -22712 3432
rect -23884 3352 -22712 3368
rect -23884 3288 -22796 3352
rect -22732 3288 -22712 3352
rect -23884 3272 -22712 3288
rect -23884 3208 -22796 3272
rect -22732 3208 -22712 3272
rect -23884 3192 -22712 3208
rect -23884 3128 -22796 3192
rect -22732 3128 -22712 3192
rect -23884 3112 -22712 3128
rect -23884 3048 -22796 3112
rect -22732 3048 -22712 3112
rect -23884 3032 -22712 3048
rect -23884 2968 -22796 3032
rect -22732 2968 -22712 3032
rect -23884 2920 -22712 2968
rect -22472 3752 -21300 3800
rect -22472 3688 -21384 3752
rect -21320 3688 -21300 3752
rect -22472 3672 -21300 3688
rect -22472 3608 -21384 3672
rect -21320 3608 -21300 3672
rect -22472 3592 -21300 3608
rect -22472 3528 -21384 3592
rect -21320 3528 -21300 3592
rect -22472 3512 -21300 3528
rect -22472 3448 -21384 3512
rect -21320 3448 -21300 3512
rect -22472 3432 -21300 3448
rect -22472 3368 -21384 3432
rect -21320 3368 -21300 3432
rect -22472 3352 -21300 3368
rect -22472 3288 -21384 3352
rect -21320 3288 -21300 3352
rect -22472 3272 -21300 3288
rect -22472 3208 -21384 3272
rect -21320 3208 -21300 3272
rect -22472 3192 -21300 3208
rect -22472 3128 -21384 3192
rect -21320 3128 -21300 3192
rect -22472 3112 -21300 3128
rect -22472 3048 -21384 3112
rect -21320 3048 -21300 3112
rect -22472 3032 -21300 3048
rect -22472 2968 -21384 3032
rect -21320 2968 -21300 3032
rect -22472 2920 -21300 2968
rect -21060 3752 -19888 3800
rect -21060 3688 -19972 3752
rect -19908 3688 -19888 3752
rect -21060 3672 -19888 3688
rect -21060 3608 -19972 3672
rect -19908 3608 -19888 3672
rect -21060 3592 -19888 3608
rect -21060 3528 -19972 3592
rect -19908 3528 -19888 3592
rect -21060 3512 -19888 3528
rect -21060 3448 -19972 3512
rect -19908 3448 -19888 3512
rect -21060 3432 -19888 3448
rect -21060 3368 -19972 3432
rect -19908 3368 -19888 3432
rect -21060 3352 -19888 3368
rect -21060 3288 -19972 3352
rect -19908 3288 -19888 3352
rect -21060 3272 -19888 3288
rect -21060 3208 -19972 3272
rect -19908 3208 -19888 3272
rect -21060 3192 -19888 3208
rect -21060 3128 -19972 3192
rect -19908 3128 -19888 3192
rect -21060 3112 -19888 3128
rect -21060 3048 -19972 3112
rect -19908 3048 -19888 3112
rect -21060 3032 -19888 3048
rect -21060 2968 -19972 3032
rect -19908 2968 -19888 3032
rect -21060 2920 -19888 2968
rect -19648 3752 -18476 3800
rect -19648 3688 -18560 3752
rect -18496 3688 -18476 3752
rect -19648 3672 -18476 3688
rect -19648 3608 -18560 3672
rect -18496 3608 -18476 3672
rect -19648 3592 -18476 3608
rect -19648 3528 -18560 3592
rect -18496 3528 -18476 3592
rect -19648 3512 -18476 3528
rect -19648 3448 -18560 3512
rect -18496 3448 -18476 3512
rect -19648 3432 -18476 3448
rect -19648 3368 -18560 3432
rect -18496 3368 -18476 3432
rect -19648 3352 -18476 3368
rect -19648 3288 -18560 3352
rect -18496 3288 -18476 3352
rect -19648 3272 -18476 3288
rect -19648 3208 -18560 3272
rect -18496 3208 -18476 3272
rect -19648 3192 -18476 3208
rect -19648 3128 -18560 3192
rect -18496 3128 -18476 3192
rect -19648 3112 -18476 3128
rect -19648 3048 -18560 3112
rect -18496 3048 -18476 3112
rect -19648 3032 -18476 3048
rect -19648 2968 -18560 3032
rect -18496 2968 -18476 3032
rect -19648 2920 -18476 2968
rect -18236 3752 -17064 3800
rect -18236 3688 -17148 3752
rect -17084 3688 -17064 3752
rect -18236 3672 -17064 3688
rect -18236 3608 -17148 3672
rect -17084 3608 -17064 3672
rect -18236 3592 -17064 3608
rect -18236 3528 -17148 3592
rect -17084 3528 -17064 3592
rect -18236 3512 -17064 3528
rect -18236 3448 -17148 3512
rect -17084 3448 -17064 3512
rect -18236 3432 -17064 3448
rect -18236 3368 -17148 3432
rect -17084 3368 -17064 3432
rect -18236 3352 -17064 3368
rect -18236 3288 -17148 3352
rect -17084 3288 -17064 3352
rect -18236 3272 -17064 3288
rect -18236 3208 -17148 3272
rect -17084 3208 -17064 3272
rect -18236 3192 -17064 3208
rect -18236 3128 -17148 3192
rect -17084 3128 -17064 3192
rect -18236 3112 -17064 3128
rect -18236 3048 -17148 3112
rect -17084 3048 -17064 3112
rect -18236 3032 -17064 3048
rect -18236 2968 -17148 3032
rect -17084 2968 -17064 3032
rect -18236 2920 -17064 2968
rect -16824 3752 -15652 3800
rect -16824 3688 -15736 3752
rect -15672 3688 -15652 3752
rect -16824 3672 -15652 3688
rect -16824 3608 -15736 3672
rect -15672 3608 -15652 3672
rect -16824 3592 -15652 3608
rect -16824 3528 -15736 3592
rect -15672 3528 -15652 3592
rect -16824 3512 -15652 3528
rect -16824 3448 -15736 3512
rect -15672 3448 -15652 3512
rect -16824 3432 -15652 3448
rect -16824 3368 -15736 3432
rect -15672 3368 -15652 3432
rect -16824 3352 -15652 3368
rect -16824 3288 -15736 3352
rect -15672 3288 -15652 3352
rect -16824 3272 -15652 3288
rect -16824 3208 -15736 3272
rect -15672 3208 -15652 3272
rect -16824 3192 -15652 3208
rect -16824 3128 -15736 3192
rect -15672 3128 -15652 3192
rect -16824 3112 -15652 3128
rect -16824 3048 -15736 3112
rect -15672 3048 -15652 3112
rect -16824 3032 -15652 3048
rect -16824 2968 -15736 3032
rect -15672 2968 -15652 3032
rect -16824 2920 -15652 2968
rect -15412 3752 -14240 3800
rect -15412 3688 -14324 3752
rect -14260 3688 -14240 3752
rect -15412 3672 -14240 3688
rect -15412 3608 -14324 3672
rect -14260 3608 -14240 3672
rect -15412 3592 -14240 3608
rect -15412 3528 -14324 3592
rect -14260 3528 -14240 3592
rect -15412 3512 -14240 3528
rect -15412 3448 -14324 3512
rect -14260 3448 -14240 3512
rect -15412 3432 -14240 3448
rect -15412 3368 -14324 3432
rect -14260 3368 -14240 3432
rect -15412 3352 -14240 3368
rect -15412 3288 -14324 3352
rect -14260 3288 -14240 3352
rect -15412 3272 -14240 3288
rect -15412 3208 -14324 3272
rect -14260 3208 -14240 3272
rect -15412 3192 -14240 3208
rect -15412 3128 -14324 3192
rect -14260 3128 -14240 3192
rect -15412 3112 -14240 3128
rect -15412 3048 -14324 3112
rect -14260 3048 -14240 3112
rect -15412 3032 -14240 3048
rect -15412 2968 -14324 3032
rect -14260 2968 -14240 3032
rect -15412 2920 -14240 2968
rect -14000 3752 -12828 3800
rect -14000 3688 -12912 3752
rect -12848 3688 -12828 3752
rect -14000 3672 -12828 3688
rect -14000 3608 -12912 3672
rect -12848 3608 -12828 3672
rect -14000 3592 -12828 3608
rect -14000 3528 -12912 3592
rect -12848 3528 -12828 3592
rect -14000 3512 -12828 3528
rect -14000 3448 -12912 3512
rect -12848 3448 -12828 3512
rect -14000 3432 -12828 3448
rect -14000 3368 -12912 3432
rect -12848 3368 -12828 3432
rect -14000 3352 -12828 3368
rect -14000 3288 -12912 3352
rect -12848 3288 -12828 3352
rect -14000 3272 -12828 3288
rect -14000 3208 -12912 3272
rect -12848 3208 -12828 3272
rect -14000 3192 -12828 3208
rect -14000 3128 -12912 3192
rect -12848 3128 -12828 3192
rect -14000 3112 -12828 3128
rect -14000 3048 -12912 3112
rect -12848 3048 -12828 3112
rect -14000 3032 -12828 3048
rect -14000 2968 -12912 3032
rect -12848 2968 -12828 3032
rect -14000 2920 -12828 2968
rect -12588 3752 -11416 3800
rect -12588 3688 -11500 3752
rect -11436 3688 -11416 3752
rect -12588 3672 -11416 3688
rect -12588 3608 -11500 3672
rect -11436 3608 -11416 3672
rect -12588 3592 -11416 3608
rect -12588 3528 -11500 3592
rect -11436 3528 -11416 3592
rect -12588 3512 -11416 3528
rect -12588 3448 -11500 3512
rect -11436 3448 -11416 3512
rect -12588 3432 -11416 3448
rect -12588 3368 -11500 3432
rect -11436 3368 -11416 3432
rect -12588 3352 -11416 3368
rect -12588 3288 -11500 3352
rect -11436 3288 -11416 3352
rect -12588 3272 -11416 3288
rect -12588 3208 -11500 3272
rect -11436 3208 -11416 3272
rect -12588 3192 -11416 3208
rect -12588 3128 -11500 3192
rect -11436 3128 -11416 3192
rect -12588 3112 -11416 3128
rect -12588 3048 -11500 3112
rect -11436 3048 -11416 3112
rect -12588 3032 -11416 3048
rect -12588 2968 -11500 3032
rect -11436 2968 -11416 3032
rect -12588 2920 -11416 2968
rect -11176 3752 -10004 3800
rect -11176 3688 -10088 3752
rect -10024 3688 -10004 3752
rect -11176 3672 -10004 3688
rect -11176 3608 -10088 3672
rect -10024 3608 -10004 3672
rect -11176 3592 -10004 3608
rect -11176 3528 -10088 3592
rect -10024 3528 -10004 3592
rect -11176 3512 -10004 3528
rect -11176 3448 -10088 3512
rect -10024 3448 -10004 3512
rect -11176 3432 -10004 3448
rect -11176 3368 -10088 3432
rect -10024 3368 -10004 3432
rect -11176 3352 -10004 3368
rect -11176 3288 -10088 3352
rect -10024 3288 -10004 3352
rect -11176 3272 -10004 3288
rect -11176 3208 -10088 3272
rect -10024 3208 -10004 3272
rect -11176 3192 -10004 3208
rect -11176 3128 -10088 3192
rect -10024 3128 -10004 3192
rect -11176 3112 -10004 3128
rect -11176 3048 -10088 3112
rect -10024 3048 -10004 3112
rect -11176 3032 -10004 3048
rect -11176 2968 -10088 3032
rect -10024 2968 -10004 3032
rect -11176 2920 -10004 2968
rect -9764 3752 -8592 3800
rect -9764 3688 -8676 3752
rect -8612 3688 -8592 3752
rect -9764 3672 -8592 3688
rect -9764 3608 -8676 3672
rect -8612 3608 -8592 3672
rect -9764 3592 -8592 3608
rect -9764 3528 -8676 3592
rect -8612 3528 -8592 3592
rect -9764 3512 -8592 3528
rect -9764 3448 -8676 3512
rect -8612 3448 -8592 3512
rect -9764 3432 -8592 3448
rect -9764 3368 -8676 3432
rect -8612 3368 -8592 3432
rect -9764 3352 -8592 3368
rect -9764 3288 -8676 3352
rect -8612 3288 -8592 3352
rect -9764 3272 -8592 3288
rect -9764 3208 -8676 3272
rect -8612 3208 -8592 3272
rect -9764 3192 -8592 3208
rect -9764 3128 -8676 3192
rect -8612 3128 -8592 3192
rect -9764 3112 -8592 3128
rect -9764 3048 -8676 3112
rect -8612 3048 -8592 3112
rect -9764 3032 -8592 3048
rect -9764 2968 -8676 3032
rect -8612 2968 -8592 3032
rect -9764 2920 -8592 2968
rect -8352 3752 -7180 3800
rect -8352 3688 -7264 3752
rect -7200 3688 -7180 3752
rect -8352 3672 -7180 3688
rect -8352 3608 -7264 3672
rect -7200 3608 -7180 3672
rect -8352 3592 -7180 3608
rect -8352 3528 -7264 3592
rect -7200 3528 -7180 3592
rect -8352 3512 -7180 3528
rect -8352 3448 -7264 3512
rect -7200 3448 -7180 3512
rect -8352 3432 -7180 3448
rect -8352 3368 -7264 3432
rect -7200 3368 -7180 3432
rect -8352 3352 -7180 3368
rect -8352 3288 -7264 3352
rect -7200 3288 -7180 3352
rect -8352 3272 -7180 3288
rect -8352 3208 -7264 3272
rect -7200 3208 -7180 3272
rect -8352 3192 -7180 3208
rect -8352 3128 -7264 3192
rect -7200 3128 -7180 3192
rect -8352 3112 -7180 3128
rect -8352 3048 -7264 3112
rect -7200 3048 -7180 3112
rect -8352 3032 -7180 3048
rect -8352 2968 -7264 3032
rect -7200 2968 -7180 3032
rect -8352 2920 -7180 2968
rect -6940 3752 -5768 3800
rect -6940 3688 -5852 3752
rect -5788 3688 -5768 3752
rect -6940 3672 -5768 3688
rect -6940 3608 -5852 3672
rect -5788 3608 -5768 3672
rect -6940 3592 -5768 3608
rect -6940 3528 -5852 3592
rect -5788 3528 -5768 3592
rect -6940 3512 -5768 3528
rect -6940 3448 -5852 3512
rect -5788 3448 -5768 3512
rect -6940 3432 -5768 3448
rect -6940 3368 -5852 3432
rect -5788 3368 -5768 3432
rect -6940 3352 -5768 3368
rect -6940 3288 -5852 3352
rect -5788 3288 -5768 3352
rect -6940 3272 -5768 3288
rect -6940 3208 -5852 3272
rect -5788 3208 -5768 3272
rect -6940 3192 -5768 3208
rect -6940 3128 -5852 3192
rect -5788 3128 -5768 3192
rect -6940 3112 -5768 3128
rect -6940 3048 -5852 3112
rect -5788 3048 -5768 3112
rect -6940 3032 -5768 3048
rect -6940 2968 -5852 3032
rect -5788 2968 -5768 3032
rect -6940 2920 -5768 2968
rect -5528 3752 -4356 3800
rect -5528 3688 -4440 3752
rect -4376 3688 -4356 3752
rect -5528 3672 -4356 3688
rect -5528 3608 -4440 3672
rect -4376 3608 -4356 3672
rect -5528 3592 -4356 3608
rect -5528 3528 -4440 3592
rect -4376 3528 -4356 3592
rect -5528 3512 -4356 3528
rect -5528 3448 -4440 3512
rect -4376 3448 -4356 3512
rect -5528 3432 -4356 3448
rect -5528 3368 -4440 3432
rect -4376 3368 -4356 3432
rect -5528 3352 -4356 3368
rect -5528 3288 -4440 3352
rect -4376 3288 -4356 3352
rect -5528 3272 -4356 3288
rect -5528 3208 -4440 3272
rect -4376 3208 -4356 3272
rect -5528 3192 -4356 3208
rect -5528 3128 -4440 3192
rect -4376 3128 -4356 3192
rect -5528 3112 -4356 3128
rect -5528 3048 -4440 3112
rect -4376 3048 -4356 3112
rect -5528 3032 -4356 3048
rect -5528 2968 -4440 3032
rect -4376 2968 -4356 3032
rect -5528 2920 -4356 2968
rect -4116 3752 -2944 3800
rect -4116 3688 -3028 3752
rect -2964 3688 -2944 3752
rect -4116 3672 -2944 3688
rect -4116 3608 -3028 3672
rect -2964 3608 -2944 3672
rect -4116 3592 -2944 3608
rect -4116 3528 -3028 3592
rect -2964 3528 -2944 3592
rect -4116 3512 -2944 3528
rect -4116 3448 -3028 3512
rect -2964 3448 -2944 3512
rect -4116 3432 -2944 3448
rect -4116 3368 -3028 3432
rect -2964 3368 -2944 3432
rect -4116 3352 -2944 3368
rect -4116 3288 -3028 3352
rect -2964 3288 -2944 3352
rect -4116 3272 -2944 3288
rect -4116 3208 -3028 3272
rect -2964 3208 -2944 3272
rect -4116 3192 -2944 3208
rect -4116 3128 -3028 3192
rect -2964 3128 -2944 3192
rect -4116 3112 -2944 3128
rect -4116 3048 -3028 3112
rect -2964 3048 -2944 3112
rect -4116 3032 -2944 3048
rect -4116 2968 -3028 3032
rect -2964 2968 -2944 3032
rect -4116 2920 -2944 2968
rect -2704 3752 -1532 3800
rect -2704 3688 -1616 3752
rect -1552 3688 -1532 3752
rect -2704 3672 -1532 3688
rect -2704 3608 -1616 3672
rect -1552 3608 -1532 3672
rect -2704 3592 -1532 3608
rect -2704 3528 -1616 3592
rect -1552 3528 -1532 3592
rect -2704 3512 -1532 3528
rect -2704 3448 -1616 3512
rect -1552 3448 -1532 3512
rect -2704 3432 -1532 3448
rect -2704 3368 -1616 3432
rect -1552 3368 -1532 3432
rect -2704 3352 -1532 3368
rect -2704 3288 -1616 3352
rect -1552 3288 -1532 3352
rect -2704 3272 -1532 3288
rect -2704 3208 -1616 3272
rect -1552 3208 -1532 3272
rect -2704 3192 -1532 3208
rect -2704 3128 -1616 3192
rect -1552 3128 -1532 3192
rect -2704 3112 -1532 3128
rect -2704 3048 -1616 3112
rect -1552 3048 -1532 3112
rect -2704 3032 -1532 3048
rect -2704 2968 -1616 3032
rect -1552 2968 -1532 3032
rect -2704 2920 -1532 2968
rect -1292 3752 -120 3800
rect -1292 3688 -204 3752
rect -140 3688 -120 3752
rect -1292 3672 -120 3688
rect -1292 3608 -204 3672
rect -140 3608 -120 3672
rect -1292 3592 -120 3608
rect -1292 3528 -204 3592
rect -140 3528 -120 3592
rect -1292 3512 -120 3528
rect -1292 3448 -204 3512
rect -140 3448 -120 3512
rect -1292 3432 -120 3448
rect -1292 3368 -204 3432
rect -140 3368 -120 3432
rect -1292 3352 -120 3368
rect -1292 3288 -204 3352
rect -140 3288 -120 3352
rect -1292 3272 -120 3288
rect -1292 3208 -204 3272
rect -140 3208 -120 3272
rect -1292 3192 -120 3208
rect -1292 3128 -204 3192
rect -140 3128 -120 3192
rect -1292 3112 -120 3128
rect -1292 3048 -204 3112
rect -140 3048 -120 3112
rect -1292 3032 -120 3048
rect -1292 2968 -204 3032
rect -140 2968 -120 3032
rect -1292 2920 -120 2968
rect 120 3752 1292 3800
rect 120 3688 1208 3752
rect 1272 3688 1292 3752
rect 120 3672 1292 3688
rect 120 3608 1208 3672
rect 1272 3608 1292 3672
rect 120 3592 1292 3608
rect 120 3528 1208 3592
rect 1272 3528 1292 3592
rect 120 3512 1292 3528
rect 120 3448 1208 3512
rect 1272 3448 1292 3512
rect 120 3432 1292 3448
rect 120 3368 1208 3432
rect 1272 3368 1292 3432
rect 120 3352 1292 3368
rect 120 3288 1208 3352
rect 1272 3288 1292 3352
rect 120 3272 1292 3288
rect 120 3208 1208 3272
rect 1272 3208 1292 3272
rect 120 3192 1292 3208
rect 120 3128 1208 3192
rect 1272 3128 1292 3192
rect 120 3112 1292 3128
rect 120 3048 1208 3112
rect 1272 3048 1292 3112
rect 120 3032 1292 3048
rect 120 2968 1208 3032
rect 1272 2968 1292 3032
rect 120 2920 1292 2968
rect 1532 3752 2704 3800
rect 1532 3688 2620 3752
rect 2684 3688 2704 3752
rect 1532 3672 2704 3688
rect 1532 3608 2620 3672
rect 2684 3608 2704 3672
rect 1532 3592 2704 3608
rect 1532 3528 2620 3592
rect 2684 3528 2704 3592
rect 1532 3512 2704 3528
rect 1532 3448 2620 3512
rect 2684 3448 2704 3512
rect 1532 3432 2704 3448
rect 1532 3368 2620 3432
rect 2684 3368 2704 3432
rect 1532 3352 2704 3368
rect 1532 3288 2620 3352
rect 2684 3288 2704 3352
rect 1532 3272 2704 3288
rect 1532 3208 2620 3272
rect 2684 3208 2704 3272
rect 1532 3192 2704 3208
rect 1532 3128 2620 3192
rect 2684 3128 2704 3192
rect 1532 3112 2704 3128
rect 1532 3048 2620 3112
rect 2684 3048 2704 3112
rect 1532 3032 2704 3048
rect 1532 2968 2620 3032
rect 2684 2968 2704 3032
rect 1532 2920 2704 2968
rect 2944 3752 4116 3800
rect 2944 3688 4032 3752
rect 4096 3688 4116 3752
rect 2944 3672 4116 3688
rect 2944 3608 4032 3672
rect 4096 3608 4116 3672
rect 2944 3592 4116 3608
rect 2944 3528 4032 3592
rect 4096 3528 4116 3592
rect 2944 3512 4116 3528
rect 2944 3448 4032 3512
rect 4096 3448 4116 3512
rect 2944 3432 4116 3448
rect 2944 3368 4032 3432
rect 4096 3368 4116 3432
rect 2944 3352 4116 3368
rect 2944 3288 4032 3352
rect 4096 3288 4116 3352
rect 2944 3272 4116 3288
rect 2944 3208 4032 3272
rect 4096 3208 4116 3272
rect 2944 3192 4116 3208
rect 2944 3128 4032 3192
rect 4096 3128 4116 3192
rect 2944 3112 4116 3128
rect 2944 3048 4032 3112
rect 4096 3048 4116 3112
rect 2944 3032 4116 3048
rect 2944 2968 4032 3032
rect 4096 2968 4116 3032
rect 2944 2920 4116 2968
rect 4356 3752 5528 3800
rect 4356 3688 5444 3752
rect 5508 3688 5528 3752
rect 4356 3672 5528 3688
rect 4356 3608 5444 3672
rect 5508 3608 5528 3672
rect 4356 3592 5528 3608
rect 4356 3528 5444 3592
rect 5508 3528 5528 3592
rect 4356 3512 5528 3528
rect 4356 3448 5444 3512
rect 5508 3448 5528 3512
rect 4356 3432 5528 3448
rect 4356 3368 5444 3432
rect 5508 3368 5528 3432
rect 4356 3352 5528 3368
rect 4356 3288 5444 3352
rect 5508 3288 5528 3352
rect 4356 3272 5528 3288
rect 4356 3208 5444 3272
rect 5508 3208 5528 3272
rect 4356 3192 5528 3208
rect 4356 3128 5444 3192
rect 5508 3128 5528 3192
rect 4356 3112 5528 3128
rect 4356 3048 5444 3112
rect 5508 3048 5528 3112
rect 4356 3032 5528 3048
rect 4356 2968 5444 3032
rect 5508 2968 5528 3032
rect 4356 2920 5528 2968
rect 5768 3752 6940 3800
rect 5768 3688 6856 3752
rect 6920 3688 6940 3752
rect 5768 3672 6940 3688
rect 5768 3608 6856 3672
rect 6920 3608 6940 3672
rect 5768 3592 6940 3608
rect 5768 3528 6856 3592
rect 6920 3528 6940 3592
rect 5768 3512 6940 3528
rect 5768 3448 6856 3512
rect 6920 3448 6940 3512
rect 5768 3432 6940 3448
rect 5768 3368 6856 3432
rect 6920 3368 6940 3432
rect 5768 3352 6940 3368
rect 5768 3288 6856 3352
rect 6920 3288 6940 3352
rect 5768 3272 6940 3288
rect 5768 3208 6856 3272
rect 6920 3208 6940 3272
rect 5768 3192 6940 3208
rect 5768 3128 6856 3192
rect 6920 3128 6940 3192
rect 5768 3112 6940 3128
rect 5768 3048 6856 3112
rect 6920 3048 6940 3112
rect 5768 3032 6940 3048
rect 5768 2968 6856 3032
rect 6920 2968 6940 3032
rect 5768 2920 6940 2968
rect 7180 3752 8352 3800
rect 7180 3688 8268 3752
rect 8332 3688 8352 3752
rect 7180 3672 8352 3688
rect 7180 3608 8268 3672
rect 8332 3608 8352 3672
rect 7180 3592 8352 3608
rect 7180 3528 8268 3592
rect 8332 3528 8352 3592
rect 7180 3512 8352 3528
rect 7180 3448 8268 3512
rect 8332 3448 8352 3512
rect 7180 3432 8352 3448
rect 7180 3368 8268 3432
rect 8332 3368 8352 3432
rect 7180 3352 8352 3368
rect 7180 3288 8268 3352
rect 8332 3288 8352 3352
rect 7180 3272 8352 3288
rect 7180 3208 8268 3272
rect 8332 3208 8352 3272
rect 7180 3192 8352 3208
rect 7180 3128 8268 3192
rect 8332 3128 8352 3192
rect 7180 3112 8352 3128
rect 7180 3048 8268 3112
rect 8332 3048 8352 3112
rect 7180 3032 8352 3048
rect 7180 2968 8268 3032
rect 8332 2968 8352 3032
rect 7180 2920 8352 2968
rect 8592 3752 9764 3800
rect 8592 3688 9680 3752
rect 9744 3688 9764 3752
rect 8592 3672 9764 3688
rect 8592 3608 9680 3672
rect 9744 3608 9764 3672
rect 8592 3592 9764 3608
rect 8592 3528 9680 3592
rect 9744 3528 9764 3592
rect 8592 3512 9764 3528
rect 8592 3448 9680 3512
rect 9744 3448 9764 3512
rect 8592 3432 9764 3448
rect 8592 3368 9680 3432
rect 9744 3368 9764 3432
rect 8592 3352 9764 3368
rect 8592 3288 9680 3352
rect 9744 3288 9764 3352
rect 8592 3272 9764 3288
rect 8592 3208 9680 3272
rect 9744 3208 9764 3272
rect 8592 3192 9764 3208
rect 8592 3128 9680 3192
rect 9744 3128 9764 3192
rect 8592 3112 9764 3128
rect 8592 3048 9680 3112
rect 9744 3048 9764 3112
rect 8592 3032 9764 3048
rect 8592 2968 9680 3032
rect 9744 2968 9764 3032
rect 8592 2920 9764 2968
rect 10004 3752 11176 3800
rect 10004 3688 11092 3752
rect 11156 3688 11176 3752
rect 10004 3672 11176 3688
rect 10004 3608 11092 3672
rect 11156 3608 11176 3672
rect 10004 3592 11176 3608
rect 10004 3528 11092 3592
rect 11156 3528 11176 3592
rect 10004 3512 11176 3528
rect 10004 3448 11092 3512
rect 11156 3448 11176 3512
rect 10004 3432 11176 3448
rect 10004 3368 11092 3432
rect 11156 3368 11176 3432
rect 10004 3352 11176 3368
rect 10004 3288 11092 3352
rect 11156 3288 11176 3352
rect 10004 3272 11176 3288
rect 10004 3208 11092 3272
rect 11156 3208 11176 3272
rect 10004 3192 11176 3208
rect 10004 3128 11092 3192
rect 11156 3128 11176 3192
rect 10004 3112 11176 3128
rect 10004 3048 11092 3112
rect 11156 3048 11176 3112
rect 10004 3032 11176 3048
rect 10004 2968 11092 3032
rect 11156 2968 11176 3032
rect 10004 2920 11176 2968
rect 11416 3752 12588 3800
rect 11416 3688 12504 3752
rect 12568 3688 12588 3752
rect 11416 3672 12588 3688
rect 11416 3608 12504 3672
rect 12568 3608 12588 3672
rect 11416 3592 12588 3608
rect 11416 3528 12504 3592
rect 12568 3528 12588 3592
rect 11416 3512 12588 3528
rect 11416 3448 12504 3512
rect 12568 3448 12588 3512
rect 11416 3432 12588 3448
rect 11416 3368 12504 3432
rect 12568 3368 12588 3432
rect 11416 3352 12588 3368
rect 11416 3288 12504 3352
rect 12568 3288 12588 3352
rect 11416 3272 12588 3288
rect 11416 3208 12504 3272
rect 12568 3208 12588 3272
rect 11416 3192 12588 3208
rect 11416 3128 12504 3192
rect 12568 3128 12588 3192
rect 11416 3112 12588 3128
rect 11416 3048 12504 3112
rect 12568 3048 12588 3112
rect 11416 3032 12588 3048
rect 11416 2968 12504 3032
rect 12568 2968 12588 3032
rect 11416 2920 12588 2968
rect 12828 3752 14000 3800
rect 12828 3688 13916 3752
rect 13980 3688 14000 3752
rect 12828 3672 14000 3688
rect 12828 3608 13916 3672
rect 13980 3608 14000 3672
rect 12828 3592 14000 3608
rect 12828 3528 13916 3592
rect 13980 3528 14000 3592
rect 12828 3512 14000 3528
rect 12828 3448 13916 3512
rect 13980 3448 14000 3512
rect 12828 3432 14000 3448
rect 12828 3368 13916 3432
rect 13980 3368 14000 3432
rect 12828 3352 14000 3368
rect 12828 3288 13916 3352
rect 13980 3288 14000 3352
rect 12828 3272 14000 3288
rect 12828 3208 13916 3272
rect 13980 3208 14000 3272
rect 12828 3192 14000 3208
rect 12828 3128 13916 3192
rect 13980 3128 14000 3192
rect 12828 3112 14000 3128
rect 12828 3048 13916 3112
rect 13980 3048 14000 3112
rect 12828 3032 14000 3048
rect 12828 2968 13916 3032
rect 13980 2968 14000 3032
rect 12828 2920 14000 2968
rect 14240 3752 15412 3800
rect 14240 3688 15328 3752
rect 15392 3688 15412 3752
rect 14240 3672 15412 3688
rect 14240 3608 15328 3672
rect 15392 3608 15412 3672
rect 14240 3592 15412 3608
rect 14240 3528 15328 3592
rect 15392 3528 15412 3592
rect 14240 3512 15412 3528
rect 14240 3448 15328 3512
rect 15392 3448 15412 3512
rect 14240 3432 15412 3448
rect 14240 3368 15328 3432
rect 15392 3368 15412 3432
rect 14240 3352 15412 3368
rect 14240 3288 15328 3352
rect 15392 3288 15412 3352
rect 14240 3272 15412 3288
rect 14240 3208 15328 3272
rect 15392 3208 15412 3272
rect 14240 3192 15412 3208
rect 14240 3128 15328 3192
rect 15392 3128 15412 3192
rect 14240 3112 15412 3128
rect 14240 3048 15328 3112
rect 15392 3048 15412 3112
rect 14240 3032 15412 3048
rect 14240 2968 15328 3032
rect 15392 2968 15412 3032
rect 14240 2920 15412 2968
rect 15652 3752 16824 3800
rect 15652 3688 16740 3752
rect 16804 3688 16824 3752
rect 15652 3672 16824 3688
rect 15652 3608 16740 3672
rect 16804 3608 16824 3672
rect 15652 3592 16824 3608
rect 15652 3528 16740 3592
rect 16804 3528 16824 3592
rect 15652 3512 16824 3528
rect 15652 3448 16740 3512
rect 16804 3448 16824 3512
rect 15652 3432 16824 3448
rect 15652 3368 16740 3432
rect 16804 3368 16824 3432
rect 15652 3352 16824 3368
rect 15652 3288 16740 3352
rect 16804 3288 16824 3352
rect 15652 3272 16824 3288
rect 15652 3208 16740 3272
rect 16804 3208 16824 3272
rect 15652 3192 16824 3208
rect 15652 3128 16740 3192
rect 16804 3128 16824 3192
rect 15652 3112 16824 3128
rect 15652 3048 16740 3112
rect 16804 3048 16824 3112
rect 15652 3032 16824 3048
rect 15652 2968 16740 3032
rect 16804 2968 16824 3032
rect 15652 2920 16824 2968
rect 17064 3752 18236 3800
rect 17064 3688 18152 3752
rect 18216 3688 18236 3752
rect 17064 3672 18236 3688
rect 17064 3608 18152 3672
rect 18216 3608 18236 3672
rect 17064 3592 18236 3608
rect 17064 3528 18152 3592
rect 18216 3528 18236 3592
rect 17064 3512 18236 3528
rect 17064 3448 18152 3512
rect 18216 3448 18236 3512
rect 17064 3432 18236 3448
rect 17064 3368 18152 3432
rect 18216 3368 18236 3432
rect 17064 3352 18236 3368
rect 17064 3288 18152 3352
rect 18216 3288 18236 3352
rect 17064 3272 18236 3288
rect 17064 3208 18152 3272
rect 18216 3208 18236 3272
rect 17064 3192 18236 3208
rect 17064 3128 18152 3192
rect 18216 3128 18236 3192
rect 17064 3112 18236 3128
rect 17064 3048 18152 3112
rect 18216 3048 18236 3112
rect 17064 3032 18236 3048
rect 17064 2968 18152 3032
rect 18216 2968 18236 3032
rect 17064 2920 18236 2968
rect 18476 3752 19648 3800
rect 18476 3688 19564 3752
rect 19628 3688 19648 3752
rect 18476 3672 19648 3688
rect 18476 3608 19564 3672
rect 19628 3608 19648 3672
rect 18476 3592 19648 3608
rect 18476 3528 19564 3592
rect 19628 3528 19648 3592
rect 18476 3512 19648 3528
rect 18476 3448 19564 3512
rect 19628 3448 19648 3512
rect 18476 3432 19648 3448
rect 18476 3368 19564 3432
rect 19628 3368 19648 3432
rect 18476 3352 19648 3368
rect 18476 3288 19564 3352
rect 19628 3288 19648 3352
rect 18476 3272 19648 3288
rect 18476 3208 19564 3272
rect 19628 3208 19648 3272
rect 18476 3192 19648 3208
rect 18476 3128 19564 3192
rect 19628 3128 19648 3192
rect 18476 3112 19648 3128
rect 18476 3048 19564 3112
rect 19628 3048 19648 3112
rect 18476 3032 19648 3048
rect 18476 2968 19564 3032
rect 19628 2968 19648 3032
rect 18476 2920 19648 2968
rect 19888 3752 21060 3800
rect 19888 3688 20976 3752
rect 21040 3688 21060 3752
rect 19888 3672 21060 3688
rect 19888 3608 20976 3672
rect 21040 3608 21060 3672
rect 19888 3592 21060 3608
rect 19888 3528 20976 3592
rect 21040 3528 21060 3592
rect 19888 3512 21060 3528
rect 19888 3448 20976 3512
rect 21040 3448 21060 3512
rect 19888 3432 21060 3448
rect 19888 3368 20976 3432
rect 21040 3368 21060 3432
rect 19888 3352 21060 3368
rect 19888 3288 20976 3352
rect 21040 3288 21060 3352
rect 19888 3272 21060 3288
rect 19888 3208 20976 3272
rect 21040 3208 21060 3272
rect 19888 3192 21060 3208
rect 19888 3128 20976 3192
rect 21040 3128 21060 3192
rect 19888 3112 21060 3128
rect 19888 3048 20976 3112
rect 21040 3048 21060 3112
rect 19888 3032 21060 3048
rect 19888 2968 20976 3032
rect 21040 2968 21060 3032
rect 19888 2920 21060 2968
rect 21300 3752 22472 3800
rect 21300 3688 22388 3752
rect 22452 3688 22472 3752
rect 21300 3672 22472 3688
rect 21300 3608 22388 3672
rect 22452 3608 22472 3672
rect 21300 3592 22472 3608
rect 21300 3528 22388 3592
rect 22452 3528 22472 3592
rect 21300 3512 22472 3528
rect 21300 3448 22388 3512
rect 22452 3448 22472 3512
rect 21300 3432 22472 3448
rect 21300 3368 22388 3432
rect 22452 3368 22472 3432
rect 21300 3352 22472 3368
rect 21300 3288 22388 3352
rect 22452 3288 22472 3352
rect 21300 3272 22472 3288
rect 21300 3208 22388 3272
rect 22452 3208 22472 3272
rect 21300 3192 22472 3208
rect 21300 3128 22388 3192
rect 22452 3128 22472 3192
rect 21300 3112 22472 3128
rect 21300 3048 22388 3112
rect 22452 3048 22472 3112
rect 21300 3032 22472 3048
rect 21300 2968 22388 3032
rect 22452 2968 22472 3032
rect 21300 2920 22472 2968
rect 22712 3752 23884 3800
rect 22712 3688 23800 3752
rect 23864 3688 23884 3752
rect 22712 3672 23884 3688
rect 22712 3608 23800 3672
rect 23864 3608 23884 3672
rect 22712 3592 23884 3608
rect 22712 3528 23800 3592
rect 23864 3528 23884 3592
rect 22712 3512 23884 3528
rect 22712 3448 23800 3512
rect 23864 3448 23884 3512
rect 22712 3432 23884 3448
rect 22712 3368 23800 3432
rect 23864 3368 23884 3432
rect 22712 3352 23884 3368
rect 22712 3288 23800 3352
rect 23864 3288 23884 3352
rect 22712 3272 23884 3288
rect 22712 3208 23800 3272
rect 23864 3208 23884 3272
rect 22712 3192 23884 3208
rect 22712 3128 23800 3192
rect 23864 3128 23884 3192
rect 22712 3112 23884 3128
rect 22712 3048 23800 3112
rect 23864 3048 23884 3112
rect 22712 3032 23884 3048
rect 22712 2968 23800 3032
rect 23864 2968 23884 3032
rect 22712 2920 23884 2968
rect -23884 2632 -22712 2680
rect -23884 2568 -22796 2632
rect -22732 2568 -22712 2632
rect -23884 2552 -22712 2568
rect -23884 2488 -22796 2552
rect -22732 2488 -22712 2552
rect -23884 2472 -22712 2488
rect -23884 2408 -22796 2472
rect -22732 2408 -22712 2472
rect -23884 2392 -22712 2408
rect -23884 2328 -22796 2392
rect -22732 2328 -22712 2392
rect -23884 2312 -22712 2328
rect -23884 2248 -22796 2312
rect -22732 2248 -22712 2312
rect -23884 2232 -22712 2248
rect -23884 2168 -22796 2232
rect -22732 2168 -22712 2232
rect -23884 2152 -22712 2168
rect -23884 2088 -22796 2152
rect -22732 2088 -22712 2152
rect -23884 2072 -22712 2088
rect -23884 2008 -22796 2072
rect -22732 2008 -22712 2072
rect -23884 1992 -22712 2008
rect -23884 1928 -22796 1992
rect -22732 1928 -22712 1992
rect -23884 1912 -22712 1928
rect -23884 1848 -22796 1912
rect -22732 1848 -22712 1912
rect -23884 1800 -22712 1848
rect -22472 2632 -21300 2680
rect -22472 2568 -21384 2632
rect -21320 2568 -21300 2632
rect -22472 2552 -21300 2568
rect -22472 2488 -21384 2552
rect -21320 2488 -21300 2552
rect -22472 2472 -21300 2488
rect -22472 2408 -21384 2472
rect -21320 2408 -21300 2472
rect -22472 2392 -21300 2408
rect -22472 2328 -21384 2392
rect -21320 2328 -21300 2392
rect -22472 2312 -21300 2328
rect -22472 2248 -21384 2312
rect -21320 2248 -21300 2312
rect -22472 2232 -21300 2248
rect -22472 2168 -21384 2232
rect -21320 2168 -21300 2232
rect -22472 2152 -21300 2168
rect -22472 2088 -21384 2152
rect -21320 2088 -21300 2152
rect -22472 2072 -21300 2088
rect -22472 2008 -21384 2072
rect -21320 2008 -21300 2072
rect -22472 1992 -21300 2008
rect -22472 1928 -21384 1992
rect -21320 1928 -21300 1992
rect -22472 1912 -21300 1928
rect -22472 1848 -21384 1912
rect -21320 1848 -21300 1912
rect -22472 1800 -21300 1848
rect -21060 2632 -19888 2680
rect -21060 2568 -19972 2632
rect -19908 2568 -19888 2632
rect -21060 2552 -19888 2568
rect -21060 2488 -19972 2552
rect -19908 2488 -19888 2552
rect -21060 2472 -19888 2488
rect -21060 2408 -19972 2472
rect -19908 2408 -19888 2472
rect -21060 2392 -19888 2408
rect -21060 2328 -19972 2392
rect -19908 2328 -19888 2392
rect -21060 2312 -19888 2328
rect -21060 2248 -19972 2312
rect -19908 2248 -19888 2312
rect -21060 2232 -19888 2248
rect -21060 2168 -19972 2232
rect -19908 2168 -19888 2232
rect -21060 2152 -19888 2168
rect -21060 2088 -19972 2152
rect -19908 2088 -19888 2152
rect -21060 2072 -19888 2088
rect -21060 2008 -19972 2072
rect -19908 2008 -19888 2072
rect -21060 1992 -19888 2008
rect -21060 1928 -19972 1992
rect -19908 1928 -19888 1992
rect -21060 1912 -19888 1928
rect -21060 1848 -19972 1912
rect -19908 1848 -19888 1912
rect -21060 1800 -19888 1848
rect -19648 2632 -18476 2680
rect -19648 2568 -18560 2632
rect -18496 2568 -18476 2632
rect -19648 2552 -18476 2568
rect -19648 2488 -18560 2552
rect -18496 2488 -18476 2552
rect -19648 2472 -18476 2488
rect -19648 2408 -18560 2472
rect -18496 2408 -18476 2472
rect -19648 2392 -18476 2408
rect -19648 2328 -18560 2392
rect -18496 2328 -18476 2392
rect -19648 2312 -18476 2328
rect -19648 2248 -18560 2312
rect -18496 2248 -18476 2312
rect -19648 2232 -18476 2248
rect -19648 2168 -18560 2232
rect -18496 2168 -18476 2232
rect -19648 2152 -18476 2168
rect -19648 2088 -18560 2152
rect -18496 2088 -18476 2152
rect -19648 2072 -18476 2088
rect -19648 2008 -18560 2072
rect -18496 2008 -18476 2072
rect -19648 1992 -18476 2008
rect -19648 1928 -18560 1992
rect -18496 1928 -18476 1992
rect -19648 1912 -18476 1928
rect -19648 1848 -18560 1912
rect -18496 1848 -18476 1912
rect -19648 1800 -18476 1848
rect -18236 2632 -17064 2680
rect -18236 2568 -17148 2632
rect -17084 2568 -17064 2632
rect -18236 2552 -17064 2568
rect -18236 2488 -17148 2552
rect -17084 2488 -17064 2552
rect -18236 2472 -17064 2488
rect -18236 2408 -17148 2472
rect -17084 2408 -17064 2472
rect -18236 2392 -17064 2408
rect -18236 2328 -17148 2392
rect -17084 2328 -17064 2392
rect -18236 2312 -17064 2328
rect -18236 2248 -17148 2312
rect -17084 2248 -17064 2312
rect -18236 2232 -17064 2248
rect -18236 2168 -17148 2232
rect -17084 2168 -17064 2232
rect -18236 2152 -17064 2168
rect -18236 2088 -17148 2152
rect -17084 2088 -17064 2152
rect -18236 2072 -17064 2088
rect -18236 2008 -17148 2072
rect -17084 2008 -17064 2072
rect -18236 1992 -17064 2008
rect -18236 1928 -17148 1992
rect -17084 1928 -17064 1992
rect -18236 1912 -17064 1928
rect -18236 1848 -17148 1912
rect -17084 1848 -17064 1912
rect -18236 1800 -17064 1848
rect -16824 2632 -15652 2680
rect -16824 2568 -15736 2632
rect -15672 2568 -15652 2632
rect -16824 2552 -15652 2568
rect -16824 2488 -15736 2552
rect -15672 2488 -15652 2552
rect -16824 2472 -15652 2488
rect -16824 2408 -15736 2472
rect -15672 2408 -15652 2472
rect -16824 2392 -15652 2408
rect -16824 2328 -15736 2392
rect -15672 2328 -15652 2392
rect -16824 2312 -15652 2328
rect -16824 2248 -15736 2312
rect -15672 2248 -15652 2312
rect -16824 2232 -15652 2248
rect -16824 2168 -15736 2232
rect -15672 2168 -15652 2232
rect -16824 2152 -15652 2168
rect -16824 2088 -15736 2152
rect -15672 2088 -15652 2152
rect -16824 2072 -15652 2088
rect -16824 2008 -15736 2072
rect -15672 2008 -15652 2072
rect -16824 1992 -15652 2008
rect -16824 1928 -15736 1992
rect -15672 1928 -15652 1992
rect -16824 1912 -15652 1928
rect -16824 1848 -15736 1912
rect -15672 1848 -15652 1912
rect -16824 1800 -15652 1848
rect -15412 2632 -14240 2680
rect -15412 2568 -14324 2632
rect -14260 2568 -14240 2632
rect -15412 2552 -14240 2568
rect -15412 2488 -14324 2552
rect -14260 2488 -14240 2552
rect -15412 2472 -14240 2488
rect -15412 2408 -14324 2472
rect -14260 2408 -14240 2472
rect -15412 2392 -14240 2408
rect -15412 2328 -14324 2392
rect -14260 2328 -14240 2392
rect -15412 2312 -14240 2328
rect -15412 2248 -14324 2312
rect -14260 2248 -14240 2312
rect -15412 2232 -14240 2248
rect -15412 2168 -14324 2232
rect -14260 2168 -14240 2232
rect -15412 2152 -14240 2168
rect -15412 2088 -14324 2152
rect -14260 2088 -14240 2152
rect -15412 2072 -14240 2088
rect -15412 2008 -14324 2072
rect -14260 2008 -14240 2072
rect -15412 1992 -14240 2008
rect -15412 1928 -14324 1992
rect -14260 1928 -14240 1992
rect -15412 1912 -14240 1928
rect -15412 1848 -14324 1912
rect -14260 1848 -14240 1912
rect -15412 1800 -14240 1848
rect -14000 2632 -12828 2680
rect -14000 2568 -12912 2632
rect -12848 2568 -12828 2632
rect -14000 2552 -12828 2568
rect -14000 2488 -12912 2552
rect -12848 2488 -12828 2552
rect -14000 2472 -12828 2488
rect -14000 2408 -12912 2472
rect -12848 2408 -12828 2472
rect -14000 2392 -12828 2408
rect -14000 2328 -12912 2392
rect -12848 2328 -12828 2392
rect -14000 2312 -12828 2328
rect -14000 2248 -12912 2312
rect -12848 2248 -12828 2312
rect -14000 2232 -12828 2248
rect -14000 2168 -12912 2232
rect -12848 2168 -12828 2232
rect -14000 2152 -12828 2168
rect -14000 2088 -12912 2152
rect -12848 2088 -12828 2152
rect -14000 2072 -12828 2088
rect -14000 2008 -12912 2072
rect -12848 2008 -12828 2072
rect -14000 1992 -12828 2008
rect -14000 1928 -12912 1992
rect -12848 1928 -12828 1992
rect -14000 1912 -12828 1928
rect -14000 1848 -12912 1912
rect -12848 1848 -12828 1912
rect -14000 1800 -12828 1848
rect -12588 2632 -11416 2680
rect -12588 2568 -11500 2632
rect -11436 2568 -11416 2632
rect -12588 2552 -11416 2568
rect -12588 2488 -11500 2552
rect -11436 2488 -11416 2552
rect -12588 2472 -11416 2488
rect -12588 2408 -11500 2472
rect -11436 2408 -11416 2472
rect -12588 2392 -11416 2408
rect -12588 2328 -11500 2392
rect -11436 2328 -11416 2392
rect -12588 2312 -11416 2328
rect -12588 2248 -11500 2312
rect -11436 2248 -11416 2312
rect -12588 2232 -11416 2248
rect -12588 2168 -11500 2232
rect -11436 2168 -11416 2232
rect -12588 2152 -11416 2168
rect -12588 2088 -11500 2152
rect -11436 2088 -11416 2152
rect -12588 2072 -11416 2088
rect -12588 2008 -11500 2072
rect -11436 2008 -11416 2072
rect -12588 1992 -11416 2008
rect -12588 1928 -11500 1992
rect -11436 1928 -11416 1992
rect -12588 1912 -11416 1928
rect -12588 1848 -11500 1912
rect -11436 1848 -11416 1912
rect -12588 1800 -11416 1848
rect -11176 2632 -10004 2680
rect -11176 2568 -10088 2632
rect -10024 2568 -10004 2632
rect -11176 2552 -10004 2568
rect -11176 2488 -10088 2552
rect -10024 2488 -10004 2552
rect -11176 2472 -10004 2488
rect -11176 2408 -10088 2472
rect -10024 2408 -10004 2472
rect -11176 2392 -10004 2408
rect -11176 2328 -10088 2392
rect -10024 2328 -10004 2392
rect -11176 2312 -10004 2328
rect -11176 2248 -10088 2312
rect -10024 2248 -10004 2312
rect -11176 2232 -10004 2248
rect -11176 2168 -10088 2232
rect -10024 2168 -10004 2232
rect -11176 2152 -10004 2168
rect -11176 2088 -10088 2152
rect -10024 2088 -10004 2152
rect -11176 2072 -10004 2088
rect -11176 2008 -10088 2072
rect -10024 2008 -10004 2072
rect -11176 1992 -10004 2008
rect -11176 1928 -10088 1992
rect -10024 1928 -10004 1992
rect -11176 1912 -10004 1928
rect -11176 1848 -10088 1912
rect -10024 1848 -10004 1912
rect -11176 1800 -10004 1848
rect -9764 2632 -8592 2680
rect -9764 2568 -8676 2632
rect -8612 2568 -8592 2632
rect -9764 2552 -8592 2568
rect -9764 2488 -8676 2552
rect -8612 2488 -8592 2552
rect -9764 2472 -8592 2488
rect -9764 2408 -8676 2472
rect -8612 2408 -8592 2472
rect -9764 2392 -8592 2408
rect -9764 2328 -8676 2392
rect -8612 2328 -8592 2392
rect -9764 2312 -8592 2328
rect -9764 2248 -8676 2312
rect -8612 2248 -8592 2312
rect -9764 2232 -8592 2248
rect -9764 2168 -8676 2232
rect -8612 2168 -8592 2232
rect -9764 2152 -8592 2168
rect -9764 2088 -8676 2152
rect -8612 2088 -8592 2152
rect -9764 2072 -8592 2088
rect -9764 2008 -8676 2072
rect -8612 2008 -8592 2072
rect -9764 1992 -8592 2008
rect -9764 1928 -8676 1992
rect -8612 1928 -8592 1992
rect -9764 1912 -8592 1928
rect -9764 1848 -8676 1912
rect -8612 1848 -8592 1912
rect -9764 1800 -8592 1848
rect -8352 2632 -7180 2680
rect -8352 2568 -7264 2632
rect -7200 2568 -7180 2632
rect -8352 2552 -7180 2568
rect -8352 2488 -7264 2552
rect -7200 2488 -7180 2552
rect -8352 2472 -7180 2488
rect -8352 2408 -7264 2472
rect -7200 2408 -7180 2472
rect -8352 2392 -7180 2408
rect -8352 2328 -7264 2392
rect -7200 2328 -7180 2392
rect -8352 2312 -7180 2328
rect -8352 2248 -7264 2312
rect -7200 2248 -7180 2312
rect -8352 2232 -7180 2248
rect -8352 2168 -7264 2232
rect -7200 2168 -7180 2232
rect -8352 2152 -7180 2168
rect -8352 2088 -7264 2152
rect -7200 2088 -7180 2152
rect -8352 2072 -7180 2088
rect -8352 2008 -7264 2072
rect -7200 2008 -7180 2072
rect -8352 1992 -7180 2008
rect -8352 1928 -7264 1992
rect -7200 1928 -7180 1992
rect -8352 1912 -7180 1928
rect -8352 1848 -7264 1912
rect -7200 1848 -7180 1912
rect -8352 1800 -7180 1848
rect -6940 2632 -5768 2680
rect -6940 2568 -5852 2632
rect -5788 2568 -5768 2632
rect -6940 2552 -5768 2568
rect -6940 2488 -5852 2552
rect -5788 2488 -5768 2552
rect -6940 2472 -5768 2488
rect -6940 2408 -5852 2472
rect -5788 2408 -5768 2472
rect -6940 2392 -5768 2408
rect -6940 2328 -5852 2392
rect -5788 2328 -5768 2392
rect -6940 2312 -5768 2328
rect -6940 2248 -5852 2312
rect -5788 2248 -5768 2312
rect -6940 2232 -5768 2248
rect -6940 2168 -5852 2232
rect -5788 2168 -5768 2232
rect -6940 2152 -5768 2168
rect -6940 2088 -5852 2152
rect -5788 2088 -5768 2152
rect -6940 2072 -5768 2088
rect -6940 2008 -5852 2072
rect -5788 2008 -5768 2072
rect -6940 1992 -5768 2008
rect -6940 1928 -5852 1992
rect -5788 1928 -5768 1992
rect -6940 1912 -5768 1928
rect -6940 1848 -5852 1912
rect -5788 1848 -5768 1912
rect -6940 1800 -5768 1848
rect -5528 2632 -4356 2680
rect -5528 2568 -4440 2632
rect -4376 2568 -4356 2632
rect -5528 2552 -4356 2568
rect -5528 2488 -4440 2552
rect -4376 2488 -4356 2552
rect -5528 2472 -4356 2488
rect -5528 2408 -4440 2472
rect -4376 2408 -4356 2472
rect -5528 2392 -4356 2408
rect -5528 2328 -4440 2392
rect -4376 2328 -4356 2392
rect -5528 2312 -4356 2328
rect -5528 2248 -4440 2312
rect -4376 2248 -4356 2312
rect -5528 2232 -4356 2248
rect -5528 2168 -4440 2232
rect -4376 2168 -4356 2232
rect -5528 2152 -4356 2168
rect -5528 2088 -4440 2152
rect -4376 2088 -4356 2152
rect -5528 2072 -4356 2088
rect -5528 2008 -4440 2072
rect -4376 2008 -4356 2072
rect -5528 1992 -4356 2008
rect -5528 1928 -4440 1992
rect -4376 1928 -4356 1992
rect -5528 1912 -4356 1928
rect -5528 1848 -4440 1912
rect -4376 1848 -4356 1912
rect -5528 1800 -4356 1848
rect -4116 2632 -2944 2680
rect -4116 2568 -3028 2632
rect -2964 2568 -2944 2632
rect -4116 2552 -2944 2568
rect -4116 2488 -3028 2552
rect -2964 2488 -2944 2552
rect -4116 2472 -2944 2488
rect -4116 2408 -3028 2472
rect -2964 2408 -2944 2472
rect -4116 2392 -2944 2408
rect -4116 2328 -3028 2392
rect -2964 2328 -2944 2392
rect -4116 2312 -2944 2328
rect -4116 2248 -3028 2312
rect -2964 2248 -2944 2312
rect -4116 2232 -2944 2248
rect -4116 2168 -3028 2232
rect -2964 2168 -2944 2232
rect -4116 2152 -2944 2168
rect -4116 2088 -3028 2152
rect -2964 2088 -2944 2152
rect -4116 2072 -2944 2088
rect -4116 2008 -3028 2072
rect -2964 2008 -2944 2072
rect -4116 1992 -2944 2008
rect -4116 1928 -3028 1992
rect -2964 1928 -2944 1992
rect -4116 1912 -2944 1928
rect -4116 1848 -3028 1912
rect -2964 1848 -2944 1912
rect -4116 1800 -2944 1848
rect -2704 2632 -1532 2680
rect -2704 2568 -1616 2632
rect -1552 2568 -1532 2632
rect -2704 2552 -1532 2568
rect -2704 2488 -1616 2552
rect -1552 2488 -1532 2552
rect -2704 2472 -1532 2488
rect -2704 2408 -1616 2472
rect -1552 2408 -1532 2472
rect -2704 2392 -1532 2408
rect -2704 2328 -1616 2392
rect -1552 2328 -1532 2392
rect -2704 2312 -1532 2328
rect -2704 2248 -1616 2312
rect -1552 2248 -1532 2312
rect -2704 2232 -1532 2248
rect -2704 2168 -1616 2232
rect -1552 2168 -1532 2232
rect -2704 2152 -1532 2168
rect -2704 2088 -1616 2152
rect -1552 2088 -1532 2152
rect -2704 2072 -1532 2088
rect -2704 2008 -1616 2072
rect -1552 2008 -1532 2072
rect -2704 1992 -1532 2008
rect -2704 1928 -1616 1992
rect -1552 1928 -1532 1992
rect -2704 1912 -1532 1928
rect -2704 1848 -1616 1912
rect -1552 1848 -1532 1912
rect -2704 1800 -1532 1848
rect -1292 2632 -120 2680
rect -1292 2568 -204 2632
rect -140 2568 -120 2632
rect -1292 2552 -120 2568
rect -1292 2488 -204 2552
rect -140 2488 -120 2552
rect -1292 2472 -120 2488
rect -1292 2408 -204 2472
rect -140 2408 -120 2472
rect -1292 2392 -120 2408
rect -1292 2328 -204 2392
rect -140 2328 -120 2392
rect -1292 2312 -120 2328
rect -1292 2248 -204 2312
rect -140 2248 -120 2312
rect -1292 2232 -120 2248
rect -1292 2168 -204 2232
rect -140 2168 -120 2232
rect -1292 2152 -120 2168
rect -1292 2088 -204 2152
rect -140 2088 -120 2152
rect -1292 2072 -120 2088
rect -1292 2008 -204 2072
rect -140 2008 -120 2072
rect -1292 1992 -120 2008
rect -1292 1928 -204 1992
rect -140 1928 -120 1992
rect -1292 1912 -120 1928
rect -1292 1848 -204 1912
rect -140 1848 -120 1912
rect -1292 1800 -120 1848
rect 120 2632 1292 2680
rect 120 2568 1208 2632
rect 1272 2568 1292 2632
rect 120 2552 1292 2568
rect 120 2488 1208 2552
rect 1272 2488 1292 2552
rect 120 2472 1292 2488
rect 120 2408 1208 2472
rect 1272 2408 1292 2472
rect 120 2392 1292 2408
rect 120 2328 1208 2392
rect 1272 2328 1292 2392
rect 120 2312 1292 2328
rect 120 2248 1208 2312
rect 1272 2248 1292 2312
rect 120 2232 1292 2248
rect 120 2168 1208 2232
rect 1272 2168 1292 2232
rect 120 2152 1292 2168
rect 120 2088 1208 2152
rect 1272 2088 1292 2152
rect 120 2072 1292 2088
rect 120 2008 1208 2072
rect 1272 2008 1292 2072
rect 120 1992 1292 2008
rect 120 1928 1208 1992
rect 1272 1928 1292 1992
rect 120 1912 1292 1928
rect 120 1848 1208 1912
rect 1272 1848 1292 1912
rect 120 1800 1292 1848
rect 1532 2632 2704 2680
rect 1532 2568 2620 2632
rect 2684 2568 2704 2632
rect 1532 2552 2704 2568
rect 1532 2488 2620 2552
rect 2684 2488 2704 2552
rect 1532 2472 2704 2488
rect 1532 2408 2620 2472
rect 2684 2408 2704 2472
rect 1532 2392 2704 2408
rect 1532 2328 2620 2392
rect 2684 2328 2704 2392
rect 1532 2312 2704 2328
rect 1532 2248 2620 2312
rect 2684 2248 2704 2312
rect 1532 2232 2704 2248
rect 1532 2168 2620 2232
rect 2684 2168 2704 2232
rect 1532 2152 2704 2168
rect 1532 2088 2620 2152
rect 2684 2088 2704 2152
rect 1532 2072 2704 2088
rect 1532 2008 2620 2072
rect 2684 2008 2704 2072
rect 1532 1992 2704 2008
rect 1532 1928 2620 1992
rect 2684 1928 2704 1992
rect 1532 1912 2704 1928
rect 1532 1848 2620 1912
rect 2684 1848 2704 1912
rect 1532 1800 2704 1848
rect 2944 2632 4116 2680
rect 2944 2568 4032 2632
rect 4096 2568 4116 2632
rect 2944 2552 4116 2568
rect 2944 2488 4032 2552
rect 4096 2488 4116 2552
rect 2944 2472 4116 2488
rect 2944 2408 4032 2472
rect 4096 2408 4116 2472
rect 2944 2392 4116 2408
rect 2944 2328 4032 2392
rect 4096 2328 4116 2392
rect 2944 2312 4116 2328
rect 2944 2248 4032 2312
rect 4096 2248 4116 2312
rect 2944 2232 4116 2248
rect 2944 2168 4032 2232
rect 4096 2168 4116 2232
rect 2944 2152 4116 2168
rect 2944 2088 4032 2152
rect 4096 2088 4116 2152
rect 2944 2072 4116 2088
rect 2944 2008 4032 2072
rect 4096 2008 4116 2072
rect 2944 1992 4116 2008
rect 2944 1928 4032 1992
rect 4096 1928 4116 1992
rect 2944 1912 4116 1928
rect 2944 1848 4032 1912
rect 4096 1848 4116 1912
rect 2944 1800 4116 1848
rect 4356 2632 5528 2680
rect 4356 2568 5444 2632
rect 5508 2568 5528 2632
rect 4356 2552 5528 2568
rect 4356 2488 5444 2552
rect 5508 2488 5528 2552
rect 4356 2472 5528 2488
rect 4356 2408 5444 2472
rect 5508 2408 5528 2472
rect 4356 2392 5528 2408
rect 4356 2328 5444 2392
rect 5508 2328 5528 2392
rect 4356 2312 5528 2328
rect 4356 2248 5444 2312
rect 5508 2248 5528 2312
rect 4356 2232 5528 2248
rect 4356 2168 5444 2232
rect 5508 2168 5528 2232
rect 4356 2152 5528 2168
rect 4356 2088 5444 2152
rect 5508 2088 5528 2152
rect 4356 2072 5528 2088
rect 4356 2008 5444 2072
rect 5508 2008 5528 2072
rect 4356 1992 5528 2008
rect 4356 1928 5444 1992
rect 5508 1928 5528 1992
rect 4356 1912 5528 1928
rect 4356 1848 5444 1912
rect 5508 1848 5528 1912
rect 4356 1800 5528 1848
rect 5768 2632 6940 2680
rect 5768 2568 6856 2632
rect 6920 2568 6940 2632
rect 5768 2552 6940 2568
rect 5768 2488 6856 2552
rect 6920 2488 6940 2552
rect 5768 2472 6940 2488
rect 5768 2408 6856 2472
rect 6920 2408 6940 2472
rect 5768 2392 6940 2408
rect 5768 2328 6856 2392
rect 6920 2328 6940 2392
rect 5768 2312 6940 2328
rect 5768 2248 6856 2312
rect 6920 2248 6940 2312
rect 5768 2232 6940 2248
rect 5768 2168 6856 2232
rect 6920 2168 6940 2232
rect 5768 2152 6940 2168
rect 5768 2088 6856 2152
rect 6920 2088 6940 2152
rect 5768 2072 6940 2088
rect 5768 2008 6856 2072
rect 6920 2008 6940 2072
rect 5768 1992 6940 2008
rect 5768 1928 6856 1992
rect 6920 1928 6940 1992
rect 5768 1912 6940 1928
rect 5768 1848 6856 1912
rect 6920 1848 6940 1912
rect 5768 1800 6940 1848
rect 7180 2632 8352 2680
rect 7180 2568 8268 2632
rect 8332 2568 8352 2632
rect 7180 2552 8352 2568
rect 7180 2488 8268 2552
rect 8332 2488 8352 2552
rect 7180 2472 8352 2488
rect 7180 2408 8268 2472
rect 8332 2408 8352 2472
rect 7180 2392 8352 2408
rect 7180 2328 8268 2392
rect 8332 2328 8352 2392
rect 7180 2312 8352 2328
rect 7180 2248 8268 2312
rect 8332 2248 8352 2312
rect 7180 2232 8352 2248
rect 7180 2168 8268 2232
rect 8332 2168 8352 2232
rect 7180 2152 8352 2168
rect 7180 2088 8268 2152
rect 8332 2088 8352 2152
rect 7180 2072 8352 2088
rect 7180 2008 8268 2072
rect 8332 2008 8352 2072
rect 7180 1992 8352 2008
rect 7180 1928 8268 1992
rect 8332 1928 8352 1992
rect 7180 1912 8352 1928
rect 7180 1848 8268 1912
rect 8332 1848 8352 1912
rect 7180 1800 8352 1848
rect 8592 2632 9764 2680
rect 8592 2568 9680 2632
rect 9744 2568 9764 2632
rect 8592 2552 9764 2568
rect 8592 2488 9680 2552
rect 9744 2488 9764 2552
rect 8592 2472 9764 2488
rect 8592 2408 9680 2472
rect 9744 2408 9764 2472
rect 8592 2392 9764 2408
rect 8592 2328 9680 2392
rect 9744 2328 9764 2392
rect 8592 2312 9764 2328
rect 8592 2248 9680 2312
rect 9744 2248 9764 2312
rect 8592 2232 9764 2248
rect 8592 2168 9680 2232
rect 9744 2168 9764 2232
rect 8592 2152 9764 2168
rect 8592 2088 9680 2152
rect 9744 2088 9764 2152
rect 8592 2072 9764 2088
rect 8592 2008 9680 2072
rect 9744 2008 9764 2072
rect 8592 1992 9764 2008
rect 8592 1928 9680 1992
rect 9744 1928 9764 1992
rect 8592 1912 9764 1928
rect 8592 1848 9680 1912
rect 9744 1848 9764 1912
rect 8592 1800 9764 1848
rect 10004 2632 11176 2680
rect 10004 2568 11092 2632
rect 11156 2568 11176 2632
rect 10004 2552 11176 2568
rect 10004 2488 11092 2552
rect 11156 2488 11176 2552
rect 10004 2472 11176 2488
rect 10004 2408 11092 2472
rect 11156 2408 11176 2472
rect 10004 2392 11176 2408
rect 10004 2328 11092 2392
rect 11156 2328 11176 2392
rect 10004 2312 11176 2328
rect 10004 2248 11092 2312
rect 11156 2248 11176 2312
rect 10004 2232 11176 2248
rect 10004 2168 11092 2232
rect 11156 2168 11176 2232
rect 10004 2152 11176 2168
rect 10004 2088 11092 2152
rect 11156 2088 11176 2152
rect 10004 2072 11176 2088
rect 10004 2008 11092 2072
rect 11156 2008 11176 2072
rect 10004 1992 11176 2008
rect 10004 1928 11092 1992
rect 11156 1928 11176 1992
rect 10004 1912 11176 1928
rect 10004 1848 11092 1912
rect 11156 1848 11176 1912
rect 10004 1800 11176 1848
rect 11416 2632 12588 2680
rect 11416 2568 12504 2632
rect 12568 2568 12588 2632
rect 11416 2552 12588 2568
rect 11416 2488 12504 2552
rect 12568 2488 12588 2552
rect 11416 2472 12588 2488
rect 11416 2408 12504 2472
rect 12568 2408 12588 2472
rect 11416 2392 12588 2408
rect 11416 2328 12504 2392
rect 12568 2328 12588 2392
rect 11416 2312 12588 2328
rect 11416 2248 12504 2312
rect 12568 2248 12588 2312
rect 11416 2232 12588 2248
rect 11416 2168 12504 2232
rect 12568 2168 12588 2232
rect 11416 2152 12588 2168
rect 11416 2088 12504 2152
rect 12568 2088 12588 2152
rect 11416 2072 12588 2088
rect 11416 2008 12504 2072
rect 12568 2008 12588 2072
rect 11416 1992 12588 2008
rect 11416 1928 12504 1992
rect 12568 1928 12588 1992
rect 11416 1912 12588 1928
rect 11416 1848 12504 1912
rect 12568 1848 12588 1912
rect 11416 1800 12588 1848
rect 12828 2632 14000 2680
rect 12828 2568 13916 2632
rect 13980 2568 14000 2632
rect 12828 2552 14000 2568
rect 12828 2488 13916 2552
rect 13980 2488 14000 2552
rect 12828 2472 14000 2488
rect 12828 2408 13916 2472
rect 13980 2408 14000 2472
rect 12828 2392 14000 2408
rect 12828 2328 13916 2392
rect 13980 2328 14000 2392
rect 12828 2312 14000 2328
rect 12828 2248 13916 2312
rect 13980 2248 14000 2312
rect 12828 2232 14000 2248
rect 12828 2168 13916 2232
rect 13980 2168 14000 2232
rect 12828 2152 14000 2168
rect 12828 2088 13916 2152
rect 13980 2088 14000 2152
rect 12828 2072 14000 2088
rect 12828 2008 13916 2072
rect 13980 2008 14000 2072
rect 12828 1992 14000 2008
rect 12828 1928 13916 1992
rect 13980 1928 14000 1992
rect 12828 1912 14000 1928
rect 12828 1848 13916 1912
rect 13980 1848 14000 1912
rect 12828 1800 14000 1848
rect 14240 2632 15412 2680
rect 14240 2568 15328 2632
rect 15392 2568 15412 2632
rect 14240 2552 15412 2568
rect 14240 2488 15328 2552
rect 15392 2488 15412 2552
rect 14240 2472 15412 2488
rect 14240 2408 15328 2472
rect 15392 2408 15412 2472
rect 14240 2392 15412 2408
rect 14240 2328 15328 2392
rect 15392 2328 15412 2392
rect 14240 2312 15412 2328
rect 14240 2248 15328 2312
rect 15392 2248 15412 2312
rect 14240 2232 15412 2248
rect 14240 2168 15328 2232
rect 15392 2168 15412 2232
rect 14240 2152 15412 2168
rect 14240 2088 15328 2152
rect 15392 2088 15412 2152
rect 14240 2072 15412 2088
rect 14240 2008 15328 2072
rect 15392 2008 15412 2072
rect 14240 1992 15412 2008
rect 14240 1928 15328 1992
rect 15392 1928 15412 1992
rect 14240 1912 15412 1928
rect 14240 1848 15328 1912
rect 15392 1848 15412 1912
rect 14240 1800 15412 1848
rect 15652 2632 16824 2680
rect 15652 2568 16740 2632
rect 16804 2568 16824 2632
rect 15652 2552 16824 2568
rect 15652 2488 16740 2552
rect 16804 2488 16824 2552
rect 15652 2472 16824 2488
rect 15652 2408 16740 2472
rect 16804 2408 16824 2472
rect 15652 2392 16824 2408
rect 15652 2328 16740 2392
rect 16804 2328 16824 2392
rect 15652 2312 16824 2328
rect 15652 2248 16740 2312
rect 16804 2248 16824 2312
rect 15652 2232 16824 2248
rect 15652 2168 16740 2232
rect 16804 2168 16824 2232
rect 15652 2152 16824 2168
rect 15652 2088 16740 2152
rect 16804 2088 16824 2152
rect 15652 2072 16824 2088
rect 15652 2008 16740 2072
rect 16804 2008 16824 2072
rect 15652 1992 16824 2008
rect 15652 1928 16740 1992
rect 16804 1928 16824 1992
rect 15652 1912 16824 1928
rect 15652 1848 16740 1912
rect 16804 1848 16824 1912
rect 15652 1800 16824 1848
rect 17064 2632 18236 2680
rect 17064 2568 18152 2632
rect 18216 2568 18236 2632
rect 17064 2552 18236 2568
rect 17064 2488 18152 2552
rect 18216 2488 18236 2552
rect 17064 2472 18236 2488
rect 17064 2408 18152 2472
rect 18216 2408 18236 2472
rect 17064 2392 18236 2408
rect 17064 2328 18152 2392
rect 18216 2328 18236 2392
rect 17064 2312 18236 2328
rect 17064 2248 18152 2312
rect 18216 2248 18236 2312
rect 17064 2232 18236 2248
rect 17064 2168 18152 2232
rect 18216 2168 18236 2232
rect 17064 2152 18236 2168
rect 17064 2088 18152 2152
rect 18216 2088 18236 2152
rect 17064 2072 18236 2088
rect 17064 2008 18152 2072
rect 18216 2008 18236 2072
rect 17064 1992 18236 2008
rect 17064 1928 18152 1992
rect 18216 1928 18236 1992
rect 17064 1912 18236 1928
rect 17064 1848 18152 1912
rect 18216 1848 18236 1912
rect 17064 1800 18236 1848
rect 18476 2632 19648 2680
rect 18476 2568 19564 2632
rect 19628 2568 19648 2632
rect 18476 2552 19648 2568
rect 18476 2488 19564 2552
rect 19628 2488 19648 2552
rect 18476 2472 19648 2488
rect 18476 2408 19564 2472
rect 19628 2408 19648 2472
rect 18476 2392 19648 2408
rect 18476 2328 19564 2392
rect 19628 2328 19648 2392
rect 18476 2312 19648 2328
rect 18476 2248 19564 2312
rect 19628 2248 19648 2312
rect 18476 2232 19648 2248
rect 18476 2168 19564 2232
rect 19628 2168 19648 2232
rect 18476 2152 19648 2168
rect 18476 2088 19564 2152
rect 19628 2088 19648 2152
rect 18476 2072 19648 2088
rect 18476 2008 19564 2072
rect 19628 2008 19648 2072
rect 18476 1992 19648 2008
rect 18476 1928 19564 1992
rect 19628 1928 19648 1992
rect 18476 1912 19648 1928
rect 18476 1848 19564 1912
rect 19628 1848 19648 1912
rect 18476 1800 19648 1848
rect 19888 2632 21060 2680
rect 19888 2568 20976 2632
rect 21040 2568 21060 2632
rect 19888 2552 21060 2568
rect 19888 2488 20976 2552
rect 21040 2488 21060 2552
rect 19888 2472 21060 2488
rect 19888 2408 20976 2472
rect 21040 2408 21060 2472
rect 19888 2392 21060 2408
rect 19888 2328 20976 2392
rect 21040 2328 21060 2392
rect 19888 2312 21060 2328
rect 19888 2248 20976 2312
rect 21040 2248 21060 2312
rect 19888 2232 21060 2248
rect 19888 2168 20976 2232
rect 21040 2168 21060 2232
rect 19888 2152 21060 2168
rect 19888 2088 20976 2152
rect 21040 2088 21060 2152
rect 19888 2072 21060 2088
rect 19888 2008 20976 2072
rect 21040 2008 21060 2072
rect 19888 1992 21060 2008
rect 19888 1928 20976 1992
rect 21040 1928 21060 1992
rect 19888 1912 21060 1928
rect 19888 1848 20976 1912
rect 21040 1848 21060 1912
rect 19888 1800 21060 1848
rect 21300 2632 22472 2680
rect 21300 2568 22388 2632
rect 22452 2568 22472 2632
rect 21300 2552 22472 2568
rect 21300 2488 22388 2552
rect 22452 2488 22472 2552
rect 21300 2472 22472 2488
rect 21300 2408 22388 2472
rect 22452 2408 22472 2472
rect 21300 2392 22472 2408
rect 21300 2328 22388 2392
rect 22452 2328 22472 2392
rect 21300 2312 22472 2328
rect 21300 2248 22388 2312
rect 22452 2248 22472 2312
rect 21300 2232 22472 2248
rect 21300 2168 22388 2232
rect 22452 2168 22472 2232
rect 21300 2152 22472 2168
rect 21300 2088 22388 2152
rect 22452 2088 22472 2152
rect 21300 2072 22472 2088
rect 21300 2008 22388 2072
rect 22452 2008 22472 2072
rect 21300 1992 22472 2008
rect 21300 1928 22388 1992
rect 22452 1928 22472 1992
rect 21300 1912 22472 1928
rect 21300 1848 22388 1912
rect 22452 1848 22472 1912
rect 21300 1800 22472 1848
rect 22712 2632 23884 2680
rect 22712 2568 23800 2632
rect 23864 2568 23884 2632
rect 22712 2552 23884 2568
rect 22712 2488 23800 2552
rect 23864 2488 23884 2552
rect 22712 2472 23884 2488
rect 22712 2408 23800 2472
rect 23864 2408 23884 2472
rect 22712 2392 23884 2408
rect 22712 2328 23800 2392
rect 23864 2328 23884 2392
rect 22712 2312 23884 2328
rect 22712 2248 23800 2312
rect 23864 2248 23884 2312
rect 22712 2232 23884 2248
rect 22712 2168 23800 2232
rect 23864 2168 23884 2232
rect 22712 2152 23884 2168
rect 22712 2088 23800 2152
rect 23864 2088 23884 2152
rect 22712 2072 23884 2088
rect 22712 2008 23800 2072
rect 23864 2008 23884 2072
rect 22712 1992 23884 2008
rect 22712 1928 23800 1992
rect 23864 1928 23884 1992
rect 22712 1912 23884 1928
rect 22712 1848 23800 1912
rect 23864 1848 23884 1912
rect 22712 1800 23884 1848
rect -23884 1512 -22712 1560
rect -23884 1448 -22796 1512
rect -22732 1448 -22712 1512
rect -23884 1432 -22712 1448
rect -23884 1368 -22796 1432
rect -22732 1368 -22712 1432
rect -23884 1352 -22712 1368
rect -23884 1288 -22796 1352
rect -22732 1288 -22712 1352
rect -23884 1272 -22712 1288
rect -23884 1208 -22796 1272
rect -22732 1208 -22712 1272
rect -23884 1192 -22712 1208
rect -23884 1128 -22796 1192
rect -22732 1128 -22712 1192
rect -23884 1112 -22712 1128
rect -23884 1048 -22796 1112
rect -22732 1048 -22712 1112
rect -23884 1032 -22712 1048
rect -23884 968 -22796 1032
rect -22732 968 -22712 1032
rect -23884 952 -22712 968
rect -23884 888 -22796 952
rect -22732 888 -22712 952
rect -23884 872 -22712 888
rect -23884 808 -22796 872
rect -22732 808 -22712 872
rect -23884 792 -22712 808
rect -23884 728 -22796 792
rect -22732 728 -22712 792
rect -23884 680 -22712 728
rect -22472 1512 -21300 1560
rect -22472 1448 -21384 1512
rect -21320 1448 -21300 1512
rect -22472 1432 -21300 1448
rect -22472 1368 -21384 1432
rect -21320 1368 -21300 1432
rect -22472 1352 -21300 1368
rect -22472 1288 -21384 1352
rect -21320 1288 -21300 1352
rect -22472 1272 -21300 1288
rect -22472 1208 -21384 1272
rect -21320 1208 -21300 1272
rect -22472 1192 -21300 1208
rect -22472 1128 -21384 1192
rect -21320 1128 -21300 1192
rect -22472 1112 -21300 1128
rect -22472 1048 -21384 1112
rect -21320 1048 -21300 1112
rect -22472 1032 -21300 1048
rect -22472 968 -21384 1032
rect -21320 968 -21300 1032
rect -22472 952 -21300 968
rect -22472 888 -21384 952
rect -21320 888 -21300 952
rect -22472 872 -21300 888
rect -22472 808 -21384 872
rect -21320 808 -21300 872
rect -22472 792 -21300 808
rect -22472 728 -21384 792
rect -21320 728 -21300 792
rect -22472 680 -21300 728
rect -21060 1512 -19888 1560
rect -21060 1448 -19972 1512
rect -19908 1448 -19888 1512
rect -21060 1432 -19888 1448
rect -21060 1368 -19972 1432
rect -19908 1368 -19888 1432
rect -21060 1352 -19888 1368
rect -21060 1288 -19972 1352
rect -19908 1288 -19888 1352
rect -21060 1272 -19888 1288
rect -21060 1208 -19972 1272
rect -19908 1208 -19888 1272
rect -21060 1192 -19888 1208
rect -21060 1128 -19972 1192
rect -19908 1128 -19888 1192
rect -21060 1112 -19888 1128
rect -21060 1048 -19972 1112
rect -19908 1048 -19888 1112
rect -21060 1032 -19888 1048
rect -21060 968 -19972 1032
rect -19908 968 -19888 1032
rect -21060 952 -19888 968
rect -21060 888 -19972 952
rect -19908 888 -19888 952
rect -21060 872 -19888 888
rect -21060 808 -19972 872
rect -19908 808 -19888 872
rect -21060 792 -19888 808
rect -21060 728 -19972 792
rect -19908 728 -19888 792
rect -21060 680 -19888 728
rect -19648 1512 -18476 1560
rect -19648 1448 -18560 1512
rect -18496 1448 -18476 1512
rect -19648 1432 -18476 1448
rect -19648 1368 -18560 1432
rect -18496 1368 -18476 1432
rect -19648 1352 -18476 1368
rect -19648 1288 -18560 1352
rect -18496 1288 -18476 1352
rect -19648 1272 -18476 1288
rect -19648 1208 -18560 1272
rect -18496 1208 -18476 1272
rect -19648 1192 -18476 1208
rect -19648 1128 -18560 1192
rect -18496 1128 -18476 1192
rect -19648 1112 -18476 1128
rect -19648 1048 -18560 1112
rect -18496 1048 -18476 1112
rect -19648 1032 -18476 1048
rect -19648 968 -18560 1032
rect -18496 968 -18476 1032
rect -19648 952 -18476 968
rect -19648 888 -18560 952
rect -18496 888 -18476 952
rect -19648 872 -18476 888
rect -19648 808 -18560 872
rect -18496 808 -18476 872
rect -19648 792 -18476 808
rect -19648 728 -18560 792
rect -18496 728 -18476 792
rect -19648 680 -18476 728
rect -18236 1512 -17064 1560
rect -18236 1448 -17148 1512
rect -17084 1448 -17064 1512
rect -18236 1432 -17064 1448
rect -18236 1368 -17148 1432
rect -17084 1368 -17064 1432
rect -18236 1352 -17064 1368
rect -18236 1288 -17148 1352
rect -17084 1288 -17064 1352
rect -18236 1272 -17064 1288
rect -18236 1208 -17148 1272
rect -17084 1208 -17064 1272
rect -18236 1192 -17064 1208
rect -18236 1128 -17148 1192
rect -17084 1128 -17064 1192
rect -18236 1112 -17064 1128
rect -18236 1048 -17148 1112
rect -17084 1048 -17064 1112
rect -18236 1032 -17064 1048
rect -18236 968 -17148 1032
rect -17084 968 -17064 1032
rect -18236 952 -17064 968
rect -18236 888 -17148 952
rect -17084 888 -17064 952
rect -18236 872 -17064 888
rect -18236 808 -17148 872
rect -17084 808 -17064 872
rect -18236 792 -17064 808
rect -18236 728 -17148 792
rect -17084 728 -17064 792
rect -18236 680 -17064 728
rect -16824 1512 -15652 1560
rect -16824 1448 -15736 1512
rect -15672 1448 -15652 1512
rect -16824 1432 -15652 1448
rect -16824 1368 -15736 1432
rect -15672 1368 -15652 1432
rect -16824 1352 -15652 1368
rect -16824 1288 -15736 1352
rect -15672 1288 -15652 1352
rect -16824 1272 -15652 1288
rect -16824 1208 -15736 1272
rect -15672 1208 -15652 1272
rect -16824 1192 -15652 1208
rect -16824 1128 -15736 1192
rect -15672 1128 -15652 1192
rect -16824 1112 -15652 1128
rect -16824 1048 -15736 1112
rect -15672 1048 -15652 1112
rect -16824 1032 -15652 1048
rect -16824 968 -15736 1032
rect -15672 968 -15652 1032
rect -16824 952 -15652 968
rect -16824 888 -15736 952
rect -15672 888 -15652 952
rect -16824 872 -15652 888
rect -16824 808 -15736 872
rect -15672 808 -15652 872
rect -16824 792 -15652 808
rect -16824 728 -15736 792
rect -15672 728 -15652 792
rect -16824 680 -15652 728
rect -15412 1512 -14240 1560
rect -15412 1448 -14324 1512
rect -14260 1448 -14240 1512
rect -15412 1432 -14240 1448
rect -15412 1368 -14324 1432
rect -14260 1368 -14240 1432
rect -15412 1352 -14240 1368
rect -15412 1288 -14324 1352
rect -14260 1288 -14240 1352
rect -15412 1272 -14240 1288
rect -15412 1208 -14324 1272
rect -14260 1208 -14240 1272
rect -15412 1192 -14240 1208
rect -15412 1128 -14324 1192
rect -14260 1128 -14240 1192
rect -15412 1112 -14240 1128
rect -15412 1048 -14324 1112
rect -14260 1048 -14240 1112
rect -15412 1032 -14240 1048
rect -15412 968 -14324 1032
rect -14260 968 -14240 1032
rect -15412 952 -14240 968
rect -15412 888 -14324 952
rect -14260 888 -14240 952
rect -15412 872 -14240 888
rect -15412 808 -14324 872
rect -14260 808 -14240 872
rect -15412 792 -14240 808
rect -15412 728 -14324 792
rect -14260 728 -14240 792
rect -15412 680 -14240 728
rect -14000 1512 -12828 1560
rect -14000 1448 -12912 1512
rect -12848 1448 -12828 1512
rect -14000 1432 -12828 1448
rect -14000 1368 -12912 1432
rect -12848 1368 -12828 1432
rect -14000 1352 -12828 1368
rect -14000 1288 -12912 1352
rect -12848 1288 -12828 1352
rect -14000 1272 -12828 1288
rect -14000 1208 -12912 1272
rect -12848 1208 -12828 1272
rect -14000 1192 -12828 1208
rect -14000 1128 -12912 1192
rect -12848 1128 -12828 1192
rect -14000 1112 -12828 1128
rect -14000 1048 -12912 1112
rect -12848 1048 -12828 1112
rect -14000 1032 -12828 1048
rect -14000 968 -12912 1032
rect -12848 968 -12828 1032
rect -14000 952 -12828 968
rect -14000 888 -12912 952
rect -12848 888 -12828 952
rect -14000 872 -12828 888
rect -14000 808 -12912 872
rect -12848 808 -12828 872
rect -14000 792 -12828 808
rect -14000 728 -12912 792
rect -12848 728 -12828 792
rect -14000 680 -12828 728
rect -12588 1512 -11416 1560
rect -12588 1448 -11500 1512
rect -11436 1448 -11416 1512
rect -12588 1432 -11416 1448
rect -12588 1368 -11500 1432
rect -11436 1368 -11416 1432
rect -12588 1352 -11416 1368
rect -12588 1288 -11500 1352
rect -11436 1288 -11416 1352
rect -12588 1272 -11416 1288
rect -12588 1208 -11500 1272
rect -11436 1208 -11416 1272
rect -12588 1192 -11416 1208
rect -12588 1128 -11500 1192
rect -11436 1128 -11416 1192
rect -12588 1112 -11416 1128
rect -12588 1048 -11500 1112
rect -11436 1048 -11416 1112
rect -12588 1032 -11416 1048
rect -12588 968 -11500 1032
rect -11436 968 -11416 1032
rect -12588 952 -11416 968
rect -12588 888 -11500 952
rect -11436 888 -11416 952
rect -12588 872 -11416 888
rect -12588 808 -11500 872
rect -11436 808 -11416 872
rect -12588 792 -11416 808
rect -12588 728 -11500 792
rect -11436 728 -11416 792
rect -12588 680 -11416 728
rect -11176 1512 -10004 1560
rect -11176 1448 -10088 1512
rect -10024 1448 -10004 1512
rect -11176 1432 -10004 1448
rect -11176 1368 -10088 1432
rect -10024 1368 -10004 1432
rect -11176 1352 -10004 1368
rect -11176 1288 -10088 1352
rect -10024 1288 -10004 1352
rect -11176 1272 -10004 1288
rect -11176 1208 -10088 1272
rect -10024 1208 -10004 1272
rect -11176 1192 -10004 1208
rect -11176 1128 -10088 1192
rect -10024 1128 -10004 1192
rect -11176 1112 -10004 1128
rect -11176 1048 -10088 1112
rect -10024 1048 -10004 1112
rect -11176 1032 -10004 1048
rect -11176 968 -10088 1032
rect -10024 968 -10004 1032
rect -11176 952 -10004 968
rect -11176 888 -10088 952
rect -10024 888 -10004 952
rect -11176 872 -10004 888
rect -11176 808 -10088 872
rect -10024 808 -10004 872
rect -11176 792 -10004 808
rect -11176 728 -10088 792
rect -10024 728 -10004 792
rect -11176 680 -10004 728
rect -9764 1512 -8592 1560
rect -9764 1448 -8676 1512
rect -8612 1448 -8592 1512
rect -9764 1432 -8592 1448
rect -9764 1368 -8676 1432
rect -8612 1368 -8592 1432
rect -9764 1352 -8592 1368
rect -9764 1288 -8676 1352
rect -8612 1288 -8592 1352
rect -9764 1272 -8592 1288
rect -9764 1208 -8676 1272
rect -8612 1208 -8592 1272
rect -9764 1192 -8592 1208
rect -9764 1128 -8676 1192
rect -8612 1128 -8592 1192
rect -9764 1112 -8592 1128
rect -9764 1048 -8676 1112
rect -8612 1048 -8592 1112
rect -9764 1032 -8592 1048
rect -9764 968 -8676 1032
rect -8612 968 -8592 1032
rect -9764 952 -8592 968
rect -9764 888 -8676 952
rect -8612 888 -8592 952
rect -9764 872 -8592 888
rect -9764 808 -8676 872
rect -8612 808 -8592 872
rect -9764 792 -8592 808
rect -9764 728 -8676 792
rect -8612 728 -8592 792
rect -9764 680 -8592 728
rect -8352 1512 -7180 1560
rect -8352 1448 -7264 1512
rect -7200 1448 -7180 1512
rect -8352 1432 -7180 1448
rect -8352 1368 -7264 1432
rect -7200 1368 -7180 1432
rect -8352 1352 -7180 1368
rect -8352 1288 -7264 1352
rect -7200 1288 -7180 1352
rect -8352 1272 -7180 1288
rect -8352 1208 -7264 1272
rect -7200 1208 -7180 1272
rect -8352 1192 -7180 1208
rect -8352 1128 -7264 1192
rect -7200 1128 -7180 1192
rect -8352 1112 -7180 1128
rect -8352 1048 -7264 1112
rect -7200 1048 -7180 1112
rect -8352 1032 -7180 1048
rect -8352 968 -7264 1032
rect -7200 968 -7180 1032
rect -8352 952 -7180 968
rect -8352 888 -7264 952
rect -7200 888 -7180 952
rect -8352 872 -7180 888
rect -8352 808 -7264 872
rect -7200 808 -7180 872
rect -8352 792 -7180 808
rect -8352 728 -7264 792
rect -7200 728 -7180 792
rect -8352 680 -7180 728
rect -6940 1512 -5768 1560
rect -6940 1448 -5852 1512
rect -5788 1448 -5768 1512
rect -6940 1432 -5768 1448
rect -6940 1368 -5852 1432
rect -5788 1368 -5768 1432
rect -6940 1352 -5768 1368
rect -6940 1288 -5852 1352
rect -5788 1288 -5768 1352
rect -6940 1272 -5768 1288
rect -6940 1208 -5852 1272
rect -5788 1208 -5768 1272
rect -6940 1192 -5768 1208
rect -6940 1128 -5852 1192
rect -5788 1128 -5768 1192
rect -6940 1112 -5768 1128
rect -6940 1048 -5852 1112
rect -5788 1048 -5768 1112
rect -6940 1032 -5768 1048
rect -6940 968 -5852 1032
rect -5788 968 -5768 1032
rect -6940 952 -5768 968
rect -6940 888 -5852 952
rect -5788 888 -5768 952
rect -6940 872 -5768 888
rect -6940 808 -5852 872
rect -5788 808 -5768 872
rect -6940 792 -5768 808
rect -6940 728 -5852 792
rect -5788 728 -5768 792
rect -6940 680 -5768 728
rect -5528 1512 -4356 1560
rect -5528 1448 -4440 1512
rect -4376 1448 -4356 1512
rect -5528 1432 -4356 1448
rect -5528 1368 -4440 1432
rect -4376 1368 -4356 1432
rect -5528 1352 -4356 1368
rect -5528 1288 -4440 1352
rect -4376 1288 -4356 1352
rect -5528 1272 -4356 1288
rect -5528 1208 -4440 1272
rect -4376 1208 -4356 1272
rect -5528 1192 -4356 1208
rect -5528 1128 -4440 1192
rect -4376 1128 -4356 1192
rect -5528 1112 -4356 1128
rect -5528 1048 -4440 1112
rect -4376 1048 -4356 1112
rect -5528 1032 -4356 1048
rect -5528 968 -4440 1032
rect -4376 968 -4356 1032
rect -5528 952 -4356 968
rect -5528 888 -4440 952
rect -4376 888 -4356 952
rect -5528 872 -4356 888
rect -5528 808 -4440 872
rect -4376 808 -4356 872
rect -5528 792 -4356 808
rect -5528 728 -4440 792
rect -4376 728 -4356 792
rect -5528 680 -4356 728
rect -4116 1512 -2944 1560
rect -4116 1448 -3028 1512
rect -2964 1448 -2944 1512
rect -4116 1432 -2944 1448
rect -4116 1368 -3028 1432
rect -2964 1368 -2944 1432
rect -4116 1352 -2944 1368
rect -4116 1288 -3028 1352
rect -2964 1288 -2944 1352
rect -4116 1272 -2944 1288
rect -4116 1208 -3028 1272
rect -2964 1208 -2944 1272
rect -4116 1192 -2944 1208
rect -4116 1128 -3028 1192
rect -2964 1128 -2944 1192
rect -4116 1112 -2944 1128
rect -4116 1048 -3028 1112
rect -2964 1048 -2944 1112
rect -4116 1032 -2944 1048
rect -4116 968 -3028 1032
rect -2964 968 -2944 1032
rect -4116 952 -2944 968
rect -4116 888 -3028 952
rect -2964 888 -2944 952
rect -4116 872 -2944 888
rect -4116 808 -3028 872
rect -2964 808 -2944 872
rect -4116 792 -2944 808
rect -4116 728 -3028 792
rect -2964 728 -2944 792
rect -4116 680 -2944 728
rect -2704 1512 -1532 1560
rect -2704 1448 -1616 1512
rect -1552 1448 -1532 1512
rect -2704 1432 -1532 1448
rect -2704 1368 -1616 1432
rect -1552 1368 -1532 1432
rect -2704 1352 -1532 1368
rect -2704 1288 -1616 1352
rect -1552 1288 -1532 1352
rect -2704 1272 -1532 1288
rect -2704 1208 -1616 1272
rect -1552 1208 -1532 1272
rect -2704 1192 -1532 1208
rect -2704 1128 -1616 1192
rect -1552 1128 -1532 1192
rect -2704 1112 -1532 1128
rect -2704 1048 -1616 1112
rect -1552 1048 -1532 1112
rect -2704 1032 -1532 1048
rect -2704 968 -1616 1032
rect -1552 968 -1532 1032
rect -2704 952 -1532 968
rect -2704 888 -1616 952
rect -1552 888 -1532 952
rect -2704 872 -1532 888
rect -2704 808 -1616 872
rect -1552 808 -1532 872
rect -2704 792 -1532 808
rect -2704 728 -1616 792
rect -1552 728 -1532 792
rect -2704 680 -1532 728
rect -1292 1512 -120 1560
rect -1292 1448 -204 1512
rect -140 1448 -120 1512
rect -1292 1432 -120 1448
rect -1292 1368 -204 1432
rect -140 1368 -120 1432
rect -1292 1352 -120 1368
rect -1292 1288 -204 1352
rect -140 1288 -120 1352
rect -1292 1272 -120 1288
rect -1292 1208 -204 1272
rect -140 1208 -120 1272
rect -1292 1192 -120 1208
rect -1292 1128 -204 1192
rect -140 1128 -120 1192
rect -1292 1112 -120 1128
rect -1292 1048 -204 1112
rect -140 1048 -120 1112
rect -1292 1032 -120 1048
rect -1292 968 -204 1032
rect -140 968 -120 1032
rect -1292 952 -120 968
rect -1292 888 -204 952
rect -140 888 -120 952
rect -1292 872 -120 888
rect -1292 808 -204 872
rect -140 808 -120 872
rect -1292 792 -120 808
rect -1292 728 -204 792
rect -140 728 -120 792
rect -1292 680 -120 728
rect 120 1512 1292 1560
rect 120 1448 1208 1512
rect 1272 1448 1292 1512
rect 120 1432 1292 1448
rect 120 1368 1208 1432
rect 1272 1368 1292 1432
rect 120 1352 1292 1368
rect 120 1288 1208 1352
rect 1272 1288 1292 1352
rect 120 1272 1292 1288
rect 120 1208 1208 1272
rect 1272 1208 1292 1272
rect 120 1192 1292 1208
rect 120 1128 1208 1192
rect 1272 1128 1292 1192
rect 120 1112 1292 1128
rect 120 1048 1208 1112
rect 1272 1048 1292 1112
rect 120 1032 1292 1048
rect 120 968 1208 1032
rect 1272 968 1292 1032
rect 120 952 1292 968
rect 120 888 1208 952
rect 1272 888 1292 952
rect 120 872 1292 888
rect 120 808 1208 872
rect 1272 808 1292 872
rect 120 792 1292 808
rect 120 728 1208 792
rect 1272 728 1292 792
rect 120 680 1292 728
rect 1532 1512 2704 1560
rect 1532 1448 2620 1512
rect 2684 1448 2704 1512
rect 1532 1432 2704 1448
rect 1532 1368 2620 1432
rect 2684 1368 2704 1432
rect 1532 1352 2704 1368
rect 1532 1288 2620 1352
rect 2684 1288 2704 1352
rect 1532 1272 2704 1288
rect 1532 1208 2620 1272
rect 2684 1208 2704 1272
rect 1532 1192 2704 1208
rect 1532 1128 2620 1192
rect 2684 1128 2704 1192
rect 1532 1112 2704 1128
rect 1532 1048 2620 1112
rect 2684 1048 2704 1112
rect 1532 1032 2704 1048
rect 1532 968 2620 1032
rect 2684 968 2704 1032
rect 1532 952 2704 968
rect 1532 888 2620 952
rect 2684 888 2704 952
rect 1532 872 2704 888
rect 1532 808 2620 872
rect 2684 808 2704 872
rect 1532 792 2704 808
rect 1532 728 2620 792
rect 2684 728 2704 792
rect 1532 680 2704 728
rect 2944 1512 4116 1560
rect 2944 1448 4032 1512
rect 4096 1448 4116 1512
rect 2944 1432 4116 1448
rect 2944 1368 4032 1432
rect 4096 1368 4116 1432
rect 2944 1352 4116 1368
rect 2944 1288 4032 1352
rect 4096 1288 4116 1352
rect 2944 1272 4116 1288
rect 2944 1208 4032 1272
rect 4096 1208 4116 1272
rect 2944 1192 4116 1208
rect 2944 1128 4032 1192
rect 4096 1128 4116 1192
rect 2944 1112 4116 1128
rect 2944 1048 4032 1112
rect 4096 1048 4116 1112
rect 2944 1032 4116 1048
rect 2944 968 4032 1032
rect 4096 968 4116 1032
rect 2944 952 4116 968
rect 2944 888 4032 952
rect 4096 888 4116 952
rect 2944 872 4116 888
rect 2944 808 4032 872
rect 4096 808 4116 872
rect 2944 792 4116 808
rect 2944 728 4032 792
rect 4096 728 4116 792
rect 2944 680 4116 728
rect 4356 1512 5528 1560
rect 4356 1448 5444 1512
rect 5508 1448 5528 1512
rect 4356 1432 5528 1448
rect 4356 1368 5444 1432
rect 5508 1368 5528 1432
rect 4356 1352 5528 1368
rect 4356 1288 5444 1352
rect 5508 1288 5528 1352
rect 4356 1272 5528 1288
rect 4356 1208 5444 1272
rect 5508 1208 5528 1272
rect 4356 1192 5528 1208
rect 4356 1128 5444 1192
rect 5508 1128 5528 1192
rect 4356 1112 5528 1128
rect 4356 1048 5444 1112
rect 5508 1048 5528 1112
rect 4356 1032 5528 1048
rect 4356 968 5444 1032
rect 5508 968 5528 1032
rect 4356 952 5528 968
rect 4356 888 5444 952
rect 5508 888 5528 952
rect 4356 872 5528 888
rect 4356 808 5444 872
rect 5508 808 5528 872
rect 4356 792 5528 808
rect 4356 728 5444 792
rect 5508 728 5528 792
rect 4356 680 5528 728
rect 5768 1512 6940 1560
rect 5768 1448 6856 1512
rect 6920 1448 6940 1512
rect 5768 1432 6940 1448
rect 5768 1368 6856 1432
rect 6920 1368 6940 1432
rect 5768 1352 6940 1368
rect 5768 1288 6856 1352
rect 6920 1288 6940 1352
rect 5768 1272 6940 1288
rect 5768 1208 6856 1272
rect 6920 1208 6940 1272
rect 5768 1192 6940 1208
rect 5768 1128 6856 1192
rect 6920 1128 6940 1192
rect 5768 1112 6940 1128
rect 5768 1048 6856 1112
rect 6920 1048 6940 1112
rect 5768 1032 6940 1048
rect 5768 968 6856 1032
rect 6920 968 6940 1032
rect 5768 952 6940 968
rect 5768 888 6856 952
rect 6920 888 6940 952
rect 5768 872 6940 888
rect 5768 808 6856 872
rect 6920 808 6940 872
rect 5768 792 6940 808
rect 5768 728 6856 792
rect 6920 728 6940 792
rect 5768 680 6940 728
rect 7180 1512 8352 1560
rect 7180 1448 8268 1512
rect 8332 1448 8352 1512
rect 7180 1432 8352 1448
rect 7180 1368 8268 1432
rect 8332 1368 8352 1432
rect 7180 1352 8352 1368
rect 7180 1288 8268 1352
rect 8332 1288 8352 1352
rect 7180 1272 8352 1288
rect 7180 1208 8268 1272
rect 8332 1208 8352 1272
rect 7180 1192 8352 1208
rect 7180 1128 8268 1192
rect 8332 1128 8352 1192
rect 7180 1112 8352 1128
rect 7180 1048 8268 1112
rect 8332 1048 8352 1112
rect 7180 1032 8352 1048
rect 7180 968 8268 1032
rect 8332 968 8352 1032
rect 7180 952 8352 968
rect 7180 888 8268 952
rect 8332 888 8352 952
rect 7180 872 8352 888
rect 7180 808 8268 872
rect 8332 808 8352 872
rect 7180 792 8352 808
rect 7180 728 8268 792
rect 8332 728 8352 792
rect 7180 680 8352 728
rect 8592 1512 9764 1560
rect 8592 1448 9680 1512
rect 9744 1448 9764 1512
rect 8592 1432 9764 1448
rect 8592 1368 9680 1432
rect 9744 1368 9764 1432
rect 8592 1352 9764 1368
rect 8592 1288 9680 1352
rect 9744 1288 9764 1352
rect 8592 1272 9764 1288
rect 8592 1208 9680 1272
rect 9744 1208 9764 1272
rect 8592 1192 9764 1208
rect 8592 1128 9680 1192
rect 9744 1128 9764 1192
rect 8592 1112 9764 1128
rect 8592 1048 9680 1112
rect 9744 1048 9764 1112
rect 8592 1032 9764 1048
rect 8592 968 9680 1032
rect 9744 968 9764 1032
rect 8592 952 9764 968
rect 8592 888 9680 952
rect 9744 888 9764 952
rect 8592 872 9764 888
rect 8592 808 9680 872
rect 9744 808 9764 872
rect 8592 792 9764 808
rect 8592 728 9680 792
rect 9744 728 9764 792
rect 8592 680 9764 728
rect 10004 1512 11176 1560
rect 10004 1448 11092 1512
rect 11156 1448 11176 1512
rect 10004 1432 11176 1448
rect 10004 1368 11092 1432
rect 11156 1368 11176 1432
rect 10004 1352 11176 1368
rect 10004 1288 11092 1352
rect 11156 1288 11176 1352
rect 10004 1272 11176 1288
rect 10004 1208 11092 1272
rect 11156 1208 11176 1272
rect 10004 1192 11176 1208
rect 10004 1128 11092 1192
rect 11156 1128 11176 1192
rect 10004 1112 11176 1128
rect 10004 1048 11092 1112
rect 11156 1048 11176 1112
rect 10004 1032 11176 1048
rect 10004 968 11092 1032
rect 11156 968 11176 1032
rect 10004 952 11176 968
rect 10004 888 11092 952
rect 11156 888 11176 952
rect 10004 872 11176 888
rect 10004 808 11092 872
rect 11156 808 11176 872
rect 10004 792 11176 808
rect 10004 728 11092 792
rect 11156 728 11176 792
rect 10004 680 11176 728
rect 11416 1512 12588 1560
rect 11416 1448 12504 1512
rect 12568 1448 12588 1512
rect 11416 1432 12588 1448
rect 11416 1368 12504 1432
rect 12568 1368 12588 1432
rect 11416 1352 12588 1368
rect 11416 1288 12504 1352
rect 12568 1288 12588 1352
rect 11416 1272 12588 1288
rect 11416 1208 12504 1272
rect 12568 1208 12588 1272
rect 11416 1192 12588 1208
rect 11416 1128 12504 1192
rect 12568 1128 12588 1192
rect 11416 1112 12588 1128
rect 11416 1048 12504 1112
rect 12568 1048 12588 1112
rect 11416 1032 12588 1048
rect 11416 968 12504 1032
rect 12568 968 12588 1032
rect 11416 952 12588 968
rect 11416 888 12504 952
rect 12568 888 12588 952
rect 11416 872 12588 888
rect 11416 808 12504 872
rect 12568 808 12588 872
rect 11416 792 12588 808
rect 11416 728 12504 792
rect 12568 728 12588 792
rect 11416 680 12588 728
rect 12828 1512 14000 1560
rect 12828 1448 13916 1512
rect 13980 1448 14000 1512
rect 12828 1432 14000 1448
rect 12828 1368 13916 1432
rect 13980 1368 14000 1432
rect 12828 1352 14000 1368
rect 12828 1288 13916 1352
rect 13980 1288 14000 1352
rect 12828 1272 14000 1288
rect 12828 1208 13916 1272
rect 13980 1208 14000 1272
rect 12828 1192 14000 1208
rect 12828 1128 13916 1192
rect 13980 1128 14000 1192
rect 12828 1112 14000 1128
rect 12828 1048 13916 1112
rect 13980 1048 14000 1112
rect 12828 1032 14000 1048
rect 12828 968 13916 1032
rect 13980 968 14000 1032
rect 12828 952 14000 968
rect 12828 888 13916 952
rect 13980 888 14000 952
rect 12828 872 14000 888
rect 12828 808 13916 872
rect 13980 808 14000 872
rect 12828 792 14000 808
rect 12828 728 13916 792
rect 13980 728 14000 792
rect 12828 680 14000 728
rect 14240 1512 15412 1560
rect 14240 1448 15328 1512
rect 15392 1448 15412 1512
rect 14240 1432 15412 1448
rect 14240 1368 15328 1432
rect 15392 1368 15412 1432
rect 14240 1352 15412 1368
rect 14240 1288 15328 1352
rect 15392 1288 15412 1352
rect 14240 1272 15412 1288
rect 14240 1208 15328 1272
rect 15392 1208 15412 1272
rect 14240 1192 15412 1208
rect 14240 1128 15328 1192
rect 15392 1128 15412 1192
rect 14240 1112 15412 1128
rect 14240 1048 15328 1112
rect 15392 1048 15412 1112
rect 14240 1032 15412 1048
rect 14240 968 15328 1032
rect 15392 968 15412 1032
rect 14240 952 15412 968
rect 14240 888 15328 952
rect 15392 888 15412 952
rect 14240 872 15412 888
rect 14240 808 15328 872
rect 15392 808 15412 872
rect 14240 792 15412 808
rect 14240 728 15328 792
rect 15392 728 15412 792
rect 14240 680 15412 728
rect 15652 1512 16824 1560
rect 15652 1448 16740 1512
rect 16804 1448 16824 1512
rect 15652 1432 16824 1448
rect 15652 1368 16740 1432
rect 16804 1368 16824 1432
rect 15652 1352 16824 1368
rect 15652 1288 16740 1352
rect 16804 1288 16824 1352
rect 15652 1272 16824 1288
rect 15652 1208 16740 1272
rect 16804 1208 16824 1272
rect 15652 1192 16824 1208
rect 15652 1128 16740 1192
rect 16804 1128 16824 1192
rect 15652 1112 16824 1128
rect 15652 1048 16740 1112
rect 16804 1048 16824 1112
rect 15652 1032 16824 1048
rect 15652 968 16740 1032
rect 16804 968 16824 1032
rect 15652 952 16824 968
rect 15652 888 16740 952
rect 16804 888 16824 952
rect 15652 872 16824 888
rect 15652 808 16740 872
rect 16804 808 16824 872
rect 15652 792 16824 808
rect 15652 728 16740 792
rect 16804 728 16824 792
rect 15652 680 16824 728
rect 17064 1512 18236 1560
rect 17064 1448 18152 1512
rect 18216 1448 18236 1512
rect 17064 1432 18236 1448
rect 17064 1368 18152 1432
rect 18216 1368 18236 1432
rect 17064 1352 18236 1368
rect 17064 1288 18152 1352
rect 18216 1288 18236 1352
rect 17064 1272 18236 1288
rect 17064 1208 18152 1272
rect 18216 1208 18236 1272
rect 17064 1192 18236 1208
rect 17064 1128 18152 1192
rect 18216 1128 18236 1192
rect 17064 1112 18236 1128
rect 17064 1048 18152 1112
rect 18216 1048 18236 1112
rect 17064 1032 18236 1048
rect 17064 968 18152 1032
rect 18216 968 18236 1032
rect 17064 952 18236 968
rect 17064 888 18152 952
rect 18216 888 18236 952
rect 17064 872 18236 888
rect 17064 808 18152 872
rect 18216 808 18236 872
rect 17064 792 18236 808
rect 17064 728 18152 792
rect 18216 728 18236 792
rect 17064 680 18236 728
rect 18476 1512 19648 1560
rect 18476 1448 19564 1512
rect 19628 1448 19648 1512
rect 18476 1432 19648 1448
rect 18476 1368 19564 1432
rect 19628 1368 19648 1432
rect 18476 1352 19648 1368
rect 18476 1288 19564 1352
rect 19628 1288 19648 1352
rect 18476 1272 19648 1288
rect 18476 1208 19564 1272
rect 19628 1208 19648 1272
rect 18476 1192 19648 1208
rect 18476 1128 19564 1192
rect 19628 1128 19648 1192
rect 18476 1112 19648 1128
rect 18476 1048 19564 1112
rect 19628 1048 19648 1112
rect 18476 1032 19648 1048
rect 18476 968 19564 1032
rect 19628 968 19648 1032
rect 18476 952 19648 968
rect 18476 888 19564 952
rect 19628 888 19648 952
rect 18476 872 19648 888
rect 18476 808 19564 872
rect 19628 808 19648 872
rect 18476 792 19648 808
rect 18476 728 19564 792
rect 19628 728 19648 792
rect 18476 680 19648 728
rect 19888 1512 21060 1560
rect 19888 1448 20976 1512
rect 21040 1448 21060 1512
rect 19888 1432 21060 1448
rect 19888 1368 20976 1432
rect 21040 1368 21060 1432
rect 19888 1352 21060 1368
rect 19888 1288 20976 1352
rect 21040 1288 21060 1352
rect 19888 1272 21060 1288
rect 19888 1208 20976 1272
rect 21040 1208 21060 1272
rect 19888 1192 21060 1208
rect 19888 1128 20976 1192
rect 21040 1128 21060 1192
rect 19888 1112 21060 1128
rect 19888 1048 20976 1112
rect 21040 1048 21060 1112
rect 19888 1032 21060 1048
rect 19888 968 20976 1032
rect 21040 968 21060 1032
rect 19888 952 21060 968
rect 19888 888 20976 952
rect 21040 888 21060 952
rect 19888 872 21060 888
rect 19888 808 20976 872
rect 21040 808 21060 872
rect 19888 792 21060 808
rect 19888 728 20976 792
rect 21040 728 21060 792
rect 19888 680 21060 728
rect 21300 1512 22472 1560
rect 21300 1448 22388 1512
rect 22452 1448 22472 1512
rect 21300 1432 22472 1448
rect 21300 1368 22388 1432
rect 22452 1368 22472 1432
rect 21300 1352 22472 1368
rect 21300 1288 22388 1352
rect 22452 1288 22472 1352
rect 21300 1272 22472 1288
rect 21300 1208 22388 1272
rect 22452 1208 22472 1272
rect 21300 1192 22472 1208
rect 21300 1128 22388 1192
rect 22452 1128 22472 1192
rect 21300 1112 22472 1128
rect 21300 1048 22388 1112
rect 22452 1048 22472 1112
rect 21300 1032 22472 1048
rect 21300 968 22388 1032
rect 22452 968 22472 1032
rect 21300 952 22472 968
rect 21300 888 22388 952
rect 22452 888 22472 952
rect 21300 872 22472 888
rect 21300 808 22388 872
rect 22452 808 22472 872
rect 21300 792 22472 808
rect 21300 728 22388 792
rect 22452 728 22472 792
rect 21300 680 22472 728
rect 22712 1512 23884 1560
rect 22712 1448 23800 1512
rect 23864 1448 23884 1512
rect 22712 1432 23884 1448
rect 22712 1368 23800 1432
rect 23864 1368 23884 1432
rect 22712 1352 23884 1368
rect 22712 1288 23800 1352
rect 23864 1288 23884 1352
rect 22712 1272 23884 1288
rect 22712 1208 23800 1272
rect 23864 1208 23884 1272
rect 22712 1192 23884 1208
rect 22712 1128 23800 1192
rect 23864 1128 23884 1192
rect 22712 1112 23884 1128
rect 22712 1048 23800 1112
rect 23864 1048 23884 1112
rect 22712 1032 23884 1048
rect 22712 968 23800 1032
rect 23864 968 23884 1032
rect 22712 952 23884 968
rect 22712 888 23800 952
rect 23864 888 23884 952
rect 22712 872 23884 888
rect 22712 808 23800 872
rect 23864 808 23884 872
rect 22712 792 23884 808
rect 22712 728 23800 792
rect 23864 728 23884 792
rect 22712 680 23884 728
rect -23884 392 -22712 440
rect -23884 328 -22796 392
rect -22732 328 -22712 392
rect -23884 312 -22712 328
rect -23884 248 -22796 312
rect -22732 248 -22712 312
rect -23884 232 -22712 248
rect -23884 168 -22796 232
rect -22732 168 -22712 232
rect -23884 152 -22712 168
rect -23884 88 -22796 152
rect -22732 88 -22712 152
rect -23884 72 -22712 88
rect -23884 8 -22796 72
rect -22732 8 -22712 72
rect -23884 -8 -22712 8
rect -23884 -72 -22796 -8
rect -22732 -72 -22712 -8
rect -23884 -88 -22712 -72
rect -23884 -152 -22796 -88
rect -22732 -152 -22712 -88
rect -23884 -168 -22712 -152
rect -23884 -232 -22796 -168
rect -22732 -232 -22712 -168
rect -23884 -248 -22712 -232
rect -23884 -312 -22796 -248
rect -22732 -312 -22712 -248
rect -23884 -328 -22712 -312
rect -23884 -392 -22796 -328
rect -22732 -392 -22712 -328
rect -23884 -440 -22712 -392
rect -22472 392 -21300 440
rect -22472 328 -21384 392
rect -21320 328 -21300 392
rect -22472 312 -21300 328
rect -22472 248 -21384 312
rect -21320 248 -21300 312
rect -22472 232 -21300 248
rect -22472 168 -21384 232
rect -21320 168 -21300 232
rect -22472 152 -21300 168
rect -22472 88 -21384 152
rect -21320 88 -21300 152
rect -22472 72 -21300 88
rect -22472 8 -21384 72
rect -21320 8 -21300 72
rect -22472 -8 -21300 8
rect -22472 -72 -21384 -8
rect -21320 -72 -21300 -8
rect -22472 -88 -21300 -72
rect -22472 -152 -21384 -88
rect -21320 -152 -21300 -88
rect -22472 -168 -21300 -152
rect -22472 -232 -21384 -168
rect -21320 -232 -21300 -168
rect -22472 -248 -21300 -232
rect -22472 -312 -21384 -248
rect -21320 -312 -21300 -248
rect -22472 -328 -21300 -312
rect -22472 -392 -21384 -328
rect -21320 -392 -21300 -328
rect -22472 -440 -21300 -392
rect -21060 392 -19888 440
rect -21060 328 -19972 392
rect -19908 328 -19888 392
rect -21060 312 -19888 328
rect -21060 248 -19972 312
rect -19908 248 -19888 312
rect -21060 232 -19888 248
rect -21060 168 -19972 232
rect -19908 168 -19888 232
rect -21060 152 -19888 168
rect -21060 88 -19972 152
rect -19908 88 -19888 152
rect -21060 72 -19888 88
rect -21060 8 -19972 72
rect -19908 8 -19888 72
rect -21060 -8 -19888 8
rect -21060 -72 -19972 -8
rect -19908 -72 -19888 -8
rect -21060 -88 -19888 -72
rect -21060 -152 -19972 -88
rect -19908 -152 -19888 -88
rect -21060 -168 -19888 -152
rect -21060 -232 -19972 -168
rect -19908 -232 -19888 -168
rect -21060 -248 -19888 -232
rect -21060 -312 -19972 -248
rect -19908 -312 -19888 -248
rect -21060 -328 -19888 -312
rect -21060 -392 -19972 -328
rect -19908 -392 -19888 -328
rect -21060 -440 -19888 -392
rect -19648 392 -18476 440
rect -19648 328 -18560 392
rect -18496 328 -18476 392
rect -19648 312 -18476 328
rect -19648 248 -18560 312
rect -18496 248 -18476 312
rect -19648 232 -18476 248
rect -19648 168 -18560 232
rect -18496 168 -18476 232
rect -19648 152 -18476 168
rect -19648 88 -18560 152
rect -18496 88 -18476 152
rect -19648 72 -18476 88
rect -19648 8 -18560 72
rect -18496 8 -18476 72
rect -19648 -8 -18476 8
rect -19648 -72 -18560 -8
rect -18496 -72 -18476 -8
rect -19648 -88 -18476 -72
rect -19648 -152 -18560 -88
rect -18496 -152 -18476 -88
rect -19648 -168 -18476 -152
rect -19648 -232 -18560 -168
rect -18496 -232 -18476 -168
rect -19648 -248 -18476 -232
rect -19648 -312 -18560 -248
rect -18496 -312 -18476 -248
rect -19648 -328 -18476 -312
rect -19648 -392 -18560 -328
rect -18496 -392 -18476 -328
rect -19648 -440 -18476 -392
rect -18236 392 -17064 440
rect -18236 328 -17148 392
rect -17084 328 -17064 392
rect -18236 312 -17064 328
rect -18236 248 -17148 312
rect -17084 248 -17064 312
rect -18236 232 -17064 248
rect -18236 168 -17148 232
rect -17084 168 -17064 232
rect -18236 152 -17064 168
rect -18236 88 -17148 152
rect -17084 88 -17064 152
rect -18236 72 -17064 88
rect -18236 8 -17148 72
rect -17084 8 -17064 72
rect -18236 -8 -17064 8
rect -18236 -72 -17148 -8
rect -17084 -72 -17064 -8
rect -18236 -88 -17064 -72
rect -18236 -152 -17148 -88
rect -17084 -152 -17064 -88
rect -18236 -168 -17064 -152
rect -18236 -232 -17148 -168
rect -17084 -232 -17064 -168
rect -18236 -248 -17064 -232
rect -18236 -312 -17148 -248
rect -17084 -312 -17064 -248
rect -18236 -328 -17064 -312
rect -18236 -392 -17148 -328
rect -17084 -392 -17064 -328
rect -18236 -440 -17064 -392
rect -16824 392 -15652 440
rect -16824 328 -15736 392
rect -15672 328 -15652 392
rect -16824 312 -15652 328
rect -16824 248 -15736 312
rect -15672 248 -15652 312
rect -16824 232 -15652 248
rect -16824 168 -15736 232
rect -15672 168 -15652 232
rect -16824 152 -15652 168
rect -16824 88 -15736 152
rect -15672 88 -15652 152
rect -16824 72 -15652 88
rect -16824 8 -15736 72
rect -15672 8 -15652 72
rect -16824 -8 -15652 8
rect -16824 -72 -15736 -8
rect -15672 -72 -15652 -8
rect -16824 -88 -15652 -72
rect -16824 -152 -15736 -88
rect -15672 -152 -15652 -88
rect -16824 -168 -15652 -152
rect -16824 -232 -15736 -168
rect -15672 -232 -15652 -168
rect -16824 -248 -15652 -232
rect -16824 -312 -15736 -248
rect -15672 -312 -15652 -248
rect -16824 -328 -15652 -312
rect -16824 -392 -15736 -328
rect -15672 -392 -15652 -328
rect -16824 -440 -15652 -392
rect -15412 392 -14240 440
rect -15412 328 -14324 392
rect -14260 328 -14240 392
rect -15412 312 -14240 328
rect -15412 248 -14324 312
rect -14260 248 -14240 312
rect -15412 232 -14240 248
rect -15412 168 -14324 232
rect -14260 168 -14240 232
rect -15412 152 -14240 168
rect -15412 88 -14324 152
rect -14260 88 -14240 152
rect -15412 72 -14240 88
rect -15412 8 -14324 72
rect -14260 8 -14240 72
rect -15412 -8 -14240 8
rect -15412 -72 -14324 -8
rect -14260 -72 -14240 -8
rect -15412 -88 -14240 -72
rect -15412 -152 -14324 -88
rect -14260 -152 -14240 -88
rect -15412 -168 -14240 -152
rect -15412 -232 -14324 -168
rect -14260 -232 -14240 -168
rect -15412 -248 -14240 -232
rect -15412 -312 -14324 -248
rect -14260 -312 -14240 -248
rect -15412 -328 -14240 -312
rect -15412 -392 -14324 -328
rect -14260 -392 -14240 -328
rect -15412 -440 -14240 -392
rect -14000 392 -12828 440
rect -14000 328 -12912 392
rect -12848 328 -12828 392
rect -14000 312 -12828 328
rect -14000 248 -12912 312
rect -12848 248 -12828 312
rect -14000 232 -12828 248
rect -14000 168 -12912 232
rect -12848 168 -12828 232
rect -14000 152 -12828 168
rect -14000 88 -12912 152
rect -12848 88 -12828 152
rect -14000 72 -12828 88
rect -14000 8 -12912 72
rect -12848 8 -12828 72
rect -14000 -8 -12828 8
rect -14000 -72 -12912 -8
rect -12848 -72 -12828 -8
rect -14000 -88 -12828 -72
rect -14000 -152 -12912 -88
rect -12848 -152 -12828 -88
rect -14000 -168 -12828 -152
rect -14000 -232 -12912 -168
rect -12848 -232 -12828 -168
rect -14000 -248 -12828 -232
rect -14000 -312 -12912 -248
rect -12848 -312 -12828 -248
rect -14000 -328 -12828 -312
rect -14000 -392 -12912 -328
rect -12848 -392 -12828 -328
rect -14000 -440 -12828 -392
rect -12588 392 -11416 440
rect -12588 328 -11500 392
rect -11436 328 -11416 392
rect -12588 312 -11416 328
rect -12588 248 -11500 312
rect -11436 248 -11416 312
rect -12588 232 -11416 248
rect -12588 168 -11500 232
rect -11436 168 -11416 232
rect -12588 152 -11416 168
rect -12588 88 -11500 152
rect -11436 88 -11416 152
rect -12588 72 -11416 88
rect -12588 8 -11500 72
rect -11436 8 -11416 72
rect -12588 -8 -11416 8
rect -12588 -72 -11500 -8
rect -11436 -72 -11416 -8
rect -12588 -88 -11416 -72
rect -12588 -152 -11500 -88
rect -11436 -152 -11416 -88
rect -12588 -168 -11416 -152
rect -12588 -232 -11500 -168
rect -11436 -232 -11416 -168
rect -12588 -248 -11416 -232
rect -12588 -312 -11500 -248
rect -11436 -312 -11416 -248
rect -12588 -328 -11416 -312
rect -12588 -392 -11500 -328
rect -11436 -392 -11416 -328
rect -12588 -440 -11416 -392
rect -11176 392 -10004 440
rect -11176 328 -10088 392
rect -10024 328 -10004 392
rect -11176 312 -10004 328
rect -11176 248 -10088 312
rect -10024 248 -10004 312
rect -11176 232 -10004 248
rect -11176 168 -10088 232
rect -10024 168 -10004 232
rect -11176 152 -10004 168
rect -11176 88 -10088 152
rect -10024 88 -10004 152
rect -11176 72 -10004 88
rect -11176 8 -10088 72
rect -10024 8 -10004 72
rect -11176 -8 -10004 8
rect -11176 -72 -10088 -8
rect -10024 -72 -10004 -8
rect -11176 -88 -10004 -72
rect -11176 -152 -10088 -88
rect -10024 -152 -10004 -88
rect -11176 -168 -10004 -152
rect -11176 -232 -10088 -168
rect -10024 -232 -10004 -168
rect -11176 -248 -10004 -232
rect -11176 -312 -10088 -248
rect -10024 -312 -10004 -248
rect -11176 -328 -10004 -312
rect -11176 -392 -10088 -328
rect -10024 -392 -10004 -328
rect -11176 -440 -10004 -392
rect -9764 392 -8592 440
rect -9764 328 -8676 392
rect -8612 328 -8592 392
rect -9764 312 -8592 328
rect -9764 248 -8676 312
rect -8612 248 -8592 312
rect -9764 232 -8592 248
rect -9764 168 -8676 232
rect -8612 168 -8592 232
rect -9764 152 -8592 168
rect -9764 88 -8676 152
rect -8612 88 -8592 152
rect -9764 72 -8592 88
rect -9764 8 -8676 72
rect -8612 8 -8592 72
rect -9764 -8 -8592 8
rect -9764 -72 -8676 -8
rect -8612 -72 -8592 -8
rect -9764 -88 -8592 -72
rect -9764 -152 -8676 -88
rect -8612 -152 -8592 -88
rect -9764 -168 -8592 -152
rect -9764 -232 -8676 -168
rect -8612 -232 -8592 -168
rect -9764 -248 -8592 -232
rect -9764 -312 -8676 -248
rect -8612 -312 -8592 -248
rect -9764 -328 -8592 -312
rect -9764 -392 -8676 -328
rect -8612 -392 -8592 -328
rect -9764 -440 -8592 -392
rect -8352 392 -7180 440
rect -8352 328 -7264 392
rect -7200 328 -7180 392
rect -8352 312 -7180 328
rect -8352 248 -7264 312
rect -7200 248 -7180 312
rect -8352 232 -7180 248
rect -8352 168 -7264 232
rect -7200 168 -7180 232
rect -8352 152 -7180 168
rect -8352 88 -7264 152
rect -7200 88 -7180 152
rect -8352 72 -7180 88
rect -8352 8 -7264 72
rect -7200 8 -7180 72
rect -8352 -8 -7180 8
rect -8352 -72 -7264 -8
rect -7200 -72 -7180 -8
rect -8352 -88 -7180 -72
rect -8352 -152 -7264 -88
rect -7200 -152 -7180 -88
rect -8352 -168 -7180 -152
rect -8352 -232 -7264 -168
rect -7200 -232 -7180 -168
rect -8352 -248 -7180 -232
rect -8352 -312 -7264 -248
rect -7200 -312 -7180 -248
rect -8352 -328 -7180 -312
rect -8352 -392 -7264 -328
rect -7200 -392 -7180 -328
rect -8352 -440 -7180 -392
rect -6940 392 -5768 440
rect -6940 328 -5852 392
rect -5788 328 -5768 392
rect -6940 312 -5768 328
rect -6940 248 -5852 312
rect -5788 248 -5768 312
rect -6940 232 -5768 248
rect -6940 168 -5852 232
rect -5788 168 -5768 232
rect -6940 152 -5768 168
rect -6940 88 -5852 152
rect -5788 88 -5768 152
rect -6940 72 -5768 88
rect -6940 8 -5852 72
rect -5788 8 -5768 72
rect -6940 -8 -5768 8
rect -6940 -72 -5852 -8
rect -5788 -72 -5768 -8
rect -6940 -88 -5768 -72
rect -6940 -152 -5852 -88
rect -5788 -152 -5768 -88
rect -6940 -168 -5768 -152
rect -6940 -232 -5852 -168
rect -5788 -232 -5768 -168
rect -6940 -248 -5768 -232
rect -6940 -312 -5852 -248
rect -5788 -312 -5768 -248
rect -6940 -328 -5768 -312
rect -6940 -392 -5852 -328
rect -5788 -392 -5768 -328
rect -6940 -440 -5768 -392
rect -5528 392 -4356 440
rect -5528 328 -4440 392
rect -4376 328 -4356 392
rect -5528 312 -4356 328
rect -5528 248 -4440 312
rect -4376 248 -4356 312
rect -5528 232 -4356 248
rect -5528 168 -4440 232
rect -4376 168 -4356 232
rect -5528 152 -4356 168
rect -5528 88 -4440 152
rect -4376 88 -4356 152
rect -5528 72 -4356 88
rect -5528 8 -4440 72
rect -4376 8 -4356 72
rect -5528 -8 -4356 8
rect -5528 -72 -4440 -8
rect -4376 -72 -4356 -8
rect -5528 -88 -4356 -72
rect -5528 -152 -4440 -88
rect -4376 -152 -4356 -88
rect -5528 -168 -4356 -152
rect -5528 -232 -4440 -168
rect -4376 -232 -4356 -168
rect -5528 -248 -4356 -232
rect -5528 -312 -4440 -248
rect -4376 -312 -4356 -248
rect -5528 -328 -4356 -312
rect -5528 -392 -4440 -328
rect -4376 -392 -4356 -328
rect -5528 -440 -4356 -392
rect -4116 392 -2944 440
rect -4116 328 -3028 392
rect -2964 328 -2944 392
rect -4116 312 -2944 328
rect -4116 248 -3028 312
rect -2964 248 -2944 312
rect -4116 232 -2944 248
rect -4116 168 -3028 232
rect -2964 168 -2944 232
rect -4116 152 -2944 168
rect -4116 88 -3028 152
rect -2964 88 -2944 152
rect -4116 72 -2944 88
rect -4116 8 -3028 72
rect -2964 8 -2944 72
rect -4116 -8 -2944 8
rect -4116 -72 -3028 -8
rect -2964 -72 -2944 -8
rect -4116 -88 -2944 -72
rect -4116 -152 -3028 -88
rect -2964 -152 -2944 -88
rect -4116 -168 -2944 -152
rect -4116 -232 -3028 -168
rect -2964 -232 -2944 -168
rect -4116 -248 -2944 -232
rect -4116 -312 -3028 -248
rect -2964 -312 -2944 -248
rect -4116 -328 -2944 -312
rect -4116 -392 -3028 -328
rect -2964 -392 -2944 -328
rect -4116 -440 -2944 -392
rect -2704 392 -1532 440
rect -2704 328 -1616 392
rect -1552 328 -1532 392
rect -2704 312 -1532 328
rect -2704 248 -1616 312
rect -1552 248 -1532 312
rect -2704 232 -1532 248
rect -2704 168 -1616 232
rect -1552 168 -1532 232
rect -2704 152 -1532 168
rect -2704 88 -1616 152
rect -1552 88 -1532 152
rect -2704 72 -1532 88
rect -2704 8 -1616 72
rect -1552 8 -1532 72
rect -2704 -8 -1532 8
rect -2704 -72 -1616 -8
rect -1552 -72 -1532 -8
rect -2704 -88 -1532 -72
rect -2704 -152 -1616 -88
rect -1552 -152 -1532 -88
rect -2704 -168 -1532 -152
rect -2704 -232 -1616 -168
rect -1552 -232 -1532 -168
rect -2704 -248 -1532 -232
rect -2704 -312 -1616 -248
rect -1552 -312 -1532 -248
rect -2704 -328 -1532 -312
rect -2704 -392 -1616 -328
rect -1552 -392 -1532 -328
rect -2704 -440 -1532 -392
rect -1292 392 -120 440
rect -1292 328 -204 392
rect -140 328 -120 392
rect -1292 312 -120 328
rect -1292 248 -204 312
rect -140 248 -120 312
rect -1292 232 -120 248
rect -1292 168 -204 232
rect -140 168 -120 232
rect -1292 152 -120 168
rect -1292 88 -204 152
rect -140 88 -120 152
rect -1292 72 -120 88
rect -1292 8 -204 72
rect -140 8 -120 72
rect -1292 -8 -120 8
rect -1292 -72 -204 -8
rect -140 -72 -120 -8
rect -1292 -88 -120 -72
rect -1292 -152 -204 -88
rect -140 -152 -120 -88
rect -1292 -168 -120 -152
rect -1292 -232 -204 -168
rect -140 -232 -120 -168
rect -1292 -248 -120 -232
rect -1292 -312 -204 -248
rect -140 -312 -120 -248
rect -1292 -328 -120 -312
rect -1292 -392 -204 -328
rect -140 -392 -120 -328
rect -1292 -440 -120 -392
rect 120 392 1292 440
rect 120 328 1208 392
rect 1272 328 1292 392
rect 120 312 1292 328
rect 120 248 1208 312
rect 1272 248 1292 312
rect 120 232 1292 248
rect 120 168 1208 232
rect 1272 168 1292 232
rect 120 152 1292 168
rect 120 88 1208 152
rect 1272 88 1292 152
rect 120 72 1292 88
rect 120 8 1208 72
rect 1272 8 1292 72
rect 120 -8 1292 8
rect 120 -72 1208 -8
rect 1272 -72 1292 -8
rect 120 -88 1292 -72
rect 120 -152 1208 -88
rect 1272 -152 1292 -88
rect 120 -168 1292 -152
rect 120 -232 1208 -168
rect 1272 -232 1292 -168
rect 120 -248 1292 -232
rect 120 -312 1208 -248
rect 1272 -312 1292 -248
rect 120 -328 1292 -312
rect 120 -392 1208 -328
rect 1272 -392 1292 -328
rect 120 -440 1292 -392
rect 1532 392 2704 440
rect 1532 328 2620 392
rect 2684 328 2704 392
rect 1532 312 2704 328
rect 1532 248 2620 312
rect 2684 248 2704 312
rect 1532 232 2704 248
rect 1532 168 2620 232
rect 2684 168 2704 232
rect 1532 152 2704 168
rect 1532 88 2620 152
rect 2684 88 2704 152
rect 1532 72 2704 88
rect 1532 8 2620 72
rect 2684 8 2704 72
rect 1532 -8 2704 8
rect 1532 -72 2620 -8
rect 2684 -72 2704 -8
rect 1532 -88 2704 -72
rect 1532 -152 2620 -88
rect 2684 -152 2704 -88
rect 1532 -168 2704 -152
rect 1532 -232 2620 -168
rect 2684 -232 2704 -168
rect 1532 -248 2704 -232
rect 1532 -312 2620 -248
rect 2684 -312 2704 -248
rect 1532 -328 2704 -312
rect 1532 -392 2620 -328
rect 2684 -392 2704 -328
rect 1532 -440 2704 -392
rect 2944 392 4116 440
rect 2944 328 4032 392
rect 4096 328 4116 392
rect 2944 312 4116 328
rect 2944 248 4032 312
rect 4096 248 4116 312
rect 2944 232 4116 248
rect 2944 168 4032 232
rect 4096 168 4116 232
rect 2944 152 4116 168
rect 2944 88 4032 152
rect 4096 88 4116 152
rect 2944 72 4116 88
rect 2944 8 4032 72
rect 4096 8 4116 72
rect 2944 -8 4116 8
rect 2944 -72 4032 -8
rect 4096 -72 4116 -8
rect 2944 -88 4116 -72
rect 2944 -152 4032 -88
rect 4096 -152 4116 -88
rect 2944 -168 4116 -152
rect 2944 -232 4032 -168
rect 4096 -232 4116 -168
rect 2944 -248 4116 -232
rect 2944 -312 4032 -248
rect 4096 -312 4116 -248
rect 2944 -328 4116 -312
rect 2944 -392 4032 -328
rect 4096 -392 4116 -328
rect 2944 -440 4116 -392
rect 4356 392 5528 440
rect 4356 328 5444 392
rect 5508 328 5528 392
rect 4356 312 5528 328
rect 4356 248 5444 312
rect 5508 248 5528 312
rect 4356 232 5528 248
rect 4356 168 5444 232
rect 5508 168 5528 232
rect 4356 152 5528 168
rect 4356 88 5444 152
rect 5508 88 5528 152
rect 4356 72 5528 88
rect 4356 8 5444 72
rect 5508 8 5528 72
rect 4356 -8 5528 8
rect 4356 -72 5444 -8
rect 5508 -72 5528 -8
rect 4356 -88 5528 -72
rect 4356 -152 5444 -88
rect 5508 -152 5528 -88
rect 4356 -168 5528 -152
rect 4356 -232 5444 -168
rect 5508 -232 5528 -168
rect 4356 -248 5528 -232
rect 4356 -312 5444 -248
rect 5508 -312 5528 -248
rect 4356 -328 5528 -312
rect 4356 -392 5444 -328
rect 5508 -392 5528 -328
rect 4356 -440 5528 -392
rect 5768 392 6940 440
rect 5768 328 6856 392
rect 6920 328 6940 392
rect 5768 312 6940 328
rect 5768 248 6856 312
rect 6920 248 6940 312
rect 5768 232 6940 248
rect 5768 168 6856 232
rect 6920 168 6940 232
rect 5768 152 6940 168
rect 5768 88 6856 152
rect 6920 88 6940 152
rect 5768 72 6940 88
rect 5768 8 6856 72
rect 6920 8 6940 72
rect 5768 -8 6940 8
rect 5768 -72 6856 -8
rect 6920 -72 6940 -8
rect 5768 -88 6940 -72
rect 5768 -152 6856 -88
rect 6920 -152 6940 -88
rect 5768 -168 6940 -152
rect 5768 -232 6856 -168
rect 6920 -232 6940 -168
rect 5768 -248 6940 -232
rect 5768 -312 6856 -248
rect 6920 -312 6940 -248
rect 5768 -328 6940 -312
rect 5768 -392 6856 -328
rect 6920 -392 6940 -328
rect 5768 -440 6940 -392
rect 7180 392 8352 440
rect 7180 328 8268 392
rect 8332 328 8352 392
rect 7180 312 8352 328
rect 7180 248 8268 312
rect 8332 248 8352 312
rect 7180 232 8352 248
rect 7180 168 8268 232
rect 8332 168 8352 232
rect 7180 152 8352 168
rect 7180 88 8268 152
rect 8332 88 8352 152
rect 7180 72 8352 88
rect 7180 8 8268 72
rect 8332 8 8352 72
rect 7180 -8 8352 8
rect 7180 -72 8268 -8
rect 8332 -72 8352 -8
rect 7180 -88 8352 -72
rect 7180 -152 8268 -88
rect 8332 -152 8352 -88
rect 7180 -168 8352 -152
rect 7180 -232 8268 -168
rect 8332 -232 8352 -168
rect 7180 -248 8352 -232
rect 7180 -312 8268 -248
rect 8332 -312 8352 -248
rect 7180 -328 8352 -312
rect 7180 -392 8268 -328
rect 8332 -392 8352 -328
rect 7180 -440 8352 -392
rect 8592 392 9764 440
rect 8592 328 9680 392
rect 9744 328 9764 392
rect 8592 312 9764 328
rect 8592 248 9680 312
rect 9744 248 9764 312
rect 8592 232 9764 248
rect 8592 168 9680 232
rect 9744 168 9764 232
rect 8592 152 9764 168
rect 8592 88 9680 152
rect 9744 88 9764 152
rect 8592 72 9764 88
rect 8592 8 9680 72
rect 9744 8 9764 72
rect 8592 -8 9764 8
rect 8592 -72 9680 -8
rect 9744 -72 9764 -8
rect 8592 -88 9764 -72
rect 8592 -152 9680 -88
rect 9744 -152 9764 -88
rect 8592 -168 9764 -152
rect 8592 -232 9680 -168
rect 9744 -232 9764 -168
rect 8592 -248 9764 -232
rect 8592 -312 9680 -248
rect 9744 -312 9764 -248
rect 8592 -328 9764 -312
rect 8592 -392 9680 -328
rect 9744 -392 9764 -328
rect 8592 -440 9764 -392
rect 10004 392 11176 440
rect 10004 328 11092 392
rect 11156 328 11176 392
rect 10004 312 11176 328
rect 10004 248 11092 312
rect 11156 248 11176 312
rect 10004 232 11176 248
rect 10004 168 11092 232
rect 11156 168 11176 232
rect 10004 152 11176 168
rect 10004 88 11092 152
rect 11156 88 11176 152
rect 10004 72 11176 88
rect 10004 8 11092 72
rect 11156 8 11176 72
rect 10004 -8 11176 8
rect 10004 -72 11092 -8
rect 11156 -72 11176 -8
rect 10004 -88 11176 -72
rect 10004 -152 11092 -88
rect 11156 -152 11176 -88
rect 10004 -168 11176 -152
rect 10004 -232 11092 -168
rect 11156 -232 11176 -168
rect 10004 -248 11176 -232
rect 10004 -312 11092 -248
rect 11156 -312 11176 -248
rect 10004 -328 11176 -312
rect 10004 -392 11092 -328
rect 11156 -392 11176 -328
rect 10004 -440 11176 -392
rect 11416 392 12588 440
rect 11416 328 12504 392
rect 12568 328 12588 392
rect 11416 312 12588 328
rect 11416 248 12504 312
rect 12568 248 12588 312
rect 11416 232 12588 248
rect 11416 168 12504 232
rect 12568 168 12588 232
rect 11416 152 12588 168
rect 11416 88 12504 152
rect 12568 88 12588 152
rect 11416 72 12588 88
rect 11416 8 12504 72
rect 12568 8 12588 72
rect 11416 -8 12588 8
rect 11416 -72 12504 -8
rect 12568 -72 12588 -8
rect 11416 -88 12588 -72
rect 11416 -152 12504 -88
rect 12568 -152 12588 -88
rect 11416 -168 12588 -152
rect 11416 -232 12504 -168
rect 12568 -232 12588 -168
rect 11416 -248 12588 -232
rect 11416 -312 12504 -248
rect 12568 -312 12588 -248
rect 11416 -328 12588 -312
rect 11416 -392 12504 -328
rect 12568 -392 12588 -328
rect 11416 -440 12588 -392
rect 12828 392 14000 440
rect 12828 328 13916 392
rect 13980 328 14000 392
rect 12828 312 14000 328
rect 12828 248 13916 312
rect 13980 248 14000 312
rect 12828 232 14000 248
rect 12828 168 13916 232
rect 13980 168 14000 232
rect 12828 152 14000 168
rect 12828 88 13916 152
rect 13980 88 14000 152
rect 12828 72 14000 88
rect 12828 8 13916 72
rect 13980 8 14000 72
rect 12828 -8 14000 8
rect 12828 -72 13916 -8
rect 13980 -72 14000 -8
rect 12828 -88 14000 -72
rect 12828 -152 13916 -88
rect 13980 -152 14000 -88
rect 12828 -168 14000 -152
rect 12828 -232 13916 -168
rect 13980 -232 14000 -168
rect 12828 -248 14000 -232
rect 12828 -312 13916 -248
rect 13980 -312 14000 -248
rect 12828 -328 14000 -312
rect 12828 -392 13916 -328
rect 13980 -392 14000 -328
rect 12828 -440 14000 -392
rect 14240 392 15412 440
rect 14240 328 15328 392
rect 15392 328 15412 392
rect 14240 312 15412 328
rect 14240 248 15328 312
rect 15392 248 15412 312
rect 14240 232 15412 248
rect 14240 168 15328 232
rect 15392 168 15412 232
rect 14240 152 15412 168
rect 14240 88 15328 152
rect 15392 88 15412 152
rect 14240 72 15412 88
rect 14240 8 15328 72
rect 15392 8 15412 72
rect 14240 -8 15412 8
rect 14240 -72 15328 -8
rect 15392 -72 15412 -8
rect 14240 -88 15412 -72
rect 14240 -152 15328 -88
rect 15392 -152 15412 -88
rect 14240 -168 15412 -152
rect 14240 -232 15328 -168
rect 15392 -232 15412 -168
rect 14240 -248 15412 -232
rect 14240 -312 15328 -248
rect 15392 -312 15412 -248
rect 14240 -328 15412 -312
rect 14240 -392 15328 -328
rect 15392 -392 15412 -328
rect 14240 -440 15412 -392
rect 15652 392 16824 440
rect 15652 328 16740 392
rect 16804 328 16824 392
rect 15652 312 16824 328
rect 15652 248 16740 312
rect 16804 248 16824 312
rect 15652 232 16824 248
rect 15652 168 16740 232
rect 16804 168 16824 232
rect 15652 152 16824 168
rect 15652 88 16740 152
rect 16804 88 16824 152
rect 15652 72 16824 88
rect 15652 8 16740 72
rect 16804 8 16824 72
rect 15652 -8 16824 8
rect 15652 -72 16740 -8
rect 16804 -72 16824 -8
rect 15652 -88 16824 -72
rect 15652 -152 16740 -88
rect 16804 -152 16824 -88
rect 15652 -168 16824 -152
rect 15652 -232 16740 -168
rect 16804 -232 16824 -168
rect 15652 -248 16824 -232
rect 15652 -312 16740 -248
rect 16804 -312 16824 -248
rect 15652 -328 16824 -312
rect 15652 -392 16740 -328
rect 16804 -392 16824 -328
rect 15652 -440 16824 -392
rect 17064 392 18236 440
rect 17064 328 18152 392
rect 18216 328 18236 392
rect 17064 312 18236 328
rect 17064 248 18152 312
rect 18216 248 18236 312
rect 17064 232 18236 248
rect 17064 168 18152 232
rect 18216 168 18236 232
rect 17064 152 18236 168
rect 17064 88 18152 152
rect 18216 88 18236 152
rect 17064 72 18236 88
rect 17064 8 18152 72
rect 18216 8 18236 72
rect 17064 -8 18236 8
rect 17064 -72 18152 -8
rect 18216 -72 18236 -8
rect 17064 -88 18236 -72
rect 17064 -152 18152 -88
rect 18216 -152 18236 -88
rect 17064 -168 18236 -152
rect 17064 -232 18152 -168
rect 18216 -232 18236 -168
rect 17064 -248 18236 -232
rect 17064 -312 18152 -248
rect 18216 -312 18236 -248
rect 17064 -328 18236 -312
rect 17064 -392 18152 -328
rect 18216 -392 18236 -328
rect 17064 -440 18236 -392
rect 18476 392 19648 440
rect 18476 328 19564 392
rect 19628 328 19648 392
rect 18476 312 19648 328
rect 18476 248 19564 312
rect 19628 248 19648 312
rect 18476 232 19648 248
rect 18476 168 19564 232
rect 19628 168 19648 232
rect 18476 152 19648 168
rect 18476 88 19564 152
rect 19628 88 19648 152
rect 18476 72 19648 88
rect 18476 8 19564 72
rect 19628 8 19648 72
rect 18476 -8 19648 8
rect 18476 -72 19564 -8
rect 19628 -72 19648 -8
rect 18476 -88 19648 -72
rect 18476 -152 19564 -88
rect 19628 -152 19648 -88
rect 18476 -168 19648 -152
rect 18476 -232 19564 -168
rect 19628 -232 19648 -168
rect 18476 -248 19648 -232
rect 18476 -312 19564 -248
rect 19628 -312 19648 -248
rect 18476 -328 19648 -312
rect 18476 -392 19564 -328
rect 19628 -392 19648 -328
rect 18476 -440 19648 -392
rect 19888 392 21060 440
rect 19888 328 20976 392
rect 21040 328 21060 392
rect 19888 312 21060 328
rect 19888 248 20976 312
rect 21040 248 21060 312
rect 19888 232 21060 248
rect 19888 168 20976 232
rect 21040 168 21060 232
rect 19888 152 21060 168
rect 19888 88 20976 152
rect 21040 88 21060 152
rect 19888 72 21060 88
rect 19888 8 20976 72
rect 21040 8 21060 72
rect 19888 -8 21060 8
rect 19888 -72 20976 -8
rect 21040 -72 21060 -8
rect 19888 -88 21060 -72
rect 19888 -152 20976 -88
rect 21040 -152 21060 -88
rect 19888 -168 21060 -152
rect 19888 -232 20976 -168
rect 21040 -232 21060 -168
rect 19888 -248 21060 -232
rect 19888 -312 20976 -248
rect 21040 -312 21060 -248
rect 19888 -328 21060 -312
rect 19888 -392 20976 -328
rect 21040 -392 21060 -328
rect 19888 -440 21060 -392
rect 21300 392 22472 440
rect 21300 328 22388 392
rect 22452 328 22472 392
rect 21300 312 22472 328
rect 21300 248 22388 312
rect 22452 248 22472 312
rect 21300 232 22472 248
rect 21300 168 22388 232
rect 22452 168 22472 232
rect 21300 152 22472 168
rect 21300 88 22388 152
rect 22452 88 22472 152
rect 21300 72 22472 88
rect 21300 8 22388 72
rect 22452 8 22472 72
rect 21300 -8 22472 8
rect 21300 -72 22388 -8
rect 22452 -72 22472 -8
rect 21300 -88 22472 -72
rect 21300 -152 22388 -88
rect 22452 -152 22472 -88
rect 21300 -168 22472 -152
rect 21300 -232 22388 -168
rect 22452 -232 22472 -168
rect 21300 -248 22472 -232
rect 21300 -312 22388 -248
rect 22452 -312 22472 -248
rect 21300 -328 22472 -312
rect 21300 -392 22388 -328
rect 22452 -392 22472 -328
rect 21300 -440 22472 -392
rect 22712 392 23884 440
rect 22712 328 23800 392
rect 23864 328 23884 392
rect 22712 312 23884 328
rect 22712 248 23800 312
rect 23864 248 23884 312
rect 22712 232 23884 248
rect 22712 168 23800 232
rect 23864 168 23884 232
rect 22712 152 23884 168
rect 22712 88 23800 152
rect 23864 88 23884 152
rect 22712 72 23884 88
rect 22712 8 23800 72
rect 23864 8 23884 72
rect 22712 -8 23884 8
rect 22712 -72 23800 -8
rect 23864 -72 23884 -8
rect 22712 -88 23884 -72
rect 22712 -152 23800 -88
rect 23864 -152 23884 -88
rect 22712 -168 23884 -152
rect 22712 -232 23800 -168
rect 23864 -232 23884 -168
rect 22712 -248 23884 -232
rect 22712 -312 23800 -248
rect 23864 -312 23884 -248
rect 22712 -328 23884 -312
rect 22712 -392 23800 -328
rect 23864 -392 23884 -328
rect 22712 -440 23884 -392
rect -23884 -728 -22712 -680
rect -23884 -792 -22796 -728
rect -22732 -792 -22712 -728
rect -23884 -808 -22712 -792
rect -23884 -872 -22796 -808
rect -22732 -872 -22712 -808
rect -23884 -888 -22712 -872
rect -23884 -952 -22796 -888
rect -22732 -952 -22712 -888
rect -23884 -968 -22712 -952
rect -23884 -1032 -22796 -968
rect -22732 -1032 -22712 -968
rect -23884 -1048 -22712 -1032
rect -23884 -1112 -22796 -1048
rect -22732 -1112 -22712 -1048
rect -23884 -1128 -22712 -1112
rect -23884 -1192 -22796 -1128
rect -22732 -1192 -22712 -1128
rect -23884 -1208 -22712 -1192
rect -23884 -1272 -22796 -1208
rect -22732 -1272 -22712 -1208
rect -23884 -1288 -22712 -1272
rect -23884 -1352 -22796 -1288
rect -22732 -1352 -22712 -1288
rect -23884 -1368 -22712 -1352
rect -23884 -1432 -22796 -1368
rect -22732 -1432 -22712 -1368
rect -23884 -1448 -22712 -1432
rect -23884 -1512 -22796 -1448
rect -22732 -1512 -22712 -1448
rect -23884 -1560 -22712 -1512
rect -22472 -728 -21300 -680
rect -22472 -792 -21384 -728
rect -21320 -792 -21300 -728
rect -22472 -808 -21300 -792
rect -22472 -872 -21384 -808
rect -21320 -872 -21300 -808
rect -22472 -888 -21300 -872
rect -22472 -952 -21384 -888
rect -21320 -952 -21300 -888
rect -22472 -968 -21300 -952
rect -22472 -1032 -21384 -968
rect -21320 -1032 -21300 -968
rect -22472 -1048 -21300 -1032
rect -22472 -1112 -21384 -1048
rect -21320 -1112 -21300 -1048
rect -22472 -1128 -21300 -1112
rect -22472 -1192 -21384 -1128
rect -21320 -1192 -21300 -1128
rect -22472 -1208 -21300 -1192
rect -22472 -1272 -21384 -1208
rect -21320 -1272 -21300 -1208
rect -22472 -1288 -21300 -1272
rect -22472 -1352 -21384 -1288
rect -21320 -1352 -21300 -1288
rect -22472 -1368 -21300 -1352
rect -22472 -1432 -21384 -1368
rect -21320 -1432 -21300 -1368
rect -22472 -1448 -21300 -1432
rect -22472 -1512 -21384 -1448
rect -21320 -1512 -21300 -1448
rect -22472 -1560 -21300 -1512
rect -21060 -728 -19888 -680
rect -21060 -792 -19972 -728
rect -19908 -792 -19888 -728
rect -21060 -808 -19888 -792
rect -21060 -872 -19972 -808
rect -19908 -872 -19888 -808
rect -21060 -888 -19888 -872
rect -21060 -952 -19972 -888
rect -19908 -952 -19888 -888
rect -21060 -968 -19888 -952
rect -21060 -1032 -19972 -968
rect -19908 -1032 -19888 -968
rect -21060 -1048 -19888 -1032
rect -21060 -1112 -19972 -1048
rect -19908 -1112 -19888 -1048
rect -21060 -1128 -19888 -1112
rect -21060 -1192 -19972 -1128
rect -19908 -1192 -19888 -1128
rect -21060 -1208 -19888 -1192
rect -21060 -1272 -19972 -1208
rect -19908 -1272 -19888 -1208
rect -21060 -1288 -19888 -1272
rect -21060 -1352 -19972 -1288
rect -19908 -1352 -19888 -1288
rect -21060 -1368 -19888 -1352
rect -21060 -1432 -19972 -1368
rect -19908 -1432 -19888 -1368
rect -21060 -1448 -19888 -1432
rect -21060 -1512 -19972 -1448
rect -19908 -1512 -19888 -1448
rect -21060 -1560 -19888 -1512
rect -19648 -728 -18476 -680
rect -19648 -792 -18560 -728
rect -18496 -792 -18476 -728
rect -19648 -808 -18476 -792
rect -19648 -872 -18560 -808
rect -18496 -872 -18476 -808
rect -19648 -888 -18476 -872
rect -19648 -952 -18560 -888
rect -18496 -952 -18476 -888
rect -19648 -968 -18476 -952
rect -19648 -1032 -18560 -968
rect -18496 -1032 -18476 -968
rect -19648 -1048 -18476 -1032
rect -19648 -1112 -18560 -1048
rect -18496 -1112 -18476 -1048
rect -19648 -1128 -18476 -1112
rect -19648 -1192 -18560 -1128
rect -18496 -1192 -18476 -1128
rect -19648 -1208 -18476 -1192
rect -19648 -1272 -18560 -1208
rect -18496 -1272 -18476 -1208
rect -19648 -1288 -18476 -1272
rect -19648 -1352 -18560 -1288
rect -18496 -1352 -18476 -1288
rect -19648 -1368 -18476 -1352
rect -19648 -1432 -18560 -1368
rect -18496 -1432 -18476 -1368
rect -19648 -1448 -18476 -1432
rect -19648 -1512 -18560 -1448
rect -18496 -1512 -18476 -1448
rect -19648 -1560 -18476 -1512
rect -18236 -728 -17064 -680
rect -18236 -792 -17148 -728
rect -17084 -792 -17064 -728
rect -18236 -808 -17064 -792
rect -18236 -872 -17148 -808
rect -17084 -872 -17064 -808
rect -18236 -888 -17064 -872
rect -18236 -952 -17148 -888
rect -17084 -952 -17064 -888
rect -18236 -968 -17064 -952
rect -18236 -1032 -17148 -968
rect -17084 -1032 -17064 -968
rect -18236 -1048 -17064 -1032
rect -18236 -1112 -17148 -1048
rect -17084 -1112 -17064 -1048
rect -18236 -1128 -17064 -1112
rect -18236 -1192 -17148 -1128
rect -17084 -1192 -17064 -1128
rect -18236 -1208 -17064 -1192
rect -18236 -1272 -17148 -1208
rect -17084 -1272 -17064 -1208
rect -18236 -1288 -17064 -1272
rect -18236 -1352 -17148 -1288
rect -17084 -1352 -17064 -1288
rect -18236 -1368 -17064 -1352
rect -18236 -1432 -17148 -1368
rect -17084 -1432 -17064 -1368
rect -18236 -1448 -17064 -1432
rect -18236 -1512 -17148 -1448
rect -17084 -1512 -17064 -1448
rect -18236 -1560 -17064 -1512
rect -16824 -728 -15652 -680
rect -16824 -792 -15736 -728
rect -15672 -792 -15652 -728
rect -16824 -808 -15652 -792
rect -16824 -872 -15736 -808
rect -15672 -872 -15652 -808
rect -16824 -888 -15652 -872
rect -16824 -952 -15736 -888
rect -15672 -952 -15652 -888
rect -16824 -968 -15652 -952
rect -16824 -1032 -15736 -968
rect -15672 -1032 -15652 -968
rect -16824 -1048 -15652 -1032
rect -16824 -1112 -15736 -1048
rect -15672 -1112 -15652 -1048
rect -16824 -1128 -15652 -1112
rect -16824 -1192 -15736 -1128
rect -15672 -1192 -15652 -1128
rect -16824 -1208 -15652 -1192
rect -16824 -1272 -15736 -1208
rect -15672 -1272 -15652 -1208
rect -16824 -1288 -15652 -1272
rect -16824 -1352 -15736 -1288
rect -15672 -1352 -15652 -1288
rect -16824 -1368 -15652 -1352
rect -16824 -1432 -15736 -1368
rect -15672 -1432 -15652 -1368
rect -16824 -1448 -15652 -1432
rect -16824 -1512 -15736 -1448
rect -15672 -1512 -15652 -1448
rect -16824 -1560 -15652 -1512
rect -15412 -728 -14240 -680
rect -15412 -792 -14324 -728
rect -14260 -792 -14240 -728
rect -15412 -808 -14240 -792
rect -15412 -872 -14324 -808
rect -14260 -872 -14240 -808
rect -15412 -888 -14240 -872
rect -15412 -952 -14324 -888
rect -14260 -952 -14240 -888
rect -15412 -968 -14240 -952
rect -15412 -1032 -14324 -968
rect -14260 -1032 -14240 -968
rect -15412 -1048 -14240 -1032
rect -15412 -1112 -14324 -1048
rect -14260 -1112 -14240 -1048
rect -15412 -1128 -14240 -1112
rect -15412 -1192 -14324 -1128
rect -14260 -1192 -14240 -1128
rect -15412 -1208 -14240 -1192
rect -15412 -1272 -14324 -1208
rect -14260 -1272 -14240 -1208
rect -15412 -1288 -14240 -1272
rect -15412 -1352 -14324 -1288
rect -14260 -1352 -14240 -1288
rect -15412 -1368 -14240 -1352
rect -15412 -1432 -14324 -1368
rect -14260 -1432 -14240 -1368
rect -15412 -1448 -14240 -1432
rect -15412 -1512 -14324 -1448
rect -14260 -1512 -14240 -1448
rect -15412 -1560 -14240 -1512
rect -14000 -728 -12828 -680
rect -14000 -792 -12912 -728
rect -12848 -792 -12828 -728
rect -14000 -808 -12828 -792
rect -14000 -872 -12912 -808
rect -12848 -872 -12828 -808
rect -14000 -888 -12828 -872
rect -14000 -952 -12912 -888
rect -12848 -952 -12828 -888
rect -14000 -968 -12828 -952
rect -14000 -1032 -12912 -968
rect -12848 -1032 -12828 -968
rect -14000 -1048 -12828 -1032
rect -14000 -1112 -12912 -1048
rect -12848 -1112 -12828 -1048
rect -14000 -1128 -12828 -1112
rect -14000 -1192 -12912 -1128
rect -12848 -1192 -12828 -1128
rect -14000 -1208 -12828 -1192
rect -14000 -1272 -12912 -1208
rect -12848 -1272 -12828 -1208
rect -14000 -1288 -12828 -1272
rect -14000 -1352 -12912 -1288
rect -12848 -1352 -12828 -1288
rect -14000 -1368 -12828 -1352
rect -14000 -1432 -12912 -1368
rect -12848 -1432 -12828 -1368
rect -14000 -1448 -12828 -1432
rect -14000 -1512 -12912 -1448
rect -12848 -1512 -12828 -1448
rect -14000 -1560 -12828 -1512
rect -12588 -728 -11416 -680
rect -12588 -792 -11500 -728
rect -11436 -792 -11416 -728
rect -12588 -808 -11416 -792
rect -12588 -872 -11500 -808
rect -11436 -872 -11416 -808
rect -12588 -888 -11416 -872
rect -12588 -952 -11500 -888
rect -11436 -952 -11416 -888
rect -12588 -968 -11416 -952
rect -12588 -1032 -11500 -968
rect -11436 -1032 -11416 -968
rect -12588 -1048 -11416 -1032
rect -12588 -1112 -11500 -1048
rect -11436 -1112 -11416 -1048
rect -12588 -1128 -11416 -1112
rect -12588 -1192 -11500 -1128
rect -11436 -1192 -11416 -1128
rect -12588 -1208 -11416 -1192
rect -12588 -1272 -11500 -1208
rect -11436 -1272 -11416 -1208
rect -12588 -1288 -11416 -1272
rect -12588 -1352 -11500 -1288
rect -11436 -1352 -11416 -1288
rect -12588 -1368 -11416 -1352
rect -12588 -1432 -11500 -1368
rect -11436 -1432 -11416 -1368
rect -12588 -1448 -11416 -1432
rect -12588 -1512 -11500 -1448
rect -11436 -1512 -11416 -1448
rect -12588 -1560 -11416 -1512
rect -11176 -728 -10004 -680
rect -11176 -792 -10088 -728
rect -10024 -792 -10004 -728
rect -11176 -808 -10004 -792
rect -11176 -872 -10088 -808
rect -10024 -872 -10004 -808
rect -11176 -888 -10004 -872
rect -11176 -952 -10088 -888
rect -10024 -952 -10004 -888
rect -11176 -968 -10004 -952
rect -11176 -1032 -10088 -968
rect -10024 -1032 -10004 -968
rect -11176 -1048 -10004 -1032
rect -11176 -1112 -10088 -1048
rect -10024 -1112 -10004 -1048
rect -11176 -1128 -10004 -1112
rect -11176 -1192 -10088 -1128
rect -10024 -1192 -10004 -1128
rect -11176 -1208 -10004 -1192
rect -11176 -1272 -10088 -1208
rect -10024 -1272 -10004 -1208
rect -11176 -1288 -10004 -1272
rect -11176 -1352 -10088 -1288
rect -10024 -1352 -10004 -1288
rect -11176 -1368 -10004 -1352
rect -11176 -1432 -10088 -1368
rect -10024 -1432 -10004 -1368
rect -11176 -1448 -10004 -1432
rect -11176 -1512 -10088 -1448
rect -10024 -1512 -10004 -1448
rect -11176 -1560 -10004 -1512
rect -9764 -728 -8592 -680
rect -9764 -792 -8676 -728
rect -8612 -792 -8592 -728
rect -9764 -808 -8592 -792
rect -9764 -872 -8676 -808
rect -8612 -872 -8592 -808
rect -9764 -888 -8592 -872
rect -9764 -952 -8676 -888
rect -8612 -952 -8592 -888
rect -9764 -968 -8592 -952
rect -9764 -1032 -8676 -968
rect -8612 -1032 -8592 -968
rect -9764 -1048 -8592 -1032
rect -9764 -1112 -8676 -1048
rect -8612 -1112 -8592 -1048
rect -9764 -1128 -8592 -1112
rect -9764 -1192 -8676 -1128
rect -8612 -1192 -8592 -1128
rect -9764 -1208 -8592 -1192
rect -9764 -1272 -8676 -1208
rect -8612 -1272 -8592 -1208
rect -9764 -1288 -8592 -1272
rect -9764 -1352 -8676 -1288
rect -8612 -1352 -8592 -1288
rect -9764 -1368 -8592 -1352
rect -9764 -1432 -8676 -1368
rect -8612 -1432 -8592 -1368
rect -9764 -1448 -8592 -1432
rect -9764 -1512 -8676 -1448
rect -8612 -1512 -8592 -1448
rect -9764 -1560 -8592 -1512
rect -8352 -728 -7180 -680
rect -8352 -792 -7264 -728
rect -7200 -792 -7180 -728
rect -8352 -808 -7180 -792
rect -8352 -872 -7264 -808
rect -7200 -872 -7180 -808
rect -8352 -888 -7180 -872
rect -8352 -952 -7264 -888
rect -7200 -952 -7180 -888
rect -8352 -968 -7180 -952
rect -8352 -1032 -7264 -968
rect -7200 -1032 -7180 -968
rect -8352 -1048 -7180 -1032
rect -8352 -1112 -7264 -1048
rect -7200 -1112 -7180 -1048
rect -8352 -1128 -7180 -1112
rect -8352 -1192 -7264 -1128
rect -7200 -1192 -7180 -1128
rect -8352 -1208 -7180 -1192
rect -8352 -1272 -7264 -1208
rect -7200 -1272 -7180 -1208
rect -8352 -1288 -7180 -1272
rect -8352 -1352 -7264 -1288
rect -7200 -1352 -7180 -1288
rect -8352 -1368 -7180 -1352
rect -8352 -1432 -7264 -1368
rect -7200 -1432 -7180 -1368
rect -8352 -1448 -7180 -1432
rect -8352 -1512 -7264 -1448
rect -7200 -1512 -7180 -1448
rect -8352 -1560 -7180 -1512
rect -6940 -728 -5768 -680
rect -6940 -792 -5852 -728
rect -5788 -792 -5768 -728
rect -6940 -808 -5768 -792
rect -6940 -872 -5852 -808
rect -5788 -872 -5768 -808
rect -6940 -888 -5768 -872
rect -6940 -952 -5852 -888
rect -5788 -952 -5768 -888
rect -6940 -968 -5768 -952
rect -6940 -1032 -5852 -968
rect -5788 -1032 -5768 -968
rect -6940 -1048 -5768 -1032
rect -6940 -1112 -5852 -1048
rect -5788 -1112 -5768 -1048
rect -6940 -1128 -5768 -1112
rect -6940 -1192 -5852 -1128
rect -5788 -1192 -5768 -1128
rect -6940 -1208 -5768 -1192
rect -6940 -1272 -5852 -1208
rect -5788 -1272 -5768 -1208
rect -6940 -1288 -5768 -1272
rect -6940 -1352 -5852 -1288
rect -5788 -1352 -5768 -1288
rect -6940 -1368 -5768 -1352
rect -6940 -1432 -5852 -1368
rect -5788 -1432 -5768 -1368
rect -6940 -1448 -5768 -1432
rect -6940 -1512 -5852 -1448
rect -5788 -1512 -5768 -1448
rect -6940 -1560 -5768 -1512
rect -5528 -728 -4356 -680
rect -5528 -792 -4440 -728
rect -4376 -792 -4356 -728
rect -5528 -808 -4356 -792
rect -5528 -872 -4440 -808
rect -4376 -872 -4356 -808
rect -5528 -888 -4356 -872
rect -5528 -952 -4440 -888
rect -4376 -952 -4356 -888
rect -5528 -968 -4356 -952
rect -5528 -1032 -4440 -968
rect -4376 -1032 -4356 -968
rect -5528 -1048 -4356 -1032
rect -5528 -1112 -4440 -1048
rect -4376 -1112 -4356 -1048
rect -5528 -1128 -4356 -1112
rect -5528 -1192 -4440 -1128
rect -4376 -1192 -4356 -1128
rect -5528 -1208 -4356 -1192
rect -5528 -1272 -4440 -1208
rect -4376 -1272 -4356 -1208
rect -5528 -1288 -4356 -1272
rect -5528 -1352 -4440 -1288
rect -4376 -1352 -4356 -1288
rect -5528 -1368 -4356 -1352
rect -5528 -1432 -4440 -1368
rect -4376 -1432 -4356 -1368
rect -5528 -1448 -4356 -1432
rect -5528 -1512 -4440 -1448
rect -4376 -1512 -4356 -1448
rect -5528 -1560 -4356 -1512
rect -4116 -728 -2944 -680
rect -4116 -792 -3028 -728
rect -2964 -792 -2944 -728
rect -4116 -808 -2944 -792
rect -4116 -872 -3028 -808
rect -2964 -872 -2944 -808
rect -4116 -888 -2944 -872
rect -4116 -952 -3028 -888
rect -2964 -952 -2944 -888
rect -4116 -968 -2944 -952
rect -4116 -1032 -3028 -968
rect -2964 -1032 -2944 -968
rect -4116 -1048 -2944 -1032
rect -4116 -1112 -3028 -1048
rect -2964 -1112 -2944 -1048
rect -4116 -1128 -2944 -1112
rect -4116 -1192 -3028 -1128
rect -2964 -1192 -2944 -1128
rect -4116 -1208 -2944 -1192
rect -4116 -1272 -3028 -1208
rect -2964 -1272 -2944 -1208
rect -4116 -1288 -2944 -1272
rect -4116 -1352 -3028 -1288
rect -2964 -1352 -2944 -1288
rect -4116 -1368 -2944 -1352
rect -4116 -1432 -3028 -1368
rect -2964 -1432 -2944 -1368
rect -4116 -1448 -2944 -1432
rect -4116 -1512 -3028 -1448
rect -2964 -1512 -2944 -1448
rect -4116 -1560 -2944 -1512
rect -2704 -728 -1532 -680
rect -2704 -792 -1616 -728
rect -1552 -792 -1532 -728
rect -2704 -808 -1532 -792
rect -2704 -872 -1616 -808
rect -1552 -872 -1532 -808
rect -2704 -888 -1532 -872
rect -2704 -952 -1616 -888
rect -1552 -952 -1532 -888
rect -2704 -968 -1532 -952
rect -2704 -1032 -1616 -968
rect -1552 -1032 -1532 -968
rect -2704 -1048 -1532 -1032
rect -2704 -1112 -1616 -1048
rect -1552 -1112 -1532 -1048
rect -2704 -1128 -1532 -1112
rect -2704 -1192 -1616 -1128
rect -1552 -1192 -1532 -1128
rect -2704 -1208 -1532 -1192
rect -2704 -1272 -1616 -1208
rect -1552 -1272 -1532 -1208
rect -2704 -1288 -1532 -1272
rect -2704 -1352 -1616 -1288
rect -1552 -1352 -1532 -1288
rect -2704 -1368 -1532 -1352
rect -2704 -1432 -1616 -1368
rect -1552 -1432 -1532 -1368
rect -2704 -1448 -1532 -1432
rect -2704 -1512 -1616 -1448
rect -1552 -1512 -1532 -1448
rect -2704 -1560 -1532 -1512
rect -1292 -728 -120 -680
rect -1292 -792 -204 -728
rect -140 -792 -120 -728
rect -1292 -808 -120 -792
rect -1292 -872 -204 -808
rect -140 -872 -120 -808
rect -1292 -888 -120 -872
rect -1292 -952 -204 -888
rect -140 -952 -120 -888
rect -1292 -968 -120 -952
rect -1292 -1032 -204 -968
rect -140 -1032 -120 -968
rect -1292 -1048 -120 -1032
rect -1292 -1112 -204 -1048
rect -140 -1112 -120 -1048
rect -1292 -1128 -120 -1112
rect -1292 -1192 -204 -1128
rect -140 -1192 -120 -1128
rect -1292 -1208 -120 -1192
rect -1292 -1272 -204 -1208
rect -140 -1272 -120 -1208
rect -1292 -1288 -120 -1272
rect -1292 -1352 -204 -1288
rect -140 -1352 -120 -1288
rect -1292 -1368 -120 -1352
rect -1292 -1432 -204 -1368
rect -140 -1432 -120 -1368
rect -1292 -1448 -120 -1432
rect -1292 -1512 -204 -1448
rect -140 -1512 -120 -1448
rect -1292 -1560 -120 -1512
rect 120 -728 1292 -680
rect 120 -792 1208 -728
rect 1272 -792 1292 -728
rect 120 -808 1292 -792
rect 120 -872 1208 -808
rect 1272 -872 1292 -808
rect 120 -888 1292 -872
rect 120 -952 1208 -888
rect 1272 -952 1292 -888
rect 120 -968 1292 -952
rect 120 -1032 1208 -968
rect 1272 -1032 1292 -968
rect 120 -1048 1292 -1032
rect 120 -1112 1208 -1048
rect 1272 -1112 1292 -1048
rect 120 -1128 1292 -1112
rect 120 -1192 1208 -1128
rect 1272 -1192 1292 -1128
rect 120 -1208 1292 -1192
rect 120 -1272 1208 -1208
rect 1272 -1272 1292 -1208
rect 120 -1288 1292 -1272
rect 120 -1352 1208 -1288
rect 1272 -1352 1292 -1288
rect 120 -1368 1292 -1352
rect 120 -1432 1208 -1368
rect 1272 -1432 1292 -1368
rect 120 -1448 1292 -1432
rect 120 -1512 1208 -1448
rect 1272 -1512 1292 -1448
rect 120 -1560 1292 -1512
rect 1532 -728 2704 -680
rect 1532 -792 2620 -728
rect 2684 -792 2704 -728
rect 1532 -808 2704 -792
rect 1532 -872 2620 -808
rect 2684 -872 2704 -808
rect 1532 -888 2704 -872
rect 1532 -952 2620 -888
rect 2684 -952 2704 -888
rect 1532 -968 2704 -952
rect 1532 -1032 2620 -968
rect 2684 -1032 2704 -968
rect 1532 -1048 2704 -1032
rect 1532 -1112 2620 -1048
rect 2684 -1112 2704 -1048
rect 1532 -1128 2704 -1112
rect 1532 -1192 2620 -1128
rect 2684 -1192 2704 -1128
rect 1532 -1208 2704 -1192
rect 1532 -1272 2620 -1208
rect 2684 -1272 2704 -1208
rect 1532 -1288 2704 -1272
rect 1532 -1352 2620 -1288
rect 2684 -1352 2704 -1288
rect 1532 -1368 2704 -1352
rect 1532 -1432 2620 -1368
rect 2684 -1432 2704 -1368
rect 1532 -1448 2704 -1432
rect 1532 -1512 2620 -1448
rect 2684 -1512 2704 -1448
rect 1532 -1560 2704 -1512
rect 2944 -728 4116 -680
rect 2944 -792 4032 -728
rect 4096 -792 4116 -728
rect 2944 -808 4116 -792
rect 2944 -872 4032 -808
rect 4096 -872 4116 -808
rect 2944 -888 4116 -872
rect 2944 -952 4032 -888
rect 4096 -952 4116 -888
rect 2944 -968 4116 -952
rect 2944 -1032 4032 -968
rect 4096 -1032 4116 -968
rect 2944 -1048 4116 -1032
rect 2944 -1112 4032 -1048
rect 4096 -1112 4116 -1048
rect 2944 -1128 4116 -1112
rect 2944 -1192 4032 -1128
rect 4096 -1192 4116 -1128
rect 2944 -1208 4116 -1192
rect 2944 -1272 4032 -1208
rect 4096 -1272 4116 -1208
rect 2944 -1288 4116 -1272
rect 2944 -1352 4032 -1288
rect 4096 -1352 4116 -1288
rect 2944 -1368 4116 -1352
rect 2944 -1432 4032 -1368
rect 4096 -1432 4116 -1368
rect 2944 -1448 4116 -1432
rect 2944 -1512 4032 -1448
rect 4096 -1512 4116 -1448
rect 2944 -1560 4116 -1512
rect 4356 -728 5528 -680
rect 4356 -792 5444 -728
rect 5508 -792 5528 -728
rect 4356 -808 5528 -792
rect 4356 -872 5444 -808
rect 5508 -872 5528 -808
rect 4356 -888 5528 -872
rect 4356 -952 5444 -888
rect 5508 -952 5528 -888
rect 4356 -968 5528 -952
rect 4356 -1032 5444 -968
rect 5508 -1032 5528 -968
rect 4356 -1048 5528 -1032
rect 4356 -1112 5444 -1048
rect 5508 -1112 5528 -1048
rect 4356 -1128 5528 -1112
rect 4356 -1192 5444 -1128
rect 5508 -1192 5528 -1128
rect 4356 -1208 5528 -1192
rect 4356 -1272 5444 -1208
rect 5508 -1272 5528 -1208
rect 4356 -1288 5528 -1272
rect 4356 -1352 5444 -1288
rect 5508 -1352 5528 -1288
rect 4356 -1368 5528 -1352
rect 4356 -1432 5444 -1368
rect 5508 -1432 5528 -1368
rect 4356 -1448 5528 -1432
rect 4356 -1512 5444 -1448
rect 5508 -1512 5528 -1448
rect 4356 -1560 5528 -1512
rect 5768 -728 6940 -680
rect 5768 -792 6856 -728
rect 6920 -792 6940 -728
rect 5768 -808 6940 -792
rect 5768 -872 6856 -808
rect 6920 -872 6940 -808
rect 5768 -888 6940 -872
rect 5768 -952 6856 -888
rect 6920 -952 6940 -888
rect 5768 -968 6940 -952
rect 5768 -1032 6856 -968
rect 6920 -1032 6940 -968
rect 5768 -1048 6940 -1032
rect 5768 -1112 6856 -1048
rect 6920 -1112 6940 -1048
rect 5768 -1128 6940 -1112
rect 5768 -1192 6856 -1128
rect 6920 -1192 6940 -1128
rect 5768 -1208 6940 -1192
rect 5768 -1272 6856 -1208
rect 6920 -1272 6940 -1208
rect 5768 -1288 6940 -1272
rect 5768 -1352 6856 -1288
rect 6920 -1352 6940 -1288
rect 5768 -1368 6940 -1352
rect 5768 -1432 6856 -1368
rect 6920 -1432 6940 -1368
rect 5768 -1448 6940 -1432
rect 5768 -1512 6856 -1448
rect 6920 -1512 6940 -1448
rect 5768 -1560 6940 -1512
rect 7180 -728 8352 -680
rect 7180 -792 8268 -728
rect 8332 -792 8352 -728
rect 7180 -808 8352 -792
rect 7180 -872 8268 -808
rect 8332 -872 8352 -808
rect 7180 -888 8352 -872
rect 7180 -952 8268 -888
rect 8332 -952 8352 -888
rect 7180 -968 8352 -952
rect 7180 -1032 8268 -968
rect 8332 -1032 8352 -968
rect 7180 -1048 8352 -1032
rect 7180 -1112 8268 -1048
rect 8332 -1112 8352 -1048
rect 7180 -1128 8352 -1112
rect 7180 -1192 8268 -1128
rect 8332 -1192 8352 -1128
rect 7180 -1208 8352 -1192
rect 7180 -1272 8268 -1208
rect 8332 -1272 8352 -1208
rect 7180 -1288 8352 -1272
rect 7180 -1352 8268 -1288
rect 8332 -1352 8352 -1288
rect 7180 -1368 8352 -1352
rect 7180 -1432 8268 -1368
rect 8332 -1432 8352 -1368
rect 7180 -1448 8352 -1432
rect 7180 -1512 8268 -1448
rect 8332 -1512 8352 -1448
rect 7180 -1560 8352 -1512
rect 8592 -728 9764 -680
rect 8592 -792 9680 -728
rect 9744 -792 9764 -728
rect 8592 -808 9764 -792
rect 8592 -872 9680 -808
rect 9744 -872 9764 -808
rect 8592 -888 9764 -872
rect 8592 -952 9680 -888
rect 9744 -952 9764 -888
rect 8592 -968 9764 -952
rect 8592 -1032 9680 -968
rect 9744 -1032 9764 -968
rect 8592 -1048 9764 -1032
rect 8592 -1112 9680 -1048
rect 9744 -1112 9764 -1048
rect 8592 -1128 9764 -1112
rect 8592 -1192 9680 -1128
rect 9744 -1192 9764 -1128
rect 8592 -1208 9764 -1192
rect 8592 -1272 9680 -1208
rect 9744 -1272 9764 -1208
rect 8592 -1288 9764 -1272
rect 8592 -1352 9680 -1288
rect 9744 -1352 9764 -1288
rect 8592 -1368 9764 -1352
rect 8592 -1432 9680 -1368
rect 9744 -1432 9764 -1368
rect 8592 -1448 9764 -1432
rect 8592 -1512 9680 -1448
rect 9744 -1512 9764 -1448
rect 8592 -1560 9764 -1512
rect 10004 -728 11176 -680
rect 10004 -792 11092 -728
rect 11156 -792 11176 -728
rect 10004 -808 11176 -792
rect 10004 -872 11092 -808
rect 11156 -872 11176 -808
rect 10004 -888 11176 -872
rect 10004 -952 11092 -888
rect 11156 -952 11176 -888
rect 10004 -968 11176 -952
rect 10004 -1032 11092 -968
rect 11156 -1032 11176 -968
rect 10004 -1048 11176 -1032
rect 10004 -1112 11092 -1048
rect 11156 -1112 11176 -1048
rect 10004 -1128 11176 -1112
rect 10004 -1192 11092 -1128
rect 11156 -1192 11176 -1128
rect 10004 -1208 11176 -1192
rect 10004 -1272 11092 -1208
rect 11156 -1272 11176 -1208
rect 10004 -1288 11176 -1272
rect 10004 -1352 11092 -1288
rect 11156 -1352 11176 -1288
rect 10004 -1368 11176 -1352
rect 10004 -1432 11092 -1368
rect 11156 -1432 11176 -1368
rect 10004 -1448 11176 -1432
rect 10004 -1512 11092 -1448
rect 11156 -1512 11176 -1448
rect 10004 -1560 11176 -1512
rect 11416 -728 12588 -680
rect 11416 -792 12504 -728
rect 12568 -792 12588 -728
rect 11416 -808 12588 -792
rect 11416 -872 12504 -808
rect 12568 -872 12588 -808
rect 11416 -888 12588 -872
rect 11416 -952 12504 -888
rect 12568 -952 12588 -888
rect 11416 -968 12588 -952
rect 11416 -1032 12504 -968
rect 12568 -1032 12588 -968
rect 11416 -1048 12588 -1032
rect 11416 -1112 12504 -1048
rect 12568 -1112 12588 -1048
rect 11416 -1128 12588 -1112
rect 11416 -1192 12504 -1128
rect 12568 -1192 12588 -1128
rect 11416 -1208 12588 -1192
rect 11416 -1272 12504 -1208
rect 12568 -1272 12588 -1208
rect 11416 -1288 12588 -1272
rect 11416 -1352 12504 -1288
rect 12568 -1352 12588 -1288
rect 11416 -1368 12588 -1352
rect 11416 -1432 12504 -1368
rect 12568 -1432 12588 -1368
rect 11416 -1448 12588 -1432
rect 11416 -1512 12504 -1448
rect 12568 -1512 12588 -1448
rect 11416 -1560 12588 -1512
rect 12828 -728 14000 -680
rect 12828 -792 13916 -728
rect 13980 -792 14000 -728
rect 12828 -808 14000 -792
rect 12828 -872 13916 -808
rect 13980 -872 14000 -808
rect 12828 -888 14000 -872
rect 12828 -952 13916 -888
rect 13980 -952 14000 -888
rect 12828 -968 14000 -952
rect 12828 -1032 13916 -968
rect 13980 -1032 14000 -968
rect 12828 -1048 14000 -1032
rect 12828 -1112 13916 -1048
rect 13980 -1112 14000 -1048
rect 12828 -1128 14000 -1112
rect 12828 -1192 13916 -1128
rect 13980 -1192 14000 -1128
rect 12828 -1208 14000 -1192
rect 12828 -1272 13916 -1208
rect 13980 -1272 14000 -1208
rect 12828 -1288 14000 -1272
rect 12828 -1352 13916 -1288
rect 13980 -1352 14000 -1288
rect 12828 -1368 14000 -1352
rect 12828 -1432 13916 -1368
rect 13980 -1432 14000 -1368
rect 12828 -1448 14000 -1432
rect 12828 -1512 13916 -1448
rect 13980 -1512 14000 -1448
rect 12828 -1560 14000 -1512
rect 14240 -728 15412 -680
rect 14240 -792 15328 -728
rect 15392 -792 15412 -728
rect 14240 -808 15412 -792
rect 14240 -872 15328 -808
rect 15392 -872 15412 -808
rect 14240 -888 15412 -872
rect 14240 -952 15328 -888
rect 15392 -952 15412 -888
rect 14240 -968 15412 -952
rect 14240 -1032 15328 -968
rect 15392 -1032 15412 -968
rect 14240 -1048 15412 -1032
rect 14240 -1112 15328 -1048
rect 15392 -1112 15412 -1048
rect 14240 -1128 15412 -1112
rect 14240 -1192 15328 -1128
rect 15392 -1192 15412 -1128
rect 14240 -1208 15412 -1192
rect 14240 -1272 15328 -1208
rect 15392 -1272 15412 -1208
rect 14240 -1288 15412 -1272
rect 14240 -1352 15328 -1288
rect 15392 -1352 15412 -1288
rect 14240 -1368 15412 -1352
rect 14240 -1432 15328 -1368
rect 15392 -1432 15412 -1368
rect 14240 -1448 15412 -1432
rect 14240 -1512 15328 -1448
rect 15392 -1512 15412 -1448
rect 14240 -1560 15412 -1512
rect 15652 -728 16824 -680
rect 15652 -792 16740 -728
rect 16804 -792 16824 -728
rect 15652 -808 16824 -792
rect 15652 -872 16740 -808
rect 16804 -872 16824 -808
rect 15652 -888 16824 -872
rect 15652 -952 16740 -888
rect 16804 -952 16824 -888
rect 15652 -968 16824 -952
rect 15652 -1032 16740 -968
rect 16804 -1032 16824 -968
rect 15652 -1048 16824 -1032
rect 15652 -1112 16740 -1048
rect 16804 -1112 16824 -1048
rect 15652 -1128 16824 -1112
rect 15652 -1192 16740 -1128
rect 16804 -1192 16824 -1128
rect 15652 -1208 16824 -1192
rect 15652 -1272 16740 -1208
rect 16804 -1272 16824 -1208
rect 15652 -1288 16824 -1272
rect 15652 -1352 16740 -1288
rect 16804 -1352 16824 -1288
rect 15652 -1368 16824 -1352
rect 15652 -1432 16740 -1368
rect 16804 -1432 16824 -1368
rect 15652 -1448 16824 -1432
rect 15652 -1512 16740 -1448
rect 16804 -1512 16824 -1448
rect 15652 -1560 16824 -1512
rect 17064 -728 18236 -680
rect 17064 -792 18152 -728
rect 18216 -792 18236 -728
rect 17064 -808 18236 -792
rect 17064 -872 18152 -808
rect 18216 -872 18236 -808
rect 17064 -888 18236 -872
rect 17064 -952 18152 -888
rect 18216 -952 18236 -888
rect 17064 -968 18236 -952
rect 17064 -1032 18152 -968
rect 18216 -1032 18236 -968
rect 17064 -1048 18236 -1032
rect 17064 -1112 18152 -1048
rect 18216 -1112 18236 -1048
rect 17064 -1128 18236 -1112
rect 17064 -1192 18152 -1128
rect 18216 -1192 18236 -1128
rect 17064 -1208 18236 -1192
rect 17064 -1272 18152 -1208
rect 18216 -1272 18236 -1208
rect 17064 -1288 18236 -1272
rect 17064 -1352 18152 -1288
rect 18216 -1352 18236 -1288
rect 17064 -1368 18236 -1352
rect 17064 -1432 18152 -1368
rect 18216 -1432 18236 -1368
rect 17064 -1448 18236 -1432
rect 17064 -1512 18152 -1448
rect 18216 -1512 18236 -1448
rect 17064 -1560 18236 -1512
rect 18476 -728 19648 -680
rect 18476 -792 19564 -728
rect 19628 -792 19648 -728
rect 18476 -808 19648 -792
rect 18476 -872 19564 -808
rect 19628 -872 19648 -808
rect 18476 -888 19648 -872
rect 18476 -952 19564 -888
rect 19628 -952 19648 -888
rect 18476 -968 19648 -952
rect 18476 -1032 19564 -968
rect 19628 -1032 19648 -968
rect 18476 -1048 19648 -1032
rect 18476 -1112 19564 -1048
rect 19628 -1112 19648 -1048
rect 18476 -1128 19648 -1112
rect 18476 -1192 19564 -1128
rect 19628 -1192 19648 -1128
rect 18476 -1208 19648 -1192
rect 18476 -1272 19564 -1208
rect 19628 -1272 19648 -1208
rect 18476 -1288 19648 -1272
rect 18476 -1352 19564 -1288
rect 19628 -1352 19648 -1288
rect 18476 -1368 19648 -1352
rect 18476 -1432 19564 -1368
rect 19628 -1432 19648 -1368
rect 18476 -1448 19648 -1432
rect 18476 -1512 19564 -1448
rect 19628 -1512 19648 -1448
rect 18476 -1560 19648 -1512
rect 19888 -728 21060 -680
rect 19888 -792 20976 -728
rect 21040 -792 21060 -728
rect 19888 -808 21060 -792
rect 19888 -872 20976 -808
rect 21040 -872 21060 -808
rect 19888 -888 21060 -872
rect 19888 -952 20976 -888
rect 21040 -952 21060 -888
rect 19888 -968 21060 -952
rect 19888 -1032 20976 -968
rect 21040 -1032 21060 -968
rect 19888 -1048 21060 -1032
rect 19888 -1112 20976 -1048
rect 21040 -1112 21060 -1048
rect 19888 -1128 21060 -1112
rect 19888 -1192 20976 -1128
rect 21040 -1192 21060 -1128
rect 19888 -1208 21060 -1192
rect 19888 -1272 20976 -1208
rect 21040 -1272 21060 -1208
rect 19888 -1288 21060 -1272
rect 19888 -1352 20976 -1288
rect 21040 -1352 21060 -1288
rect 19888 -1368 21060 -1352
rect 19888 -1432 20976 -1368
rect 21040 -1432 21060 -1368
rect 19888 -1448 21060 -1432
rect 19888 -1512 20976 -1448
rect 21040 -1512 21060 -1448
rect 19888 -1560 21060 -1512
rect 21300 -728 22472 -680
rect 21300 -792 22388 -728
rect 22452 -792 22472 -728
rect 21300 -808 22472 -792
rect 21300 -872 22388 -808
rect 22452 -872 22472 -808
rect 21300 -888 22472 -872
rect 21300 -952 22388 -888
rect 22452 -952 22472 -888
rect 21300 -968 22472 -952
rect 21300 -1032 22388 -968
rect 22452 -1032 22472 -968
rect 21300 -1048 22472 -1032
rect 21300 -1112 22388 -1048
rect 22452 -1112 22472 -1048
rect 21300 -1128 22472 -1112
rect 21300 -1192 22388 -1128
rect 22452 -1192 22472 -1128
rect 21300 -1208 22472 -1192
rect 21300 -1272 22388 -1208
rect 22452 -1272 22472 -1208
rect 21300 -1288 22472 -1272
rect 21300 -1352 22388 -1288
rect 22452 -1352 22472 -1288
rect 21300 -1368 22472 -1352
rect 21300 -1432 22388 -1368
rect 22452 -1432 22472 -1368
rect 21300 -1448 22472 -1432
rect 21300 -1512 22388 -1448
rect 22452 -1512 22472 -1448
rect 21300 -1560 22472 -1512
rect 22712 -728 23884 -680
rect 22712 -792 23800 -728
rect 23864 -792 23884 -728
rect 22712 -808 23884 -792
rect 22712 -872 23800 -808
rect 23864 -872 23884 -808
rect 22712 -888 23884 -872
rect 22712 -952 23800 -888
rect 23864 -952 23884 -888
rect 22712 -968 23884 -952
rect 22712 -1032 23800 -968
rect 23864 -1032 23884 -968
rect 22712 -1048 23884 -1032
rect 22712 -1112 23800 -1048
rect 23864 -1112 23884 -1048
rect 22712 -1128 23884 -1112
rect 22712 -1192 23800 -1128
rect 23864 -1192 23884 -1128
rect 22712 -1208 23884 -1192
rect 22712 -1272 23800 -1208
rect 23864 -1272 23884 -1208
rect 22712 -1288 23884 -1272
rect 22712 -1352 23800 -1288
rect 23864 -1352 23884 -1288
rect 22712 -1368 23884 -1352
rect 22712 -1432 23800 -1368
rect 23864 -1432 23884 -1368
rect 22712 -1448 23884 -1432
rect 22712 -1512 23800 -1448
rect 23864 -1512 23884 -1448
rect 22712 -1560 23884 -1512
rect -23884 -1848 -22712 -1800
rect -23884 -1912 -22796 -1848
rect -22732 -1912 -22712 -1848
rect -23884 -1928 -22712 -1912
rect -23884 -1992 -22796 -1928
rect -22732 -1992 -22712 -1928
rect -23884 -2008 -22712 -1992
rect -23884 -2072 -22796 -2008
rect -22732 -2072 -22712 -2008
rect -23884 -2088 -22712 -2072
rect -23884 -2152 -22796 -2088
rect -22732 -2152 -22712 -2088
rect -23884 -2168 -22712 -2152
rect -23884 -2232 -22796 -2168
rect -22732 -2232 -22712 -2168
rect -23884 -2248 -22712 -2232
rect -23884 -2312 -22796 -2248
rect -22732 -2312 -22712 -2248
rect -23884 -2328 -22712 -2312
rect -23884 -2392 -22796 -2328
rect -22732 -2392 -22712 -2328
rect -23884 -2408 -22712 -2392
rect -23884 -2472 -22796 -2408
rect -22732 -2472 -22712 -2408
rect -23884 -2488 -22712 -2472
rect -23884 -2552 -22796 -2488
rect -22732 -2552 -22712 -2488
rect -23884 -2568 -22712 -2552
rect -23884 -2632 -22796 -2568
rect -22732 -2632 -22712 -2568
rect -23884 -2680 -22712 -2632
rect -22472 -1848 -21300 -1800
rect -22472 -1912 -21384 -1848
rect -21320 -1912 -21300 -1848
rect -22472 -1928 -21300 -1912
rect -22472 -1992 -21384 -1928
rect -21320 -1992 -21300 -1928
rect -22472 -2008 -21300 -1992
rect -22472 -2072 -21384 -2008
rect -21320 -2072 -21300 -2008
rect -22472 -2088 -21300 -2072
rect -22472 -2152 -21384 -2088
rect -21320 -2152 -21300 -2088
rect -22472 -2168 -21300 -2152
rect -22472 -2232 -21384 -2168
rect -21320 -2232 -21300 -2168
rect -22472 -2248 -21300 -2232
rect -22472 -2312 -21384 -2248
rect -21320 -2312 -21300 -2248
rect -22472 -2328 -21300 -2312
rect -22472 -2392 -21384 -2328
rect -21320 -2392 -21300 -2328
rect -22472 -2408 -21300 -2392
rect -22472 -2472 -21384 -2408
rect -21320 -2472 -21300 -2408
rect -22472 -2488 -21300 -2472
rect -22472 -2552 -21384 -2488
rect -21320 -2552 -21300 -2488
rect -22472 -2568 -21300 -2552
rect -22472 -2632 -21384 -2568
rect -21320 -2632 -21300 -2568
rect -22472 -2680 -21300 -2632
rect -21060 -1848 -19888 -1800
rect -21060 -1912 -19972 -1848
rect -19908 -1912 -19888 -1848
rect -21060 -1928 -19888 -1912
rect -21060 -1992 -19972 -1928
rect -19908 -1992 -19888 -1928
rect -21060 -2008 -19888 -1992
rect -21060 -2072 -19972 -2008
rect -19908 -2072 -19888 -2008
rect -21060 -2088 -19888 -2072
rect -21060 -2152 -19972 -2088
rect -19908 -2152 -19888 -2088
rect -21060 -2168 -19888 -2152
rect -21060 -2232 -19972 -2168
rect -19908 -2232 -19888 -2168
rect -21060 -2248 -19888 -2232
rect -21060 -2312 -19972 -2248
rect -19908 -2312 -19888 -2248
rect -21060 -2328 -19888 -2312
rect -21060 -2392 -19972 -2328
rect -19908 -2392 -19888 -2328
rect -21060 -2408 -19888 -2392
rect -21060 -2472 -19972 -2408
rect -19908 -2472 -19888 -2408
rect -21060 -2488 -19888 -2472
rect -21060 -2552 -19972 -2488
rect -19908 -2552 -19888 -2488
rect -21060 -2568 -19888 -2552
rect -21060 -2632 -19972 -2568
rect -19908 -2632 -19888 -2568
rect -21060 -2680 -19888 -2632
rect -19648 -1848 -18476 -1800
rect -19648 -1912 -18560 -1848
rect -18496 -1912 -18476 -1848
rect -19648 -1928 -18476 -1912
rect -19648 -1992 -18560 -1928
rect -18496 -1992 -18476 -1928
rect -19648 -2008 -18476 -1992
rect -19648 -2072 -18560 -2008
rect -18496 -2072 -18476 -2008
rect -19648 -2088 -18476 -2072
rect -19648 -2152 -18560 -2088
rect -18496 -2152 -18476 -2088
rect -19648 -2168 -18476 -2152
rect -19648 -2232 -18560 -2168
rect -18496 -2232 -18476 -2168
rect -19648 -2248 -18476 -2232
rect -19648 -2312 -18560 -2248
rect -18496 -2312 -18476 -2248
rect -19648 -2328 -18476 -2312
rect -19648 -2392 -18560 -2328
rect -18496 -2392 -18476 -2328
rect -19648 -2408 -18476 -2392
rect -19648 -2472 -18560 -2408
rect -18496 -2472 -18476 -2408
rect -19648 -2488 -18476 -2472
rect -19648 -2552 -18560 -2488
rect -18496 -2552 -18476 -2488
rect -19648 -2568 -18476 -2552
rect -19648 -2632 -18560 -2568
rect -18496 -2632 -18476 -2568
rect -19648 -2680 -18476 -2632
rect -18236 -1848 -17064 -1800
rect -18236 -1912 -17148 -1848
rect -17084 -1912 -17064 -1848
rect -18236 -1928 -17064 -1912
rect -18236 -1992 -17148 -1928
rect -17084 -1992 -17064 -1928
rect -18236 -2008 -17064 -1992
rect -18236 -2072 -17148 -2008
rect -17084 -2072 -17064 -2008
rect -18236 -2088 -17064 -2072
rect -18236 -2152 -17148 -2088
rect -17084 -2152 -17064 -2088
rect -18236 -2168 -17064 -2152
rect -18236 -2232 -17148 -2168
rect -17084 -2232 -17064 -2168
rect -18236 -2248 -17064 -2232
rect -18236 -2312 -17148 -2248
rect -17084 -2312 -17064 -2248
rect -18236 -2328 -17064 -2312
rect -18236 -2392 -17148 -2328
rect -17084 -2392 -17064 -2328
rect -18236 -2408 -17064 -2392
rect -18236 -2472 -17148 -2408
rect -17084 -2472 -17064 -2408
rect -18236 -2488 -17064 -2472
rect -18236 -2552 -17148 -2488
rect -17084 -2552 -17064 -2488
rect -18236 -2568 -17064 -2552
rect -18236 -2632 -17148 -2568
rect -17084 -2632 -17064 -2568
rect -18236 -2680 -17064 -2632
rect -16824 -1848 -15652 -1800
rect -16824 -1912 -15736 -1848
rect -15672 -1912 -15652 -1848
rect -16824 -1928 -15652 -1912
rect -16824 -1992 -15736 -1928
rect -15672 -1992 -15652 -1928
rect -16824 -2008 -15652 -1992
rect -16824 -2072 -15736 -2008
rect -15672 -2072 -15652 -2008
rect -16824 -2088 -15652 -2072
rect -16824 -2152 -15736 -2088
rect -15672 -2152 -15652 -2088
rect -16824 -2168 -15652 -2152
rect -16824 -2232 -15736 -2168
rect -15672 -2232 -15652 -2168
rect -16824 -2248 -15652 -2232
rect -16824 -2312 -15736 -2248
rect -15672 -2312 -15652 -2248
rect -16824 -2328 -15652 -2312
rect -16824 -2392 -15736 -2328
rect -15672 -2392 -15652 -2328
rect -16824 -2408 -15652 -2392
rect -16824 -2472 -15736 -2408
rect -15672 -2472 -15652 -2408
rect -16824 -2488 -15652 -2472
rect -16824 -2552 -15736 -2488
rect -15672 -2552 -15652 -2488
rect -16824 -2568 -15652 -2552
rect -16824 -2632 -15736 -2568
rect -15672 -2632 -15652 -2568
rect -16824 -2680 -15652 -2632
rect -15412 -1848 -14240 -1800
rect -15412 -1912 -14324 -1848
rect -14260 -1912 -14240 -1848
rect -15412 -1928 -14240 -1912
rect -15412 -1992 -14324 -1928
rect -14260 -1992 -14240 -1928
rect -15412 -2008 -14240 -1992
rect -15412 -2072 -14324 -2008
rect -14260 -2072 -14240 -2008
rect -15412 -2088 -14240 -2072
rect -15412 -2152 -14324 -2088
rect -14260 -2152 -14240 -2088
rect -15412 -2168 -14240 -2152
rect -15412 -2232 -14324 -2168
rect -14260 -2232 -14240 -2168
rect -15412 -2248 -14240 -2232
rect -15412 -2312 -14324 -2248
rect -14260 -2312 -14240 -2248
rect -15412 -2328 -14240 -2312
rect -15412 -2392 -14324 -2328
rect -14260 -2392 -14240 -2328
rect -15412 -2408 -14240 -2392
rect -15412 -2472 -14324 -2408
rect -14260 -2472 -14240 -2408
rect -15412 -2488 -14240 -2472
rect -15412 -2552 -14324 -2488
rect -14260 -2552 -14240 -2488
rect -15412 -2568 -14240 -2552
rect -15412 -2632 -14324 -2568
rect -14260 -2632 -14240 -2568
rect -15412 -2680 -14240 -2632
rect -14000 -1848 -12828 -1800
rect -14000 -1912 -12912 -1848
rect -12848 -1912 -12828 -1848
rect -14000 -1928 -12828 -1912
rect -14000 -1992 -12912 -1928
rect -12848 -1992 -12828 -1928
rect -14000 -2008 -12828 -1992
rect -14000 -2072 -12912 -2008
rect -12848 -2072 -12828 -2008
rect -14000 -2088 -12828 -2072
rect -14000 -2152 -12912 -2088
rect -12848 -2152 -12828 -2088
rect -14000 -2168 -12828 -2152
rect -14000 -2232 -12912 -2168
rect -12848 -2232 -12828 -2168
rect -14000 -2248 -12828 -2232
rect -14000 -2312 -12912 -2248
rect -12848 -2312 -12828 -2248
rect -14000 -2328 -12828 -2312
rect -14000 -2392 -12912 -2328
rect -12848 -2392 -12828 -2328
rect -14000 -2408 -12828 -2392
rect -14000 -2472 -12912 -2408
rect -12848 -2472 -12828 -2408
rect -14000 -2488 -12828 -2472
rect -14000 -2552 -12912 -2488
rect -12848 -2552 -12828 -2488
rect -14000 -2568 -12828 -2552
rect -14000 -2632 -12912 -2568
rect -12848 -2632 -12828 -2568
rect -14000 -2680 -12828 -2632
rect -12588 -1848 -11416 -1800
rect -12588 -1912 -11500 -1848
rect -11436 -1912 -11416 -1848
rect -12588 -1928 -11416 -1912
rect -12588 -1992 -11500 -1928
rect -11436 -1992 -11416 -1928
rect -12588 -2008 -11416 -1992
rect -12588 -2072 -11500 -2008
rect -11436 -2072 -11416 -2008
rect -12588 -2088 -11416 -2072
rect -12588 -2152 -11500 -2088
rect -11436 -2152 -11416 -2088
rect -12588 -2168 -11416 -2152
rect -12588 -2232 -11500 -2168
rect -11436 -2232 -11416 -2168
rect -12588 -2248 -11416 -2232
rect -12588 -2312 -11500 -2248
rect -11436 -2312 -11416 -2248
rect -12588 -2328 -11416 -2312
rect -12588 -2392 -11500 -2328
rect -11436 -2392 -11416 -2328
rect -12588 -2408 -11416 -2392
rect -12588 -2472 -11500 -2408
rect -11436 -2472 -11416 -2408
rect -12588 -2488 -11416 -2472
rect -12588 -2552 -11500 -2488
rect -11436 -2552 -11416 -2488
rect -12588 -2568 -11416 -2552
rect -12588 -2632 -11500 -2568
rect -11436 -2632 -11416 -2568
rect -12588 -2680 -11416 -2632
rect -11176 -1848 -10004 -1800
rect -11176 -1912 -10088 -1848
rect -10024 -1912 -10004 -1848
rect -11176 -1928 -10004 -1912
rect -11176 -1992 -10088 -1928
rect -10024 -1992 -10004 -1928
rect -11176 -2008 -10004 -1992
rect -11176 -2072 -10088 -2008
rect -10024 -2072 -10004 -2008
rect -11176 -2088 -10004 -2072
rect -11176 -2152 -10088 -2088
rect -10024 -2152 -10004 -2088
rect -11176 -2168 -10004 -2152
rect -11176 -2232 -10088 -2168
rect -10024 -2232 -10004 -2168
rect -11176 -2248 -10004 -2232
rect -11176 -2312 -10088 -2248
rect -10024 -2312 -10004 -2248
rect -11176 -2328 -10004 -2312
rect -11176 -2392 -10088 -2328
rect -10024 -2392 -10004 -2328
rect -11176 -2408 -10004 -2392
rect -11176 -2472 -10088 -2408
rect -10024 -2472 -10004 -2408
rect -11176 -2488 -10004 -2472
rect -11176 -2552 -10088 -2488
rect -10024 -2552 -10004 -2488
rect -11176 -2568 -10004 -2552
rect -11176 -2632 -10088 -2568
rect -10024 -2632 -10004 -2568
rect -11176 -2680 -10004 -2632
rect -9764 -1848 -8592 -1800
rect -9764 -1912 -8676 -1848
rect -8612 -1912 -8592 -1848
rect -9764 -1928 -8592 -1912
rect -9764 -1992 -8676 -1928
rect -8612 -1992 -8592 -1928
rect -9764 -2008 -8592 -1992
rect -9764 -2072 -8676 -2008
rect -8612 -2072 -8592 -2008
rect -9764 -2088 -8592 -2072
rect -9764 -2152 -8676 -2088
rect -8612 -2152 -8592 -2088
rect -9764 -2168 -8592 -2152
rect -9764 -2232 -8676 -2168
rect -8612 -2232 -8592 -2168
rect -9764 -2248 -8592 -2232
rect -9764 -2312 -8676 -2248
rect -8612 -2312 -8592 -2248
rect -9764 -2328 -8592 -2312
rect -9764 -2392 -8676 -2328
rect -8612 -2392 -8592 -2328
rect -9764 -2408 -8592 -2392
rect -9764 -2472 -8676 -2408
rect -8612 -2472 -8592 -2408
rect -9764 -2488 -8592 -2472
rect -9764 -2552 -8676 -2488
rect -8612 -2552 -8592 -2488
rect -9764 -2568 -8592 -2552
rect -9764 -2632 -8676 -2568
rect -8612 -2632 -8592 -2568
rect -9764 -2680 -8592 -2632
rect -8352 -1848 -7180 -1800
rect -8352 -1912 -7264 -1848
rect -7200 -1912 -7180 -1848
rect -8352 -1928 -7180 -1912
rect -8352 -1992 -7264 -1928
rect -7200 -1992 -7180 -1928
rect -8352 -2008 -7180 -1992
rect -8352 -2072 -7264 -2008
rect -7200 -2072 -7180 -2008
rect -8352 -2088 -7180 -2072
rect -8352 -2152 -7264 -2088
rect -7200 -2152 -7180 -2088
rect -8352 -2168 -7180 -2152
rect -8352 -2232 -7264 -2168
rect -7200 -2232 -7180 -2168
rect -8352 -2248 -7180 -2232
rect -8352 -2312 -7264 -2248
rect -7200 -2312 -7180 -2248
rect -8352 -2328 -7180 -2312
rect -8352 -2392 -7264 -2328
rect -7200 -2392 -7180 -2328
rect -8352 -2408 -7180 -2392
rect -8352 -2472 -7264 -2408
rect -7200 -2472 -7180 -2408
rect -8352 -2488 -7180 -2472
rect -8352 -2552 -7264 -2488
rect -7200 -2552 -7180 -2488
rect -8352 -2568 -7180 -2552
rect -8352 -2632 -7264 -2568
rect -7200 -2632 -7180 -2568
rect -8352 -2680 -7180 -2632
rect -6940 -1848 -5768 -1800
rect -6940 -1912 -5852 -1848
rect -5788 -1912 -5768 -1848
rect -6940 -1928 -5768 -1912
rect -6940 -1992 -5852 -1928
rect -5788 -1992 -5768 -1928
rect -6940 -2008 -5768 -1992
rect -6940 -2072 -5852 -2008
rect -5788 -2072 -5768 -2008
rect -6940 -2088 -5768 -2072
rect -6940 -2152 -5852 -2088
rect -5788 -2152 -5768 -2088
rect -6940 -2168 -5768 -2152
rect -6940 -2232 -5852 -2168
rect -5788 -2232 -5768 -2168
rect -6940 -2248 -5768 -2232
rect -6940 -2312 -5852 -2248
rect -5788 -2312 -5768 -2248
rect -6940 -2328 -5768 -2312
rect -6940 -2392 -5852 -2328
rect -5788 -2392 -5768 -2328
rect -6940 -2408 -5768 -2392
rect -6940 -2472 -5852 -2408
rect -5788 -2472 -5768 -2408
rect -6940 -2488 -5768 -2472
rect -6940 -2552 -5852 -2488
rect -5788 -2552 -5768 -2488
rect -6940 -2568 -5768 -2552
rect -6940 -2632 -5852 -2568
rect -5788 -2632 -5768 -2568
rect -6940 -2680 -5768 -2632
rect -5528 -1848 -4356 -1800
rect -5528 -1912 -4440 -1848
rect -4376 -1912 -4356 -1848
rect -5528 -1928 -4356 -1912
rect -5528 -1992 -4440 -1928
rect -4376 -1992 -4356 -1928
rect -5528 -2008 -4356 -1992
rect -5528 -2072 -4440 -2008
rect -4376 -2072 -4356 -2008
rect -5528 -2088 -4356 -2072
rect -5528 -2152 -4440 -2088
rect -4376 -2152 -4356 -2088
rect -5528 -2168 -4356 -2152
rect -5528 -2232 -4440 -2168
rect -4376 -2232 -4356 -2168
rect -5528 -2248 -4356 -2232
rect -5528 -2312 -4440 -2248
rect -4376 -2312 -4356 -2248
rect -5528 -2328 -4356 -2312
rect -5528 -2392 -4440 -2328
rect -4376 -2392 -4356 -2328
rect -5528 -2408 -4356 -2392
rect -5528 -2472 -4440 -2408
rect -4376 -2472 -4356 -2408
rect -5528 -2488 -4356 -2472
rect -5528 -2552 -4440 -2488
rect -4376 -2552 -4356 -2488
rect -5528 -2568 -4356 -2552
rect -5528 -2632 -4440 -2568
rect -4376 -2632 -4356 -2568
rect -5528 -2680 -4356 -2632
rect -4116 -1848 -2944 -1800
rect -4116 -1912 -3028 -1848
rect -2964 -1912 -2944 -1848
rect -4116 -1928 -2944 -1912
rect -4116 -1992 -3028 -1928
rect -2964 -1992 -2944 -1928
rect -4116 -2008 -2944 -1992
rect -4116 -2072 -3028 -2008
rect -2964 -2072 -2944 -2008
rect -4116 -2088 -2944 -2072
rect -4116 -2152 -3028 -2088
rect -2964 -2152 -2944 -2088
rect -4116 -2168 -2944 -2152
rect -4116 -2232 -3028 -2168
rect -2964 -2232 -2944 -2168
rect -4116 -2248 -2944 -2232
rect -4116 -2312 -3028 -2248
rect -2964 -2312 -2944 -2248
rect -4116 -2328 -2944 -2312
rect -4116 -2392 -3028 -2328
rect -2964 -2392 -2944 -2328
rect -4116 -2408 -2944 -2392
rect -4116 -2472 -3028 -2408
rect -2964 -2472 -2944 -2408
rect -4116 -2488 -2944 -2472
rect -4116 -2552 -3028 -2488
rect -2964 -2552 -2944 -2488
rect -4116 -2568 -2944 -2552
rect -4116 -2632 -3028 -2568
rect -2964 -2632 -2944 -2568
rect -4116 -2680 -2944 -2632
rect -2704 -1848 -1532 -1800
rect -2704 -1912 -1616 -1848
rect -1552 -1912 -1532 -1848
rect -2704 -1928 -1532 -1912
rect -2704 -1992 -1616 -1928
rect -1552 -1992 -1532 -1928
rect -2704 -2008 -1532 -1992
rect -2704 -2072 -1616 -2008
rect -1552 -2072 -1532 -2008
rect -2704 -2088 -1532 -2072
rect -2704 -2152 -1616 -2088
rect -1552 -2152 -1532 -2088
rect -2704 -2168 -1532 -2152
rect -2704 -2232 -1616 -2168
rect -1552 -2232 -1532 -2168
rect -2704 -2248 -1532 -2232
rect -2704 -2312 -1616 -2248
rect -1552 -2312 -1532 -2248
rect -2704 -2328 -1532 -2312
rect -2704 -2392 -1616 -2328
rect -1552 -2392 -1532 -2328
rect -2704 -2408 -1532 -2392
rect -2704 -2472 -1616 -2408
rect -1552 -2472 -1532 -2408
rect -2704 -2488 -1532 -2472
rect -2704 -2552 -1616 -2488
rect -1552 -2552 -1532 -2488
rect -2704 -2568 -1532 -2552
rect -2704 -2632 -1616 -2568
rect -1552 -2632 -1532 -2568
rect -2704 -2680 -1532 -2632
rect -1292 -1848 -120 -1800
rect -1292 -1912 -204 -1848
rect -140 -1912 -120 -1848
rect -1292 -1928 -120 -1912
rect -1292 -1992 -204 -1928
rect -140 -1992 -120 -1928
rect -1292 -2008 -120 -1992
rect -1292 -2072 -204 -2008
rect -140 -2072 -120 -2008
rect -1292 -2088 -120 -2072
rect -1292 -2152 -204 -2088
rect -140 -2152 -120 -2088
rect -1292 -2168 -120 -2152
rect -1292 -2232 -204 -2168
rect -140 -2232 -120 -2168
rect -1292 -2248 -120 -2232
rect -1292 -2312 -204 -2248
rect -140 -2312 -120 -2248
rect -1292 -2328 -120 -2312
rect -1292 -2392 -204 -2328
rect -140 -2392 -120 -2328
rect -1292 -2408 -120 -2392
rect -1292 -2472 -204 -2408
rect -140 -2472 -120 -2408
rect -1292 -2488 -120 -2472
rect -1292 -2552 -204 -2488
rect -140 -2552 -120 -2488
rect -1292 -2568 -120 -2552
rect -1292 -2632 -204 -2568
rect -140 -2632 -120 -2568
rect -1292 -2680 -120 -2632
rect 120 -1848 1292 -1800
rect 120 -1912 1208 -1848
rect 1272 -1912 1292 -1848
rect 120 -1928 1292 -1912
rect 120 -1992 1208 -1928
rect 1272 -1992 1292 -1928
rect 120 -2008 1292 -1992
rect 120 -2072 1208 -2008
rect 1272 -2072 1292 -2008
rect 120 -2088 1292 -2072
rect 120 -2152 1208 -2088
rect 1272 -2152 1292 -2088
rect 120 -2168 1292 -2152
rect 120 -2232 1208 -2168
rect 1272 -2232 1292 -2168
rect 120 -2248 1292 -2232
rect 120 -2312 1208 -2248
rect 1272 -2312 1292 -2248
rect 120 -2328 1292 -2312
rect 120 -2392 1208 -2328
rect 1272 -2392 1292 -2328
rect 120 -2408 1292 -2392
rect 120 -2472 1208 -2408
rect 1272 -2472 1292 -2408
rect 120 -2488 1292 -2472
rect 120 -2552 1208 -2488
rect 1272 -2552 1292 -2488
rect 120 -2568 1292 -2552
rect 120 -2632 1208 -2568
rect 1272 -2632 1292 -2568
rect 120 -2680 1292 -2632
rect 1532 -1848 2704 -1800
rect 1532 -1912 2620 -1848
rect 2684 -1912 2704 -1848
rect 1532 -1928 2704 -1912
rect 1532 -1992 2620 -1928
rect 2684 -1992 2704 -1928
rect 1532 -2008 2704 -1992
rect 1532 -2072 2620 -2008
rect 2684 -2072 2704 -2008
rect 1532 -2088 2704 -2072
rect 1532 -2152 2620 -2088
rect 2684 -2152 2704 -2088
rect 1532 -2168 2704 -2152
rect 1532 -2232 2620 -2168
rect 2684 -2232 2704 -2168
rect 1532 -2248 2704 -2232
rect 1532 -2312 2620 -2248
rect 2684 -2312 2704 -2248
rect 1532 -2328 2704 -2312
rect 1532 -2392 2620 -2328
rect 2684 -2392 2704 -2328
rect 1532 -2408 2704 -2392
rect 1532 -2472 2620 -2408
rect 2684 -2472 2704 -2408
rect 1532 -2488 2704 -2472
rect 1532 -2552 2620 -2488
rect 2684 -2552 2704 -2488
rect 1532 -2568 2704 -2552
rect 1532 -2632 2620 -2568
rect 2684 -2632 2704 -2568
rect 1532 -2680 2704 -2632
rect 2944 -1848 4116 -1800
rect 2944 -1912 4032 -1848
rect 4096 -1912 4116 -1848
rect 2944 -1928 4116 -1912
rect 2944 -1992 4032 -1928
rect 4096 -1992 4116 -1928
rect 2944 -2008 4116 -1992
rect 2944 -2072 4032 -2008
rect 4096 -2072 4116 -2008
rect 2944 -2088 4116 -2072
rect 2944 -2152 4032 -2088
rect 4096 -2152 4116 -2088
rect 2944 -2168 4116 -2152
rect 2944 -2232 4032 -2168
rect 4096 -2232 4116 -2168
rect 2944 -2248 4116 -2232
rect 2944 -2312 4032 -2248
rect 4096 -2312 4116 -2248
rect 2944 -2328 4116 -2312
rect 2944 -2392 4032 -2328
rect 4096 -2392 4116 -2328
rect 2944 -2408 4116 -2392
rect 2944 -2472 4032 -2408
rect 4096 -2472 4116 -2408
rect 2944 -2488 4116 -2472
rect 2944 -2552 4032 -2488
rect 4096 -2552 4116 -2488
rect 2944 -2568 4116 -2552
rect 2944 -2632 4032 -2568
rect 4096 -2632 4116 -2568
rect 2944 -2680 4116 -2632
rect 4356 -1848 5528 -1800
rect 4356 -1912 5444 -1848
rect 5508 -1912 5528 -1848
rect 4356 -1928 5528 -1912
rect 4356 -1992 5444 -1928
rect 5508 -1992 5528 -1928
rect 4356 -2008 5528 -1992
rect 4356 -2072 5444 -2008
rect 5508 -2072 5528 -2008
rect 4356 -2088 5528 -2072
rect 4356 -2152 5444 -2088
rect 5508 -2152 5528 -2088
rect 4356 -2168 5528 -2152
rect 4356 -2232 5444 -2168
rect 5508 -2232 5528 -2168
rect 4356 -2248 5528 -2232
rect 4356 -2312 5444 -2248
rect 5508 -2312 5528 -2248
rect 4356 -2328 5528 -2312
rect 4356 -2392 5444 -2328
rect 5508 -2392 5528 -2328
rect 4356 -2408 5528 -2392
rect 4356 -2472 5444 -2408
rect 5508 -2472 5528 -2408
rect 4356 -2488 5528 -2472
rect 4356 -2552 5444 -2488
rect 5508 -2552 5528 -2488
rect 4356 -2568 5528 -2552
rect 4356 -2632 5444 -2568
rect 5508 -2632 5528 -2568
rect 4356 -2680 5528 -2632
rect 5768 -1848 6940 -1800
rect 5768 -1912 6856 -1848
rect 6920 -1912 6940 -1848
rect 5768 -1928 6940 -1912
rect 5768 -1992 6856 -1928
rect 6920 -1992 6940 -1928
rect 5768 -2008 6940 -1992
rect 5768 -2072 6856 -2008
rect 6920 -2072 6940 -2008
rect 5768 -2088 6940 -2072
rect 5768 -2152 6856 -2088
rect 6920 -2152 6940 -2088
rect 5768 -2168 6940 -2152
rect 5768 -2232 6856 -2168
rect 6920 -2232 6940 -2168
rect 5768 -2248 6940 -2232
rect 5768 -2312 6856 -2248
rect 6920 -2312 6940 -2248
rect 5768 -2328 6940 -2312
rect 5768 -2392 6856 -2328
rect 6920 -2392 6940 -2328
rect 5768 -2408 6940 -2392
rect 5768 -2472 6856 -2408
rect 6920 -2472 6940 -2408
rect 5768 -2488 6940 -2472
rect 5768 -2552 6856 -2488
rect 6920 -2552 6940 -2488
rect 5768 -2568 6940 -2552
rect 5768 -2632 6856 -2568
rect 6920 -2632 6940 -2568
rect 5768 -2680 6940 -2632
rect 7180 -1848 8352 -1800
rect 7180 -1912 8268 -1848
rect 8332 -1912 8352 -1848
rect 7180 -1928 8352 -1912
rect 7180 -1992 8268 -1928
rect 8332 -1992 8352 -1928
rect 7180 -2008 8352 -1992
rect 7180 -2072 8268 -2008
rect 8332 -2072 8352 -2008
rect 7180 -2088 8352 -2072
rect 7180 -2152 8268 -2088
rect 8332 -2152 8352 -2088
rect 7180 -2168 8352 -2152
rect 7180 -2232 8268 -2168
rect 8332 -2232 8352 -2168
rect 7180 -2248 8352 -2232
rect 7180 -2312 8268 -2248
rect 8332 -2312 8352 -2248
rect 7180 -2328 8352 -2312
rect 7180 -2392 8268 -2328
rect 8332 -2392 8352 -2328
rect 7180 -2408 8352 -2392
rect 7180 -2472 8268 -2408
rect 8332 -2472 8352 -2408
rect 7180 -2488 8352 -2472
rect 7180 -2552 8268 -2488
rect 8332 -2552 8352 -2488
rect 7180 -2568 8352 -2552
rect 7180 -2632 8268 -2568
rect 8332 -2632 8352 -2568
rect 7180 -2680 8352 -2632
rect 8592 -1848 9764 -1800
rect 8592 -1912 9680 -1848
rect 9744 -1912 9764 -1848
rect 8592 -1928 9764 -1912
rect 8592 -1992 9680 -1928
rect 9744 -1992 9764 -1928
rect 8592 -2008 9764 -1992
rect 8592 -2072 9680 -2008
rect 9744 -2072 9764 -2008
rect 8592 -2088 9764 -2072
rect 8592 -2152 9680 -2088
rect 9744 -2152 9764 -2088
rect 8592 -2168 9764 -2152
rect 8592 -2232 9680 -2168
rect 9744 -2232 9764 -2168
rect 8592 -2248 9764 -2232
rect 8592 -2312 9680 -2248
rect 9744 -2312 9764 -2248
rect 8592 -2328 9764 -2312
rect 8592 -2392 9680 -2328
rect 9744 -2392 9764 -2328
rect 8592 -2408 9764 -2392
rect 8592 -2472 9680 -2408
rect 9744 -2472 9764 -2408
rect 8592 -2488 9764 -2472
rect 8592 -2552 9680 -2488
rect 9744 -2552 9764 -2488
rect 8592 -2568 9764 -2552
rect 8592 -2632 9680 -2568
rect 9744 -2632 9764 -2568
rect 8592 -2680 9764 -2632
rect 10004 -1848 11176 -1800
rect 10004 -1912 11092 -1848
rect 11156 -1912 11176 -1848
rect 10004 -1928 11176 -1912
rect 10004 -1992 11092 -1928
rect 11156 -1992 11176 -1928
rect 10004 -2008 11176 -1992
rect 10004 -2072 11092 -2008
rect 11156 -2072 11176 -2008
rect 10004 -2088 11176 -2072
rect 10004 -2152 11092 -2088
rect 11156 -2152 11176 -2088
rect 10004 -2168 11176 -2152
rect 10004 -2232 11092 -2168
rect 11156 -2232 11176 -2168
rect 10004 -2248 11176 -2232
rect 10004 -2312 11092 -2248
rect 11156 -2312 11176 -2248
rect 10004 -2328 11176 -2312
rect 10004 -2392 11092 -2328
rect 11156 -2392 11176 -2328
rect 10004 -2408 11176 -2392
rect 10004 -2472 11092 -2408
rect 11156 -2472 11176 -2408
rect 10004 -2488 11176 -2472
rect 10004 -2552 11092 -2488
rect 11156 -2552 11176 -2488
rect 10004 -2568 11176 -2552
rect 10004 -2632 11092 -2568
rect 11156 -2632 11176 -2568
rect 10004 -2680 11176 -2632
rect 11416 -1848 12588 -1800
rect 11416 -1912 12504 -1848
rect 12568 -1912 12588 -1848
rect 11416 -1928 12588 -1912
rect 11416 -1992 12504 -1928
rect 12568 -1992 12588 -1928
rect 11416 -2008 12588 -1992
rect 11416 -2072 12504 -2008
rect 12568 -2072 12588 -2008
rect 11416 -2088 12588 -2072
rect 11416 -2152 12504 -2088
rect 12568 -2152 12588 -2088
rect 11416 -2168 12588 -2152
rect 11416 -2232 12504 -2168
rect 12568 -2232 12588 -2168
rect 11416 -2248 12588 -2232
rect 11416 -2312 12504 -2248
rect 12568 -2312 12588 -2248
rect 11416 -2328 12588 -2312
rect 11416 -2392 12504 -2328
rect 12568 -2392 12588 -2328
rect 11416 -2408 12588 -2392
rect 11416 -2472 12504 -2408
rect 12568 -2472 12588 -2408
rect 11416 -2488 12588 -2472
rect 11416 -2552 12504 -2488
rect 12568 -2552 12588 -2488
rect 11416 -2568 12588 -2552
rect 11416 -2632 12504 -2568
rect 12568 -2632 12588 -2568
rect 11416 -2680 12588 -2632
rect 12828 -1848 14000 -1800
rect 12828 -1912 13916 -1848
rect 13980 -1912 14000 -1848
rect 12828 -1928 14000 -1912
rect 12828 -1992 13916 -1928
rect 13980 -1992 14000 -1928
rect 12828 -2008 14000 -1992
rect 12828 -2072 13916 -2008
rect 13980 -2072 14000 -2008
rect 12828 -2088 14000 -2072
rect 12828 -2152 13916 -2088
rect 13980 -2152 14000 -2088
rect 12828 -2168 14000 -2152
rect 12828 -2232 13916 -2168
rect 13980 -2232 14000 -2168
rect 12828 -2248 14000 -2232
rect 12828 -2312 13916 -2248
rect 13980 -2312 14000 -2248
rect 12828 -2328 14000 -2312
rect 12828 -2392 13916 -2328
rect 13980 -2392 14000 -2328
rect 12828 -2408 14000 -2392
rect 12828 -2472 13916 -2408
rect 13980 -2472 14000 -2408
rect 12828 -2488 14000 -2472
rect 12828 -2552 13916 -2488
rect 13980 -2552 14000 -2488
rect 12828 -2568 14000 -2552
rect 12828 -2632 13916 -2568
rect 13980 -2632 14000 -2568
rect 12828 -2680 14000 -2632
rect 14240 -1848 15412 -1800
rect 14240 -1912 15328 -1848
rect 15392 -1912 15412 -1848
rect 14240 -1928 15412 -1912
rect 14240 -1992 15328 -1928
rect 15392 -1992 15412 -1928
rect 14240 -2008 15412 -1992
rect 14240 -2072 15328 -2008
rect 15392 -2072 15412 -2008
rect 14240 -2088 15412 -2072
rect 14240 -2152 15328 -2088
rect 15392 -2152 15412 -2088
rect 14240 -2168 15412 -2152
rect 14240 -2232 15328 -2168
rect 15392 -2232 15412 -2168
rect 14240 -2248 15412 -2232
rect 14240 -2312 15328 -2248
rect 15392 -2312 15412 -2248
rect 14240 -2328 15412 -2312
rect 14240 -2392 15328 -2328
rect 15392 -2392 15412 -2328
rect 14240 -2408 15412 -2392
rect 14240 -2472 15328 -2408
rect 15392 -2472 15412 -2408
rect 14240 -2488 15412 -2472
rect 14240 -2552 15328 -2488
rect 15392 -2552 15412 -2488
rect 14240 -2568 15412 -2552
rect 14240 -2632 15328 -2568
rect 15392 -2632 15412 -2568
rect 14240 -2680 15412 -2632
rect 15652 -1848 16824 -1800
rect 15652 -1912 16740 -1848
rect 16804 -1912 16824 -1848
rect 15652 -1928 16824 -1912
rect 15652 -1992 16740 -1928
rect 16804 -1992 16824 -1928
rect 15652 -2008 16824 -1992
rect 15652 -2072 16740 -2008
rect 16804 -2072 16824 -2008
rect 15652 -2088 16824 -2072
rect 15652 -2152 16740 -2088
rect 16804 -2152 16824 -2088
rect 15652 -2168 16824 -2152
rect 15652 -2232 16740 -2168
rect 16804 -2232 16824 -2168
rect 15652 -2248 16824 -2232
rect 15652 -2312 16740 -2248
rect 16804 -2312 16824 -2248
rect 15652 -2328 16824 -2312
rect 15652 -2392 16740 -2328
rect 16804 -2392 16824 -2328
rect 15652 -2408 16824 -2392
rect 15652 -2472 16740 -2408
rect 16804 -2472 16824 -2408
rect 15652 -2488 16824 -2472
rect 15652 -2552 16740 -2488
rect 16804 -2552 16824 -2488
rect 15652 -2568 16824 -2552
rect 15652 -2632 16740 -2568
rect 16804 -2632 16824 -2568
rect 15652 -2680 16824 -2632
rect 17064 -1848 18236 -1800
rect 17064 -1912 18152 -1848
rect 18216 -1912 18236 -1848
rect 17064 -1928 18236 -1912
rect 17064 -1992 18152 -1928
rect 18216 -1992 18236 -1928
rect 17064 -2008 18236 -1992
rect 17064 -2072 18152 -2008
rect 18216 -2072 18236 -2008
rect 17064 -2088 18236 -2072
rect 17064 -2152 18152 -2088
rect 18216 -2152 18236 -2088
rect 17064 -2168 18236 -2152
rect 17064 -2232 18152 -2168
rect 18216 -2232 18236 -2168
rect 17064 -2248 18236 -2232
rect 17064 -2312 18152 -2248
rect 18216 -2312 18236 -2248
rect 17064 -2328 18236 -2312
rect 17064 -2392 18152 -2328
rect 18216 -2392 18236 -2328
rect 17064 -2408 18236 -2392
rect 17064 -2472 18152 -2408
rect 18216 -2472 18236 -2408
rect 17064 -2488 18236 -2472
rect 17064 -2552 18152 -2488
rect 18216 -2552 18236 -2488
rect 17064 -2568 18236 -2552
rect 17064 -2632 18152 -2568
rect 18216 -2632 18236 -2568
rect 17064 -2680 18236 -2632
rect 18476 -1848 19648 -1800
rect 18476 -1912 19564 -1848
rect 19628 -1912 19648 -1848
rect 18476 -1928 19648 -1912
rect 18476 -1992 19564 -1928
rect 19628 -1992 19648 -1928
rect 18476 -2008 19648 -1992
rect 18476 -2072 19564 -2008
rect 19628 -2072 19648 -2008
rect 18476 -2088 19648 -2072
rect 18476 -2152 19564 -2088
rect 19628 -2152 19648 -2088
rect 18476 -2168 19648 -2152
rect 18476 -2232 19564 -2168
rect 19628 -2232 19648 -2168
rect 18476 -2248 19648 -2232
rect 18476 -2312 19564 -2248
rect 19628 -2312 19648 -2248
rect 18476 -2328 19648 -2312
rect 18476 -2392 19564 -2328
rect 19628 -2392 19648 -2328
rect 18476 -2408 19648 -2392
rect 18476 -2472 19564 -2408
rect 19628 -2472 19648 -2408
rect 18476 -2488 19648 -2472
rect 18476 -2552 19564 -2488
rect 19628 -2552 19648 -2488
rect 18476 -2568 19648 -2552
rect 18476 -2632 19564 -2568
rect 19628 -2632 19648 -2568
rect 18476 -2680 19648 -2632
rect 19888 -1848 21060 -1800
rect 19888 -1912 20976 -1848
rect 21040 -1912 21060 -1848
rect 19888 -1928 21060 -1912
rect 19888 -1992 20976 -1928
rect 21040 -1992 21060 -1928
rect 19888 -2008 21060 -1992
rect 19888 -2072 20976 -2008
rect 21040 -2072 21060 -2008
rect 19888 -2088 21060 -2072
rect 19888 -2152 20976 -2088
rect 21040 -2152 21060 -2088
rect 19888 -2168 21060 -2152
rect 19888 -2232 20976 -2168
rect 21040 -2232 21060 -2168
rect 19888 -2248 21060 -2232
rect 19888 -2312 20976 -2248
rect 21040 -2312 21060 -2248
rect 19888 -2328 21060 -2312
rect 19888 -2392 20976 -2328
rect 21040 -2392 21060 -2328
rect 19888 -2408 21060 -2392
rect 19888 -2472 20976 -2408
rect 21040 -2472 21060 -2408
rect 19888 -2488 21060 -2472
rect 19888 -2552 20976 -2488
rect 21040 -2552 21060 -2488
rect 19888 -2568 21060 -2552
rect 19888 -2632 20976 -2568
rect 21040 -2632 21060 -2568
rect 19888 -2680 21060 -2632
rect 21300 -1848 22472 -1800
rect 21300 -1912 22388 -1848
rect 22452 -1912 22472 -1848
rect 21300 -1928 22472 -1912
rect 21300 -1992 22388 -1928
rect 22452 -1992 22472 -1928
rect 21300 -2008 22472 -1992
rect 21300 -2072 22388 -2008
rect 22452 -2072 22472 -2008
rect 21300 -2088 22472 -2072
rect 21300 -2152 22388 -2088
rect 22452 -2152 22472 -2088
rect 21300 -2168 22472 -2152
rect 21300 -2232 22388 -2168
rect 22452 -2232 22472 -2168
rect 21300 -2248 22472 -2232
rect 21300 -2312 22388 -2248
rect 22452 -2312 22472 -2248
rect 21300 -2328 22472 -2312
rect 21300 -2392 22388 -2328
rect 22452 -2392 22472 -2328
rect 21300 -2408 22472 -2392
rect 21300 -2472 22388 -2408
rect 22452 -2472 22472 -2408
rect 21300 -2488 22472 -2472
rect 21300 -2552 22388 -2488
rect 22452 -2552 22472 -2488
rect 21300 -2568 22472 -2552
rect 21300 -2632 22388 -2568
rect 22452 -2632 22472 -2568
rect 21300 -2680 22472 -2632
rect 22712 -1848 23884 -1800
rect 22712 -1912 23800 -1848
rect 23864 -1912 23884 -1848
rect 22712 -1928 23884 -1912
rect 22712 -1992 23800 -1928
rect 23864 -1992 23884 -1928
rect 22712 -2008 23884 -1992
rect 22712 -2072 23800 -2008
rect 23864 -2072 23884 -2008
rect 22712 -2088 23884 -2072
rect 22712 -2152 23800 -2088
rect 23864 -2152 23884 -2088
rect 22712 -2168 23884 -2152
rect 22712 -2232 23800 -2168
rect 23864 -2232 23884 -2168
rect 22712 -2248 23884 -2232
rect 22712 -2312 23800 -2248
rect 23864 -2312 23884 -2248
rect 22712 -2328 23884 -2312
rect 22712 -2392 23800 -2328
rect 23864 -2392 23884 -2328
rect 22712 -2408 23884 -2392
rect 22712 -2472 23800 -2408
rect 23864 -2472 23884 -2408
rect 22712 -2488 23884 -2472
rect 22712 -2552 23800 -2488
rect 23864 -2552 23884 -2488
rect 22712 -2568 23884 -2552
rect 22712 -2632 23800 -2568
rect 23864 -2632 23884 -2568
rect 22712 -2680 23884 -2632
rect -23884 -2968 -22712 -2920
rect -23884 -3032 -22796 -2968
rect -22732 -3032 -22712 -2968
rect -23884 -3048 -22712 -3032
rect -23884 -3112 -22796 -3048
rect -22732 -3112 -22712 -3048
rect -23884 -3128 -22712 -3112
rect -23884 -3192 -22796 -3128
rect -22732 -3192 -22712 -3128
rect -23884 -3208 -22712 -3192
rect -23884 -3272 -22796 -3208
rect -22732 -3272 -22712 -3208
rect -23884 -3288 -22712 -3272
rect -23884 -3352 -22796 -3288
rect -22732 -3352 -22712 -3288
rect -23884 -3368 -22712 -3352
rect -23884 -3432 -22796 -3368
rect -22732 -3432 -22712 -3368
rect -23884 -3448 -22712 -3432
rect -23884 -3512 -22796 -3448
rect -22732 -3512 -22712 -3448
rect -23884 -3528 -22712 -3512
rect -23884 -3592 -22796 -3528
rect -22732 -3592 -22712 -3528
rect -23884 -3608 -22712 -3592
rect -23884 -3672 -22796 -3608
rect -22732 -3672 -22712 -3608
rect -23884 -3688 -22712 -3672
rect -23884 -3752 -22796 -3688
rect -22732 -3752 -22712 -3688
rect -23884 -3800 -22712 -3752
rect -22472 -2968 -21300 -2920
rect -22472 -3032 -21384 -2968
rect -21320 -3032 -21300 -2968
rect -22472 -3048 -21300 -3032
rect -22472 -3112 -21384 -3048
rect -21320 -3112 -21300 -3048
rect -22472 -3128 -21300 -3112
rect -22472 -3192 -21384 -3128
rect -21320 -3192 -21300 -3128
rect -22472 -3208 -21300 -3192
rect -22472 -3272 -21384 -3208
rect -21320 -3272 -21300 -3208
rect -22472 -3288 -21300 -3272
rect -22472 -3352 -21384 -3288
rect -21320 -3352 -21300 -3288
rect -22472 -3368 -21300 -3352
rect -22472 -3432 -21384 -3368
rect -21320 -3432 -21300 -3368
rect -22472 -3448 -21300 -3432
rect -22472 -3512 -21384 -3448
rect -21320 -3512 -21300 -3448
rect -22472 -3528 -21300 -3512
rect -22472 -3592 -21384 -3528
rect -21320 -3592 -21300 -3528
rect -22472 -3608 -21300 -3592
rect -22472 -3672 -21384 -3608
rect -21320 -3672 -21300 -3608
rect -22472 -3688 -21300 -3672
rect -22472 -3752 -21384 -3688
rect -21320 -3752 -21300 -3688
rect -22472 -3800 -21300 -3752
rect -21060 -2968 -19888 -2920
rect -21060 -3032 -19972 -2968
rect -19908 -3032 -19888 -2968
rect -21060 -3048 -19888 -3032
rect -21060 -3112 -19972 -3048
rect -19908 -3112 -19888 -3048
rect -21060 -3128 -19888 -3112
rect -21060 -3192 -19972 -3128
rect -19908 -3192 -19888 -3128
rect -21060 -3208 -19888 -3192
rect -21060 -3272 -19972 -3208
rect -19908 -3272 -19888 -3208
rect -21060 -3288 -19888 -3272
rect -21060 -3352 -19972 -3288
rect -19908 -3352 -19888 -3288
rect -21060 -3368 -19888 -3352
rect -21060 -3432 -19972 -3368
rect -19908 -3432 -19888 -3368
rect -21060 -3448 -19888 -3432
rect -21060 -3512 -19972 -3448
rect -19908 -3512 -19888 -3448
rect -21060 -3528 -19888 -3512
rect -21060 -3592 -19972 -3528
rect -19908 -3592 -19888 -3528
rect -21060 -3608 -19888 -3592
rect -21060 -3672 -19972 -3608
rect -19908 -3672 -19888 -3608
rect -21060 -3688 -19888 -3672
rect -21060 -3752 -19972 -3688
rect -19908 -3752 -19888 -3688
rect -21060 -3800 -19888 -3752
rect -19648 -2968 -18476 -2920
rect -19648 -3032 -18560 -2968
rect -18496 -3032 -18476 -2968
rect -19648 -3048 -18476 -3032
rect -19648 -3112 -18560 -3048
rect -18496 -3112 -18476 -3048
rect -19648 -3128 -18476 -3112
rect -19648 -3192 -18560 -3128
rect -18496 -3192 -18476 -3128
rect -19648 -3208 -18476 -3192
rect -19648 -3272 -18560 -3208
rect -18496 -3272 -18476 -3208
rect -19648 -3288 -18476 -3272
rect -19648 -3352 -18560 -3288
rect -18496 -3352 -18476 -3288
rect -19648 -3368 -18476 -3352
rect -19648 -3432 -18560 -3368
rect -18496 -3432 -18476 -3368
rect -19648 -3448 -18476 -3432
rect -19648 -3512 -18560 -3448
rect -18496 -3512 -18476 -3448
rect -19648 -3528 -18476 -3512
rect -19648 -3592 -18560 -3528
rect -18496 -3592 -18476 -3528
rect -19648 -3608 -18476 -3592
rect -19648 -3672 -18560 -3608
rect -18496 -3672 -18476 -3608
rect -19648 -3688 -18476 -3672
rect -19648 -3752 -18560 -3688
rect -18496 -3752 -18476 -3688
rect -19648 -3800 -18476 -3752
rect -18236 -2968 -17064 -2920
rect -18236 -3032 -17148 -2968
rect -17084 -3032 -17064 -2968
rect -18236 -3048 -17064 -3032
rect -18236 -3112 -17148 -3048
rect -17084 -3112 -17064 -3048
rect -18236 -3128 -17064 -3112
rect -18236 -3192 -17148 -3128
rect -17084 -3192 -17064 -3128
rect -18236 -3208 -17064 -3192
rect -18236 -3272 -17148 -3208
rect -17084 -3272 -17064 -3208
rect -18236 -3288 -17064 -3272
rect -18236 -3352 -17148 -3288
rect -17084 -3352 -17064 -3288
rect -18236 -3368 -17064 -3352
rect -18236 -3432 -17148 -3368
rect -17084 -3432 -17064 -3368
rect -18236 -3448 -17064 -3432
rect -18236 -3512 -17148 -3448
rect -17084 -3512 -17064 -3448
rect -18236 -3528 -17064 -3512
rect -18236 -3592 -17148 -3528
rect -17084 -3592 -17064 -3528
rect -18236 -3608 -17064 -3592
rect -18236 -3672 -17148 -3608
rect -17084 -3672 -17064 -3608
rect -18236 -3688 -17064 -3672
rect -18236 -3752 -17148 -3688
rect -17084 -3752 -17064 -3688
rect -18236 -3800 -17064 -3752
rect -16824 -2968 -15652 -2920
rect -16824 -3032 -15736 -2968
rect -15672 -3032 -15652 -2968
rect -16824 -3048 -15652 -3032
rect -16824 -3112 -15736 -3048
rect -15672 -3112 -15652 -3048
rect -16824 -3128 -15652 -3112
rect -16824 -3192 -15736 -3128
rect -15672 -3192 -15652 -3128
rect -16824 -3208 -15652 -3192
rect -16824 -3272 -15736 -3208
rect -15672 -3272 -15652 -3208
rect -16824 -3288 -15652 -3272
rect -16824 -3352 -15736 -3288
rect -15672 -3352 -15652 -3288
rect -16824 -3368 -15652 -3352
rect -16824 -3432 -15736 -3368
rect -15672 -3432 -15652 -3368
rect -16824 -3448 -15652 -3432
rect -16824 -3512 -15736 -3448
rect -15672 -3512 -15652 -3448
rect -16824 -3528 -15652 -3512
rect -16824 -3592 -15736 -3528
rect -15672 -3592 -15652 -3528
rect -16824 -3608 -15652 -3592
rect -16824 -3672 -15736 -3608
rect -15672 -3672 -15652 -3608
rect -16824 -3688 -15652 -3672
rect -16824 -3752 -15736 -3688
rect -15672 -3752 -15652 -3688
rect -16824 -3800 -15652 -3752
rect -15412 -2968 -14240 -2920
rect -15412 -3032 -14324 -2968
rect -14260 -3032 -14240 -2968
rect -15412 -3048 -14240 -3032
rect -15412 -3112 -14324 -3048
rect -14260 -3112 -14240 -3048
rect -15412 -3128 -14240 -3112
rect -15412 -3192 -14324 -3128
rect -14260 -3192 -14240 -3128
rect -15412 -3208 -14240 -3192
rect -15412 -3272 -14324 -3208
rect -14260 -3272 -14240 -3208
rect -15412 -3288 -14240 -3272
rect -15412 -3352 -14324 -3288
rect -14260 -3352 -14240 -3288
rect -15412 -3368 -14240 -3352
rect -15412 -3432 -14324 -3368
rect -14260 -3432 -14240 -3368
rect -15412 -3448 -14240 -3432
rect -15412 -3512 -14324 -3448
rect -14260 -3512 -14240 -3448
rect -15412 -3528 -14240 -3512
rect -15412 -3592 -14324 -3528
rect -14260 -3592 -14240 -3528
rect -15412 -3608 -14240 -3592
rect -15412 -3672 -14324 -3608
rect -14260 -3672 -14240 -3608
rect -15412 -3688 -14240 -3672
rect -15412 -3752 -14324 -3688
rect -14260 -3752 -14240 -3688
rect -15412 -3800 -14240 -3752
rect -14000 -2968 -12828 -2920
rect -14000 -3032 -12912 -2968
rect -12848 -3032 -12828 -2968
rect -14000 -3048 -12828 -3032
rect -14000 -3112 -12912 -3048
rect -12848 -3112 -12828 -3048
rect -14000 -3128 -12828 -3112
rect -14000 -3192 -12912 -3128
rect -12848 -3192 -12828 -3128
rect -14000 -3208 -12828 -3192
rect -14000 -3272 -12912 -3208
rect -12848 -3272 -12828 -3208
rect -14000 -3288 -12828 -3272
rect -14000 -3352 -12912 -3288
rect -12848 -3352 -12828 -3288
rect -14000 -3368 -12828 -3352
rect -14000 -3432 -12912 -3368
rect -12848 -3432 -12828 -3368
rect -14000 -3448 -12828 -3432
rect -14000 -3512 -12912 -3448
rect -12848 -3512 -12828 -3448
rect -14000 -3528 -12828 -3512
rect -14000 -3592 -12912 -3528
rect -12848 -3592 -12828 -3528
rect -14000 -3608 -12828 -3592
rect -14000 -3672 -12912 -3608
rect -12848 -3672 -12828 -3608
rect -14000 -3688 -12828 -3672
rect -14000 -3752 -12912 -3688
rect -12848 -3752 -12828 -3688
rect -14000 -3800 -12828 -3752
rect -12588 -2968 -11416 -2920
rect -12588 -3032 -11500 -2968
rect -11436 -3032 -11416 -2968
rect -12588 -3048 -11416 -3032
rect -12588 -3112 -11500 -3048
rect -11436 -3112 -11416 -3048
rect -12588 -3128 -11416 -3112
rect -12588 -3192 -11500 -3128
rect -11436 -3192 -11416 -3128
rect -12588 -3208 -11416 -3192
rect -12588 -3272 -11500 -3208
rect -11436 -3272 -11416 -3208
rect -12588 -3288 -11416 -3272
rect -12588 -3352 -11500 -3288
rect -11436 -3352 -11416 -3288
rect -12588 -3368 -11416 -3352
rect -12588 -3432 -11500 -3368
rect -11436 -3432 -11416 -3368
rect -12588 -3448 -11416 -3432
rect -12588 -3512 -11500 -3448
rect -11436 -3512 -11416 -3448
rect -12588 -3528 -11416 -3512
rect -12588 -3592 -11500 -3528
rect -11436 -3592 -11416 -3528
rect -12588 -3608 -11416 -3592
rect -12588 -3672 -11500 -3608
rect -11436 -3672 -11416 -3608
rect -12588 -3688 -11416 -3672
rect -12588 -3752 -11500 -3688
rect -11436 -3752 -11416 -3688
rect -12588 -3800 -11416 -3752
rect -11176 -2968 -10004 -2920
rect -11176 -3032 -10088 -2968
rect -10024 -3032 -10004 -2968
rect -11176 -3048 -10004 -3032
rect -11176 -3112 -10088 -3048
rect -10024 -3112 -10004 -3048
rect -11176 -3128 -10004 -3112
rect -11176 -3192 -10088 -3128
rect -10024 -3192 -10004 -3128
rect -11176 -3208 -10004 -3192
rect -11176 -3272 -10088 -3208
rect -10024 -3272 -10004 -3208
rect -11176 -3288 -10004 -3272
rect -11176 -3352 -10088 -3288
rect -10024 -3352 -10004 -3288
rect -11176 -3368 -10004 -3352
rect -11176 -3432 -10088 -3368
rect -10024 -3432 -10004 -3368
rect -11176 -3448 -10004 -3432
rect -11176 -3512 -10088 -3448
rect -10024 -3512 -10004 -3448
rect -11176 -3528 -10004 -3512
rect -11176 -3592 -10088 -3528
rect -10024 -3592 -10004 -3528
rect -11176 -3608 -10004 -3592
rect -11176 -3672 -10088 -3608
rect -10024 -3672 -10004 -3608
rect -11176 -3688 -10004 -3672
rect -11176 -3752 -10088 -3688
rect -10024 -3752 -10004 -3688
rect -11176 -3800 -10004 -3752
rect -9764 -2968 -8592 -2920
rect -9764 -3032 -8676 -2968
rect -8612 -3032 -8592 -2968
rect -9764 -3048 -8592 -3032
rect -9764 -3112 -8676 -3048
rect -8612 -3112 -8592 -3048
rect -9764 -3128 -8592 -3112
rect -9764 -3192 -8676 -3128
rect -8612 -3192 -8592 -3128
rect -9764 -3208 -8592 -3192
rect -9764 -3272 -8676 -3208
rect -8612 -3272 -8592 -3208
rect -9764 -3288 -8592 -3272
rect -9764 -3352 -8676 -3288
rect -8612 -3352 -8592 -3288
rect -9764 -3368 -8592 -3352
rect -9764 -3432 -8676 -3368
rect -8612 -3432 -8592 -3368
rect -9764 -3448 -8592 -3432
rect -9764 -3512 -8676 -3448
rect -8612 -3512 -8592 -3448
rect -9764 -3528 -8592 -3512
rect -9764 -3592 -8676 -3528
rect -8612 -3592 -8592 -3528
rect -9764 -3608 -8592 -3592
rect -9764 -3672 -8676 -3608
rect -8612 -3672 -8592 -3608
rect -9764 -3688 -8592 -3672
rect -9764 -3752 -8676 -3688
rect -8612 -3752 -8592 -3688
rect -9764 -3800 -8592 -3752
rect -8352 -2968 -7180 -2920
rect -8352 -3032 -7264 -2968
rect -7200 -3032 -7180 -2968
rect -8352 -3048 -7180 -3032
rect -8352 -3112 -7264 -3048
rect -7200 -3112 -7180 -3048
rect -8352 -3128 -7180 -3112
rect -8352 -3192 -7264 -3128
rect -7200 -3192 -7180 -3128
rect -8352 -3208 -7180 -3192
rect -8352 -3272 -7264 -3208
rect -7200 -3272 -7180 -3208
rect -8352 -3288 -7180 -3272
rect -8352 -3352 -7264 -3288
rect -7200 -3352 -7180 -3288
rect -8352 -3368 -7180 -3352
rect -8352 -3432 -7264 -3368
rect -7200 -3432 -7180 -3368
rect -8352 -3448 -7180 -3432
rect -8352 -3512 -7264 -3448
rect -7200 -3512 -7180 -3448
rect -8352 -3528 -7180 -3512
rect -8352 -3592 -7264 -3528
rect -7200 -3592 -7180 -3528
rect -8352 -3608 -7180 -3592
rect -8352 -3672 -7264 -3608
rect -7200 -3672 -7180 -3608
rect -8352 -3688 -7180 -3672
rect -8352 -3752 -7264 -3688
rect -7200 -3752 -7180 -3688
rect -8352 -3800 -7180 -3752
rect -6940 -2968 -5768 -2920
rect -6940 -3032 -5852 -2968
rect -5788 -3032 -5768 -2968
rect -6940 -3048 -5768 -3032
rect -6940 -3112 -5852 -3048
rect -5788 -3112 -5768 -3048
rect -6940 -3128 -5768 -3112
rect -6940 -3192 -5852 -3128
rect -5788 -3192 -5768 -3128
rect -6940 -3208 -5768 -3192
rect -6940 -3272 -5852 -3208
rect -5788 -3272 -5768 -3208
rect -6940 -3288 -5768 -3272
rect -6940 -3352 -5852 -3288
rect -5788 -3352 -5768 -3288
rect -6940 -3368 -5768 -3352
rect -6940 -3432 -5852 -3368
rect -5788 -3432 -5768 -3368
rect -6940 -3448 -5768 -3432
rect -6940 -3512 -5852 -3448
rect -5788 -3512 -5768 -3448
rect -6940 -3528 -5768 -3512
rect -6940 -3592 -5852 -3528
rect -5788 -3592 -5768 -3528
rect -6940 -3608 -5768 -3592
rect -6940 -3672 -5852 -3608
rect -5788 -3672 -5768 -3608
rect -6940 -3688 -5768 -3672
rect -6940 -3752 -5852 -3688
rect -5788 -3752 -5768 -3688
rect -6940 -3800 -5768 -3752
rect -5528 -2968 -4356 -2920
rect -5528 -3032 -4440 -2968
rect -4376 -3032 -4356 -2968
rect -5528 -3048 -4356 -3032
rect -5528 -3112 -4440 -3048
rect -4376 -3112 -4356 -3048
rect -5528 -3128 -4356 -3112
rect -5528 -3192 -4440 -3128
rect -4376 -3192 -4356 -3128
rect -5528 -3208 -4356 -3192
rect -5528 -3272 -4440 -3208
rect -4376 -3272 -4356 -3208
rect -5528 -3288 -4356 -3272
rect -5528 -3352 -4440 -3288
rect -4376 -3352 -4356 -3288
rect -5528 -3368 -4356 -3352
rect -5528 -3432 -4440 -3368
rect -4376 -3432 -4356 -3368
rect -5528 -3448 -4356 -3432
rect -5528 -3512 -4440 -3448
rect -4376 -3512 -4356 -3448
rect -5528 -3528 -4356 -3512
rect -5528 -3592 -4440 -3528
rect -4376 -3592 -4356 -3528
rect -5528 -3608 -4356 -3592
rect -5528 -3672 -4440 -3608
rect -4376 -3672 -4356 -3608
rect -5528 -3688 -4356 -3672
rect -5528 -3752 -4440 -3688
rect -4376 -3752 -4356 -3688
rect -5528 -3800 -4356 -3752
rect -4116 -2968 -2944 -2920
rect -4116 -3032 -3028 -2968
rect -2964 -3032 -2944 -2968
rect -4116 -3048 -2944 -3032
rect -4116 -3112 -3028 -3048
rect -2964 -3112 -2944 -3048
rect -4116 -3128 -2944 -3112
rect -4116 -3192 -3028 -3128
rect -2964 -3192 -2944 -3128
rect -4116 -3208 -2944 -3192
rect -4116 -3272 -3028 -3208
rect -2964 -3272 -2944 -3208
rect -4116 -3288 -2944 -3272
rect -4116 -3352 -3028 -3288
rect -2964 -3352 -2944 -3288
rect -4116 -3368 -2944 -3352
rect -4116 -3432 -3028 -3368
rect -2964 -3432 -2944 -3368
rect -4116 -3448 -2944 -3432
rect -4116 -3512 -3028 -3448
rect -2964 -3512 -2944 -3448
rect -4116 -3528 -2944 -3512
rect -4116 -3592 -3028 -3528
rect -2964 -3592 -2944 -3528
rect -4116 -3608 -2944 -3592
rect -4116 -3672 -3028 -3608
rect -2964 -3672 -2944 -3608
rect -4116 -3688 -2944 -3672
rect -4116 -3752 -3028 -3688
rect -2964 -3752 -2944 -3688
rect -4116 -3800 -2944 -3752
rect -2704 -2968 -1532 -2920
rect -2704 -3032 -1616 -2968
rect -1552 -3032 -1532 -2968
rect -2704 -3048 -1532 -3032
rect -2704 -3112 -1616 -3048
rect -1552 -3112 -1532 -3048
rect -2704 -3128 -1532 -3112
rect -2704 -3192 -1616 -3128
rect -1552 -3192 -1532 -3128
rect -2704 -3208 -1532 -3192
rect -2704 -3272 -1616 -3208
rect -1552 -3272 -1532 -3208
rect -2704 -3288 -1532 -3272
rect -2704 -3352 -1616 -3288
rect -1552 -3352 -1532 -3288
rect -2704 -3368 -1532 -3352
rect -2704 -3432 -1616 -3368
rect -1552 -3432 -1532 -3368
rect -2704 -3448 -1532 -3432
rect -2704 -3512 -1616 -3448
rect -1552 -3512 -1532 -3448
rect -2704 -3528 -1532 -3512
rect -2704 -3592 -1616 -3528
rect -1552 -3592 -1532 -3528
rect -2704 -3608 -1532 -3592
rect -2704 -3672 -1616 -3608
rect -1552 -3672 -1532 -3608
rect -2704 -3688 -1532 -3672
rect -2704 -3752 -1616 -3688
rect -1552 -3752 -1532 -3688
rect -2704 -3800 -1532 -3752
rect -1292 -2968 -120 -2920
rect -1292 -3032 -204 -2968
rect -140 -3032 -120 -2968
rect -1292 -3048 -120 -3032
rect -1292 -3112 -204 -3048
rect -140 -3112 -120 -3048
rect -1292 -3128 -120 -3112
rect -1292 -3192 -204 -3128
rect -140 -3192 -120 -3128
rect -1292 -3208 -120 -3192
rect -1292 -3272 -204 -3208
rect -140 -3272 -120 -3208
rect -1292 -3288 -120 -3272
rect -1292 -3352 -204 -3288
rect -140 -3352 -120 -3288
rect -1292 -3368 -120 -3352
rect -1292 -3432 -204 -3368
rect -140 -3432 -120 -3368
rect -1292 -3448 -120 -3432
rect -1292 -3512 -204 -3448
rect -140 -3512 -120 -3448
rect -1292 -3528 -120 -3512
rect -1292 -3592 -204 -3528
rect -140 -3592 -120 -3528
rect -1292 -3608 -120 -3592
rect -1292 -3672 -204 -3608
rect -140 -3672 -120 -3608
rect -1292 -3688 -120 -3672
rect -1292 -3752 -204 -3688
rect -140 -3752 -120 -3688
rect -1292 -3800 -120 -3752
rect 120 -2968 1292 -2920
rect 120 -3032 1208 -2968
rect 1272 -3032 1292 -2968
rect 120 -3048 1292 -3032
rect 120 -3112 1208 -3048
rect 1272 -3112 1292 -3048
rect 120 -3128 1292 -3112
rect 120 -3192 1208 -3128
rect 1272 -3192 1292 -3128
rect 120 -3208 1292 -3192
rect 120 -3272 1208 -3208
rect 1272 -3272 1292 -3208
rect 120 -3288 1292 -3272
rect 120 -3352 1208 -3288
rect 1272 -3352 1292 -3288
rect 120 -3368 1292 -3352
rect 120 -3432 1208 -3368
rect 1272 -3432 1292 -3368
rect 120 -3448 1292 -3432
rect 120 -3512 1208 -3448
rect 1272 -3512 1292 -3448
rect 120 -3528 1292 -3512
rect 120 -3592 1208 -3528
rect 1272 -3592 1292 -3528
rect 120 -3608 1292 -3592
rect 120 -3672 1208 -3608
rect 1272 -3672 1292 -3608
rect 120 -3688 1292 -3672
rect 120 -3752 1208 -3688
rect 1272 -3752 1292 -3688
rect 120 -3800 1292 -3752
rect 1532 -2968 2704 -2920
rect 1532 -3032 2620 -2968
rect 2684 -3032 2704 -2968
rect 1532 -3048 2704 -3032
rect 1532 -3112 2620 -3048
rect 2684 -3112 2704 -3048
rect 1532 -3128 2704 -3112
rect 1532 -3192 2620 -3128
rect 2684 -3192 2704 -3128
rect 1532 -3208 2704 -3192
rect 1532 -3272 2620 -3208
rect 2684 -3272 2704 -3208
rect 1532 -3288 2704 -3272
rect 1532 -3352 2620 -3288
rect 2684 -3352 2704 -3288
rect 1532 -3368 2704 -3352
rect 1532 -3432 2620 -3368
rect 2684 -3432 2704 -3368
rect 1532 -3448 2704 -3432
rect 1532 -3512 2620 -3448
rect 2684 -3512 2704 -3448
rect 1532 -3528 2704 -3512
rect 1532 -3592 2620 -3528
rect 2684 -3592 2704 -3528
rect 1532 -3608 2704 -3592
rect 1532 -3672 2620 -3608
rect 2684 -3672 2704 -3608
rect 1532 -3688 2704 -3672
rect 1532 -3752 2620 -3688
rect 2684 -3752 2704 -3688
rect 1532 -3800 2704 -3752
rect 2944 -2968 4116 -2920
rect 2944 -3032 4032 -2968
rect 4096 -3032 4116 -2968
rect 2944 -3048 4116 -3032
rect 2944 -3112 4032 -3048
rect 4096 -3112 4116 -3048
rect 2944 -3128 4116 -3112
rect 2944 -3192 4032 -3128
rect 4096 -3192 4116 -3128
rect 2944 -3208 4116 -3192
rect 2944 -3272 4032 -3208
rect 4096 -3272 4116 -3208
rect 2944 -3288 4116 -3272
rect 2944 -3352 4032 -3288
rect 4096 -3352 4116 -3288
rect 2944 -3368 4116 -3352
rect 2944 -3432 4032 -3368
rect 4096 -3432 4116 -3368
rect 2944 -3448 4116 -3432
rect 2944 -3512 4032 -3448
rect 4096 -3512 4116 -3448
rect 2944 -3528 4116 -3512
rect 2944 -3592 4032 -3528
rect 4096 -3592 4116 -3528
rect 2944 -3608 4116 -3592
rect 2944 -3672 4032 -3608
rect 4096 -3672 4116 -3608
rect 2944 -3688 4116 -3672
rect 2944 -3752 4032 -3688
rect 4096 -3752 4116 -3688
rect 2944 -3800 4116 -3752
rect 4356 -2968 5528 -2920
rect 4356 -3032 5444 -2968
rect 5508 -3032 5528 -2968
rect 4356 -3048 5528 -3032
rect 4356 -3112 5444 -3048
rect 5508 -3112 5528 -3048
rect 4356 -3128 5528 -3112
rect 4356 -3192 5444 -3128
rect 5508 -3192 5528 -3128
rect 4356 -3208 5528 -3192
rect 4356 -3272 5444 -3208
rect 5508 -3272 5528 -3208
rect 4356 -3288 5528 -3272
rect 4356 -3352 5444 -3288
rect 5508 -3352 5528 -3288
rect 4356 -3368 5528 -3352
rect 4356 -3432 5444 -3368
rect 5508 -3432 5528 -3368
rect 4356 -3448 5528 -3432
rect 4356 -3512 5444 -3448
rect 5508 -3512 5528 -3448
rect 4356 -3528 5528 -3512
rect 4356 -3592 5444 -3528
rect 5508 -3592 5528 -3528
rect 4356 -3608 5528 -3592
rect 4356 -3672 5444 -3608
rect 5508 -3672 5528 -3608
rect 4356 -3688 5528 -3672
rect 4356 -3752 5444 -3688
rect 5508 -3752 5528 -3688
rect 4356 -3800 5528 -3752
rect 5768 -2968 6940 -2920
rect 5768 -3032 6856 -2968
rect 6920 -3032 6940 -2968
rect 5768 -3048 6940 -3032
rect 5768 -3112 6856 -3048
rect 6920 -3112 6940 -3048
rect 5768 -3128 6940 -3112
rect 5768 -3192 6856 -3128
rect 6920 -3192 6940 -3128
rect 5768 -3208 6940 -3192
rect 5768 -3272 6856 -3208
rect 6920 -3272 6940 -3208
rect 5768 -3288 6940 -3272
rect 5768 -3352 6856 -3288
rect 6920 -3352 6940 -3288
rect 5768 -3368 6940 -3352
rect 5768 -3432 6856 -3368
rect 6920 -3432 6940 -3368
rect 5768 -3448 6940 -3432
rect 5768 -3512 6856 -3448
rect 6920 -3512 6940 -3448
rect 5768 -3528 6940 -3512
rect 5768 -3592 6856 -3528
rect 6920 -3592 6940 -3528
rect 5768 -3608 6940 -3592
rect 5768 -3672 6856 -3608
rect 6920 -3672 6940 -3608
rect 5768 -3688 6940 -3672
rect 5768 -3752 6856 -3688
rect 6920 -3752 6940 -3688
rect 5768 -3800 6940 -3752
rect 7180 -2968 8352 -2920
rect 7180 -3032 8268 -2968
rect 8332 -3032 8352 -2968
rect 7180 -3048 8352 -3032
rect 7180 -3112 8268 -3048
rect 8332 -3112 8352 -3048
rect 7180 -3128 8352 -3112
rect 7180 -3192 8268 -3128
rect 8332 -3192 8352 -3128
rect 7180 -3208 8352 -3192
rect 7180 -3272 8268 -3208
rect 8332 -3272 8352 -3208
rect 7180 -3288 8352 -3272
rect 7180 -3352 8268 -3288
rect 8332 -3352 8352 -3288
rect 7180 -3368 8352 -3352
rect 7180 -3432 8268 -3368
rect 8332 -3432 8352 -3368
rect 7180 -3448 8352 -3432
rect 7180 -3512 8268 -3448
rect 8332 -3512 8352 -3448
rect 7180 -3528 8352 -3512
rect 7180 -3592 8268 -3528
rect 8332 -3592 8352 -3528
rect 7180 -3608 8352 -3592
rect 7180 -3672 8268 -3608
rect 8332 -3672 8352 -3608
rect 7180 -3688 8352 -3672
rect 7180 -3752 8268 -3688
rect 8332 -3752 8352 -3688
rect 7180 -3800 8352 -3752
rect 8592 -2968 9764 -2920
rect 8592 -3032 9680 -2968
rect 9744 -3032 9764 -2968
rect 8592 -3048 9764 -3032
rect 8592 -3112 9680 -3048
rect 9744 -3112 9764 -3048
rect 8592 -3128 9764 -3112
rect 8592 -3192 9680 -3128
rect 9744 -3192 9764 -3128
rect 8592 -3208 9764 -3192
rect 8592 -3272 9680 -3208
rect 9744 -3272 9764 -3208
rect 8592 -3288 9764 -3272
rect 8592 -3352 9680 -3288
rect 9744 -3352 9764 -3288
rect 8592 -3368 9764 -3352
rect 8592 -3432 9680 -3368
rect 9744 -3432 9764 -3368
rect 8592 -3448 9764 -3432
rect 8592 -3512 9680 -3448
rect 9744 -3512 9764 -3448
rect 8592 -3528 9764 -3512
rect 8592 -3592 9680 -3528
rect 9744 -3592 9764 -3528
rect 8592 -3608 9764 -3592
rect 8592 -3672 9680 -3608
rect 9744 -3672 9764 -3608
rect 8592 -3688 9764 -3672
rect 8592 -3752 9680 -3688
rect 9744 -3752 9764 -3688
rect 8592 -3800 9764 -3752
rect 10004 -2968 11176 -2920
rect 10004 -3032 11092 -2968
rect 11156 -3032 11176 -2968
rect 10004 -3048 11176 -3032
rect 10004 -3112 11092 -3048
rect 11156 -3112 11176 -3048
rect 10004 -3128 11176 -3112
rect 10004 -3192 11092 -3128
rect 11156 -3192 11176 -3128
rect 10004 -3208 11176 -3192
rect 10004 -3272 11092 -3208
rect 11156 -3272 11176 -3208
rect 10004 -3288 11176 -3272
rect 10004 -3352 11092 -3288
rect 11156 -3352 11176 -3288
rect 10004 -3368 11176 -3352
rect 10004 -3432 11092 -3368
rect 11156 -3432 11176 -3368
rect 10004 -3448 11176 -3432
rect 10004 -3512 11092 -3448
rect 11156 -3512 11176 -3448
rect 10004 -3528 11176 -3512
rect 10004 -3592 11092 -3528
rect 11156 -3592 11176 -3528
rect 10004 -3608 11176 -3592
rect 10004 -3672 11092 -3608
rect 11156 -3672 11176 -3608
rect 10004 -3688 11176 -3672
rect 10004 -3752 11092 -3688
rect 11156 -3752 11176 -3688
rect 10004 -3800 11176 -3752
rect 11416 -2968 12588 -2920
rect 11416 -3032 12504 -2968
rect 12568 -3032 12588 -2968
rect 11416 -3048 12588 -3032
rect 11416 -3112 12504 -3048
rect 12568 -3112 12588 -3048
rect 11416 -3128 12588 -3112
rect 11416 -3192 12504 -3128
rect 12568 -3192 12588 -3128
rect 11416 -3208 12588 -3192
rect 11416 -3272 12504 -3208
rect 12568 -3272 12588 -3208
rect 11416 -3288 12588 -3272
rect 11416 -3352 12504 -3288
rect 12568 -3352 12588 -3288
rect 11416 -3368 12588 -3352
rect 11416 -3432 12504 -3368
rect 12568 -3432 12588 -3368
rect 11416 -3448 12588 -3432
rect 11416 -3512 12504 -3448
rect 12568 -3512 12588 -3448
rect 11416 -3528 12588 -3512
rect 11416 -3592 12504 -3528
rect 12568 -3592 12588 -3528
rect 11416 -3608 12588 -3592
rect 11416 -3672 12504 -3608
rect 12568 -3672 12588 -3608
rect 11416 -3688 12588 -3672
rect 11416 -3752 12504 -3688
rect 12568 -3752 12588 -3688
rect 11416 -3800 12588 -3752
rect 12828 -2968 14000 -2920
rect 12828 -3032 13916 -2968
rect 13980 -3032 14000 -2968
rect 12828 -3048 14000 -3032
rect 12828 -3112 13916 -3048
rect 13980 -3112 14000 -3048
rect 12828 -3128 14000 -3112
rect 12828 -3192 13916 -3128
rect 13980 -3192 14000 -3128
rect 12828 -3208 14000 -3192
rect 12828 -3272 13916 -3208
rect 13980 -3272 14000 -3208
rect 12828 -3288 14000 -3272
rect 12828 -3352 13916 -3288
rect 13980 -3352 14000 -3288
rect 12828 -3368 14000 -3352
rect 12828 -3432 13916 -3368
rect 13980 -3432 14000 -3368
rect 12828 -3448 14000 -3432
rect 12828 -3512 13916 -3448
rect 13980 -3512 14000 -3448
rect 12828 -3528 14000 -3512
rect 12828 -3592 13916 -3528
rect 13980 -3592 14000 -3528
rect 12828 -3608 14000 -3592
rect 12828 -3672 13916 -3608
rect 13980 -3672 14000 -3608
rect 12828 -3688 14000 -3672
rect 12828 -3752 13916 -3688
rect 13980 -3752 14000 -3688
rect 12828 -3800 14000 -3752
rect 14240 -2968 15412 -2920
rect 14240 -3032 15328 -2968
rect 15392 -3032 15412 -2968
rect 14240 -3048 15412 -3032
rect 14240 -3112 15328 -3048
rect 15392 -3112 15412 -3048
rect 14240 -3128 15412 -3112
rect 14240 -3192 15328 -3128
rect 15392 -3192 15412 -3128
rect 14240 -3208 15412 -3192
rect 14240 -3272 15328 -3208
rect 15392 -3272 15412 -3208
rect 14240 -3288 15412 -3272
rect 14240 -3352 15328 -3288
rect 15392 -3352 15412 -3288
rect 14240 -3368 15412 -3352
rect 14240 -3432 15328 -3368
rect 15392 -3432 15412 -3368
rect 14240 -3448 15412 -3432
rect 14240 -3512 15328 -3448
rect 15392 -3512 15412 -3448
rect 14240 -3528 15412 -3512
rect 14240 -3592 15328 -3528
rect 15392 -3592 15412 -3528
rect 14240 -3608 15412 -3592
rect 14240 -3672 15328 -3608
rect 15392 -3672 15412 -3608
rect 14240 -3688 15412 -3672
rect 14240 -3752 15328 -3688
rect 15392 -3752 15412 -3688
rect 14240 -3800 15412 -3752
rect 15652 -2968 16824 -2920
rect 15652 -3032 16740 -2968
rect 16804 -3032 16824 -2968
rect 15652 -3048 16824 -3032
rect 15652 -3112 16740 -3048
rect 16804 -3112 16824 -3048
rect 15652 -3128 16824 -3112
rect 15652 -3192 16740 -3128
rect 16804 -3192 16824 -3128
rect 15652 -3208 16824 -3192
rect 15652 -3272 16740 -3208
rect 16804 -3272 16824 -3208
rect 15652 -3288 16824 -3272
rect 15652 -3352 16740 -3288
rect 16804 -3352 16824 -3288
rect 15652 -3368 16824 -3352
rect 15652 -3432 16740 -3368
rect 16804 -3432 16824 -3368
rect 15652 -3448 16824 -3432
rect 15652 -3512 16740 -3448
rect 16804 -3512 16824 -3448
rect 15652 -3528 16824 -3512
rect 15652 -3592 16740 -3528
rect 16804 -3592 16824 -3528
rect 15652 -3608 16824 -3592
rect 15652 -3672 16740 -3608
rect 16804 -3672 16824 -3608
rect 15652 -3688 16824 -3672
rect 15652 -3752 16740 -3688
rect 16804 -3752 16824 -3688
rect 15652 -3800 16824 -3752
rect 17064 -2968 18236 -2920
rect 17064 -3032 18152 -2968
rect 18216 -3032 18236 -2968
rect 17064 -3048 18236 -3032
rect 17064 -3112 18152 -3048
rect 18216 -3112 18236 -3048
rect 17064 -3128 18236 -3112
rect 17064 -3192 18152 -3128
rect 18216 -3192 18236 -3128
rect 17064 -3208 18236 -3192
rect 17064 -3272 18152 -3208
rect 18216 -3272 18236 -3208
rect 17064 -3288 18236 -3272
rect 17064 -3352 18152 -3288
rect 18216 -3352 18236 -3288
rect 17064 -3368 18236 -3352
rect 17064 -3432 18152 -3368
rect 18216 -3432 18236 -3368
rect 17064 -3448 18236 -3432
rect 17064 -3512 18152 -3448
rect 18216 -3512 18236 -3448
rect 17064 -3528 18236 -3512
rect 17064 -3592 18152 -3528
rect 18216 -3592 18236 -3528
rect 17064 -3608 18236 -3592
rect 17064 -3672 18152 -3608
rect 18216 -3672 18236 -3608
rect 17064 -3688 18236 -3672
rect 17064 -3752 18152 -3688
rect 18216 -3752 18236 -3688
rect 17064 -3800 18236 -3752
rect 18476 -2968 19648 -2920
rect 18476 -3032 19564 -2968
rect 19628 -3032 19648 -2968
rect 18476 -3048 19648 -3032
rect 18476 -3112 19564 -3048
rect 19628 -3112 19648 -3048
rect 18476 -3128 19648 -3112
rect 18476 -3192 19564 -3128
rect 19628 -3192 19648 -3128
rect 18476 -3208 19648 -3192
rect 18476 -3272 19564 -3208
rect 19628 -3272 19648 -3208
rect 18476 -3288 19648 -3272
rect 18476 -3352 19564 -3288
rect 19628 -3352 19648 -3288
rect 18476 -3368 19648 -3352
rect 18476 -3432 19564 -3368
rect 19628 -3432 19648 -3368
rect 18476 -3448 19648 -3432
rect 18476 -3512 19564 -3448
rect 19628 -3512 19648 -3448
rect 18476 -3528 19648 -3512
rect 18476 -3592 19564 -3528
rect 19628 -3592 19648 -3528
rect 18476 -3608 19648 -3592
rect 18476 -3672 19564 -3608
rect 19628 -3672 19648 -3608
rect 18476 -3688 19648 -3672
rect 18476 -3752 19564 -3688
rect 19628 -3752 19648 -3688
rect 18476 -3800 19648 -3752
rect 19888 -2968 21060 -2920
rect 19888 -3032 20976 -2968
rect 21040 -3032 21060 -2968
rect 19888 -3048 21060 -3032
rect 19888 -3112 20976 -3048
rect 21040 -3112 21060 -3048
rect 19888 -3128 21060 -3112
rect 19888 -3192 20976 -3128
rect 21040 -3192 21060 -3128
rect 19888 -3208 21060 -3192
rect 19888 -3272 20976 -3208
rect 21040 -3272 21060 -3208
rect 19888 -3288 21060 -3272
rect 19888 -3352 20976 -3288
rect 21040 -3352 21060 -3288
rect 19888 -3368 21060 -3352
rect 19888 -3432 20976 -3368
rect 21040 -3432 21060 -3368
rect 19888 -3448 21060 -3432
rect 19888 -3512 20976 -3448
rect 21040 -3512 21060 -3448
rect 19888 -3528 21060 -3512
rect 19888 -3592 20976 -3528
rect 21040 -3592 21060 -3528
rect 19888 -3608 21060 -3592
rect 19888 -3672 20976 -3608
rect 21040 -3672 21060 -3608
rect 19888 -3688 21060 -3672
rect 19888 -3752 20976 -3688
rect 21040 -3752 21060 -3688
rect 19888 -3800 21060 -3752
rect 21300 -2968 22472 -2920
rect 21300 -3032 22388 -2968
rect 22452 -3032 22472 -2968
rect 21300 -3048 22472 -3032
rect 21300 -3112 22388 -3048
rect 22452 -3112 22472 -3048
rect 21300 -3128 22472 -3112
rect 21300 -3192 22388 -3128
rect 22452 -3192 22472 -3128
rect 21300 -3208 22472 -3192
rect 21300 -3272 22388 -3208
rect 22452 -3272 22472 -3208
rect 21300 -3288 22472 -3272
rect 21300 -3352 22388 -3288
rect 22452 -3352 22472 -3288
rect 21300 -3368 22472 -3352
rect 21300 -3432 22388 -3368
rect 22452 -3432 22472 -3368
rect 21300 -3448 22472 -3432
rect 21300 -3512 22388 -3448
rect 22452 -3512 22472 -3448
rect 21300 -3528 22472 -3512
rect 21300 -3592 22388 -3528
rect 22452 -3592 22472 -3528
rect 21300 -3608 22472 -3592
rect 21300 -3672 22388 -3608
rect 22452 -3672 22472 -3608
rect 21300 -3688 22472 -3672
rect 21300 -3752 22388 -3688
rect 22452 -3752 22472 -3688
rect 21300 -3800 22472 -3752
rect 22712 -2968 23884 -2920
rect 22712 -3032 23800 -2968
rect 23864 -3032 23884 -2968
rect 22712 -3048 23884 -3032
rect 22712 -3112 23800 -3048
rect 23864 -3112 23884 -3048
rect 22712 -3128 23884 -3112
rect 22712 -3192 23800 -3128
rect 23864 -3192 23884 -3128
rect 22712 -3208 23884 -3192
rect 22712 -3272 23800 -3208
rect 23864 -3272 23884 -3208
rect 22712 -3288 23884 -3272
rect 22712 -3352 23800 -3288
rect 23864 -3352 23884 -3288
rect 22712 -3368 23884 -3352
rect 22712 -3432 23800 -3368
rect 23864 -3432 23884 -3368
rect 22712 -3448 23884 -3432
rect 22712 -3512 23800 -3448
rect 23864 -3512 23884 -3448
rect 22712 -3528 23884 -3512
rect 22712 -3592 23800 -3528
rect 23864 -3592 23884 -3528
rect 22712 -3608 23884 -3592
rect 22712 -3672 23800 -3608
rect 23864 -3672 23884 -3608
rect 22712 -3688 23884 -3672
rect 22712 -3752 23800 -3688
rect 23864 -3752 23884 -3688
rect 22712 -3800 23884 -3752
rect -23884 -4088 -22712 -4040
rect -23884 -4152 -22796 -4088
rect -22732 -4152 -22712 -4088
rect -23884 -4168 -22712 -4152
rect -23884 -4232 -22796 -4168
rect -22732 -4232 -22712 -4168
rect -23884 -4248 -22712 -4232
rect -23884 -4312 -22796 -4248
rect -22732 -4312 -22712 -4248
rect -23884 -4328 -22712 -4312
rect -23884 -4392 -22796 -4328
rect -22732 -4392 -22712 -4328
rect -23884 -4408 -22712 -4392
rect -23884 -4472 -22796 -4408
rect -22732 -4472 -22712 -4408
rect -23884 -4488 -22712 -4472
rect -23884 -4552 -22796 -4488
rect -22732 -4552 -22712 -4488
rect -23884 -4568 -22712 -4552
rect -23884 -4632 -22796 -4568
rect -22732 -4632 -22712 -4568
rect -23884 -4648 -22712 -4632
rect -23884 -4712 -22796 -4648
rect -22732 -4712 -22712 -4648
rect -23884 -4728 -22712 -4712
rect -23884 -4792 -22796 -4728
rect -22732 -4792 -22712 -4728
rect -23884 -4808 -22712 -4792
rect -23884 -4872 -22796 -4808
rect -22732 -4872 -22712 -4808
rect -23884 -4920 -22712 -4872
rect -22472 -4088 -21300 -4040
rect -22472 -4152 -21384 -4088
rect -21320 -4152 -21300 -4088
rect -22472 -4168 -21300 -4152
rect -22472 -4232 -21384 -4168
rect -21320 -4232 -21300 -4168
rect -22472 -4248 -21300 -4232
rect -22472 -4312 -21384 -4248
rect -21320 -4312 -21300 -4248
rect -22472 -4328 -21300 -4312
rect -22472 -4392 -21384 -4328
rect -21320 -4392 -21300 -4328
rect -22472 -4408 -21300 -4392
rect -22472 -4472 -21384 -4408
rect -21320 -4472 -21300 -4408
rect -22472 -4488 -21300 -4472
rect -22472 -4552 -21384 -4488
rect -21320 -4552 -21300 -4488
rect -22472 -4568 -21300 -4552
rect -22472 -4632 -21384 -4568
rect -21320 -4632 -21300 -4568
rect -22472 -4648 -21300 -4632
rect -22472 -4712 -21384 -4648
rect -21320 -4712 -21300 -4648
rect -22472 -4728 -21300 -4712
rect -22472 -4792 -21384 -4728
rect -21320 -4792 -21300 -4728
rect -22472 -4808 -21300 -4792
rect -22472 -4872 -21384 -4808
rect -21320 -4872 -21300 -4808
rect -22472 -4920 -21300 -4872
rect -21060 -4088 -19888 -4040
rect -21060 -4152 -19972 -4088
rect -19908 -4152 -19888 -4088
rect -21060 -4168 -19888 -4152
rect -21060 -4232 -19972 -4168
rect -19908 -4232 -19888 -4168
rect -21060 -4248 -19888 -4232
rect -21060 -4312 -19972 -4248
rect -19908 -4312 -19888 -4248
rect -21060 -4328 -19888 -4312
rect -21060 -4392 -19972 -4328
rect -19908 -4392 -19888 -4328
rect -21060 -4408 -19888 -4392
rect -21060 -4472 -19972 -4408
rect -19908 -4472 -19888 -4408
rect -21060 -4488 -19888 -4472
rect -21060 -4552 -19972 -4488
rect -19908 -4552 -19888 -4488
rect -21060 -4568 -19888 -4552
rect -21060 -4632 -19972 -4568
rect -19908 -4632 -19888 -4568
rect -21060 -4648 -19888 -4632
rect -21060 -4712 -19972 -4648
rect -19908 -4712 -19888 -4648
rect -21060 -4728 -19888 -4712
rect -21060 -4792 -19972 -4728
rect -19908 -4792 -19888 -4728
rect -21060 -4808 -19888 -4792
rect -21060 -4872 -19972 -4808
rect -19908 -4872 -19888 -4808
rect -21060 -4920 -19888 -4872
rect -19648 -4088 -18476 -4040
rect -19648 -4152 -18560 -4088
rect -18496 -4152 -18476 -4088
rect -19648 -4168 -18476 -4152
rect -19648 -4232 -18560 -4168
rect -18496 -4232 -18476 -4168
rect -19648 -4248 -18476 -4232
rect -19648 -4312 -18560 -4248
rect -18496 -4312 -18476 -4248
rect -19648 -4328 -18476 -4312
rect -19648 -4392 -18560 -4328
rect -18496 -4392 -18476 -4328
rect -19648 -4408 -18476 -4392
rect -19648 -4472 -18560 -4408
rect -18496 -4472 -18476 -4408
rect -19648 -4488 -18476 -4472
rect -19648 -4552 -18560 -4488
rect -18496 -4552 -18476 -4488
rect -19648 -4568 -18476 -4552
rect -19648 -4632 -18560 -4568
rect -18496 -4632 -18476 -4568
rect -19648 -4648 -18476 -4632
rect -19648 -4712 -18560 -4648
rect -18496 -4712 -18476 -4648
rect -19648 -4728 -18476 -4712
rect -19648 -4792 -18560 -4728
rect -18496 -4792 -18476 -4728
rect -19648 -4808 -18476 -4792
rect -19648 -4872 -18560 -4808
rect -18496 -4872 -18476 -4808
rect -19648 -4920 -18476 -4872
rect -18236 -4088 -17064 -4040
rect -18236 -4152 -17148 -4088
rect -17084 -4152 -17064 -4088
rect -18236 -4168 -17064 -4152
rect -18236 -4232 -17148 -4168
rect -17084 -4232 -17064 -4168
rect -18236 -4248 -17064 -4232
rect -18236 -4312 -17148 -4248
rect -17084 -4312 -17064 -4248
rect -18236 -4328 -17064 -4312
rect -18236 -4392 -17148 -4328
rect -17084 -4392 -17064 -4328
rect -18236 -4408 -17064 -4392
rect -18236 -4472 -17148 -4408
rect -17084 -4472 -17064 -4408
rect -18236 -4488 -17064 -4472
rect -18236 -4552 -17148 -4488
rect -17084 -4552 -17064 -4488
rect -18236 -4568 -17064 -4552
rect -18236 -4632 -17148 -4568
rect -17084 -4632 -17064 -4568
rect -18236 -4648 -17064 -4632
rect -18236 -4712 -17148 -4648
rect -17084 -4712 -17064 -4648
rect -18236 -4728 -17064 -4712
rect -18236 -4792 -17148 -4728
rect -17084 -4792 -17064 -4728
rect -18236 -4808 -17064 -4792
rect -18236 -4872 -17148 -4808
rect -17084 -4872 -17064 -4808
rect -18236 -4920 -17064 -4872
rect -16824 -4088 -15652 -4040
rect -16824 -4152 -15736 -4088
rect -15672 -4152 -15652 -4088
rect -16824 -4168 -15652 -4152
rect -16824 -4232 -15736 -4168
rect -15672 -4232 -15652 -4168
rect -16824 -4248 -15652 -4232
rect -16824 -4312 -15736 -4248
rect -15672 -4312 -15652 -4248
rect -16824 -4328 -15652 -4312
rect -16824 -4392 -15736 -4328
rect -15672 -4392 -15652 -4328
rect -16824 -4408 -15652 -4392
rect -16824 -4472 -15736 -4408
rect -15672 -4472 -15652 -4408
rect -16824 -4488 -15652 -4472
rect -16824 -4552 -15736 -4488
rect -15672 -4552 -15652 -4488
rect -16824 -4568 -15652 -4552
rect -16824 -4632 -15736 -4568
rect -15672 -4632 -15652 -4568
rect -16824 -4648 -15652 -4632
rect -16824 -4712 -15736 -4648
rect -15672 -4712 -15652 -4648
rect -16824 -4728 -15652 -4712
rect -16824 -4792 -15736 -4728
rect -15672 -4792 -15652 -4728
rect -16824 -4808 -15652 -4792
rect -16824 -4872 -15736 -4808
rect -15672 -4872 -15652 -4808
rect -16824 -4920 -15652 -4872
rect -15412 -4088 -14240 -4040
rect -15412 -4152 -14324 -4088
rect -14260 -4152 -14240 -4088
rect -15412 -4168 -14240 -4152
rect -15412 -4232 -14324 -4168
rect -14260 -4232 -14240 -4168
rect -15412 -4248 -14240 -4232
rect -15412 -4312 -14324 -4248
rect -14260 -4312 -14240 -4248
rect -15412 -4328 -14240 -4312
rect -15412 -4392 -14324 -4328
rect -14260 -4392 -14240 -4328
rect -15412 -4408 -14240 -4392
rect -15412 -4472 -14324 -4408
rect -14260 -4472 -14240 -4408
rect -15412 -4488 -14240 -4472
rect -15412 -4552 -14324 -4488
rect -14260 -4552 -14240 -4488
rect -15412 -4568 -14240 -4552
rect -15412 -4632 -14324 -4568
rect -14260 -4632 -14240 -4568
rect -15412 -4648 -14240 -4632
rect -15412 -4712 -14324 -4648
rect -14260 -4712 -14240 -4648
rect -15412 -4728 -14240 -4712
rect -15412 -4792 -14324 -4728
rect -14260 -4792 -14240 -4728
rect -15412 -4808 -14240 -4792
rect -15412 -4872 -14324 -4808
rect -14260 -4872 -14240 -4808
rect -15412 -4920 -14240 -4872
rect -14000 -4088 -12828 -4040
rect -14000 -4152 -12912 -4088
rect -12848 -4152 -12828 -4088
rect -14000 -4168 -12828 -4152
rect -14000 -4232 -12912 -4168
rect -12848 -4232 -12828 -4168
rect -14000 -4248 -12828 -4232
rect -14000 -4312 -12912 -4248
rect -12848 -4312 -12828 -4248
rect -14000 -4328 -12828 -4312
rect -14000 -4392 -12912 -4328
rect -12848 -4392 -12828 -4328
rect -14000 -4408 -12828 -4392
rect -14000 -4472 -12912 -4408
rect -12848 -4472 -12828 -4408
rect -14000 -4488 -12828 -4472
rect -14000 -4552 -12912 -4488
rect -12848 -4552 -12828 -4488
rect -14000 -4568 -12828 -4552
rect -14000 -4632 -12912 -4568
rect -12848 -4632 -12828 -4568
rect -14000 -4648 -12828 -4632
rect -14000 -4712 -12912 -4648
rect -12848 -4712 -12828 -4648
rect -14000 -4728 -12828 -4712
rect -14000 -4792 -12912 -4728
rect -12848 -4792 -12828 -4728
rect -14000 -4808 -12828 -4792
rect -14000 -4872 -12912 -4808
rect -12848 -4872 -12828 -4808
rect -14000 -4920 -12828 -4872
rect -12588 -4088 -11416 -4040
rect -12588 -4152 -11500 -4088
rect -11436 -4152 -11416 -4088
rect -12588 -4168 -11416 -4152
rect -12588 -4232 -11500 -4168
rect -11436 -4232 -11416 -4168
rect -12588 -4248 -11416 -4232
rect -12588 -4312 -11500 -4248
rect -11436 -4312 -11416 -4248
rect -12588 -4328 -11416 -4312
rect -12588 -4392 -11500 -4328
rect -11436 -4392 -11416 -4328
rect -12588 -4408 -11416 -4392
rect -12588 -4472 -11500 -4408
rect -11436 -4472 -11416 -4408
rect -12588 -4488 -11416 -4472
rect -12588 -4552 -11500 -4488
rect -11436 -4552 -11416 -4488
rect -12588 -4568 -11416 -4552
rect -12588 -4632 -11500 -4568
rect -11436 -4632 -11416 -4568
rect -12588 -4648 -11416 -4632
rect -12588 -4712 -11500 -4648
rect -11436 -4712 -11416 -4648
rect -12588 -4728 -11416 -4712
rect -12588 -4792 -11500 -4728
rect -11436 -4792 -11416 -4728
rect -12588 -4808 -11416 -4792
rect -12588 -4872 -11500 -4808
rect -11436 -4872 -11416 -4808
rect -12588 -4920 -11416 -4872
rect -11176 -4088 -10004 -4040
rect -11176 -4152 -10088 -4088
rect -10024 -4152 -10004 -4088
rect -11176 -4168 -10004 -4152
rect -11176 -4232 -10088 -4168
rect -10024 -4232 -10004 -4168
rect -11176 -4248 -10004 -4232
rect -11176 -4312 -10088 -4248
rect -10024 -4312 -10004 -4248
rect -11176 -4328 -10004 -4312
rect -11176 -4392 -10088 -4328
rect -10024 -4392 -10004 -4328
rect -11176 -4408 -10004 -4392
rect -11176 -4472 -10088 -4408
rect -10024 -4472 -10004 -4408
rect -11176 -4488 -10004 -4472
rect -11176 -4552 -10088 -4488
rect -10024 -4552 -10004 -4488
rect -11176 -4568 -10004 -4552
rect -11176 -4632 -10088 -4568
rect -10024 -4632 -10004 -4568
rect -11176 -4648 -10004 -4632
rect -11176 -4712 -10088 -4648
rect -10024 -4712 -10004 -4648
rect -11176 -4728 -10004 -4712
rect -11176 -4792 -10088 -4728
rect -10024 -4792 -10004 -4728
rect -11176 -4808 -10004 -4792
rect -11176 -4872 -10088 -4808
rect -10024 -4872 -10004 -4808
rect -11176 -4920 -10004 -4872
rect -9764 -4088 -8592 -4040
rect -9764 -4152 -8676 -4088
rect -8612 -4152 -8592 -4088
rect -9764 -4168 -8592 -4152
rect -9764 -4232 -8676 -4168
rect -8612 -4232 -8592 -4168
rect -9764 -4248 -8592 -4232
rect -9764 -4312 -8676 -4248
rect -8612 -4312 -8592 -4248
rect -9764 -4328 -8592 -4312
rect -9764 -4392 -8676 -4328
rect -8612 -4392 -8592 -4328
rect -9764 -4408 -8592 -4392
rect -9764 -4472 -8676 -4408
rect -8612 -4472 -8592 -4408
rect -9764 -4488 -8592 -4472
rect -9764 -4552 -8676 -4488
rect -8612 -4552 -8592 -4488
rect -9764 -4568 -8592 -4552
rect -9764 -4632 -8676 -4568
rect -8612 -4632 -8592 -4568
rect -9764 -4648 -8592 -4632
rect -9764 -4712 -8676 -4648
rect -8612 -4712 -8592 -4648
rect -9764 -4728 -8592 -4712
rect -9764 -4792 -8676 -4728
rect -8612 -4792 -8592 -4728
rect -9764 -4808 -8592 -4792
rect -9764 -4872 -8676 -4808
rect -8612 -4872 -8592 -4808
rect -9764 -4920 -8592 -4872
rect -8352 -4088 -7180 -4040
rect -8352 -4152 -7264 -4088
rect -7200 -4152 -7180 -4088
rect -8352 -4168 -7180 -4152
rect -8352 -4232 -7264 -4168
rect -7200 -4232 -7180 -4168
rect -8352 -4248 -7180 -4232
rect -8352 -4312 -7264 -4248
rect -7200 -4312 -7180 -4248
rect -8352 -4328 -7180 -4312
rect -8352 -4392 -7264 -4328
rect -7200 -4392 -7180 -4328
rect -8352 -4408 -7180 -4392
rect -8352 -4472 -7264 -4408
rect -7200 -4472 -7180 -4408
rect -8352 -4488 -7180 -4472
rect -8352 -4552 -7264 -4488
rect -7200 -4552 -7180 -4488
rect -8352 -4568 -7180 -4552
rect -8352 -4632 -7264 -4568
rect -7200 -4632 -7180 -4568
rect -8352 -4648 -7180 -4632
rect -8352 -4712 -7264 -4648
rect -7200 -4712 -7180 -4648
rect -8352 -4728 -7180 -4712
rect -8352 -4792 -7264 -4728
rect -7200 -4792 -7180 -4728
rect -8352 -4808 -7180 -4792
rect -8352 -4872 -7264 -4808
rect -7200 -4872 -7180 -4808
rect -8352 -4920 -7180 -4872
rect -6940 -4088 -5768 -4040
rect -6940 -4152 -5852 -4088
rect -5788 -4152 -5768 -4088
rect -6940 -4168 -5768 -4152
rect -6940 -4232 -5852 -4168
rect -5788 -4232 -5768 -4168
rect -6940 -4248 -5768 -4232
rect -6940 -4312 -5852 -4248
rect -5788 -4312 -5768 -4248
rect -6940 -4328 -5768 -4312
rect -6940 -4392 -5852 -4328
rect -5788 -4392 -5768 -4328
rect -6940 -4408 -5768 -4392
rect -6940 -4472 -5852 -4408
rect -5788 -4472 -5768 -4408
rect -6940 -4488 -5768 -4472
rect -6940 -4552 -5852 -4488
rect -5788 -4552 -5768 -4488
rect -6940 -4568 -5768 -4552
rect -6940 -4632 -5852 -4568
rect -5788 -4632 -5768 -4568
rect -6940 -4648 -5768 -4632
rect -6940 -4712 -5852 -4648
rect -5788 -4712 -5768 -4648
rect -6940 -4728 -5768 -4712
rect -6940 -4792 -5852 -4728
rect -5788 -4792 -5768 -4728
rect -6940 -4808 -5768 -4792
rect -6940 -4872 -5852 -4808
rect -5788 -4872 -5768 -4808
rect -6940 -4920 -5768 -4872
rect -5528 -4088 -4356 -4040
rect -5528 -4152 -4440 -4088
rect -4376 -4152 -4356 -4088
rect -5528 -4168 -4356 -4152
rect -5528 -4232 -4440 -4168
rect -4376 -4232 -4356 -4168
rect -5528 -4248 -4356 -4232
rect -5528 -4312 -4440 -4248
rect -4376 -4312 -4356 -4248
rect -5528 -4328 -4356 -4312
rect -5528 -4392 -4440 -4328
rect -4376 -4392 -4356 -4328
rect -5528 -4408 -4356 -4392
rect -5528 -4472 -4440 -4408
rect -4376 -4472 -4356 -4408
rect -5528 -4488 -4356 -4472
rect -5528 -4552 -4440 -4488
rect -4376 -4552 -4356 -4488
rect -5528 -4568 -4356 -4552
rect -5528 -4632 -4440 -4568
rect -4376 -4632 -4356 -4568
rect -5528 -4648 -4356 -4632
rect -5528 -4712 -4440 -4648
rect -4376 -4712 -4356 -4648
rect -5528 -4728 -4356 -4712
rect -5528 -4792 -4440 -4728
rect -4376 -4792 -4356 -4728
rect -5528 -4808 -4356 -4792
rect -5528 -4872 -4440 -4808
rect -4376 -4872 -4356 -4808
rect -5528 -4920 -4356 -4872
rect -4116 -4088 -2944 -4040
rect -4116 -4152 -3028 -4088
rect -2964 -4152 -2944 -4088
rect -4116 -4168 -2944 -4152
rect -4116 -4232 -3028 -4168
rect -2964 -4232 -2944 -4168
rect -4116 -4248 -2944 -4232
rect -4116 -4312 -3028 -4248
rect -2964 -4312 -2944 -4248
rect -4116 -4328 -2944 -4312
rect -4116 -4392 -3028 -4328
rect -2964 -4392 -2944 -4328
rect -4116 -4408 -2944 -4392
rect -4116 -4472 -3028 -4408
rect -2964 -4472 -2944 -4408
rect -4116 -4488 -2944 -4472
rect -4116 -4552 -3028 -4488
rect -2964 -4552 -2944 -4488
rect -4116 -4568 -2944 -4552
rect -4116 -4632 -3028 -4568
rect -2964 -4632 -2944 -4568
rect -4116 -4648 -2944 -4632
rect -4116 -4712 -3028 -4648
rect -2964 -4712 -2944 -4648
rect -4116 -4728 -2944 -4712
rect -4116 -4792 -3028 -4728
rect -2964 -4792 -2944 -4728
rect -4116 -4808 -2944 -4792
rect -4116 -4872 -3028 -4808
rect -2964 -4872 -2944 -4808
rect -4116 -4920 -2944 -4872
rect -2704 -4088 -1532 -4040
rect -2704 -4152 -1616 -4088
rect -1552 -4152 -1532 -4088
rect -2704 -4168 -1532 -4152
rect -2704 -4232 -1616 -4168
rect -1552 -4232 -1532 -4168
rect -2704 -4248 -1532 -4232
rect -2704 -4312 -1616 -4248
rect -1552 -4312 -1532 -4248
rect -2704 -4328 -1532 -4312
rect -2704 -4392 -1616 -4328
rect -1552 -4392 -1532 -4328
rect -2704 -4408 -1532 -4392
rect -2704 -4472 -1616 -4408
rect -1552 -4472 -1532 -4408
rect -2704 -4488 -1532 -4472
rect -2704 -4552 -1616 -4488
rect -1552 -4552 -1532 -4488
rect -2704 -4568 -1532 -4552
rect -2704 -4632 -1616 -4568
rect -1552 -4632 -1532 -4568
rect -2704 -4648 -1532 -4632
rect -2704 -4712 -1616 -4648
rect -1552 -4712 -1532 -4648
rect -2704 -4728 -1532 -4712
rect -2704 -4792 -1616 -4728
rect -1552 -4792 -1532 -4728
rect -2704 -4808 -1532 -4792
rect -2704 -4872 -1616 -4808
rect -1552 -4872 -1532 -4808
rect -2704 -4920 -1532 -4872
rect -1292 -4088 -120 -4040
rect -1292 -4152 -204 -4088
rect -140 -4152 -120 -4088
rect -1292 -4168 -120 -4152
rect -1292 -4232 -204 -4168
rect -140 -4232 -120 -4168
rect -1292 -4248 -120 -4232
rect -1292 -4312 -204 -4248
rect -140 -4312 -120 -4248
rect -1292 -4328 -120 -4312
rect -1292 -4392 -204 -4328
rect -140 -4392 -120 -4328
rect -1292 -4408 -120 -4392
rect -1292 -4472 -204 -4408
rect -140 -4472 -120 -4408
rect -1292 -4488 -120 -4472
rect -1292 -4552 -204 -4488
rect -140 -4552 -120 -4488
rect -1292 -4568 -120 -4552
rect -1292 -4632 -204 -4568
rect -140 -4632 -120 -4568
rect -1292 -4648 -120 -4632
rect -1292 -4712 -204 -4648
rect -140 -4712 -120 -4648
rect -1292 -4728 -120 -4712
rect -1292 -4792 -204 -4728
rect -140 -4792 -120 -4728
rect -1292 -4808 -120 -4792
rect -1292 -4872 -204 -4808
rect -140 -4872 -120 -4808
rect -1292 -4920 -120 -4872
rect 120 -4088 1292 -4040
rect 120 -4152 1208 -4088
rect 1272 -4152 1292 -4088
rect 120 -4168 1292 -4152
rect 120 -4232 1208 -4168
rect 1272 -4232 1292 -4168
rect 120 -4248 1292 -4232
rect 120 -4312 1208 -4248
rect 1272 -4312 1292 -4248
rect 120 -4328 1292 -4312
rect 120 -4392 1208 -4328
rect 1272 -4392 1292 -4328
rect 120 -4408 1292 -4392
rect 120 -4472 1208 -4408
rect 1272 -4472 1292 -4408
rect 120 -4488 1292 -4472
rect 120 -4552 1208 -4488
rect 1272 -4552 1292 -4488
rect 120 -4568 1292 -4552
rect 120 -4632 1208 -4568
rect 1272 -4632 1292 -4568
rect 120 -4648 1292 -4632
rect 120 -4712 1208 -4648
rect 1272 -4712 1292 -4648
rect 120 -4728 1292 -4712
rect 120 -4792 1208 -4728
rect 1272 -4792 1292 -4728
rect 120 -4808 1292 -4792
rect 120 -4872 1208 -4808
rect 1272 -4872 1292 -4808
rect 120 -4920 1292 -4872
rect 1532 -4088 2704 -4040
rect 1532 -4152 2620 -4088
rect 2684 -4152 2704 -4088
rect 1532 -4168 2704 -4152
rect 1532 -4232 2620 -4168
rect 2684 -4232 2704 -4168
rect 1532 -4248 2704 -4232
rect 1532 -4312 2620 -4248
rect 2684 -4312 2704 -4248
rect 1532 -4328 2704 -4312
rect 1532 -4392 2620 -4328
rect 2684 -4392 2704 -4328
rect 1532 -4408 2704 -4392
rect 1532 -4472 2620 -4408
rect 2684 -4472 2704 -4408
rect 1532 -4488 2704 -4472
rect 1532 -4552 2620 -4488
rect 2684 -4552 2704 -4488
rect 1532 -4568 2704 -4552
rect 1532 -4632 2620 -4568
rect 2684 -4632 2704 -4568
rect 1532 -4648 2704 -4632
rect 1532 -4712 2620 -4648
rect 2684 -4712 2704 -4648
rect 1532 -4728 2704 -4712
rect 1532 -4792 2620 -4728
rect 2684 -4792 2704 -4728
rect 1532 -4808 2704 -4792
rect 1532 -4872 2620 -4808
rect 2684 -4872 2704 -4808
rect 1532 -4920 2704 -4872
rect 2944 -4088 4116 -4040
rect 2944 -4152 4032 -4088
rect 4096 -4152 4116 -4088
rect 2944 -4168 4116 -4152
rect 2944 -4232 4032 -4168
rect 4096 -4232 4116 -4168
rect 2944 -4248 4116 -4232
rect 2944 -4312 4032 -4248
rect 4096 -4312 4116 -4248
rect 2944 -4328 4116 -4312
rect 2944 -4392 4032 -4328
rect 4096 -4392 4116 -4328
rect 2944 -4408 4116 -4392
rect 2944 -4472 4032 -4408
rect 4096 -4472 4116 -4408
rect 2944 -4488 4116 -4472
rect 2944 -4552 4032 -4488
rect 4096 -4552 4116 -4488
rect 2944 -4568 4116 -4552
rect 2944 -4632 4032 -4568
rect 4096 -4632 4116 -4568
rect 2944 -4648 4116 -4632
rect 2944 -4712 4032 -4648
rect 4096 -4712 4116 -4648
rect 2944 -4728 4116 -4712
rect 2944 -4792 4032 -4728
rect 4096 -4792 4116 -4728
rect 2944 -4808 4116 -4792
rect 2944 -4872 4032 -4808
rect 4096 -4872 4116 -4808
rect 2944 -4920 4116 -4872
rect 4356 -4088 5528 -4040
rect 4356 -4152 5444 -4088
rect 5508 -4152 5528 -4088
rect 4356 -4168 5528 -4152
rect 4356 -4232 5444 -4168
rect 5508 -4232 5528 -4168
rect 4356 -4248 5528 -4232
rect 4356 -4312 5444 -4248
rect 5508 -4312 5528 -4248
rect 4356 -4328 5528 -4312
rect 4356 -4392 5444 -4328
rect 5508 -4392 5528 -4328
rect 4356 -4408 5528 -4392
rect 4356 -4472 5444 -4408
rect 5508 -4472 5528 -4408
rect 4356 -4488 5528 -4472
rect 4356 -4552 5444 -4488
rect 5508 -4552 5528 -4488
rect 4356 -4568 5528 -4552
rect 4356 -4632 5444 -4568
rect 5508 -4632 5528 -4568
rect 4356 -4648 5528 -4632
rect 4356 -4712 5444 -4648
rect 5508 -4712 5528 -4648
rect 4356 -4728 5528 -4712
rect 4356 -4792 5444 -4728
rect 5508 -4792 5528 -4728
rect 4356 -4808 5528 -4792
rect 4356 -4872 5444 -4808
rect 5508 -4872 5528 -4808
rect 4356 -4920 5528 -4872
rect 5768 -4088 6940 -4040
rect 5768 -4152 6856 -4088
rect 6920 -4152 6940 -4088
rect 5768 -4168 6940 -4152
rect 5768 -4232 6856 -4168
rect 6920 -4232 6940 -4168
rect 5768 -4248 6940 -4232
rect 5768 -4312 6856 -4248
rect 6920 -4312 6940 -4248
rect 5768 -4328 6940 -4312
rect 5768 -4392 6856 -4328
rect 6920 -4392 6940 -4328
rect 5768 -4408 6940 -4392
rect 5768 -4472 6856 -4408
rect 6920 -4472 6940 -4408
rect 5768 -4488 6940 -4472
rect 5768 -4552 6856 -4488
rect 6920 -4552 6940 -4488
rect 5768 -4568 6940 -4552
rect 5768 -4632 6856 -4568
rect 6920 -4632 6940 -4568
rect 5768 -4648 6940 -4632
rect 5768 -4712 6856 -4648
rect 6920 -4712 6940 -4648
rect 5768 -4728 6940 -4712
rect 5768 -4792 6856 -4728
rect 6920 -4792 6940 -4728
rect 5768 -4808 6940 -4792
rect 5768 -4872 6856 -4808
rect 6920 -4872 6940 -4808
rect 5768 -4920 6940 -4872
rect 7180 -4088 8352 -4040
rect 7180 -4152 8268 -4088
rect 8332 -4152 8352 -4088
rect 7180 -4168 8352 -4152
rect 7180 -4232 8268 -4168
rect 8332 -4232 8352 -4168
rect 7180 -4248 8352 -4232
rect 7180 -4312 8268 -4248
rect 8332 -4312 8352 -4248
rect 7180 -4328 8352 -4312
rect 7180 -4392 8268 -4328
rect 8332 -4392 8352 -4328
rect 7180 -4408 8352 -4392
rect 7180 -4472 8268 -4408
rect 8332 -4472 8352 -4408
rect 7180 -4488 8352 -4472
rect 7180 -4552 8268 -4488
rect 8332 -4552 8352 -4488
rect 7180 -4568 8352 -4552
rect 7180 -4632 8268 -4568
rect 8332 -4632 8352 -4568
rect 7180 -4648 8352 -4632
rect 7180 -4712 8268 -4648
rect 8332 -4712 8352 -4648
rect 7180 -4728 8352 -4712
rect 7180 -4792 8268 -4728
rect 8332 -4792 8352 -4728
rect 7180 -4808 8352 -4792
rect 7180 -4872 8268 -4808
rect 8332 -4872 8352 -4808
rect 7180 -4920 8352 -4872
rect 8592 -4088 9764 -4040
rect 8592 -4152 9680 -4088
rect 9744 -4152 9764 -4088
rect 8592 -4168 9764 -4152
rect 8592 -4232 9680 -4168
rect 9744 -4232 9764 -4168
rect 8592 -4248 9764 -4232
rect 8592 -4312 9680 -4248
rect 9744 -4312 9764 -4248
rect 8592 -4328 9764 -4312
rect 8592 -4392 9680 -4328
rect 9744 -4392 9764 -4328
rect 8592 -4408 9764 -4392
rect 8592 -4472 9680 -4408
rect 9744 -4472 9764 -4408
rect 8592 -4488 9764 -4472
rect 8592 -4552 9680 -4488
rect 9744 -4552 9764 -4488
rect 8592 -4568 9764 -4552
rect 8592 -4632 9680 -4568
rect 9744 -4632 9764 -4568
rect 8592 -4648 9764 -4632
rect 8592 -4712 9680 -4648
rect 9744 -4712 9764 -4648
rect 8592 -4728 9764 -4712
rect 8592 -4792 9680 -4728
rect 9744 -4792 9764 -4728
rect 8592 -4808 9764 -4792
rect 8592 -4872 9680 -4808
rect 9744 -4872 9764 -4808
rect 8592 -4920 9764 -4872
rect 10004 -4088 11176 -4040
rect 10004 -4152 11092 -4088
rect 11156 -4152 11176 -4088
rect 10004 -4168 11176 -4152
rect 10004 -4232 11092 -4168
rect 11156 -4232 11176 -4168
rect 10004 -4248 11176 -4232
rect 10004 -4312 11092 -4248
rect 11156 -4312 11176 -4248
rect 10004 -4328 11176 -4312
rect 10004 -4392 11092 -4328
rect 11156 -4392 11176 -4328
rect 10004 -4408 11176 -4392
rect 10004 -4472 11092 -4408
rect 11156 -4472 11176 -4408
rect 10004 -4488 11176 -4472
rect 10004 -4552 11092 -4488
rect 11156 -4552 11176 -4488
rect 10004 -4568 11176 -4552
rect 10004 -4632 11092 -4568
rect 11156 -4632 11176 -4568
rect 10004 -4648 11176 -4632
rect 10004 -4712 11092 -4648
rect 11156 -4712 11176 -4648
rect 10004 -4728 11176 -4712
rect 10004 -4792 11092 -4728
rect 11156 -4792 11176 -4728
rect 10004 -4808 11176 -4792
rect 10004 -4872 11092 -4808
rect 11156 -4872 11176 -4808
rect 10004 -4920 11176 -4872
rect 11416 -4088 12588 -4040
rect 11416 -4152 12504 -4088
rect 12568 -4152 12588 -4088
rect 11416 -4168 12588 -4152
rect 11416 -4232 12504 -4168
rect 12568 -4232 12588 -4168
rect 11416 -4248 12588 -4232
rect 11416 -4312 12504 -4248
rect 12568 -4312 12588 -4248
rect 11416 -4328 12588 -4312
rect 11416 -4392 12504 -4328
rect 12568 -4392 12588 -4328
rect 11416 -4408 12588 -4392
rect 11416 -4472 12504 -4408
rect 12568 -4472 12588 -4408
rect 11416 -4488 12588 -4472
rect 11416 -4552 12504 -4488
rect 12568 -4552 12588 -4488
rect 11416 -4568 12588 -4552
rect 11416 -4632 12504 -4568
rect 12568 -4632 12588 -4568
rect 11416 -4648 12588 -4632
rect 11416 -4712 12504 -4648
rect 12568 -4712 12588 -4648
rect 11416 -4728 12588 -4712
rect 11416 -4792 12504 -4728
rect 12568 -4792 12588 -4728
rect 11416 -4808 12588 -4792
rect 11416 -4872 12504 -4808
rect 12568 -4872 12588 -4808
rect 11416 -4920 12588 -4872
rect 12828 -4088 14000 -4040
rect 12828 -4152 13916 -4088
rect 13980 -4152 14000 -4088
rect 12828 -4168 14000 -4152
rect 12828 -4232 13916 -4168
rect 13980 -4232 14000 -4168
rect 12828 -4248 14000 -4232
rect 12828 -4312 13916 -4248
rect 13980 -4312 14000 -4248
rect 12828 -4328 14000 -4312
rect 12828 -4392 13916 -4328
rect 13980 -4392 14000 -4328
rect 12828 -4408 14000 -4392
rect 12828 -4472 13916 -4408
rect 13980 -4472 14000 -4408
rect 12828 -4488 14000 -4472
rect 12828 -4552 13916 -4488
rect 13980 -4552 14000 -4488
rect 12828 -4568 14000 -4552
rect 12828 -4632 13916 -4568
rect 13980 -4632 14000 -4568
rect 12828 -4648 14000 -4632
rect 12828 -4712 13916 -4648
rect 13980 -4712 14000 -4648
rect 12828 -4728 14000 -4712
rect 12828 -4792 13916 -4728
rect 13980 -4792 14000 -4728
rect 12828 -4808 14000 -4792
rect 12828 -4872 13916 -4808
rect 13980 -4872 14000 -4808
rect 12828 -4920 14000 -4872
rect 14240 -4088 15412 -4040
rect 14240 -4152 15328 -4088
rect 15392 -4152 15412 -4088
rect 14240 -4168 15412 -4152
rect 14240 -4232 15328 -4168
rect 15392 -4232 15412 -4168
rect 14240 -4248 15412 -4232
rect 14240 -4312 15328 -4248
rect 15392 -4312 15412 -4248
rect 14240 -4328 15412 -4312
rect 14240 -4392 15328 -4328
rect 15392 -4392 15412 -4328
rect 14240 -4408 15412 -4392
rect 14240 -4472 15328 -4408
rect 15392 -4472 15412 -4408
rect 14240 -4488 15412 -4472
rect 14240 -4552 15328 -4488
rect 15392 -4552 15412 -4488
rect 14240 -4568 15412 -4552
rect 14240 -4632 15328 -4568
rect 15392 -4632 15412 -4568
rect 14240 -4648 15412 -4632
rect 14240 -4712 15328 -4648
rect 15392 -4712 15412 -4648
rect 14240 -4728 15412 -4712
rect 14240 -4792 15328 -4728
rect 15392 -4792 15412 -4728
rect 14240 -4808 15412 -4792
rect 14240 -4872 15328 -4808
rect 15392 -4872 15412 -4808
rect 14240 -4920 15412 -4872
rect 15652 -4088 16824 -4040
rect 15652 -4152 16740 -4088
rect 16804 -4152 16824 -4088
rect 15652 -4168 16824 -4152
rect 15652 -4232 16740 -4168
rect 16804 -4232 16824 -4168
rect 15652 -4248 16824 -4232
rect 15652 -4312 16740 -4248
rect 16804 -4312 16824 -4248
rect 15652 -4328 16824 -4312
rect 15652 -4392 16740 -4328
rect 16804 -4392 16824 -4328
rect 15652 -4408 16824 -4392
rect 15652 -4472 16740 -4408
rect 16804 -4472 16824 -4408
rect 15652 -4488 16824 -4472
rect 15652 -4552 16740 -4488
rect 16804 -4552 16824 -4488
rect 15652 -4568 16824 -4552
rect 15652 -4632 16740 -4568
rect 16804 -4632 16824 -4568
rect 15652 -4648 16824 -4632
rect 15652 -4712 16740 -4648
rect 16804 -4712 16824 -4648
rect 15652 -4728 16824 -4712
rect 15652 -4792 16740 -4728
rect 16804 -4792 16824 -4728
rect 15652 -4808 16824 -4792
rect 15652 -4872 16740 -4808
rect 16804 -4872 16824 -4808
rect 15652 -4920 16824 -4872
rect 17064 -4088 18236 -4040
rect 17064 -4152 18152 -4088
rect 18216 -4152 18236 -4088
rect 17064 -4168 18236 -4152
rect 17064 -4232 18152 -4168
rect 18216 -4232 18236 -4168
rect 17064 -4248 18236 -4232
rect 17064 -4312 18152 -4248
rect 18216 -4312 18236 -4248
rect 17064 -4328 18236 -4312
rect 17064 -4392 18152 -4328
rect 18216 -4392 18236 -4328
rect 17064 -4408 18236 -4392
rect 17064 -4472 18152 -4408
rect 18216 -4472 18236 -4408
rect 17064 -4488 18236 -4472
rect 17064 -4552 18152 -4488
rect 18216 -4552 18236 -4488
rect 17064 -4568 18236 -4552
rect 17064 -4632 18152 -4568
rect 18216 -4632 18236 -4568
rect 17064 -4648 18236 -4632
rect 17064 -4712 18152 -4648
rect 18216 -4712 18236 -4648
rect 17064 -4728 18236 -4712
rect 17064 -4792 18152 -4728
rect 18216 -4792 18236 -4728
rect 17064 -4808 18236 -4792
rect 17064 -4872 18152 -4808
rect 18216 -4872 18236 -4808
rect 17064 -4920 18236 -4872
rect 18476 -4088 19648 -4040
rect 18476 -4152 19564 -4088
rect 19628 -4152 19648 -4088
rect 18476 -4168 19648 -4152
rect 18476 -4232 19564 -4168
rect 19628 -4232 19648 -4168
rect 18476 -4248 19648 -4232
rect 18476 -4312 19564 -4248
rect 19628 -4312 19648 -4248
rect 18476 -4328 19648 -4312
rect 18476 -4392 19564 -4328
rect 19628 -4392 19648 -4328
rect 18476 -4408 19648 -4392
rect 18476 -4472 19564 -4408
rect 19628 -4472 19648 -4408
rect 18476 -4488 19648 -4472
rect 18476 -4552 19564 -4488
rect 19628 -4552 19648 -4488
rect 18476 -4568 19648 -4552
rect 18476 -4632 19564 -4568
rect 19628 -4632 19648 -4568
rect 18476 -4648 19648 -4632
rect 18476 -4712 19564 -4648
rect 19628 -4712 19648 -4648
rect 18476 -4728 19648 -4712
rect 18476 -4792 19564 -4728
rect 19628 -4792 19648 -4728
rect 18476 -4808 19648 -4792
rect 18476 -4872 19564 -4808
rect 19628 -4872 19648 -4808
rect 18476 -4920 19648 -4872
rect 19888 -4088 21060 -4040
rect 19888 -4152 20976 -4088
rect 21040 -4152 21060 -4088
rect 19888 -4168 21060 -4152
rect 19888 -4232 20976 -4168
rect 21040 -4232 21060 -4168
rect 19888 -4248 21060 -4232
rect 19888 -4312 20976 -4248
rect 21040 -4312 21060 -4248
rect 19888 -4328 21060 -4312
rect 19888 -4392 20976 -4328
rect 21040 -4392 21060 -4328
rect 19888 -4408 21060 -4392
rect 19888 -4472 20976 -4408
rect 21040 -4472 21060 -4408
rect 19888 -4488 21060 -4472
rect 19888 -4552 20976 -4488
rect 21040 -4552 21060 -4488
rect 19888 -4568 21060 -4552
rect 19888 -4632 20976 -4568
rect 21040 -4632 21060 -4568
rect 19888 -4648 21060 -4632
rect 19888 -4712 20976 -4648
rect 21040 -4712 21060 -4648
rect 19888 -4728 21060 -4712
rect 19888 -4792 20976 -4728
rect 21040 -4792 21060 -4728
rect 19888 -4808 21060 -4792
rect 19888 -4872 20976 -4808
rect 21040 -4872 21060 -4808
rect 19888 -4920 21060 -4872
rect 21300 -4088 22472 -4040
rect 21300 -4152 22388 -4088
rect 22452 -4152 22472 -4088
rect 21300 -4168 22472 -4152
rect 21300 -4232 22388 -4168
rect 22452 -4232 22472 -4168
rect 21300 -4248 22472 -4232
rect 21300 -4312 22388 -4248
rect 22452 -4312 22472 -4248
rect 21300 -4328 22472 -4312
rect 21300 -4392 22388 -4328
rect 22452 -4392 22472 -4328
rect 21300 -4408 22472 -4392
rect 21300 -4472 22388 -4408
rect 22452 -4472 22472 -4408
rect 21300 -4488 22472 -4472
rect 21300 -4552 22388 -4488
rect 22452 -4552 22472 -4488
rect 21300 -4568 22472 -4552
rect 21300 -4632 22388 -4568
rect 22452 -4632 22472 -4568
rect 21300 -4648 22472 -4632
rect 21300 -4712 22388 -4648
rect 22452 -4712 22472 -4648
rect 21300 -4728 22472 -4712
rect 21300 -4792 22388 -4728
rect 22452 -4792 22472 -4728
rect 21300 -4808 22472 -4792
rect 21300 -4872 22388 -4808
rect 22452 -4872 22472 -4808
rect 21300 -4920 22472 -4872
rect 22712 -4088 23884 -4040
rect 22712 -4152 23800 -4088
rect 23864 -4152 23884 -4088
rect 22712 -4168 23884 -4152
rect 22712 -4232 23800 -4168
rect 23864 -4232 23884 -4168
rect 22712 -4248 23884 -4232
rect 22712 -4312 23800 -4248
rect 23864 -4312 23884 -4248
rect 22712 -4328 23884 -4312
rect 22712 -4392 23800 -4328
rect 23864 -4392 23884 -4328
rect 22712 -4408 23884 -4392
rect 22712 -4472 23800 -4408
rect 23864 -4472 23884 -4408
rect 22712 -4488 23884 -4472
rect 22712 -4552 23800 -4488
rect 23864 -4552 23884 -4488
rect 22712 -4568 23884 -4552
rect 22712 -4632 23800 -4568
rect 23864 -4632 23884 -4568
rect 22712 -4648 23884 -4632
rect 22712 -4712 23800 -4648
rect 23864 -4712 23884 -4648
rect 22712 -4728 23884 -4712
rect 22712 -4792 23800 -4728
rect 23864 -4792 23884 -4728
rect 22712 -4808 23884 -4792
rect 22712 -4872 23800 -4808
rect 23864 -4872 23884 -4808
rect 22712 -4920 23884 -4872
rect -23884 -5208 -22712 -5160
rect -23884 -5272 -22796 -5208
rect -22732 -5272 -22712 -5208
rect -23884 -5288 -22712 -5272
rect -23884 -5352 -22796 -5288
rect -22732 -5352 -22712 -5288
rect -23884 -5368 -22712 -5352
rect -23884 -5432 -22796 -5368
rect -22732 -5432 -22712 -5368
rect -23884 -5448 -22712 -5432
rect -23884 -5512 -22796 -5448
rect -22732 -5512 -22712 -5448
rect -23884 -5528 -22712 -5512
rect -23884 -5592 -22796 -5528
rect -22732 -5592 -22712 -5528
rect -23884 -5608 -22712 -5592
rect -23884 -5672 -22796 -5608
rect -22732 -5672 -22712 -5608
rect -23884 -5688 -22712 -5672
rect -23884 -5752 -22796 -5688
rect -22732 -5752 -22712 -5688
rect -23884 -5768 -22712 -5752
rect -23884 -5832 -22796 -5768
rect -22732 -5832 -22712 -5768
rect -23884 -5848 -22712 -5832
rect -23884 -5912 -22796 -5848
rect -22732 -5912 -22712 -5848
rect -23884 -5928 -22712 -5912
rect -23884 -5992 -22796 -5928
rect -22732 -5992 -22712 -5928
rect -23884 -6040 -22712 -5992
rect -22472 -5208 -21300 -5160
rect -22472 -5272 -21384 -5208
rect -21320 -5272 -21300 -5208
rect -22472 -5288 -21300 -5272
rect -22472 -5352 -21384 -5288
rect -21320 -5352 -21300 -5288
rect -22472 -5368 -21300 -5352
rect -22472 -5432 -21384 -5368
rect -21320 -5432 -21300 -5368
rect -22472 -5448 -21300 -5432
rect -22472 -5512 -21384 -5448
rect -21320 -5512 -21300 -5448
rect -22472 -5528 -21300 -5512
rect -22472 -5592 -21384 -5528
rect -21320 -5592 -21300 -5528
rect -22472 -5608 -21300 -5592
rect -22472 -5672 -21384 -5608
rect -21320 -5672 -21300 -5608
rect -22472 -5688 -21300 -5672
rect -22472 -5752 -21384 -5688
rect -21320 -5752 -21300 -5688
rect -22472 -5768 -21300 -5752
rect -22472 -5832 -21384 -5768
rect -21320 -5832 -21300 -5768
rect -22472 -5848 -21300 -5832
rect -22472 -5912 -21384 -5848
rect -21320 -5912 -21300 -5848
rect -22472 -5928 -21300 -5912
rect -22472 -5992 -21384 -5928
rect -21320 -5992 -21300 -5928
rect -22472 -6040 -21300 -5992
rect -21060 -5208 -19888 -5160
rect -21060 -5272 -19972 -5208
rect -19908 -5272 -19888 -5208
rect -21060 -5288 -19888 -5272
rect -21060 -5352 -19972 -5288
rect -19908 -5352 -19888 -5288
rect -21060 -5368 -19888 -5352
rect -21060 -5432 -19972 -5368
rect -19908 -5432 -19888 -5368
rect -21060 -5448 -19888 -5432
rect -21060 -5512 -19972 -5448
rect -19908 -5512 -19888 -5448
rect -21060 -5528 -19888 -5512
rect -21060 -5592 -19972 -5528
rect -19908 -5592 -19888 -5528
rect -21060 -5608 -19888 -5592
rect -21060 -5672 -19972 -5608
rect -19908 -5672 -19888 -5608
rect -21060 -5688 -19888 -5672
rect -21060 -5752 -19972 -5688
rect -19908 -5752 -19888 -5688
rect -21060 -5768 -19888 -5752
rect -21060 -5832 -19972 -5768
rect -19908 -5832 -19888 -5768
rect -21060 -5848 -19888 -5832
rect -21060 -5912 -19972 -5848
rect -19908 -5912 -19888 -5848
rect -21060 -5928 -19888 -5912
rect -21060 -5992 -19972 -5928
rect -19908 -5992 -19888 -5928
rect -21060 -6040 -19888 -5992
rect -19648 -5208 -18476 -5160
rect -19648 -5272 -18560 -5208
rect -18496 -5272 -18476 -5208
rect -19648 -5288 -18476 -5272
rect -19648 -5352 -18560 -5288
rect -18496 -5352 -18476 -5288
rect -19648 -5368 -18476 -5352
rect -19648 -5432 -18560 -5368
rect -18496 -5432 -18476 -5368
rect -19648 -5448 -18476 -5432
rect -19648 -5512 -18560 -5448
rect -18496 -5512 -18476 -5448
rect -19648 -5528 -18476 -5512
rect -19648 -5592 -18560 -5528
rect -18496 -5592 -18476 -5528
rect -19648 -5608 -18476 -5592
rect -19648 -5672 -18560 -5608
rect -18496 -5672 -18476 -5608
rect -19648 -5688 -18476 -5672
rect -19648 -5752 -18560 -5688
rect -18496 -5752 -18476 -5688
rect -19648 -5768 -18476 -5752
rect -19648 -5832 -18560 -5768
rect -18496 -5832 -18476 -5768
rect -19648 -5848 -18476 -5832
rect -19648 -5912 -18560 -5848
rect -18496 -5912 -18476 -5848
rect -19648 -5928 -18476 -5912
rect -19648 -5992 -18560 -5928
rect -18496 -5992 -18476 -5928
rect -19648 -6040 -18476 -5992
rect -18236 -5208 -17064 -5160
rect -18236 -5272 -17148 -5208
rect -17084 -5272 -17064 -5208
rect -18236 -5288 -17064 -5272
rect -18236 -5352 -17148 -5288
rect -17084 -5352 -17064 -5288
rect -18236 -5368 -17064 -5352
rect -18236 -5432 -17148 -5368
rect -17084 -5432 -17064 -5368
rect -18236 -5448 -17064 -5432
rect -18236 -5512 -17148 -5448
rect -17084 -5512 -17064 -5448
rect -18236 -5528 -17064 -5512
rect -18236 -5592 -17148 -5528
rect -17084 -5592 -17064 -5528
rect -18236 -5608 -17064 -5592
rect -18236 -5672 -17148 -5608
rect -17084 -5672 -17064 -5608
rect -18236 -5688 -17064 -5672
rect -18236 -5752 -17148 -5688
rect -17084 -5752 -17064 -5688
rect -18236 -5768 -17064 -5752
rect -18236 -5832 -17148 -5768
rect -17084 -5832 -17064 -5768
rect -18236 -5848 -17064 -5832
rect -18236 -5912 -17148 -5848
rect -17084 -5912 -17064 -5848
rect -18236 -5928 -17064 -5912
rect -18236 -5992 -17148 -5928
rect -17084 -5992 -17064 -5928
rect -18236 -6040 -17064 -5992
rect -16824 -5208 -15652 -5160
rect -16824 -5272 -15736 -5208
rect -15672 -5272 -15652 -5208
rect -16824 -5288 -15652 -5272
rect -16824 -5352 -15736 -5288
rect -15672 -5352 -15652 -5288
rect -16824 -5368 -15652 -5352
rect -16824 -5432 -15736 -5368
rect -15672 -5432 -15652 -5368
rect -16824 -5448 -15652 -5432
rect -16824 -5512 -15736 -5448
rect -15672 -5512 -15652 -5448
rect -16824 -5528 -15652 -5512
rect -16824 -5592 -15736 -5528
rect -15672 -5592 -15652 -5528
rect -16824 -5608 -15652 -5592
rect -16824 -5672 -15736 -5608
rect -15672 -5672 -15652 -5608
rect -16824 -5688 -15652 -5672
rect -16824 -5752 -15736 -5688
rect -15672 -5752 -15652 -5688
rect -16824 -5768 -15652 -5752
rect -16824 -5832 -15736 -5768
rect -15672 -5832 -15652 -5768
rect -16824 -5848 -15652 -5832
rect -16824 -5912 -15736 -5848
rect -15672 -5912 -15652 -5848
rect -16824 -5928 -15652 -5912
rect -16824 -5992 -15736 -5928
rect -15672 -5992 -15652 -5928
rect -16824 -6040 -15652 -5992
rect -15412 -5208 -14240 -5160
rect -15412 -5272 -14324 -5208
rect -14260 -5272 -14240 -5208
rect -15412 -5288 -14240 -5272
rect -15412 -5352 -14324 -5288
rect -14260 -5352 -14240 -5288
rect -15412 -5368 -14240 -5352
rect -15412 -5432 -14324 -5368
rect -14260 -5432 -14240 -5368
rect -15412 -5448 -14240 -5432
rect -15412 -5512 -14324 -5448
rect -14260 -5512 -14240 -5448
rect -15412 -5528 -14240 -5512
rect -15412 -5592 -14324 -5528
rect -14260 -5592 -14240 -5528
rect -15412 -5608 -14240 -5592
rect -15412 -5672 -14324 -5608
rect -14260 -5672 -14240 -5608
rect -15412 -5688 -14240 -5672
rect -15412 -5752 -14324 -5688
rect -14260 -5752 -14240 -5688
rect -15412 -5768 -14240 -5752
rect -15412 -5832 -14324 -5768
rect -14260 -5832 -14240 -5768
rect -15412 -5848 -14240 -5832
rect -15412 -5912 -14324 -5848
rect -14260 -5912 -14240 -5848
rect -15412 -5928 -14240 -5912
rect -15412 -5992 -14324 -5928
rect -14260 -5992 -14240 -5928
rect -15412 -6040 -14240 -5992
rect -14000 -5208 -12828 -5160
rect -14000 -5272 -12912 -5208
rect -12848 -5272 -12828 -5208
rect -14000 -5288 -12828 -5272
rect -14000 -5352 -12912 -5288
rect -12848 -5352 -12828 -5288
rect -14000 -5368 -12828 -5352
rect -14000 -5432 -12912 -5368
rect -12848 -5432 -12828 -5368
rect -14000 -5448 -12828 -5432
rect -14000 -5512 -12912 -5448
rect -12848 -5512 -12828 -5448
rect -14000 -5528 -12828 -5512
rect -14000 -5592 -12912 -5528
rect -12848 -5592 -12828 -5528
rect -14000 -5608 -12828 -5592
rect -14000 -5672 -12912 -5608
rect -12848 -5672 -12828 -5608
rect -14000 -5688 -12828 -5672
rect -14000 -5752 -12912 -5688
rect -12848 -5752 -12828 -5688
rect -14000 -5768 -12828 -5752
rect -14000 -5832 -12912 -5768
rect -12848 -5832 -12828 -5768
rect -14000 -5848 -12828 -5832
rect -14000 -5912 -12912 -5848
rect -12848 -5912 -12828 -5848
rect -14000 -5928 -12828 -5912
rect -14000 -5992 -12912 -5928
rect -12848 -5992 -12828 -5928
rect -14000 -6040 -12828 -5992
rect -12588 -5208 -11416 -5160
rect -12588 -5272 -11500 -5208
rect -11436 -5272 -11416 -5208
rect -12588 -5288 -11416 -5272
rect -12588 -5352 -11500 -5288
rect -11436 -5352 -11416 -5288
rect -12588 -5368 -11416 -5352
rect -12588 -5432 -11500 -5368
rect -11436 -5432 -11416 -5368
rect -12588 -5448 -11416 -5432
rect -12588 -5512 -11500 -5448
rect -11436 -5512 -11416 -5448
rect -12588 -5528 -11416 -5512
rect -12588 -5592 -11500 -5528
rect -11436 -5592 -11416 -5528
rect -12588 -5608 -11416 -5592
rect -12588 -5672 -11500 -5608
rect -11436 -5672 -11416 -5608
rect -12588 -5688 -11416 -5672
rect -12588 -5752 -11500 -5688
rect -11436 -5752 -11416 -5688
rect -12588 -5768 -11416 -5752
rect -12588 -5832 -11500 -5768
rect -11436 -5832 -11416 -5768
rect -12588 -5848 -11416 -5832
rect -12588 -5912 -11500 -5848
rect -11436 -5912 -11416 -5848
rect -12588 -5928 -11416 -5912
rect -12588 -5992 -11500 -5928
rect -11436 -5992 -11416 -5928
rect -12588 -6040 -11416 -5992
rect -11176 -5208 -10004 -5160
rect -11176 -5272 -10088 -5208
rect -10024 -5272 -10004 -5208
rect -11176 -5288 -10004 -5272
rect -11176 -5352 -10088 -5288
rect -10024 -5352 -10004 -5288
rect -11176 -5368 -10004 -5352
rect -11176 -5432 -10088 -5368
rect -10024 -5432 -10004 -5368
rect -11176 -5448 -10004 -5432
rect -11176 -5512 -10088 -5448
rect -10024 -5512 -10004 -5448
rect -11176 -5528 -10004 -5512
rect -11176 -5592 -10088 -5528
rect -10024 -5592 -10004 -5528
rect -11176 -5608 -10004 -5592
rect -11176 -5672 -10088 -5608
rect -10024 -5672 -10004 -5608
rect -11176 -5688 -10004 -5672
rect -11176 -5752 -10088 -5688
rect -10024 -5752 -10004 -5688
rect -11176 -5768 -10004 -5752
rect -11176 -5832 -10088 -5768
rect -10024 -5832 -10004 -5768
rect -11176 -5848 -10004 -5832
rect -11176 -5912 -10088 -5848
rect -10024 -5912 -10004 -5848
rect -11176 -5928 -10004 -5912
rect -11176 -5992 -10088 -5928
rect -10024 -5992 -10004 -5928
rect -11176 -6040 -10004 -5992
rect -9764 -5208 -8592 -5160
rect -9764 -5272 -8676 -5208
rect -8612 -5272 -8592 -5208
rect -9764 -5288 -8592 -5272
rect -9764 -5352 -8676 -5288
rect -8612 -5352 -8592 -5288
rect -9764 -5368 -8592 -5352
rect -9764 -5432 -8676 -5368
rect -8612 -5432 -8592 -5368
rect -9764 -5448 -8592 -5432
rect -9764 -5512 -8676 -5448
rect -8612 -5512 -8592 -5448
rect -9764 -5528 -8592 -5512
rect -9764 -5592 -8676 -5528
rect -8612 -5592 -8592 -5528
rect -9764 -5608 -8592 -5592
rect -9764 -5672 -8676 -5608
rect -8612 -5672 -8592 -5608
rect -9764 -5688 -8592 -5672
rect -9764 -5752 -8676 -5688
rect -8612 -5752 -8592 -5688
rect -9764 -5768 -8592 -5752
rect -9764 -5832 -8676 -5768
rect -8612 -5832 -8592 -5768
rect -9764 -5848 -8592 -5832
rect -9764 -5912 -8676 -5848
rect -8612 -5912 -8592 -5848
rect -9764 -5928 -8592 -5912
rect -9764 -5992 -8676 -5928
rect -8612 -5992 -8592 -5928
rect -9764 -6040 -8592 -5992
rect -8352 -5208 -7180 -5160
rect -8352 -5272 -7264 -5208
rect -7200 -5272 -7180 -5208
rect -8352 -5288 -7180 -5272
rect -8352 -5352 -7264 -5288
rect -7200 -5352 -7180 -5288
rect -8352 -5368 -7180 -5352
rect -8352 -5432 -7264 -5368
rect -7200 -5432 -7180 -5368
rect -8352 -5448 -7180 -5432
rect -8352 -5512 -7264 -5448
rect -7200 -5512 -7180 -5448
rect -8352 -5528 -7180 -5512
rect -8352 -5592 -7264 -5528
rect -7200 -5592 -7180 -5528
rect -8352 -5608 -7180 -5592
rect -8352 -5672 -7264 -5608
rect -7200 -5672 -7180 -5608
rect -8352 -5688 -7180 -5672
rect -8352 -5752 -7264 -5688
rect -7200 -5752 -7180 -5688
rect -8352 -5768 -7180 -5752
rect -8352 -5832 -7264 -5768
rect -7200 -5832 -7180 -5768
rect -8352 -5848 -7180 -5832
rect -8352 -5912 -7264 -5848
rect -7200 -5912 -7180 -5848
rect -8352 -5928 -7180 -5912
rect -8352 -5992 -7264 -5928
rect -7200 -5992 -7180 -5928
rect -8352 -6040 -7180 -5992
rect -6940 -5208 -5768 -5160
rect -6940 -5272 -5852 -5208
rect -5788 -5272 -5768 -5208
rect -6940 -5288 -5768 -5272
rect -6940 -5352 -5852 -5288
rect -5788 -5352 -5768 -5288
rect -6940 -5368 -5768 -5352
rect -6940 -5432 -5852 -5368
rect -5788 -5432 -5768 -5368
rect -6940 -5448 -5768 -5432
rect -6940 -5512 -5852 -5448
rect -5788 -5512 -5768 -5448
rect -6940 -5528 -5768 -5512
rect -6940 -5592 -5852 -5528
rect -5788 -5592 -5768 -5528
rect -6940 -5608 -5768 -5592
rect -6940 -5672 -5852 -5608
rect -5788 -5672 -5768 -5608
rect -6940 -5688 -5768 -5672
rect -6940 -5752 -5852 -5688
rect -5788 -5752 -5768 -5688
rect -6940 -5768 -5768 -5752
rect -6940 -5832 -5852 -5768
rect -5788 -5832 -5768 -5768
rect -6940 -5848 -5768 -5832
rect -6940 -5912 -5852 -5848
rect -5788 -5912 -5768 -5848
rect -6940 -5928 -5768 -5912
rect -6940 -5992 -5852 -5928
rect -5788 -5992 -5768 -5928
rect -6940 -6040 -5768 -5992
rect -5528 -5208 -4356 -5160
rect -5528 -5272 -4440 -5208
rect -4376 -5272 -4356 -5208
rect -5528 -5288 -4356 -5272
rect -5528 -5352 -4440 -5288
rect -4376 -5352 -4356 -5288
rect -5528 -5368 -4356 -5352
rect -5528 -5432 -4440 -5368
rect -4376 -5432 -4356 -5368
rect -5528 -5448 -4356 -5432
rect -5528 -5512 -4440 -5448
rect -4376 -5512 -4356 -5448
rect -5528 -5528 -4356 -5512
rect -5528 -5592 -4440 -5528
rect -4376 -5592 -4356 -5528
rect -5528 -5608 -4356 -5592
rect -5528 -5672 -4440 -5608
rect -4376 -5672 -4356 -5608
rect -5528 -5688 -4356 -5672
rect -5528 -5752 -4440 -5688
rect -4376 -5752 -4356 -5688
rect -5528 -5768 -4356 -5752
rect -5528 -5832 -4440 -5768
rect -4376 -5832 -4356 -5768
rect -5528 -5848 -4356 -5832
rect -5528 -5912 -4440 -5848
rect -4376 -5912 -4356 -5848
rect -5528 -5928 -4356 -5912
rect -5528 -5992 -4440 -5928
rect -4376 -5992 -4356 -5928
rect -5528 -6040 -4356 -5992
rect -4116 -5208 -2944 -5160
rect -4116 -5272 -3028 -5208
rect -2964 -5272 -2944 -5208
rect -4116 -5288 -2944 -5272
rect -4116 -5352 -3028 -5288
rect -2964 -5352 -2944 -5288
rect -4116 -5368 -2944 -5352
rect -4116 -5432 -3028 -5368
rect -2964 -5432 -2944 -5368
rect -4116 -5448 -2944 -5432
rect -4116 -5512 -3028 -5448
rect -2964 -5512 -2944 -5448
rect -4116 -5528 -2944 -5512
rect -4116 -5592 -3028 -5528
rect -2964 -5592 -2944 -5528
rect -4116 -5608 -2944 -5592
rect -4116 -5672 -3028 -5608
rect -2964 -5672 -2944 -5608
rect -4116 -5688 -2944 -5672
rect -4116 -5752 -3028 -5688
rect -2964 -5752 -2944 -5688
rect -4116 -5768 -2944 -5752
rect -4116 -5832 -3028 -5768
rect -2964 -5832 -2944 -5768
rect -4116 -5848 -2944 -5832
rect -4116 -5912 -3028 -5848
rect -2964 -5912 -2944 -5848
rect -4116 -5928 -2944 -5912
rect -4116 -5992 -3028 -5928
rect -2964 -5992 -2944 -5928
rect -4116 -6040 -2944 -5992
rect -2704 -5208 -1532 -5160
rect -2704 -5272 -1616 -5208
rect -1552 -5272 -1532 -5208
rect -2704 -5288 -1532 -5272
rect -2704 -5352 -1616 -5288
rect -1552 -5352 -1532 -5288
rect -2704 -5368 -1532 -5352
rect -2704 -5432 -1616 -5368
rect -1552 -5432 -1532 -5368
rect -2704 -5448 -1532 -5432
rect -2704 -5512 -1616 -5448
rect -1552 -5512 -1532 -5448
rect -2704 -5528 -1532 -5512
rect -2704 -5592 -1616 -5528
rect -1552 -5592 -1532 -5528
rect -2704 -5608 -1532 -5592
rect -2704 -5672 -1616 -5608
rect -1552 -5672 -1532 -5608
rect -2704 -5688 -1532 -5672
rect -2704 -5752 -1616 -5688
rect -1552 -5752 -1532 -5688
rect -2704 -5768 -1532 -5752
rect -2704 -5832 -1616 -5768
rect -1552 -5832 -1532 -5768
rect -2704 -5848 -1532 -5832
rect -2704 -5912 -1616 -5848
rect -1552 -5912 -1532 -5848
rect -2704 -5928 -1532 -5912
rect -2704 -5992 -1616 -5928
rect -1552 -5992 -1532 -5928
rect -2704 -6040 -1532 -5992
rect -1292 -5208 -120 -5160
rect -1292 -5272 -204 -5208
rect -140 -5272 -120 -5208
rect -1292 -5288 -120 -5272
rect -1292 -5352 -204 -5288
rect -140 -5352 -120 -5288
rect -1292 -5368 -120 -5352
rect -1292 -5432 -204 -5368
rect -140 -5432 -120 -5368
rect -1292 -5448 -120 -5432
rect -1292 -5512 -204 -5448
rect -140 -5512 -120 -5448
rect -1292 -5528 -120 -5512
rect -1292 -5592 -204 -5528
rect -140 -5592 -120 -5528
rect -1292 -5608 -120 -5592
rect -1292 -5672 -204 -5608
rect -140 -5672 -120 -5608
rect -1292 -5688 -120 -5672
rect -1292 -5752 -204 -5688
rect -140 -5752 -120 -5688
rect -1292 -5768 -120 -5752
rect -1292 -5832 -204 -5768
rect -140 -5832 -120 -5768
rect -1292 -5848 -120 -5832
rect -1292 -5912 -204 -5848
rect -140 -5912 -120 -5848
rect -1292 -5928 -120 -5912
rect -1292 -5992 -204 -5928
rect -140 -5992 -120 -5928
rect -1292 -6040 -120 -5992
rect 120 -5208 1292 -5160
rect 120 -5272 1208 -5208
rect 1272 -5272 1292 -5208
rect 120 -5288 1292 -5272
rect 120 -5352 1208 -5288
rect 1272 -5352 1292 -5288
rect 120 -5368 1292 -5352
rect 120 -5432 1208 -5368
rect 1272 -5432 1292 -5368
rect 120 -5448 1292 -5432
rect 120 -5512 1208 -5448
rect 1272 -5512 1292 -5448
rect 120 -5528 1292 -5512
rect 120 -5592 1208 -5528
rect 1272 -5592 1292 -5528
rect 120 -5608 1292 -5592
rect 120 -5672 1208 -5608
rect 1272 -5672 1292 -5608
rect 120 -5688 1292 -5672
rect 120 -5752 1208 -5688
rect 1272 -5752 1292 -5688
rect 120 -5768 1292 -5752
rect 120 -5832 1208 -5768
rect 1272 -5832 1292 -5768
rect 120 -5848 1292 -5832
rect 120 -5912 1208 -5848
rect 1272 -5912 1292 -5848
rect 120 -5928 1292 -5912
rect 120 -5992 1208 -5928
rect 1272 -5992 1292 -5928
rect 120 -6040 1292 -5992
rect 1532 -5208 2704 -5160
rect 1532 -5272 2620 -5208
rect 2684 -5272 2704 -5208
rect 1532 -5288 2704 -5272
rect 1532 -5352 2620 -5288
rect 2684 -5352 2704 -5288
rect 1532 -5368 2704 -5352
rect 1532 -5432 2620 -5368
rect 2684 -5432 2704 -5368
rect 1532 -5448 2704 -5432
rect 1532 -5512 2620 -5448
rect 2684 -5512 2704 -5448
rect 1532 -5528 2704 -5512
rect 1532 -5592 2620 -5528
rect 2684 -5592 2704 -5528
rect 1532 -5608 2704 -5592
rect 1532 -5672 2620 -5608
rect 2684 -5672 2704 -5608
rect 1532 -5688 2704 -5672
rect 1532 -5752 2620 -5688
rect 2684 -5752 2704 -5688
rect 1532 -5768 2704 -5752
rect 1532 -5832 2620 -5768
rect 2684 -5832 2704 -5768
rect 1532 -5848 2704 -5832
rect 1532 -5912 2620 -5848
rect 2684 -5912 2704 -5848
rect 1532 -5928 2704 -5912
rect 1532 -5992 2620 -5928
rect 2684 -5992 2704 -5928
rect 1532 -6040 2704 -5992
rect 2944 -5208 4116 -5160
rect 2944 -5272 4032 -5208
rect 4096 -5272 4116 -5208
rect 2944 -5288 4116 -5272
rect 2944 -5352 4032 -5288
rect 4096 -5352 4116 -5288
rect 2944 -5368 4116 -5352
rect 2944 -5432 4032 -5368
rect 4096 -5432 4116 -5368
rect 2944 -5448 4116 -5432
rect 2944 -5512 4032 -5448
rect 4096 -5512 4116 -5448
rect 2944 -5528 4116 -5512
rect 2944 -5592 4032 -5528
rect 4096 -5592 4116 -5528
rect 2944 -5608 4116 -5592
rect 2944 -5672 4032 -5608
rect 4096 -5672 4116 -5608
rect 2944 -5688 4116 -5672
rect 2944 -5752 4032 -5688
rect 4096 -5752 4116 -5688
rect 2944 -5768 4116 -5752
rect 2944 -5832 4032 -5768
rect 4096 -5832 4116 -5768
rect 2944 -5848 4116 -5832
rect 2944 -5912 4032 -5848
rect 4096 -5912 4116 -5848
rect 2944 -5928 4116 -5912
rect 2944 -5992 4032 -5928
rect 4096 -5992 4116 -5928
rect 2944 -6040 4116 -5992
rect 4356 -5208 5528 -5160
rect 4356 -5272 5444 -5208
rect 5508 -5272 5528 -5208
rect 4356 -5288 5528 -5272
rect 4356 -5352 5444 -5288
rect 5508 -5352 5528 -5288
rect 4356 -5368 5528 -5352
rect 4356 -5432 5444 -5368
rect 5508 -5432 5528 -5368
rect 4356 -5448 5528 -5432
rect 4356 -5512 5444 -5448
rect 5508 -5512 5528 -5448
rect 4356 -5528 5528 -5512
rect 4356 -5592 5444 -5528
rect 5508 -5592 5528 -5528
rect 4356 -5608 5528 -5592
rect 4356 -5672 5444 -5608
rect 5508 -5672 5528 -5608
rect 4356 -5688 5528 -5672
rect 4356 -5752 5444 -5688
rect 5508 -5752 5528 -5688
rect 4356 -5768 5528 -5752
rect 4356 -5832 5444 -5768
rect 5508 -5832 5528 -5768
rect 4356 -5848 5528 -5832
rect 4356 -5912 5444 -5848
rect 5508 -5912 5528 -5848
rect 4356 -5928 5528 -5912
rect 4356 -5992 5444 -5928
rect 5508 -5992 5528 -5928
rect 4356 -6040 5528 -5992
rect 5768 -5208 6940 -5160
rect 5768 -5272 6856 -5208
rect 6920 -5272 6940 -5208
rect 5768 -5288 6940 -5272
rect 5768 -5352 6856 -5288
rect 6920 -5352 6940 -5288
rect 5768 -5368 6940 -5352
rect 5768 -5432 6856 -5368
rect 6920 -5432 6940 -5368
rect 5768 -5448 6940 -5432
rect 5768 -5512 6856 -5448
rect 6920 -5512 6940 -5448
rect 5768 -5528 6940 -5512
rect 5768 -5592 6856 -5528
rect 6920 -5592 6940 -5528
rect 5768 -5608 6940 -5592
rect 5768 -5672 6856 -5608
rect 6920 -5672 6940 -5608
rect 5768 -5688 6940 -5672
rect 5768 -5752 6856 -5688
rect 6920 -5752 6940 -5688
rect 5768 -5768 6940 -5752
rect 5768 -5832 6856 -5768
rect 6920 -5832 6940 -5768
rect 5768 -5848 6940 -5832
rect 5768 -5912 6856 -5848
rect 6920 -5912 6940 -5848
rect 5768 -5928 6940 -5912
rect 5768 -5992 6856 -5928
rect 6920 -5992 6940 -5928
rect 5768 -6040 6940 -5992
rect 7180 -5208 8352 -5160
rect 7180 -5272 8268 -5208
rect 8332 -5272 8352 -5208
rect 7180 -5288 8352 -5272
rect 7180 -5352 8268 -5288
rect 8332 -5352 8352 -5288
rect 7180 -5368 8352 -5352
rect 7180 -5432 8268 -5368
rect 8332 -5432 8352 -5368
rect 7180 -5448 8352 -5432
rect 7180 -5512 8268 -5448
rect 8332 -5512 8352 -5448
rect 7180 -5528 8352 -5512
rect 7180 -5592 8268 -5528
rect 8332 -5592 8352 -5528
rect 7180 -5608 8352 -5592
rect 7180 -5672 8268 -5608
rect 8332 -5672 8352 -5608
rect 7180 -5688 8352 -5672
rect 7180 -5752 8268 -5688
rect 8332 -5752 8352 -5688
rect 7180 -5768 8352 -5752
rect 7180 -5832 8268 -5768
rect 8332 -5832 8352 -5768
rect 7180 -5848 8352 -5832
rect 7180 -5912 8268 -5848
rect 8332 -5912 8352 -5848
rect 7180 -5928 8352 -5912
rect 7180 -5992 8268 -5928
rect 8332 -5992 8352 -5928
rect 7180 -6040 8352 -5992
rect 8592 -5208 9764 -5160
rect 8592 -5272 9680 -5208
rect 9744 -5272 9764 -5208
rect 8592 -5288 9764 -5272
rect 8592 -5352 9680 -5288
rect 9744 -5352 9764 -5288
rect 8592 -5368 9764 -5352
rect 8592 -5432 9680 -5368
rect 9744 -5432 9764 -5368
rect 8592 -5448 9764 -5432
rect 8592 -5512 9680 -5448
rect 9744 -5512 9764 -5448
rect 8592 -5528 9764 -5512
rect 8592 -5592 9680 -5528
rect 9744 -5592 9764 -5528
rect 8592 -5608 9764 -5592
rect 8592 -5672 9680 -5608
rect 9744 -5672 9764 -5608
rect 8592 -5688 9764 -5672
rect 8592 -5752 9680 -5688
rect 9744 -5752 9764 -5688
rect 8592 -5768 9764 -5752
rect 8592 -5832 9680 -5768
rect 9744 -5832 9764 -5768
rect 8592 -5848 9764 -5832
rect 8592 -5912 9680 -5848
rect 9744 -5912 9764 -5848
rect 8592 -5928 9764 -5912
rect 8592 -5992 9680 -5928
rect 9744 -5992 9764 -5928
rect 8592 -6040 9764 -5992
rect 10004 -5208 11176 -5160
rect 10004 -5272 11092 -5208
rect 11156 -5272 11176 -5208
rect 10004 -5288 11176 -5272
rect 10004 -5352 11092 -5288
rect 11156 -5352 11176 -5288
rect 10004 -5368 11176 -5352
rect 10004 -5432 11092 -5368
rect 11156 -5432 11176 -5368
rect 10004 -5448 11176 -5432
rect 10004 -5512 11092 -5448
rect 11156 -5512 11176 -5448
rect 10004 -5528 11176 -5512
rect 10004 -5592 11092 -5528
rect 11156 -5592 11176 -5528
rect 10004 -5608 11176 -5592
rect 10004 -5672 11092 -5608
rect 11156 -5672 11176 -5608
rect 10004 -5688 11176 -5672
rect 10004 -5752 11092 -5688
rect 11156 -5752 11176 -5688
rect 10004 -5768 11176 -5752
rect 10004 -5832 11092 -5768
rect 11156 -5832 11176 -5768
rect 10004 -5848 11176 -5832
rect 10004 -5912 11092 -5848
rect 11156 -5912 11176 -5848
rect 10004 -5928 11176 -5912
rect 10004 -5992 11092 -5928
rect 11156 -5992 11176 -5928
rect 10004 -6040 11176 -5992
rect 11416 -5208 12588 -5160
rect 11416 -5272 12504 -5208
rect 12568 -5272 12588 -5208
rect 11416 -5288 12588 -5272
rect 11416 -5352 12504 -5288
rect 12568 -5352 12588 -5288
rect 11416 -5368 12588 -5352
rect 11416 -5432 12504 -5368
rect 12568 -5432 12588 -5368
rect 11416 -5448 12588 -5432
rect 11416 -5512 12504 -5448
rect 12568 -5512 12588 -5448
rect 11416 -5528 12588 -5512
rect 11416 -5592 12504 -5528
rect 12568 -5592 12588 -5528
rect 11416 -5608 12588 -5592
rect 11416 -5672 12504 -5608
rect 12568 -5672 12588 -5608
rect 11416 -5688 12588 -5672
rect 11416 -5752 12504 -5688
rect 12568 -5752 12588 -5688
rect 11416 -5768 12588 -5752
rect 11416 -5832 12504 -5768
rect 12568 -5832 12588 -5768
rect 11416 -5848 12588 -5832
rect 11416 -5912 12504 -5848
rect 12568 -5912 12588 -5848
rect 11416 -5928 12588 -5912
rect 11416 -5992 12504 -5928
rect 12568 -5992 12588 -5928
rect 11416 -6040 12588 -5992
rect 12828 -5208 14000 -5160
rect 12828 -5272 13916 -5208
rect 13980 -5272 14000 -5208
rect 12828 -5288 14000 -5272
rect 12828 -5352 13916 -5288
rect 13980 -5352 14000 -5288
rect 12828 -5368 14000 -5352
rect 12828 -5432 13916 -5368
rect 13980 -5432 14000 -5368
rect 12828 -5448 14000 -5432
rect 12828 -5512 13916 -5448
rect 13980 -5512 14000 -5448
rect 12828 -5528 14000 -5512
rect 12828 -5592 13916 -5528
rect 13980 -5592 14000 -5528
rect 12828 -5608 14000 -5592
rect 12828 -5672 13916 -5608
rect 13980 -5672 14000 -5608
rect 12828 -5688 14000 -5672
rect 12828 -5752 13916 -5688
rect 13980 -5752 14000 -5688
rect 12828 -5768 14000 -5752
rect 12828 -5832 13916 -5768
rect 13980 -5832 14000 -5768
rect 12828 -5848 14000 -5832
rect 12828 -5912 13916 -5848
rect 13980 -5912 14000 -5848
rect 12828 -5928 14000 -5912
rect 12828 -5992 13916 -5928
rect 13980 -5992 14000 -5928
rect 12828 -6040 14000 -5992
rect 14240 -5208 15412 -5160
rect 14240 -5272 15328 -5208
rect 15392 -5272 15412 -5208
rect 14240 -5288 15412 -5272
rect 14240 -5352 15328 -5288
rect 15392 -5352 15412 -5288
rect 14240 -5368 15412 -5352
rect 14240 -5432 15328 -5368
rect 15392 -5432 15412 -5368
rect 14240 -5448 15412 -5432
rect 14240 -5512 15328 -5448
rect 15392 -5512 15412 -5448
rect 14240 -5528 15412 -5512
rect 14240 -5592 15328 -5528
rect 15392 -5592 15412 -5528
rect 14240 -5608 15412 -5592
rect 14240 -5672 15328 -5608
rect 15392 -5672 15412 -5608
rect 14240 -5688 15412 -5672
rect 14240 -5752 15328 -5688
rect 15392 -5752 15412 -5688
rect 14240 -5768 15412 -5752
rect 14240 -5832 15328 -5768
rect 15392 -5832 15412 -5768
rect 14240 -5848 15412 -5832
rect 14240 -5912 15328 -5848
rect 15392 -5912 15412 -5848
rect 14240 -5928 15412 -5912
rect 14240 -5992 15328 -5928
rect 15392 -5992 15412 -5928
rect 14240 -6040 15412 -5992
rect 15652 -5208 16824 -5160
rect 15652 -5272 16740 -5208
rect 16804 -5272 16824 -5208
rect 15652 -5288 16824 -5272
rect 15652 -5352 16740 -5288
rect 16804 -5352 16824 -5288
rect 15652 -5368 16824 -5352
rect 15652 -5432 16740 -5368
rect 16804 -5432 16824 -5368
rect 15652 -5448 16824 -5432
rect 15652 -5512 16740 -5448
rect 16804 -5512 16824 -5448
rect 15652 -5528 16824 -5512
rect 15652 -5592 16740 -5528
rect 16804 -5592 16824 -5528
rect 15652 -5608 16824 -5592
rect 15652 -5672 16740 -5608
rect 16804 -5672 16824 -5608
rect 15652 -5688 16824 -5672
rect 15652 -5752 16740 -5688
rect 16804 -5752 16824 -5688
rect 15652 -5768 16824 -5752
rect 15652 -5832 16740 -5768
rect 16804 -5832 16824 -5768
rect 15652 -5848 16824 -5832
rect 15652 -5912 16740 -5848
rect 16804 -5912 16824 -5848
rect 15652 -5928 16824 -5912
rect 15652 -5992 16740 -5928
rect 16804 -5992 16824 -5928
rect 15652 -6040 16824 -5992
rect 17064 -5208 18236 -5160
rect 17064 -5272 18152 -5208
rect 18216 -5272 18236 -5208
rect 17064 -5288 18236 -5272
rect 17064 -5352 18152 -5288
rect 18216 -5352 18236 -5288
rect 17064 -5368 18236 -5352
rect 17064 -5432 18152 -5368
rect 18216 -5432 18236 -5368
rect 17064 -5448 18236 -5432
rect 17064 -5512 18152 -5448
rect 18216 -5512 18236 -5448
rect 17064 -5528 18236 -5512
rect 17064 -5592 18152 -5528
rect 18216 -5592 18236 -5528
rect 17064 -5608 18236 -5592
rect 17064 -5672 18152 -5608
rect 18216 -5672 18236 -5608
rect 17064 -5688 18236 -5672
rect 17064 -5752 18152 -5688
rect 18216 -5752 18236 -5688
rect 17064 -5768 18236 -5752
rect 17064 -5832 18152 -5768
rect 18216 -5832 18236 -5768
rect 17064 -5848 18236 -5832
rect 17064 -5912 18152 -5848
rect 18216 -5912 18236 -5848
rect 17064 -5928 18236 -5912
rect 17064 -5992 18152 -5928
rect 18216 -5992 18236 -5928
rect 17064 -6040 18236 -5992
rect 18476 -5208 19648 -5160
rect 18476 -5272 19564 -5208
rect 19628 -5272 19648 -5208
rect 18476 -5288 19648 -5272
rect 18476 -5352 19564 -5288
rect 19628 -5352 19648 -5288
rect 18476 -5368 19648 -5352
rect 18476 -5432 19564 -5368
rect 19628 -5432 19648 -5368
rect 18476 -5448 19648 -5432
rect 18476 -5512 19564 -5448
rect 19628 -5512 19648 -5448
rect 18476 -5528 19648 -5512
rect 18476 -5592 19564 -5528
rect 19628 -5592 19648 -5528
rect 18476 -5608 19648 -5592
rect 18476 -5672 19564 -5608
rect 19628 -5672 19648 -5608
rect 18476 -5688 19648 -5672
rect 18476 -5752 19564 -5688
rect 19628 -5752 19648 -5688
rect 18476 -5768 19648 -5752
rect 18476 -5832 19564 -5768
rect 19628 -5832 19648 -5768
rect 18476 -5848 19648 -5832
rect 18476 -5912 19564 -5848
rect 19628 -5912 19648 -5848
rect 18476 -5928 19648 -5912
rect 18476 -5992 19564 -5928
rect 19628 -5992 19648 -5928
rect 18476 -6040 19648 -5992
rect 19888 -5208 21060 -5160
rect 19888 -5272 20976 -5208
rect 21040 -5272 21060 -5208
rect 19888 -5288 21060 -5272
rect 19888 -5352 20976 -5288
rect 21040 -5352 21060 -5288
rect 19888 -5368 21060 -5352
rect 19888 -5432 20976 -5368
rect 21040 -5432 21060 -5368
rect 19888 -5448 21060 -5432
rect 19888 -5512 20976 -5448
rect 21040 -5512 21060 -5448
rect 19888 -5528 21060 -5512
rect 19888 -5592 20976 -5528
rect 21040 -5592 21060 -5528
rect 19888 -5608 21060 -5592
rect 19888 -5672 20976 -5608
rect 21040 -5672 21060 -5608
rect 19888 -5688 21060 -5672
rect 19888 -5752 20976 -5688
rect 21040 -5752 21060 -5688
rect 19888 -5768 21060 -5752
rect 19888 -5832 20976 -5768
rect 21040 -5832 21060 -5768
rect 19888 -5848 21060 -5832
rect 19888 -5912 20976 -5848
rect 21040 -5912 21060 -5848
rect 19888 -5928 21060 -5912
rect 19888 -5992 20976 -5928
rect 21040 -5992 21060 -5928
rect 19888 -6040 21060 -5992
rect 21300 -5208 22472 -5160
rect 21300 -5272 22388 -5208
rect 22452 -5272 22472 -5208
rect 21300 -5288 22472 -5272
rect 21300 -5352 22388 -5288
rect 22452 -5352 22472 -5288
rect 21300 -5368 22472 -5352
rect 21300 -5432 22388 -5368
rect 22452 -5432 22472 -5368
rect 21300 -5448 22472 -5432
rect 21300 -5512 22388 -5448
rect 22452 -5512 22472 -5448
rect 21300 -5528 22472 -5512
rect 21300 -5592 22388 -5528
rect 22452 -5592 22472 -5528
rect 21300 -5608 22472 -5592
rect 21300 -5672 22388 -5608
rect 22452 -5672 22472 -5608
rect 21300 -5688 22472 -5672
rect 21300 -5752 22388 -5688
rect 22452 -5752 22472 -5688
rect 21300 -5768 22472 -5752
rect 21300 -5832 22388 -5768
rect 22452 -5832 22472 -5768
rect 21300 -5848 22472 -5832
rect 21300 -5912 22388 -5848
rect 22452 -5912 22472 -5848
rect 21300 -5928 22472 -5912
rect 21300 -5992 22388 -5928
rect 22452 -5992 22472 -5928
rect 21300 -6040 22472 -5992
rect 22712 -5208 23884 -5160
rect 22712 -5272 23800 -5208
rect 23864 -5272 23884 -5208
rect 22712 -5288 23884 -5272
rect 22712 -5352 23800 -5288
rect 23864 -5352 23884 -5288
rect 22712 -5368 23884 -5352
rect 22712 -5432 23800 -5368
rect 23864 -5432 23884 -5368
rect 22712 -5448 23884 -5432
rect 22712 -5512 23800 -5448
rect 23864 -5512 23884 -5448
rect 22712 -5528 23884 -5512
rect 22712 -5592 23800 -5528
rect 23864 -5592 23884 -5528
rect 22712 -5608 23884 -5592
rect 22712 -5672 23800 -5608
rect 23864 -5672 23884 -5608
rect 22712 -5688 23884 -5672
rect 22712 -5752 23800 -5688
rect 23864 -5752 23884 -5688
rect 22712 -5768 23884 -5752
rect 22712 -5832 23800 -5768
rect 23864 -5832 23884 -5768
rect 22712 -5848 23884 -5832
rect 22712 -5912 23800 -5848
rect 23864 -5912 23884 -5848
rect 22712 -5928 23884 -5912
rect 22712 -5992 23800 -5928
rect 23864 -5992 23884 -5928
rect 22712 -6040 23884 -5992
rect -23884 -6328 -22712 -6280
rect -23884 -6392 -22796 -6328
rect -22732 -6392 -22712 -6328
rect -23884 -6408 -22712 -6392
rect -23884 -6472 -22796 -6408
rect -22732 -6472 -22712 -6408
rect -23884 -6488 -22712 -6472
rect -23884 -6552 -22796 -6488
rect -22732 -6552 -22712 -6488
rect -23884 -6568 -22712 -6552
rect -23884 -6632 -22796 -6568
rect -22732 -6632 -22712 -6568
rect -23884 -6648 -22712 -6632
rect -23884 -6712 -22796 -6648
rect -22732 -6712 -22712 -6648
rect -23884 -6728 -22712 -6712
rect -23884 -6792 -22796 -6728
rect -22732 -6792 -22712 -6728
rect -23884 -6808 -22712 -6792
rect -23884 -6872 -22796 -6808
rect -22732 -6872 -22712 -6808
rect -23884 -6888 -22712 -6872
rect -23884 -6952 -22796 -6888
rect -22732 -6952 -22712 -6888
rect -23884 -6968 -22712 -6952
rect -23884 -7032 -22796 -6968
rect -22732 -7032 -22712 -6968
rect -23884 -7048 -22712 -7032
rect -23884 -7112 -22796 -7048
rect -22732 -7112 -22712 -7048
rect -23884 -7160 -22712 -7112
rect -22472 -6328 -21300 -6280
rect -22472 -6392 -21384 -6328
rect -21320 -6392 -21300 -6328
rect -22472 -6408 -21300 -6392
rect -22472 -6472 -21384 -6408
rect -21320 -6472 -21300 -6408
rect -22472 -6488 -21300 -6472
rect -22472 -6552 -21384 -6488
rect -21320 -6552 -21300 -6488
rect -22472 -6568 -21300 -6552
rect -22472 -6632 -21384 -6568
rect -21320 -6632 -21300 -6568
rect -22472 -6648 -21300 -6632
rect -22472 -6712 -21384 -6648
rect -21320 -6712 -21300 -6648
rect -22472 -6728 -21300 -6712
rect -22472 -6792 -21384 -6728
rect -21320 -6792 -21300 -6728
rect -22472 -6808 -21300 -6792
rect -22472 -6872 -21384 -6808
rect -21320 -6872 -21300 -6808
rect -22472 -6888 -21300 -6872
rect -22472 -6952 -21384 -6888
rect -21320 -6952 -21300 -6888
rect -22472 -6968 -21300 -6952
rect -22472 -7032 -21384 -6968
rect -21320 -7032 -21300 -6968
rect -22472 -7048 -21300 -7032
rect -22472 -7112 -21384 -7048
rect -21320 -7112 -21300 -7048
rect -22472 -7160 -21300 -7112
rect -21060 -6328 -19888 -6280
rect -21060 -6392 -19972 -6328
rect -19908 -6392 -19888 -6328
rect -21060 -6408 -19888 -6392
rect -21060 -6472 -19972 -6408
rect -19908 -6472 -19888 -6408
rect -21060 -6488 -19888 -6472
rect -21060 -6552 -19972 -6488
rect -19908 -6552 -19888 -6488
rect -21060 -6568 -19888 -6552
rect -21060 -6632 -19972 -6568
rect -19908 -6632 -19888 -6568
rect -21060 -6648 -19888 -6632
rect -21060 -6712 -19972 -6648
rect -19908 -6712 -19888 -6648
rect -21060 -6728 -19888 -6712
rect -21060 -6792 -19972 -6728
rect -19908 -6792 -19888 -6728
rect -21060 -6808 -19888 -6792
rect -21060 -6872 -19972 -6808
rect -19908 -6872 -19888 -6808
rect -21060 -6888 -19888 -6872
rect -21060 -6952 -19972 -6888
rect -19908 -6952 -19888 -6888
rect -21060 -6968 -19888 -6952
rect -21060 -7032 -19972 -6968
rect -19908 -7032 -19888 -6968
rect -21060 -7048 -19888 -7032
rect -21060 -7112 -19972 -7048
rect -19908 -7112 -19888 -7048
rect -21060 -7160 -19888 -7112
rect -19648 -6328 -18476 -6280
rect -19648 -6392 -18560 -6328
rect -18496 -6392 -18476 -6328
rect -19648 -6408 -18476 -6392
rect -19648 -6472 -18560 -6408
rect -18496 -6472 -18476 -6408
rect -19648 -6488 -18476 -6472
rect -19648 -6552 -18560 -6488
rect -18496 -6552 -18476 -6488
rect -19648 -6568 -18476 -6552
rect -19648 -6632 -18560 -6568
rect -18496 -6632 -18476 -6568
rect -19648 -6648 -18476 -6632
rect -19648 -6712 -18560 -6648
rect -18496 -6712 -18476 -6648
rect -19648 -6728 -18476 -6712
rect -19648 -6792 -18560 -6728
rect -18496 -6792 -18476 -6728
rect -19648 -6808 -18476 -6792
rect -19648 -6872 -18560 -6808
rect -18496 -6872 -18476 -6808
rect -19648 -6888 -18476 -6872
rect -19648 -6952 -18560 -6888
rect -18496 -6952 -18476 -6888
rect -19648 -6968 -18476 -6952
rect -19648 -7032 -18560 -6968
rect -18496 -7032 -18476 -6968
rect -19648 -7048 -18476 -7032
rect -19648 -7112 -18560 -7048
rect -18496 -7112 -18476 -7048
rect -19648 -7160 -18476 -7112
rect -18236 -6328 -17064 -6280
rect -18236 -6392 -17148 -6328
rect -17084 -6392 -17064 -6328
rect -18236 -6408 -17064 -6392
rect -18236 -6472 -17148 -6408
rect -17084 -6472 -17064 -6408
rect -18236 -6488 -17064 -6472
rect -18236 -6552 -17148 -6488
rect -17084 -6552 -17064 -6488
rect -18236 -6568 -17064 -6552
rect -18236 -6632 -17148 -6568
rect -17084 -6632 -17064 -6568
rect -18236 -6648 -17064 -6632
rect -18236 -6712 -17148 -6648
rect -17084 -6712 -17064 -6648
rect -18236 -6728 -17064 -6712
rect -18236 -6792 -17148 -6728
rect -17084 -6792 -17064 -6728
rect -18236 -6808 -17064 -6792
rect -18236 -6872 -17148 -6808
rect -17084 -6872 -17064 -6808
rect -18236 -6888 -17064 -6872
rect -18236 -6952 -17148 -6888
rect -17084 -6952 -17064 -6888
rect -18236 -6968 -17064 -6952
rect -18236 -7032 -17148 -6968
rect -17084 -7032 -17064 -6968
rect -18236 -7048 -17064 -7032
rect -18236 -7112 -17148 -7048
rect -17084 -7112 -17064 -7048
rect -18236 -7160 -17064 -7112
rect -16824 -6328 -15652 -6280
rect -16824 -6392 -15736 -6328
rect -15672 -6392 -15652 -6328
rect -16824 -6408 -15652 -6392
rect -16824 -6472 -15736 -6408
rect -15672 -6472 -15652 -6408
rect -16824 -6488 -15652 -6472
rect -16824 -6552 -15736 -6488
rect -15672 -6552 -15652 -6488
rect -16824 -6568 -15652 -6552
rect -16824 -6632 -15736 -6568
rect -15672 -6632 -15652 -6568
rect -16824 -6648 -15652 -6632
rect -16824 -6712 -15736 -6648
rect -15672 -6712 -15652 -6648
rect -16824 -6728 -15652 -6712
rect -16824 -6792 -15736 -6728
rect -15672 -6792 -15652 -6728
rect -16824 -6808 -15652 -6792
rect -16824 -6872 -15736 -6808
rect -15672 -6872 -15652 -6808
rect -16824 -6888 -15652 -6872
rect -16824 -6952 -15736 -6888
rect -15672 -6952 -15652 -6888
rect -16824 -6968 -15652 -6952
rect -16824 -7032 -15736 -6968
rect -15672 -7032 -15652 -6968
rect -16824 -7048 -15652 -7032
rect -16824 -7112 -15736 -7048
rect -15672 -7112 -15652 -7048
rect -16824 -7160 -15652 -7112
rect -15412 -6328 -14240 -6280
rect -15412 -6392 -14324 -6328
rect -14260 -6392 -14240 -6328
rect -15412 -6408 -14240 -6392
rect -15412 -6472 -14324 -6408
rect -14260 -6472 -14240 -6408
rect -15412 -6488 -14240 -6472
rect -15412 -6552 -14324 -6488
rect -14260 -6552 -14240 -6488
rect -15412 -6568 -14240 -6552
rect -15412 -6632 -14324 -6568
rect -14260 -6632 -14240 -6568
rect -15412 -6648 -14240 -6632
rect -15412 -6712 -14324 -6648
rect -14260 -6712 -14240 -6648
rect -15412 -6728 -14240 -6712
rect -15412 -6792 -14324 -6728
rect -14260 -6792 -14240 -6728
rect -15412 -6808 -14240 -6792
rect -15412 -6872 -14324 -6808
rect -14260 -6872 -14240 -6808
rect -15412 -6888 -14240 -6872
rect -15412 -6952 -14324 -6888
rect -14260 -6952 -14240 -6888
rect -15412 -6968 -14240 -6952
rect -15412 -7032 -14324 -6968
rect -14260 -7032 -14240 -6968
rect -15412 -7048 -14240 -7032
rect -15412 -7112 -14324 -7048
rect -14260 -7112 -14240 -7048
rect -15412 -7160 -14240 -7112
rect -14000 -6328 -12828 -6280
rect -14000 -6392 -12912 -6328
rect -12848 -6392 -12828 -6328
rect -14000 -6408 -12828 -6392
rect -14000 -6472 -12912 -6408
rect -12848 -6472 -12828 -6408
rect -14000 -6488 -12828 -6472
rect -14000 -6552 -12912 -6488
rect -12848 -6552 -12828 -6488
rect -14000 -6568 -12828 -6552
rect -14000 -6632 -12912 -6568
rect -12848 -6632 -12828 -6568
rect -14000 -6648 -12828 -6632
rect -14000 -6712 -12912 -6648
rect -12848 -6712 -12828 -6648
rect -14000 -6728 -12828 -6712
rect -14000 -6792 -12912 -6728
rect -12848 -6792 -12828 -6728
rect -14000 -6808 -12828 -6792
rect -14000 -6872 -12912 -6808
rect -12848 -6872 -12828 -6808
rect -14000 -6888 -12828 -6872
rect -14000 -6952 -12912 -6888
rect -12848 -6952 -12828 -6888
rect -14000 -6968 -12828 -6952
rect -14000 -7032 -12912 -6968
rect -12848 -7032 -12828 -6968
rect -14000 -7048 -12828 -7032
rect -14000 -7112 -12912 -7048
rect -12848 -7112 -12828 -7048
rect -14000 -7160 -12828 -7112
rect -12588 -6328 -11416 -6280
rect -12588 -6392 -11500 -6328
rect -11436 -6392 -11416 -6328
rect -12588 -6408 -11416 -6392
rect -12588 -6472 -11500 -6408
rect -11436 -6472 -11416 -6408
rect -12588 -6488 -11416 -6472
rect -12588 -6552 -11500 -6488
rect -11436 -6552 -11416 -6488
rect -12588 -6568 -11416 -6552
rect -12588 -6632 -11500 -6568
rect -11436 -6632 -11416 -6568
rect -12588 -6648 -11416 -6632
rect -12588 -6712 -11500 -6648
rect -11436 -6712 -11416 -6648
rect -12588 -6728 -11416 -6712
rect -12588 -6792 -11500 -6728
rect -11436 -6792 -11416 -6728
rect -12588 -6808 -11416 -6792
rect -12588 -6872 -11500 -6808
rect -11436 -6872 -11416 -6808
rect -12588 -6888 -11416 -6872
rect -12588 -6952 -11500 -6888
rect -11436 -6952 -11416 -6888
rect -12588 -6968 -11416 -6952
rect -12588 -7032 -11500 -6968
rect -11436 -7032 -11416 -6968
rect -12588 -7048 -11416 -7032
rect -12588 -7112 -11500 -7048
rect -11436 -7112 -11416 -7048
rect -12588 -7160 -11416 -7112
rect -11176 -6328 -10004 -6280
rect -11176 -6392 -10088 -6328
rect -10024 -6392 -10004 -6328
rect -11176 -6408 -10004 -6392
rect -11176 -6472 -10088 -6408
rect -10024 -6472 -10004 -6408
rect -11176 -6488 -10004 -6472
rect -11176 -6552 -10088 -6488
rect -10024 -6552 -10004 -6488
rect -11176 -6568 -10004 -6552
rect -11176 -6632 -10088 -6568
rect -10024 -6632 -10004 -6568
rect -11176 -6648 -10004 -6632
rect -11176 -6712 -10088 -6648
rect -10024 -6712 -10004 -6648
rect -11176 -6728 -10004 -6712
rect -11176 -6792 -10088 -6728
rect -10024 -6792 -10004 -6728
rect -11176 -6808 -10004 -6792
rect -11176 -6872 -10088 -6808
rect -10024 -6872 -10004 -6808
rect -11176 -6888 -10004 -6872
rect -11176 -6952 -10088 -6888
rect -10024 -6952 -10004 -6888
rect -11176 -6968 -10004 -6952
rect -11176 -7032 -10088 -6968
rect -10024 -7032 -10004 -6968
rect -11176 -7048 -10004 -7032
rect -11176 -7112 -10088 -7048
rect -10024 -7112 -10004 -7048
rect -11176 -7160 -10004 -7112
rect -9764 -6328 -8592 -6280
rect -9764 -6392 -8676 -6328
rect -8612 -6392 -8592 -6328
rect -9764 -6408 -8592 -6392
rect -9764 -6472 -8676 -6408
rect -8612 -6472 -8592 -6408
rect -9764 -6488 -8592 -6472
rect -9764 -6552 -8676 -6488
rect -8612 -6552 -8592 -6488
rect -9764 -6568 -8592 -6552
rect -9764 -6632 -8676 -6568
rect -8612 -6632 -8592 -6568
rect -9764 -6648 -8592 -6632
rect -9764 -6712 -8676 -6648
rect -8612 -6712 -8592 -6648
rect -9764 -6728 -8592 -6712
rect -9764 -6792 -8676 -6728
rect -8612 -6792 -8592 -6728
rect -9764 -6808 -8592 -6792
rect -9764 -6872 -8676 -6808
rect -8612 -6872 -8592 -6808
rect -9764 -6888 -8592 -6872
rect -9764 -6952 -8676 -6888
rect -8612 -6952 -8592 -6888
rect -9764 -6968 -8592 -6952
rect -9764 -7032 -8676 -6968
rect -8612 -7032 -8592 -6968
rect -9764 -7048 -8592 -7032
rect -9764 -7112 -8676 -7048
rect -8612 -7112 -8592 -7048
rect -9764 -7160 -8592 -7112
rect -8352 -6328 -7180 -6280
rect -8352 -6392 -7264 -6328
rect -7200 -6392 -7180 -6328
rect -8352 -6408 -7180 -6392
rect -8352 -6472 -7264 -6408
rect -7200 -6472 -7180 -6408
rect -8352 -6488 -7180 -6472
rect -8352 -6552 -7264 -6488
rect -7200 -6552 -7180 -6488
rect -8352 -6568 -7180 -6552
rect -8352 -6632 -7264 -6568
rect -7200 -6632 -7180 -6568
rect -8352 -6648 -7180 -6632
rect -8352 -6712 -7264 -6648
rect -7200 -6712 -7180 -6648
rect -8352 -6728 -7180 -6712
rect -8352 -6792 -7264 -6728
rect -7200 -6792 -7180 -6728
rect -8352 -6808 -7180 -6792
rect -8352 -6872 -7264 -6808
rect -7200 -6872 -7180 -6808
rect -8352 -6888 -7180 -6872
rect -8352 -6952 -7264 -6888
rect -7200 -6952 -7180 -6888
rect -8352 -6968 -7180 -6952
rect -8352 -7032 -7264 -6968
rect -7200 -7032 -7180 -6968
rect -8352 -7048 -7180 -7032
rect -8352 -7112 -7264 -7048
rect -7200 -7112 -7180 -7048
rect -8352 -7160 -7180 -7112
rect -6940 -6328 -5768 -6280
rect -6940 -6392 -5852 -6328
rect -5788 -6392 -5768 -6328
rect -6940 -6408 -5768 -6392
rect -6940 -6472 -5852 -6408
rect -5788 -6472 -5768 -6408
rect -6940 -6488 -5768 -6472
rect -6940 -6552 -5852 -6488
rect -5788 -6552 -5768 -6488
rect -6940 -6568 -5768 -6552
rect -6940 -6632 -5852 -6568
rect -5788 -6632 -5768 -6568
rect -6940 -6648 -5768 -6632
rect -6940 -6712 -5852 -6648
rect -5788 -6712 -5768 -6648
rect -6940 -6728 -5768 -6712
rect -6940 -6792 -5852 -6728
rect -5788 -6792 -5768 -6728
rect -6940 -6808 -5768 -6792
rect -6940 -6872 -5852 -6808
rect -5788 -6872 -5768 -6808
rect -6940 -6888 -5768 -6872
rect -6940 -6952 -5852 -6888
rect -5788 -6952 -5768 -6888
rect -6940 -6968 -5768 -6952
rect -6940 -7032 -5852 -6968
rect -5788 -7032 -5768 -6968
rect -6940 -7048 -5768 -7032
rect -6940 -7112 -5852 -7048
rect -5788 -7112 -5768 -7048
rect -6940 -7160 -5768 -7112
rect -5528 -6328 -4356 -6280
rect -5528 -6392 -4440 -6328
rect -4376 -6392 -4356 -6328
rect -5528 -6408 -4356 -6392
rect -5528 -6472 -4440 -6408
rect -4376 -6472 -4356 -6408
rect -5528 -6488 -4356 -6472
rect -5528 -6552 -4440 -6488
rect -4376 -6552 -4356 -6488
rect -5528 -6568 -4356 -6552
rect -5528 -6632 -4440 -6568
rect -4376 -6632 -4356 -6568
rect -5528 -6648 -4356 -6632
rect -5528 -6712 -4440 -6648
rect -4376 -6712 -4356 -6648
rect -5528 -6728 -4356 -6712
rect -5528 -6792 -4440 -6728
rect -4376 -6792 -4356 -6728
rect -5528 -6808 -4356 -6792
rect -5528 -6872 -4440 -6808
rect -4376 -6872 -4356 -6808
rect -5528 -6888 -4356 -6872
rect -5528 -6952 -4440 -6888
rect -4376 -6952 -4356 -6888
rect -5528 -6968 -4356 -6952
rect -5528 -7032 -4440 -6968
rect -4376 -7032 -4356 -6968
rect -5528 -7048 -4356 -7032
rect -5528 -7112 -4440 -7048
rect -4376 -7112 -4356 -7048
rect -5528 -7160 -4356 -7112
rect -4116 -6328 -2944 -6280
rect -4116 -6392 -3028 -6328
rect -2964 -6392 -2944 -6328
rect -4116 -6408 -2944 -6392
rect -4116 -6472 -3028 -6408
rect -2964 -6472 -2944 -6408
rect -4116 -6488 -2944 -6472
rect -4116 -6552 -3028 -6488
rect -2964 -6552 -2944 -6488
rect -4116 -6568 -2944 -6552
rect -4116 -6632 -3028 -6568
rect -2964 -6632 -2944 -6568
rect -4116 -6648 -2944 -6632
rect -4116 -6712 -3028 -6648
rect -2964 -6712 -2944 -6648
rect -4116 -6728 -2944 -6712
rect -4116 -6792 -3028 -6728
rect -2964 -6792 -2944 -6728
rect -4116 -6808 -2944 -6792
rect -4116 -6872 -3028 -6808
rect -2964 -6872 -2944 -6808
rect -4116 -6888 -2944 -6872
rect -4116 -6952 -3028 -6888
rect -2964 -6952 -2944 -6888
rect -4116 -6968 -2944 -6952
rect -4116 -7032 -3028 -6968
rect -2964 -7032 -2944 -6968
rect -4116 -7048 -2944 -7032
rect -4116 -7112 -3028 -7048
rect -2964 -7112 -2944 -7048
rect -4116 -7160 -2944 -7112
rect -2704 -6328 -1532 -6280
rect -2704 -6392 -1616 -6328
rect -1552 -6392 -1532 -6328
rect -2704 -6408 -1532 -6392
rect -2704 -6472 -1616 -6408
rect -1552 -6472 -1532 -6408
rect -2704 -6488 -1532 -6472
rect -2704 -6552 -1616 -6488
rect -1552 -6552 -1532 -6488
rect -2704 -6568 -1532 -6552
rect -2704 -6632 -1616 -6568
rect -1552 -6632 -1532 -6568
rect -2704 -6648 -1532 -6632
rect -2704 -6712 -1616 -6648
rect -1552 -6712 -1532 -6648
rect -2704 -6728 -1532 -6712
rect -2704 -6792 -1616 -6728
rect -1552 -6792 -1532 -6728
rect -2704 -6808 -1532 -6792
rect -2704 -6872 -1616 -6808
rect -1552 -6872 -1532 -6808
rect -2704 -6888 -1532 -6872
rect -2704 -6952 -1616 -6888
rect -1552 -6952 -1532 -6888
rect -2704 -6968 -1532 -6952
rect -2704 -7032 -1616 -6968
rect -1552 -7032 -1532 -6968
rect -2704 -7048 -1532 -7032
rect -2704 -7112 -1616 -7048
rect -1552 -7112 -1532 -7048
rect -2704 -7160 -1532 -7112
rect -1292 -6328 -120 -6280
rect -1292 -6392 -204 -6328
rect -140 -6392 -120 -6328
rect -1292 -6408 -120 -6392
rect -1292 -6472 -204 -6408
rect -140 -6472 -120 -6408
rect -1292 -6488 -120 -6472
rect -1292 -6552 -204 -6488
rect -140 -6552 -120 -6488
rect -1292 -6568 -120 -6552
rect -1292 -6632 -204 -6568
rect -140 -6632 -120 -6568
rect -1292 -6648 -120 -6632
rect -1292 -6712 -204 -6648
rect -140 -6712 -120 -6648
rect -1292 -6728 -120 -6712
rect -1292 -6792 -204 -6728
rect -140 -6792 -120 -6728
rect -1292 -6808 -120 -6792
rect -1292 -6872 -204 -6808
rect -140 -6872 -120 -6808
rect -1292 -6888 -120 -6872
rect -1292 -6952 -204 -6888
rect -140 -6952 -120 -6888
rect -1292 -6968 -120 -6952
rect -1292 -7032 -204 -6968
rect -140 -7032 -120 -6968
rect -1292 -7048 -120 -7032
rect -1292 -7112 -204 -7048
rect -140 -7112 -120 -7048
rect -1292 -7160 -120 -7112
rect 120 -6328 1292 -6280
rect 120 -6392 1208 -6328
rect 1272 -6392 1292 -6328
rect 120 -6408 1292 -6392
rect 120 -6472 1208 -6408
rect 1272 -6472 1292 -6408
rect 120 -6488 1292 -6472
rect 120 -6552 1208 -6488
rect 1272 -6552 1292 -6488
rect 120 -6568 1292 -6552
rect 120 -6632 1208 -6568
rect 1272 -6632 1292 -6568
rect 120 -6648 1292 -6632
rect 120 -6712 1208 -6648
rect 1272 -6712 1292 -6648
rect 120 -6728 1292 -6712
rect 120 -6792 1208 -6728
rect 1272 -6792 1292 -6728
rect 120 -6808 1292 -6792
rect 120 -6872 1208 -6808
rect 1272 -6872 1292 -6808
rect 120 -6888 1292 -6872
rect 120 -6952 1208 -6888
rect 1272 -6952 1292 -6888
rect 120 -6968 1292 -6952
rect 120 -7032 1208 -6968
rect 1272 -7032 1292 -6968
rect 120 -7048 1292 -7032
rect 120 -7112 1208 -7048
rect 1272 -7112 1292 -7048
rect 120 -7160 1292 -7112
rect 1532 -6328 2704 -6280
rect 1532 -6392 2620 -6328
rect 2684 -6392 2704 -6328
rect 1532 -6408 2704 -6392
rect 1532 -6472 2620 -6408
rect 2684 -6472 2704 -6408
rect 1532 -6488 2704 -6472
rect 1532 -6552 2620 -6488
rect 2684 -6552 2704 -6488
rect 1532 -6568 2704 -6552
rect 1532 -6632 2620 -6568
rect 2684 -6632 2704 -6568
rect 1532 -6648 2704 -6632
rect 1532 -6712 2620 -6648
rect 2684 -6712 2704 -6648
rect 1532 -6728 2704 -6712
rect 1532 -6792 2620 -6728
rect 2684 -6792 2704 -6728
rect 1532 -6808 2704 -6792
rect 1532 -6872 2620 -6808
rect 2684 -6872 2704 -6808
rect 1532 -6888 2704 -6872
rect 1532 -6952 2620 -6888
rect 2684 -6952 2704 -6888
rect 1532 -6968 2704 -6952
rect 1532 -7032 2620 -6968
rect 2684 -7032 2704 -6968
rect 1532 -7048 2704 -7032
rect 1532 -7112 2620 -7048
rect 2684 -7112 2704 -7048
rect 1532 -7160 2704 -7112
rect 2944 -6328 4116 -6280
rect 2944 -6392 4032 -6328
rect 4096 -6392 4116 -6328
rect 2944 -6408 4116 -6392
rect 2944 -6472 4032 -6408
rect 4096 -6472 4116 -6408
rect 2944 -6488 4116 -6472
rect 2944 -6552 4032 -6488
rect 4096 -6552 4116 -6488
rect 2944 -6568 4116 -6552
rect 2944 -6632 4032 -6568
rect 4096 -6632 4116 -6568
rect 2944 -6648 4116 -6632
rect 2944 -6712 4032 -6648
rect 4096 -6712 4116 -6648
rect 2944 -6728 4116 -6712
rect 2944 -6792 4032 -6728
rect 4096 -6792 4116 -6728
rect 2944 -6808 4116 -6792
rect 2944 -6872 4032 -6808
rect 4096 -6872 4116 -6808
rect 2944 -6888 4116 -6872
rect 2944 -6952 4032 -6888
rect 4096 -6952 4116 -6888
rect 2944 -6968 4116 -6952
rect 2944 -7032 4032 -6968
rect 4096 -7032 4116 -6968
rect 2944 -7048 4116 -7032
rect 2944 -7112 4032 -7048
rect 4096 -7112 4116 -7048
rect 2944 -7160 4116 -7112
rect 4356 -6328 5528 -6280
rect 4356 -6392 5444 -6328
rect 5508 -6392 5528 -6328
rect 4356 -6408 5528 -6392
rect 4356 -6472 5444 -6408
rect 5508 -6472 5528 -6408
rect 4356 -6488 5528 -6472
rect 4356 -6552 5444 -6488
rect 5508 -6552 5528 -6488
rect 4356 -6568 5528 -6552
rect 4356 -6632 5444 -6568
rect 5508 -6632 5528 -6568
rect 4356 -6648 5528 -6632
rect 4356 -6712 5444 -6648
rect 5508 -6712 5528 -6648
rect 4356 -6728 5528 -6712
rect 4356 -6792 5444 -6728
rect 5508 -6792 5528 -6728
rect 4356 -6808 5528 -6792
rect 4356 -6872 5444 -6808
rect 5508 -6872 5528 -6808
rect 4356 -6888 5528 -6872
rect 4356 -6952 5444 -6888
rect 5508 -6952 5528 -6888
rect 4356 -6968 5528 -6952
rect 4356 -7032 5444 -6968
rect 5508 -7032 5528 -6968
rect 4356 -7048 5528 -7032
rect 4356 -7112 5444 -7048
rect 5508 -7112 5528 -7048
rect 4356 -7160 5528 -7112
rect 5768 -6328 6940 -6280
rect 5768 -6392 6856 -6328
rect 6920 -6392 6940 -6328
rect 5768 -6408 6940 -6392
rect 5768 -6472 6856 -6408
rect 6920 -6472 6940 -6408
rect 5768 -6488 6940 -6472
rect 5768 -6552 6856 -6488
rect 6920 -6552 6940 -6488
rect 5768 -6568 6940 -6552
rect 5768 -6632 6856 -6568
rect 6920 -6632 6940 -6568
rect 5768 -6648 6940 -6632
rect 5768 -6712 6856 -6648
rect 6920 -6712 6940 -6648
rect 5768 -6728 6940 -6712
rect 5768 -6792 6856 -6728
rect 6920 -6792 6940 -6728
rect 5768 -6808 6940 -6792
rect 5768 -6872 6856 -6808
rect 6920 -6872 6940 -6808
rect 5768 -6888 6940 -6872
rect 5768 -6952 6856 -6888
rect 6920 -6952 6940 -6888
rect 5768 -6968 6940 -6952
rect 5768 -7032 6856 -6968
rect 6920 -7032 6940 -6968
rect 5768 -7048 6940 -7032
rect 5768 -7112 6856 -7048
rect 6920 -7112 6940 -7048
rect 5768 -7160 6940 -7112
rect 7180 -6328 8352 -6280
rect 7180 -6392 8268 -6328
rect 8332 -6392 8352 -6328
rect 7180 -6408 8352 -6392
rect 7180 -6472 8268 -6408
rect 8332 -6472 8352 -6408
rect 7180 -6488 8352 -6472
rect 7180 -6552 8268 -6488
rect 8332 -6552 8352 -6488
rect 7180 -6568 8352 -6552
rect 7180 -6632 8268 -6568
rect 8332 -6632 8352 -6568
rect 7180 -6648 8352 -6632
rect 7180 -6712 8268 -6648
rect 8332 -6712 8352 -6648
rect 7180 -6728 8352 -6712
rect 7180 -6792 8268 -6728
rect 8332 -6792 8352 -6728
rect 7180 -6808 8352 -6792
rect 7180 -6872 8268 -6808
rect 8332 -6872 8352 -6808
rect 7180 -6888 8352 -6872
rect 7180 -6952 8268 -6888
rect 8332 -6952 8352 -6888
rect 7180 -6968 8352 -6952
rect 7180 -7032 8268 -6968
rect 8332 -7032 8352 -6968
rect 7180 -7048 8352 -7032
rect 7180 -7112 8268 -7048
rect 8332 -7112 8352 -7048
rect 7180 -7160 8352 -7112
rect 8592 -6328 9764 -6280
rect 8592 -6392 9680 -6328
rect 9744 -6392 9764 -6328
rect 8592 -6408 9764 -6392
rect 8592 -6472 9680 -6408
rect 9744 -6472 9764 -6408
rect 8592 -6488 9764 -6472
rect 8592 -6552 9680 -6488
rect 9744 -6552 9764 -6488
rect 8592 -6568 9764 -6552
rect 8592 -6632 9680 -6568
rect 9744 -6632 9764 -6568
rect 8592 -6648 9764 -6632
rect 8592 -6712 9680 -6648
rect 9744 -6712 9764 -6648
rect 8592 -6728 9764 -6712
rect 8592 -6792 9680 -6728
rect 9744 -6792 9764 -6728
rect 8592 -6808 9764 -6792
rect 8592 -6872 9680 -6808
rect 9744 -6872 9764 -6808
rect 8592 -6888 9764 -6872
rect 8592 -6952 9680 -6888
rect 9744 -6952 9764 -6888
rect 8592 -6968 9764 -6952
rect 8592 -7032 9680 -6968
rect 9744 -7032 9764 -6968
rect 8592 -7048 9764 -7032
rect 8592 -7112 9680 -7048
rect 9744 -7112 9764 -7048
rect 8592 -7160 9764 -7112
rect 10004 -6328 11176 -6280
rect 10004 -6392 11092 -6328
rect 11156 -6392 11176 -6328
rect 10004 -6408 11176 -6392
rect 10004 -6472 11092 -6408
rect 11156 -6472 11176 -6408
rect 10004 -6488 11176 -6472
rect 10004 -6552 11092 -6488
rect 11156 -6552 11176 -6488
rect 10004 -6568 11176 -6552
rect 10004 -6632 11092 -6568
rect 11156 -6632 11176 -6568
rect 10004 -6648 11176 -6632
rect 10004 -6712 11092 -6648
rect 11156 -6712 11176 -6648
rect 10004 -6728 11176 -6712
rect 10004 -6792 11092 -6728
rect 11156 -6792 11176 -6728
rect 10004 -6808 11176 -6792
rect 10004 -6872 11092 -6808
rect 11156 -6872 11176 -6808
rect 10004 -6888 11176 -6872
rect 10004 -6952 11092 -6888
rect 11156 -6952 11176 -6888
rect 10004 -6968 11176 -6952
rect 10004 -7032 11092 -6968
rect 11156 -7032 11176 -6968
rect 10004 -7048 11176 -7032
rect 10004 -7112 11092 -7048
rect 11156 -7112 11176 -7048
rect 10004 -7160 11176 -7112
rect 11416 -6328 12588 -6280
rect 11416 -6392 12504 -6328
rect 12568 -6392 12588 -6328
rect 11416 -6408 12588 -6392
rect 11416 -6472 12504 -6408
rect 12568 -6472 12588 -6408
rect 11416 -6488 12588 -6472
rect 11416 -6552 12504 -6488
rect 12568 -6552 12588 -6488
rect 11416 -6568 12588 -6552
rect 11416 -6632 12504 -6568
rect 12568 -6632 12588 -6568
rect 11416 -6648 12588 -6632
rect 11416 -6712 12504 -6648
rect 12568 -6712 12588 -6648
rect 11416 -6728 12588 -6712
rect 11416 -6792 12504 -6728
rect 12568 -6792 12588 -6728
rect 11416 -6808 12588 -6792
rect 11416 -6872 12504 -6808
rect 12568 -6872 12588 -6808
rect 11416 -6888 12588 -6872
rect 11416 -6952 12504 -6888
rect 12568 -6952 12588 -6888
rect 11416 -6968 12588 -6952
rect 11416 -7032 12504 -6968
rect 12568 -7032 12588 -6968
rect 11416 -7048 12588 -7032
rect 11416 -7112 12504 -7048
rect 12568 -7112 12588 -7048
rect 11416 -7160 12588 -7112
rect 12828 -6328 14000 -6280
rect 12828 -6392 13916 -6328
rect 13980 -6392 14000 -6328
rect 12828 -6408 14000 -6392
rect 12828 -6472 13916 -6408
rect 13980 -6472 14000 -6408
rect 12828 -6488 14000 -6472
rect 12828 -6552 13916 -6488
rect 13980 -6552 14000 -6488
rect 12828 -6568 14000 -6552
rect 12828 -6632 13916 -6568
rect 13980 -6632 14000 -6568
rect 12828 -6648 14000 -6632
rect 12828 -6712 13916 -6648
rect 13980 -6712 14000 -6648
rect 12828 -6728 14000 -6712
rect 12828 -6792 13916 -6728
rect 13980 -6792 14000 -6728
rect 12828 -6808 14000 -6792
rect 12828 -6872 13916 -6808
rect 13980 -6872 14000 -6808
rect 12828 -6888 14000 -6872
rect 12828 -6952 13916 -6888
rect 13980 -6952 14000 -6888
rect 12828 -6968 14000 -6952
rect 12828 -7032 13916 -6968
rect 13980 -7032 14000 -6968
rect 12828 -7048 14000 -7032
rect 12828 -7112 13916 -7048
rect 13980 -7112 14000 -7048
rect 12828 -7160 14000 -7112
rect 14240 -6328 15412 -6280
rect 14240 -6392 15328 -6328
rect 15392 -6392 15412 -6328
rect 14240 -6408 15412 -6392
rect 14240 -6472 15328 -6408
rect 15392 -6472 15412 -6408
rect 14240 -6488 15412 -6472
rect 14240 -6552 15328 -6488
rect 15392 -6552 15412 -6488
rect 14240 -6568 15412 -6552
rect 14240 -6632 15328 -6568
rect 15392 -6632 15412 -6568
rect 14240 -6648 15412 -6632
rect 14240 -6712 15328 -6648
rect 15392 -6712 15412 -6648
rect 14240 -6728 15412 -6712
rect 14240 -6792 15328 -6728
rect 15392 -6792 15412 -6728
rect 14240 -6808 15412 -6792
rect 14240 -6872 15328 -6808
rect 15392 -6872 15412 -6808
rect 14240 -6888 15412 -6872
rect 14240 -6952 15328 -6888
rect 15392 -6952 15412 -6888
rect 14240 -6968 15412 -6952
rect 14240 -7032 15328 -6968
rect 15392 -7032 15412 -6968
rect 14240 -7048 15412 -7032
rect 14240 -7112 15328 -7048
rect 15392 -7112 15412 -7048
rect 14240 -7160 15412 -7112
rect 15652 -6328 16824 -6280
rect 15652 -6392 16740 -6328
rect 16804 -6392 16824 -6328
rect 15652 -6408 16824 -6392
rect 15652 -6472 16740 -6408
rect 16804 -6472 16824 -6408
rect 15652 -6488 16824 -6472
rect 15652 -6552 16740 -6488
rect 16804 -6552 16824 -6488
rect 15652 -6568 16824 -6552
rect 15652 -6632 16740 -6568
rect 16804 -6632 16824 -6568
rect 15652 -6648 16824 -6632
rect 15652 -6712 16740 -6648
rect 16804 -6712 16824 -6648
rect 15652 -6728 16824 -6712
rect 15652 -6792 16740 -6728
rect 16804 -6792 16824 -6728
rect 15652 -6808 16824 -6792
rect 15652 -6872 16740 -6808
rect 16804 -6872 16824 -6808
rect 15652 -6888 16824 -6872
rect 15652 -6952 16740 -6888
rect 16804 -6952 16824 -6888
rect 15652 -6968 16824 -6952
rect 15652 -7032 16740 -6968
rect 16804 -7032 16824 -6968
rect 15652 -7048 16824 -7032
rect 15652 -7112 16740 -7048
rect 16804 -7112 16824 -7048
rect 15652 -7160 16824 -7112
rect 17064 -6328 18236 -6280
rect 17064 -6392 18152 -6328
rect 18216 -6392 18236 -6328
rect 17064 -6408 18236 -6392
rect 17064 -6472 18152 -6408
rect 18216 -6472 18236 -6408
rect 17064 -6488 18236 -6472
rect 17064 -6552 18152 -6488
rect 18216 -6552 18236 -6488
rect 17064 -6568 18236 -6552
rect 17064 -6632 18152 -6568
rect 18216 -6632 18236 -6568
rect 17064 -6648 18236 -6632
rect 17064 -6712 18152 -6648
rect 18216 -6712 18236 -6648
rect 17064 -6728 18236 -6712
rect 17064 -6792 18152 -6728
rect 18216 -6792 18236 -6728
rect 17064 -6808 18236 -6792
rect 17064 -6872 18152 -6808
rect 18216 -6872 18236 -6808
rect 17064 -6888 18236 -6872
rect 17064 -6952 18152 -6888
rect 18216 -6952 18236 -6888
rect 17064 -6968 18236 -6952
rect 17064 -7032 18152 -6968
rect 18216 -7032 18236 -6968
rect 17064 -7048 18236 -7032
rect 17064 -7112 18152 -7048
rect 18216 -7112 18236 -7048
rect 17064 -7160 18236 -7112
rect 18476 -6328 19648 -6280
rect 18476 -6392 19564 -6328
rect 19628 -6392 19648 -6328
rect 18476 -6408 19648 -6392
rect 18476 -6472 19564 -6408
rect 19628 -6472 19648 -6408
rect 18476 -6488 19648 -6472
rect 18476 -6552 19564 -6488
rect 19628 -6552 19648 -6488
rect 18476 -6568 19648 -6552
rect 18476 -6632 19564 -6568
rect 19628 -6632 19648 -6568
rect 18476 -6648 19648 -6632
rect 18476 -6712 19564 -6648
rect 19628 -6712 19648 -6648
rect 18476 -6728 19648 -6712
rect 18476 -6792 19564 -6728
rect 19628 -6792 19648 -6728
rect 18476 -6808 19648 -6792
rect 18476 -6872 19564 -6808
rect 19628 -6872 19648 -6808
rect 18476 -6888 19648 -6872
rect 18476 -6952 19564 -6888
rect 19628 -6952 19648 -6888
rect 18476 -6968 19648 -6952
rect 18476 -7032 19564 -6968
rect 19628 -7032 19648 -6968
rect 18476 -7048 19648 -7032
rect 18476 -7112 19564 -7048
rect 19628 -7112 19648 -7048
rect 18476 -7160 19648 -7112
rect 19888 -6328 21060 -6280
rect 19888 -6392 20976 -6328
rect 21040 -6392 21060 -6328
rect 19888 -6408 21060 -6392
rect 19888 -6472 20976 -6408
rect 21040 -6472 21060 -6408
rect 19888 -6488 21060 -6472
rect 19888 -6552 20976 -6488
rect 21040 -6552 21060 -6488
rect 19888 -6568 21060 -6552
rect 19888 -6632 20976 -6568
rect 21040 -6632 21060 -6568
rect 19888 -6648 21060 -6632
rect 19888 -6712 20976 -6648
rect 21040 -6712 21060 -6648
rect 19888 -6728 21060 -6712
rect 19888 -6792 20976 -6728
rect 21040 -6792 21060 -6728
rect 19888 -6808 21060 -6792
rect 19888 -6872 20976 -6808
rect 21040 -6872 21060 -6808
rect 19888 -6888 21060 -6872
rect 19888 -6952 20976 -6888
rect 21040 -6952 21060 -6888
rect 19888 -6968 21060 -6952
rect 19888 -7032 20976 -6968
rect 21040 -7032 21060 -6968
rect 19888 -7048 21060 -7032
rect 19888 -7112 20976 -7048
rect 21040 -7112 21060 -7048
rect 19888 -7160 21060 -7112
rect 21300 -6328 22472 -6280
rect 21300 -6392 22388 -6328
rect 22452 -6392 22472 -6328
rect 21300 -6408 22472 -6392
rect 21300 -6472 22388 -6408
rect 22452 -6472 22472 -6408
rect 21300 -6488 22472 -6472
rect 21300 -6552 22388 -6488
rect 22452 -6552 22472 -6488
rect 21300 -6568 22472 -6552
rect 21300 -6632 22388 -6568
rect 22452 -6632 22472 -6568
rect 21300 -6648 22472 -6632
rect 21300 -6712 22388 -6648
rect 22452 -6712 22472 -6648
rect 21300 -6728 22472 -6712
rect 21300 -6792 22388 -6728
rect 22452 -6792 22472 -6728
rect 21300 -6808 22472 -6792
rect 21300 -6872 22388 -6808
rect 22452 -6872 22472 -6808
rect 21300 -6888 22472 -6872
rect 21300 -6952 22388 -6888
rect 22452 -6952 22472 -6888
rect 21300 -6968 22472 -6952
rect 21300 -7032 22388 -6968
rect 22452 -7032 22472 -6968
rect 21300 -7048 22472 -7032
rect 21300 -7112 22388 -7048
rect 22452 -7112 22472 -7048
rect 21300 -7160 22472 -7112
rect 22712 -6328 23884 -6280
rect 22712 -6392 23800 -6328
rect 23864 -6392 23884 -6328
rect 22712 -6408 23884 -6392
rect 22712 -6472 23800 -6408
rect 23864 -6472 23884 -6408
rect 22712 -6488 23884 -6472
rect 22712 -6552 23800 -6488
rect 23864 -6552 23884 -6488
rect 22712 -6568 23884 -6552
rect 22712 -6632 23800 -6568
rect 23864 -6632 23884 -6568
rect 22712 -6648 23884 -6632
rect 22712 -6712 23800 -6648
rect 23864 -6712 23884 -6648
rect 22712 -6728 23884 -6712
rect 22712 -6792 23800 -6728
rect 23864 -6792 23884 -6728
rect 22712 -6808 23884 -6792
rect 22712 -6872 23800 -6808
rect 23864 -6872 23884 -6808
rect 22712 -6888 23884 -6872
rect 22712 -6952 23800 -6888
rect 23864 -6952 23884 -6888
rect 22712 -6968 23884 -6952
rect 22712 -7032 23800 -6968
rect 23864 -7032 23884 -6968
rect 22712 -7048 23884 -7032
rect 22712 -7112 23800 -7048
rect 23864 -7112 23884 -7048
rect 22712 -7160 23884 -7112
rect -23884 -7448 -22712 -7400
rect -23884 -7512 -22796 -7448
rect -22732 -7512 -22712 -7448
rect -23884 -7528 -22712 -7512
rect -23884 -7592 -22796 -7528
rect -22732 -7592 -22712 -7528
rect -23884 -7608 -22712 -7592
rect -23884 -7672 -22796 -7608
rect -22732 -7672 -22712 -7608
rect -23884 -7688 -22712 -7672
rect -23884 -7752 -22796 -7688
rect -22732 -7752 -22712 -7688
rect -23884 -7768 -22712 -7752
rect -23884 -7832 -22796 -7768
rect -22732 -7832 -22712 -7768
rect -23884 -7848 -22712 -7832
rect -23884 -7912 -22796 -7848
rect -22732 -7912 -22712 -7848
rect -23884 -7928 -22712 -7912
rect -23884 -7992 -22796 -7928
rect -22732 -7992 -22712 -7928
rect -23884 -8008 -22712 -7992
rect -23884 -8072 -22796 -8008
rect -22732 -8072 -22712 -8008
rect -23884 -8088 -22712 -8072
rect -23884 -8152 -22796 -8088
rect -22732 -8152 -22712 -8088
rect -23884 -8168 -22712 -8152
rect -23884 -8232 -22796 -8168
rect -22732 -8232 -22712 -8168
rect -23884 -8280 -22712 -8232
rect -22472 -7448 -21300 -7400
rect -22472 -7512 -21384 -7448
rect -21320 -7512 -21300 -7448
rect -22472 -7528 -21300 -7512
rect -22472 -7592 -21384 -7528
rect -21320 -7592 -21300 -7528
rect -22472 -7608 -21300 -7592
rect -22472 -7672 -21384 -7608
rect -21320 -7672 -21300 -7608
rect -22472 -7688 -21300 -7672
rect -22472 -7752 -21384 -7688
rect -21320 -7752 -21300 -7688
rect -22472 -7768 -21300 -7752
rect -22472 -7832 -21384 -7768
rect -21320 -7832 -21300 -7768
rect -22472 -7848 -21300 -7832
rect -22472 -7912 -21384 -7848
rect -21320 -7912 -21300 -7848
rect -22472 -7928 -21300 -7912
rect -22472 -7992 -21384 -7928
rect -21320 -7992 -21300 -7928
rect -22472 -8008 -21300 -7992
rect -22472 -8072 -21384 -8008
rect -21320 -8072 -21300 -8008
rect -22472 -8088 -21300 -8072
rect -22472 -8152 -21384 -8088
rect -21320 -8152 -21300 -8088
rect -22472 -8168 -21300 -8152
rect -22472 -8232 -21384 -8168
rect -21320 -8232 -21300 -8168
rect -22472 -8280 -21300 -8232
rect -21060 -7448 -19888 -7400
rect -21060 -7512 -19972 -7448
rect -19908 -7512 -19888 -7448
rect -21060 -7528 -19888 -7512
rect -21060 -7592 -19972 -7528
rect -19908 -7592 -19888 -7528
rect -21060 -7608 -19888 -7592
rect -21060 -7672 -19972 -7608
rect -19908 -7672 -19888 -7608
rect -21060 -7688 -19888 -7672
rect -21060 -7752 -19972 -7688
rect -19908 -7752 -19888 -7688
rect -21060 -7768 -19888 -7752
rect -21060 -7832 -19972 -7768
rect -19908 -7832 -19888 -7768
rect -21060 -7848 -19888 -7832
rect -21060 -7912 -19972 -7848
rect -19908 -7912 -19888 -7848
rect -21060 -7928 -19888 -7912
rect -21060 -7992 -19972 -7928
rect -19908 -7992 -19888 -7928
rect -21060 -8008 -19888 -7992
rect -21060 -8072 -19972 -8008
rect -19908 -8072 -19888 -8008
rect -21060 -8088 -19888 -8072
rect -21060 -8152 -19972 -8088
rect -19908 -8152 -19888 -8088
rect -21060 -8168 -19888 -8152
rect -21060 -8232 -19972 -8168
rect -19908 -8232 -19888 -8168
rect -21060 -8280 -19888 -8232
rect -19648 -7448 -18476 -7400
rect -19648 -7512 -18560 -7448
rect -18496 -7512 -18476 -7448
rect -19648 -7528 -18476 -7512
rect -19648 -7592 -18560 -7528
rect -18496 -7592 -18476 -7528
rect -19648 -7608 -18476 -7592
rect -19648 -7672 -18560 -7608
rect -18496 -7672 -18476 -7608
rect -19648 -7688 -18476 -7672
rect -19648 -7752 -18560 -7688
rect -18496 -7752 -18476 -7688
rect -19648 -7768 -18476 -7752
rect -19648 -7832 -18560 -7768
rect -18496 -7832 -18476 -7768
rect -19648 -7848 -18476 -7832
rect -19648 -7912 -18560 -7848
rect -18496 -7912 -18476 -7848
rect -19648 -7928 -18476 -7912
rect -19648 -7992 -18560 -7928
rect -18496 -7992 -18476 -7928
rect -19648 -8008 -18476 -7992
rect -19648 -8072 -18560 -8008
rect -18496 -8072 -18476 -8008
rect -19648 -8088 -18476 -8072
rect -19648 -8152 -18560 -8088
rect -18496 -8152 -18476 -8088
rect -19648 -8168 -18476 -8152
rect -19648 -8232 -18560 -8168
rect -18496 -8232 -18476 -8168
rect -19648 -8280 -18476 -8232
rect -18236 -7448 -17064 -7400
rect -18236 -7512 -17148 -7448
rect -17084 -7512 -17064 -7448
rect -18236 -7528 -17064 -7512
rect -18236 -7592 -17148 -7528
rect -17084 -7592 -17064 -7528
rect -18236 -7608 -17064 -7592
rect -18236 -7672 -17148 -7608
rect -17084 -7672 -17064 -7608
rect -18236 -7688 -17064 -7672
rect -18236 -7752 -17148 -7688
rect -17084 -7752 -17064 -7688
rect -18236 -7768 -17064 -7752
rect -18236 -7832 -17148 -7768
rect -17084 -7832 -17064 -7768
rect -18236 -7848 -17064 -7832
rect -18236 -7912 -17148 -7848
rect -17084 -7912 -17064 -7848
rect -18236 -7928 -17064 -7912
rect -18236 -7992 -17148 -7928
rect -17084 -7992 -17064 -7928
rect -18236 -8008 -17064 -7992
rect -18236 -8072 -17148 -8008
rect -17084 -8072 -17064 -8008
rect -18236 -8088 -17064 -8072
rect -18236 -8152 -17148 -8088
rect -17084 -8152 -17064 -8088
rect -18236 -8168 -17064 -8152
rect -18236 -8232 -17148 -8168
rect -17084 -8232 -17064 -8168
rect -18236 -8280 -17064 -8232
rect -16824 -7448 -15652 -7400
rect -16824 -7512 -15736 -7448
rect -15672 -7512 -15652 -7448
rect -16824 -7528 -15652 -7512
rect -16824 -7592 -15736 -7528
rect -15672 -7592 -15652 -7528
rect -16824 -7608 -15652 -7592
rect -16824 -7672 -15736 -7608
rect -15672 -7672 -15652 -7608
rect -16824 -7688 -15652 -7672
rect -16824 -7752 -15736 -7688
rect -15672 -7752 -15652 -7688
rect -16824 -7768 -15652 -7752
rect -16824 -7832 -15736 -7768
rect -15672 -7832 -15652 -7768
rect -16824 -7848 -15652 -7832
rect -16824 -7912 -15736 -7848
rect -15672 -7912 -15652 -7848
rect -16824 -7928 -15652 -7912
rect -16824 -7992 -15736 -7928
rect -15672 -7992 -15652 -7928
rect -16824 -8008 -15652 -7992
rect -16824 -8072 -15736 -8008
rect -15672 -8072 -15652 -8008
rect -16824 -8088 -15652 -8072
rect -16824 -8152 -15736 -8088
rect -15672 -8152 -15652 -8088
rect -16824 -8168 -15652 -8152
rect -16824 -8232 -15736 -8168
rect -15672 -8232 -15652 -8168
rect -16824 -8280 -15652 -8232
rect -15412 -7448 -14240 -7400
rect -15412 -7512 -14324 -7448
rect -14260 -7512 -14240 -7448
rect -15412 -7528 -14240 -7512
rect -15412 -7592 -14324 -7528
rect -14260 -7592 -14240 -7528
rect -15412 -7608 -14240 -7592
rect -15412 -7672 -14324 -7608
rect -14260 -7672 -14240 -7608
rect -15412 -7688 -14240 -7672
rect -15412 -7752 -14324 -7688
rect -14260 -7752 -14240 -7688
rect -15412 -7768 -14240 -7752
rect -15412 -7832 -14324 -7768
rect -14260 -7832 -14240 -7768
rect -15412 -7848 -14240 -7832
rect -15412 -7912 -14324 -7848
rect -14260 -7912 -14240 -7848
rect -15412 -7928 -14240 -7912
rect -15412 -7992 -14324 -7928
rect -14260 -7992 -14240 -7928
rect -15412 -8008 -14240 -7992
rect -15412 -8072 -14324 -8008
rect -14260 -8072 -14240 -8008
rect -15412 -8088 -14240 -8072
rect -15412 -8152 -14324 -8088
rect -14260 -8152 -14240 -8088
rect -15412 -8168 -14240 -8152
rect -15412 -8232 -14324 -8168
rect -14260 -8232 -14240 -8168
rect -15412 -8280 -14240 -8232
rect -14000 -7448 -12828 -7400
rect -14000 -7512 -12912 -7448
rect -12848 -7512 -12828 -7448
rect -14000 -7528 -12828 -7512
rect -14000 -7592 -12912 -7528
rect -12848 -7592 -12828 -7528
rect -14000 -7608 -12828 -7592
rect -14000 -7672 -12912 -7608
rect -12848 -7672 -12828 -7608
rect -14000 -7688 -12828 -7672
rect -14000 -7752 -12912 -7688
rect -12848 -7752 -12828 -7688
rect -14000 -7768 -12828 -7752
rect -14000 -7832 -12912 -7768
rect -12848 -7832 -12828 -7768
rect -14000 -7848 -12828 -7832
rect -14000 -7912 -12912 -7848
rect -12848 -7912 -12828 -7848
rect -14000 -7928 -12828 -7912
rect -14000 -7992 -12912 -7928
rect -12848 -7992 -12828 -7928
rect -14000 -8008 -12828 -7992
rect -14000 -8072 -12912 -8008
rect -12848 -8072 -12828 -8008
rect -14000 -8088 -12828 -8072
rect -14000 -8152 -12912 -8088
rect -12848 -8152 -12828 -8088
rect -14000 -8168 -12828 -8152
rect -14000 -8232 -12912 -8168
rect -12848 -8232 -12828 -8168
rect -14000 -8280 -12828 -8232
rect -12588 -7448 -11416 -7400
rect -12588 -7512 -11500 -7448
rect -11436 -7512 -11416 -7448
rect -12588 -7528 -11416 -7512
rect -12588 -7592 -11500 -7528
rect -11436 -7592 -11416 -7528
rect -12588 -7608 -11416 -7592
rect -12588 -7672 -11500 -7608
rect -11436 -7672 -11416 -7608
rect -12588 -7688 -11416 -7672
rect -12588 -7752 -11500 -7688
rect -11436 -7752 -11416 -7688
rect -12588 -7768 -11416 -7752
rect -12588 -7832 -11500 -7768
rect -11436 -7832 -11416 -7768
rect -12588 -7848 -11416 -7832
rect -12588 -7912 -11500 -7848
rect -11436 -7912 -11416 -7848
rect -12588 -7928 -11416 -7912
rect -12588 -7992 -11500 -7928
rect -11436 -7992 -11416 -7928
rect -12588 -8008 -11416 -7992
rect -12588 -8072 -11500 -8008
rect -11436 -8072 -11416 -8008
rect -12588 -8088 -11416 -8072
rect -12588 -8152 -11500 -8088
rect -11436 -8152 -11416 -8088
rect -12588 -8168 -11416 -8152
rect -12588 -8232 -11500 -8168
rect -11436 -8232 -11416 -8168
rect -12588 -8280 -11416 -8232
rect -11176 -7448 -10004 -7400
rect -11176 -7512 -10088 -7448
rect -10024 -7512 -10004 -7448
rect -11176 -7528 -10004 -7512
rect -11176 -7592 -10088 -7528
rect -10024 -7592 -10004 -7528
rect -11176 -7608 -10004 -7592
rect -11176 -7672 -10088 -7608
rect -10024 -7672 -10004 -7608
rect -11176 -7688 -10004 -7672
rect -11176 -7752 -10088 -7688
rect -10024 -7752 -10004 -7688
rect -11176 -7768 -10004 -7752
rect -11176 -7832 -10088 -7768
rect -10024 -7832 -10004 -7768
rect -11176 -7848 -10004 -7832
rect -11176 -7912 -10088 -7848
rect -10024 -7912 -10004 -7848
rect -11176 -7928 -10004 -7912
rect -11176 -7992 -10088 -7928
rect -10024 -7992 -10004 -7928
rect -11176 -8008 -10004 -7992
rect -11176 -8072 -10088 -8008
rect -10024 -8072 -10004 -8008
rect -11176 -8088 -10004 -8072
rect -11176 -8152 -10088 -8088
rect -10024 -8152 -10004 -8088
rect -11176 -8168 -10004 -8152
rect -11176 -8232 -10088 -8168
rect -10024 -8232 -10004 -8168
rect -11176 -8280 -10004 -8232
rect -9764 -7448 -8592 -7400
rect -9764 -7512 -8676 -7448
rect -8612 -7512 -8592 -7448
rect -9764 -7528 -8592 -7512
rect -9764 -7592 -8676 -7528
rect -8612 -7592 -8592 -7528
rect -9764 -7608 -8592 -7592
rect -9764 -7672 -8676 -7608
rect -8612 -7672 -8592 -7608
rect -9764 -7688 -8592 -7672
rect -9764 -7752 -8676 -7688
rect -8612 -7752 -8592 -7688
rect -9764 -7768 -8592 -7752
rect -9764 -7832 -8676 -7768
rect -8612 -7832 -8592 -7768
rect -9764 -7848 -8592 -7832
rect -9764 -7912 -8676 -7848
rect -8612 -7912 -8592 -7848
rect -9764 -7928 -8592 -7912
rect -9764 -7992 -8676 -7928
rect -8612 -7992 -8592 -7928
rect -9764 -8008 -8592 -7992
rect -9764 -8072 -8676 -8008
rect -8612 -8072 -8592 -8008
rect -9764 -8088 -8592 -8072
rect -9764 -8152 -8676 -8088
rect -8612 -8152 -8592 -8088
rect -9764 -8168 -8592 -8152
rect -9764 -8232 -8676 -8168
rect -8612 -8232 -8592 -8168
rect -9764 -8280 -8592 -8232
rect -8352 -7448 -7180 -7400
rect -8352 -7512 -7264 -7448
rect -7200 -7512 -7180 -7448
rect -8352 -7528 -7180 -7512
rect -8352 -7592 -7264 -7528
rect -7200 -7592 -7180 -7528
rect -8352 -7608 -7180 -7592
rect -8352 -7672 -7264 -7608
rect -7200 -7672 -7180 -7608
rect -8352 -7688 -7180 -7672
rect -8352 -7752 -7264 -7688
rect -7200 -7752 -7180 -7688
rect -8352 -7768 -7180 -7752
rect -8352 -7832 -7264 -7768
rect -7200 -7832 -7180 -7768
rect -8352 -7848 -7180 -7832
rect -8352 -7912 -7264 -7848
rect -7200 -7912 -7180 -7848
rect -8352 -7928 -7180 -7912
rect -8352 -7992 -7264 -7928
rect -7200 -7992 -7180 -7928
rect -8352 -8008 -7180 -7992
rect -8352 -8072 -7264 -8008
rect -7200 -8072 -7180 -8008
rect -8352 -8088 -7180 -8072
rect -8352 -8152 -7264 -8088
rect -7200 -8152 -7180 -8088
rect -8352 -8168 -7180 -8152
rect -8352 -8232 -7264 -8168
rect -7200 -8232 -7180 -8168
rect -8352 -8280 -7180 -8232
rect -6940 -7448 -5768 -7400
rect -6940 -7512 -5852 -7448
rect -5788 -7512 -5768 -7448
rect -6940 -7528 -5768 -7512
rect -6940 -7592 -5852 -7528
rect -5788 -7592 -5768 -7528
rect -6940 -7608 -5768 -7592
rect -6940 -7672 -5852 -7608
rect -5788 -7672 -5768 -7608
rect -6940 -7688 -5768 -7672
rect -6940 -7752 -5852 -7688
rect -5788 -7752 -5768 -7688
rect -6940 -7768 -5768 -7752
rect -6940 -7832 -5852 -7768
rect -5788 -7832 -5768 -7768
rect -6940 -7848 -5768 -7832
rect -6940 -7912 -5852 -7848
rect -5788 -7912 -5768 -7848
rect -6940 -7928 -5768 -7912
rect -6940 -7992 -5852 -7928
rect -5788 -7992 -5768 -7928
rect -6940 -8008 -5768 -7992
rect -6940 -8072 -5852 -8008
rect -5788 -8072 -5768 -8008
rect -6940 -8088 -5768 -8072
rect -6940 -8152 -5852 -8088
rect -5788 -8152 -5768 -8088
rect -6940 -8168 -5768 -8152
rect -6940 -8232 -5852 -8168
rect -5788 -8232 -5768 -8168
rect -6940 -8280 -5768 -8232
rect -5528 -7448 -4356 -7400
rect -5528 -7512 -4440 -7448
rect -4376 -7512 -4356 -7448
rect -5528 -7528 -4356 -7512
rect -5528 -7592 -4440 -7528
rect -4376 -7592 -4356 -7528
rect -5528 -7608 -4356 -7592
rect -5528 -7672 -4440 -7608
rect -4376 -7672 -4356 -7608
rect -5528 -7688 -4356 -7672
rect -5528 -7752 -4440 -7688
rect -4376 -7752 -4356 -7688
rect -5528 -7768 -4356 -7752
rect -5528 -7832 -4440 -7768
rect -4376 -7832 -4356 -7768
rect -5528 -7848 -4356 -7832
rect -5528 -7912 -4440 -7848
rect -4376 -7912 -4356 -7848
rect -5528 -7928 -4356 -7912
rect -5528 -7992 -4440 -7928
rect -4376 -7992 -4356 -7928
rect -5528 -8008 -4356 -7992
rect -5528 -8072 -4440 -8008
rect -4376 -8072 -4356 -8008
rect -5528 -8088 -4356 -8072
rect -5528 -8152 -4440 -8088
rect -4376 -8152 -4356 -8088
rect -5528 -8168 -4356 -8152
rect -5528 -8232 -4440 -8168
rect -4376 -8232 -4356 -8168
rect -5528 -8280 -4356 -8232
rect -4116 -7448 -2944 -7400
rect -4116 -7512 -3028 -7448
rect -2964 -7512 -2944 -7448
rect -4116 -7528 -2944 -7512
rect -4116 -7592 -3028 -7528
rect -2964 -7592 -2944 -7528
rect -4116 -7608 -2944 -7592
rect -4116 -7672 -3028 -7608
rect -2964 -7672 -2944 -7608
rect -4116 -7688 -2944 -7672
rect -4116 -7752 -3028 -7688
rect -2964 -7752 -2944 -7688
rect -4116 -7768 -2944 -7752
rect -4116 -7832 -3028 -7768
rect -2964 -7832 -2944 -7768
rect -4116 -7848 -2944 -7832
rect -4116 -7912 -3028 -7848
rect -2964 -7912 -2944 -7848
rect -4116 -7928 -2944 -7912
rect -4116 -7992 -3028 -7928
rect -2964 -7992 -2944 -7928
rect -4116 -8008 -2944 -7992
rect -4116 -8072 -3028 -8008
rect -2964 -8072 -2944 -8008
rect -4116 -8088 -2944 -8072
rect -4116 -8152 -3028 -8088
rect -2964 -8152 -2944 -8088
rect -4116 -8168 -2944 -8152
rect -4116 -8232 -3028 -8168
rect -2964 -8232 -2944 -8168
rect -4116 -8280 -2944 -8232
rect -2704 -7448 -1532 -7400
rect -2704 -7512 -1616 -7448
rect -1552 -7512 -1532 -7448
rect -2704 -7528 -1532 -7512
rect -2704 -7592 -1616 -7528
rect -1552 -7592 -1532 -7528
rect -2704 -7608 -1532 -7592
rect -2704 -7672 -1616 -7608
rect -1552 -7672 -1532 -7608
rect -2704 -7688 -1532 -7672
rect -2704 -7752 -1616 -7688
rect -1552 -7752 -1532 -7688
rect -2704 -7768 -1532 -7752
rect -2704 -7832 -1616 -7768
rect -1552 -7832 -1532 -7768
rect -2704 -7848 -1532 -7832
rect -2704 -7912 -1616 -7848
rect -1552 -7912 -1532 -7848
rect -2704 -7928 -1532 -7912
rect -2704 -7992 -1616 -7928
rect -1552 -7992 -1532 -7928
rect -2704 -8008 -1532 -7992
rect -2704 -8072 -1616 -8008
rect -1552 -8072 -1532 -8008
rect -2704 -8088 -1532 -8072
rect -2704 -8152 -1616 -8088
rect -1552 -8152 -1532 -8088
rect -2704 -8168 -1532 -8152
rect -2704 -8232 -1616 -8168
rect -1552 -8232 -1532 -8168
rect -2704 -8280 -1532 -8232
rect -1292 -7448 -120 -7400
rect -1292 -7512 -204 -7448
rect -140 -7512 -120 -7448
rect -1292 -7528 -120 -7512
rect -1292 -7592 -204 -7528
rect -140 -7592 -120 -7528
rect -1292 -7608 -120 -7592
rect -1292 -7672 -204 -7608
rect -140 -7672 -120 -7608
rect -1292 -7688 -120 -7672
rect -1292 -7752 -204 -7688
rect -140 -7752 -120 -7688
rect -1292 -7768 -120 -7752
rect -1292 -7832 -204 -7768
rect -140 -7832 -120 -7768
rect -1292 -7848 -120 -7832
rect -1292 -7912 -204 -7848
rect -140 -7912 -120 -7848
rect -1292 -7928 -120 -7912
rect -1292 -7992 -204 -7928
rect -140 -7992 -120 -7928
rect -1292 -8008 -120 -7992
rect -1292 -8072 -204 -8008
rect -140 -8072 -120 -8008
rect -1292 -8088 -120 -8072
rect -1292 -8152 -204 -8088
rect -140 -8152 -120 -8088
rect -1292 -8168 -120 -8152
rect -1292 -8232 -204 -8168
rect -140 -8232 -120 -8168
rect -1292 -8280 -120 -8232
rect 120 -7448 1292 -7400
rect 120 -7512 1208 -7448
rect 1272 -7512 1292 -7448
rect 120 -7528 1292 -7512
rect 120 -7592 1208 -7528
rect 1272 -7592 1292 -7528
rect 120 -7608 1292 -7592
rect 120 -7672 1208 -7608
rect 1272 -7672 1292 -7608
rect 120 -7688 1292 -7672
rect 120 -7752 1208 -7688
rect 1272 -7752 1292 -7688
rect 120 -7768 1292 -7752
rect 120 -7832 1208 -7768
rect 1272 -7832 1292 -7768
rect 120 -7848 1292 -7832
rect 120 -7912 1208 -7848
rect 1272 -7912 1292 -7848
rect 120 -7928 1292 -7912
rect 120 -7992 1208 -7928
rect 1272 -7992 1292 -7928
rect 120 -8008 1292 -7992
rect 120 -8072 1208 -8008
rect 1272 -8072 1292 -8008
rect 120 -8088 1292 -8072
rect 120 -8152 1208 -8088
rect 1272 -8152 1292 -8088
rect 120 -8168 1292 -8152
rect 120 -8232 1208 -8168
rect 1272 -8232 1292 -8168
rect 120 -8280 1292 -8232
rect 1532 -7448 2704 -7400
rect 1532 -7512 2620 -7448
rect 2684 -7512 2704 -7448
rect 1532 -7528 2704 -7512
rect 1532 -7592 2620 -7528
rect 2684 -7592 2704 -7528
rect 1532 -7608 2704 -7592
rect 1532 -7672 2620 -7608
rect 2684 -7672 2704 -7608
rect 1532 -7688 2704 -7672
rect 1532 -7752 2620 -7688
rect 2684 -7752 2704 -7688
rect 1532 -7768 2704 -7752
rect 1532 -7832 2620 -7768
rect 2684 -7832 2704 -7768
rect 1532 -7848 2704 -7832
rect 1532 -7912 2620 -7848
rect 2684 -7912 2704 -7848
rect 1532 -7928 2704 -7912
rect 1532 -7992 2620 -7928
rect 2684 -7992 2704 -7928
rect 1532 -8008 2704 -7992
rect 1532 -8072 2620 -8008
rect 2684 -8072 2704 -8008
rect 1532 -8088 2704 -8072
rect 1532 -8152 2620 -8088
rect 2684 -8152 2704 -8088
rect 1532 -8168 2704 -8152
rect 1532 -8232 2620 -8168
rect 2684 -8232 2704 -8168
rect 1532 -8280 2704 -8232
rect 2944 -7448 4116 -7400
rect 2944 -7512 4032 -7448
rect 4096 -7512 4116 -7448
rect 2944 -7528 4116 -7512
rect 2944 -7592 4032 -7528
rect 4096 -7592 4116 -7528
rect 2944 -7608 4116 -7592
rect 2944 -7672 4032 -7608
rect 4096 -7672 4116 -7608
rect 2944 -7688 4116 -7672
rect 2944 -7752 4032 -7688
rect 4096 -7752 4116 -7688
rect 2944 -7768 4116 -7752
rect 2944 -7832 4032 -7768
rect 4096 -7832 4116 -7768
rect 2944 -7848 4116 -7832
rect 2944 -7912 4032 -7848
rect 4096 -7912 4116 -7848
rect 2944 -7928 4116 -7912
rect 2944 -7992 4032 -7928
rect 4096 -7992 4116 -7928
rect 2944 -8008 4116 -7992
rect 2944 -8072 4032 -8008
rect 4096 -8072 4116 -8008
rect 2944 -8088 4116 -8072
rect 2944 -8152 4032 -8088
rect 4096 -8152 4116 -8088
rect 2944 -8168 4116 -8152
rect 2944 -8232 4032 -8168
rect 4096 -8232 4116 -8168
rect 2944 -8280 4116 -8232
rect 4356 -7448 5528 -7400
rect 4356 -7512 5444 -7448
rect 5508 -7512 5528 -7448
rect 4356 -7528 5528 -7512
rect 4356 -7592 5444 -7528
rect 5508 -7592 5528 -7528
rect 4356 -7608 5528 -7592
rect 4356 -7672 5444 -7608
rect 5508 -7672 5528 -7608
rect 4356 -7688 5528 -7672
rect 4356 -7752 5444 -7688
rect 5508 -7752 5528 -7688
rect 4356 -7768 5528 -7752
rect 4356 -7832 5444 -7768
rect 5508 -7832 5528 -7768
rect 4356 -7848 5528 -7832
rect 4356 -7912 5444 -7848
rect 5508 -7912 5528 -7848
rect 4356 -7928 5528 -7912
rect 4356 -7992 5444 -7928
rect 5508 -7992 5528 -7928
rect 4356 -8008 5528 -7992
rect 4356 -8072 5444 -8008
rect 5508 -8072 5528 -8008
rect 4356 -8088 5528 -8072
rect 4356 -8152 5444 -8088
rect 5508 -8152 5528 -8088
rect 4356 -8168 5528 -8152
rect 4356 -8232 5444 -8168
rect 5508 -8232 5528 -8168
rect 4356 -8280 5528 -8232
rect 5768 -7448 6940 -7400
rect 5768 -7512 6856 -7448
rect 6920 -7512 6940 -7448
rect 5768 -7528 6940 -7512
rect 5768 -7592 6856 -7528
rect 6920 -7592 6940 -7528
rect 5768 -7608 6940 -7592
rect 5768 -7672 6856 -7608
rect 6920 -7672 6940 -7608
rect 5768 -7688 6940 -7672
rect 5768 -7752 6856 -7688
rect 6920 -7752 6940 -7688
rect 5768 -7768 6940 -7752
rect 5768 -7832 6856 -7768
rect 6920 -7832 6940 -7768
rect 5768 -7848 6940 -7832
rect 5768 -7912 6856 -7848
rect 6920 -7912 6940 -7848
rect 5768 -7928 6940 -7912
rect 5768 -7992 6856 -7928
rect 6920 -7992 6940 -7928
rect 5768 -8008 6940 -7992
rect 5768 -8072 6856 -8008
rect 6920 -8072 6940 -8008
rect 5768 -8088 6940 -8072
rect 5768 -8152 6856 -8088
rect 6920 -8152 6940 -8088
rect 5768 -8168 6940 -8152
rect 5768 -8232 6856 -8168
rect 6920 -8232 6940 -8168
rect 5768 -8280 6940 -8232
rect 7180 -7448 8352 -7400
rect 7180 -7512 8268 -7448
rect 8332 -7512 8352 -7448
rect 7180 -7528 8352 -7512
rect 7180 -7592 8268 -7528
rect 8332 -7592 8352 -7528
rect 7180 -7608 8352 -7592
rect 7180 -7672 8268 -7608
rect 8332 -7672 8352 -7608
rect 7180 -7688 8352 -7672
rect 7180 -7752 8268 -7688
rect 8332 -7752 8352 -7688
rect 7180 -7768 8352 -7752
rect 7180 -7832 8268 -7768
rect 8332 -7832 8352 -7768
rect 7180 -7848 8352 -7832
rect 7180 -7912 8268 -7848
rect 8332 -7912 8352 -7848
rect 7180 -7928 8352 -7912
rect 7180 -7992 8268 -7928
rect 8332 -7992 8352 -7928
rect 7180 -8008 8352 -7992
rect 7180 -8072 8268 -8008
rect 8332 -8072 8352 -8008
rect 7180 -8088 8352 -8072
rect 7180 -8152 8268 -8088
rect 8332 -8152 8352 -8088
rect 7180 -8168 8352 -8152
rect 7180 -8232 8268 -8168
rect 8332 -8232 8352 -8168
rect 7180 -8280 8352 -8232
rect 8592 -7448 9764 -7400
rect 8592 -7512 9680 -7448
rect 9744 -7512 9764 -7448
rect 8592 -7528 9764 -7512
rect 8592 -7592 9680 -7528
rect 9744 -7592 9764 -7528
rect 8592 -7608 9764 -7592
rect 8592 -7672 9680 -7608
rect 9744 -7672 9764 -7608
rect 8592 -7688 9764 -7672
rect 8592 -7752 9680 -7688
rect 9744 -7752 9764 -7688
rect 8592 -7768 9764 -7752
rect 8592 -7832 9680 -7768
rect 9744 -7832 9764 -7768
rect 8592 -7848 9764 -7832
rect 8592 -7912 9680 -7848
rect 9744 -7912 9764 -7848
rect 8592 -7928 9764 -7912
rect 8592 -7992 9680 -7928
rect 9744 -7992 9764 -7928
rect 8592 -8008 9764 -7992
rect 8592 -8072 9680 -8008
rect 9744 -8072 9764 -8008
rect 8592 -8088 9764 -8072
rect 8592 -8152 9680 -8088
rect 9744 -8152 9764 -8088
rect 8592 -8168 9764 -8152
rect 8592 -8232 9680 -8168
rect 9744 -8232 9764 -8168
rect 8592 -8280 9764 -8232
rect 10004 -7448 11176 -7400
rect 10004 -7512 11092 -7448
rect 11156 -7512 11176 -7448
rect 10004 -7528 11176 -7512
rect 10004 -7592 11092 -7528
rect 11156 -7592 11176 -7528
rect 10004 -7608 11176 -7592
rect 10004 -7672 11092 -7608
rect 11156 -7672 11176 -7608
rect 10004 -7688 11176 -7672
rect 10004 -7752 11092 -7688
rect 11156 -7752 11176 -7688
rect 10004 -7768 11176 -7752
rect 10004 -7832 11092 -7768
rect 11156 -7832 11176 -7768
rect 10004 -7848 11176 -7832
rect 10004 -7912 11092 -7848
rect 11156 -7912 11176 -7848
rect 10004 -7928 11176 -7912
rect 10004 -7992 11092 -7928
rect 11156 -7992 11176 -7928
rect 10004 -8008 11176 -7992
rect 10004 -8072 11092 -8008
rect 11156 -8072 11176 -8008
rect 10004 -8088 11176 -8072
rect 10004 -8152 11092 -8088
rect 11156 -8152 11176 -8088
rect 10004 -8168 11176 -8152
rect 10004 -8232 11092 -8168
rect 11156 -8232 11176 -8168
rect 10004 -8280 11176 -8232
rect 11416 -7448 12588 -7400
rect 11416 -7512 12504 -7448
rect 12568 -7512 12588 -7448
rect 11416 -7528 12588 -7512
rect 11416 -7592 12504 -7528
rect 12568 -7592 12588 -7528
rect 11416 -7608 12588 -7592
rect 11416 -7672 12504 -7608
rect 12568 -7672 12588 -7608
rect 11416 -7688 12588 -7672
rect 11416 -7752 12504 -7688
rect 12568 -7752 12588 -7688
rect 11416 -7768 12588 -7752
rect 11416 -7832 12504 -7768
rect 12568 -7832 12588 -7768
rect 11416 -7848 12588 -7832
rect 11416 -7912 12504 -7848
rect 12568 -7912 12588 -7848
rect 11416 -7928 12588 -7912
rect 11416 -7992 12504 -7928
rect 12568 -7992 12588 -7928
rect 11416 -8008 12588 -7992
rect 11416 -8072 12504 -8008
rect 12568 -8072 12588 -8008
rect 11416 -8088 12588 -8072
rect 11416 -8152 12504 -8088
rect 12568 -8152 12588 -8088
rect 11416 -8168 12588 -8152
rect 11416 -8232 12504 -8168
rect 12568 -8232 12588 -8168
rect 11416 -8280 12588 -8232
rect 12828 -7448 14000 -7400
rect 12828 -7512 13916 -7448
rect 13980 -7512 14000 -7448
rect 12828 -7528 14000 -7512
rect 12828 -7592 13916 -7528
rect 13980 -7592 14000 -7528
rect 12828 -7608 14000 -7592
rect 12828 -7672 13916 -7608
rect 13980 -7672 14000 -7608
rect 12828 -7688 14000 -7672
rect 12828 -7752 13916 -7688
rect 13980 -7752 14000 -7688
rect 12828 -7768 14000 -7752
rect 12828 -7832 13916 -7768
rect 13980 -7832 14000 -7768
rect 12828 -7848 14000 -7832
rect 12828 -7912 13916 -7848
rect 13980 -7912 14000 -7848
rect 12828 -7928 14000 -7912
rect 12828 -7992 13916 -7928
rect 13980 -7992 14000 -7928
rect 12828 -8008 14000 -7992
rect 12828 -8072 13916 -8008
rect 13980 -8072 14000 -8008
rect 12828 -8088 14000 -8072
rect 12828 -8152 13916 -8088
rect 13980 -8152 14000 -8088
rect 12828 -8168 14000 -8152
rect 12828 -8232 13916 -8168
rect 13980 -8232 14000 -8168
rect 12828 -8280 14000 -8232
rect 14240 -7448 15412 -7400
rect 14240 -7512 15328 -7448
rect 15392 -7512 15412 -7448
rect 14240 -7528 15412 -7512
rect 14240 -7592 15328 -7528
rect 15392 -7592 15412 -7528
rect 14240 -7608 15412 -7592
rect 14240 -7672 15328 -7608
rect 15392 -7672 15412 -7608
rect 14240 -7688 15412 -7672
rect 14240 -7752 15328 -7688
rect 15392 -7752 15412 -7688
rect 14240 -7768 15412 -7752
rect 14240 -7832 15328 -7768
rect 15392 -7832 15412 -7768
rect 14240 -7848 15412 -7832
rect 14240 -7912 15328 -7848
rect 15392 -7912 15412 -7848
rect 14240 -7928 15412 -7912
rect 14240 -7992 15328 -7928
rect 15392 -7992 15412 -7928
rect 14240 -8008 15412 -7992
rect 14240 -8072 15328 -8008
rect 15392 -8072 15412 -8008
rect 14240 -8088 15412 -8072
rect 14240 -8152 15328 -8088
rect 15392 -8152 15412 -8088
rect 14240 -8168 15412 -8152
rect 14240 -8232 15328 -8168
rect 15392 -8232 15412 -8168
rect 14240 -8280 15412 -8232
rect 15652 -7448 16824 -7400
rect 15652 -7512 16740 -7448
rect 16804 -7512 16824 -7448
rect 15652 -7528 16824 -7512
rect 15652 -7592 16740 -7528
rect 16804 -7592 16824 -7528
rect 15652 -7608 16824 -7592
rect 15652 -7672 16740 -7608
rect 16804 -7672 16824 -7608
rect 15652 -7688 16824 -7672
rect 15652 -7752 16740 -7688
rect 16804 -7752 16824 -7688
rect 15652 -7768 16824 -7752
rect 15652 -7832 16740 -7768
rect 16804 -7832 16824 -7768
rect 15652 -7848 16824 -7832
rect 15652 -7912 16740 -7848
rect 16804 -7912 16824 -7848
rect 15652 -7928 16824 -7912
rect 15652 -7992 16740 -7928
rect 16804 -7992 16824 -7928
rect 15652 -8008 16824 -7992
rect 15652 -8072 16740 -8008
rect 16804 -8072 16824 -8008
rect 15652 -8088 16824 -8072
rect 15652 -8152 16740 -8088
rect 16804 -8152 16824 -8088
rect 15652 -8168 16824 -8152
rect 15652 -8232 16740 -8168
rect 16804 -8232 16824 -8168
rect 15652 -8280 16824 -8232
rect 17064 -7448 18236 -7400
rect 17064 -7512 18152 -7448
rect 18216 -7512 18236 -7448
rect 17064 -7528 18236 -7512
rect 17064 -7592 18152 -7528
rect 18216 -7592 18236 -7528
rect 17064 -7608 18236 -7592
rect 17064 -7672 18152 -7608
rect 18216 -7672 18236 -7608
rect 17064 -7688 18236 -7672
rect 17064 -7752 18152 -7688
rect 18216 -7752 18236 -7688
rect 17064 -7768 18236 -7752
rect 17064 -7832 18152 -7768
rect 18216 -7832 18236 -7768
rect 17064 -7848 18236 -7832
rect 17064 -7912 18152 -7848
rect 18216 -7912 18236 -7848
rect 17064 -7928 18236 -7912
rect 17064 -7992 18152 -7928
rect 18216 -7992 18236 -7928
rect 17064 -8008 18236 -7992
rect 17064 -8072 18152 -8008
rect 18216 -8072 18236 -8008
rect 17064 -8088 18236 -8072
rect 17064 -8152 18152 -8088
rect 18216 -8152 18236 -8088
rect 17064 -8168 18236 -8152
rect 17064 -8232 18152 -8168
rect 18216 -8232 18236 -8168
rect 17064 -8280 18236 -8232
rect 18476 -7448 19648 -7400
rect 18476 -7512 19564 -7448
rect 19628 -7512 19648 -7448
rect 18476 -7528 19648 -7512
rect 18476 -7592 19564 -7528
rect 19628 -7592 19648 -7528
rect 18476 -7608 19648 -7592
rect 18476 -7672 19564 -7608
rect 19628 -7672 19648 -7608
rect 18476 -7688 19648 -7672
rect 18476 -7752 19564 -7688
rect 19628 -7752 19648 -7688
rect 18476 -7768 19648 -7752
rect 18476 -7832 19564 -7768
rect 19628 -7832 19648 -7768
rect 18476 -7848 19648 -7832
rect 18476 -7912 19564 -7848
rect 19628 -7912 19648 -7848
rect 18476 -7928 19648 -7912
rect 18476 -7992 19564 -7928
rect 19628 -7992 19648 -7928
rect 18476 -8008 19648 -7992
rect 18476 -8072 19564 -8008
rect 19628 -8072 19648 -8008
rect 18476 -8088 19648 -8072
rect 18476 -8152 19564 -8088
rect 19628 -8152 19648 -8088
rect 18476 -8168 19648 -8152
rect 18476 -8232 19564 -8168
rect 19628 -8232 19648 -8168
rect 18476 -8280 19648 -8232
rect 19888 -7448 21060 -7400
rect 19888 -7512 20976 -7448
rect 21040 -7512 21060 -7448
rect 19888 -7528 21060 -7512
rect 19888 -7592 20976 -7528
rect 21040 -7592 21060 -7528
rect 19888 -7608 21060 -7592
rect 19888 -7672 20976 -7608
rect 21040 -7672 21060 -7608
rect 19888 -7688 21060 -7672
rect 19888 -7752 20976 -7688
rect 21040 -7752 21060 -7688
rect 19888 -7768 21060 -7752
rect 19888 -7832 20976 -7768
rect 21040 -7832 21060 -7768
rect 19888 -7848 21060 -7832
rect 19888 -7912 20976 -7848
rect 21040 -7912 21060 -7848
rect 19888 -7928 21060 -7912
rect 19888 -7992 20976 -7928
rect 21040 -7992 21060 -7928
rect 19888 -8008 21060 -7992
rect 19888 -8072 20976 -8008
rect 21040 -8072 21060 -8008
rect 19888 -8088 21060 -8072
rect 19888 -8152 20976 -8088
rect 21040 -8152 21060 -8088
rect 19888 -8168 21060 -8152
rect 19888 -8232 20976 -8168
rect 21040 -8232 21060 -8168
rect 19888 -8280 21060 -8232
rect 21300 -7448 22472 -7400
rect 21300 -7512 22388 -7448
rect 22452 -7512 22472 -7448
rect 21300 -7528 22472 -7512
rect 21300 -7592 22388 -7528
rect 22452 -7592 22472 -7528
rect 21300 -7608 22472 -7592
rect 21300 -7672 22388 -7608
rect 22452 -7672 22472 -7608
rect 21300 -7688 22472 -7672
rect 21300 -7752 22388 -7688
rect 22452 -7752 22472 -7688
rect 21300 -7768 22472 -7752
rect 21300 -7832 22388 -7768
rect 22452 -7832 22472 -7768
rect 21300 -7848 22472 -7832
rect 21300 -7912 22388 -7848
rect 22452 -7912 22472 -7848
rect 21300 -7928 22472 -7912
rect 21300 -7992 22388 -7928
rect 22452 -7992 22472 -7928
rect 21300 -8008 22472 -7992
rect 21300 -8072 22388 -8008
rect 22452 -8072 22472 -8008
rect 21300 -8088 22472 -8072
rect 21300 -8152 22388 -8088
rect 22452 -8152 22472 -8088
rect 21300 -8168 22472 -8152
rect 21300 -8232 22388 -8168
rect 22452 -8232 22472 -8168
rect 21300 -8280 22472 -8232
rect 22712 -7448 23884 -7400
rect 22712 -7512 23800 -7448
rect 23864 -7512 23884 -7448
rect 22712 -7528 23884 -7512
rect 22712 -7592 23800 -7528
rect 23864 -7592 23884 -7528
rect 22712 -7608 23884 -7592
rect 22712 -7672 23800 -7608
rect 23864 -7672 23884 -7608
rect 22712 -7688 23884 -7672
rect 22712 -7752 23800 -7688
rect 23864 -7752 23884 -7688
rect 22712 -7768 23884 -7752
rect 22712 -7832 23800 -7768
rect 23864 -7832 23884 -7768
rect 22712 -7848 23884 -7832
rect 22712 -7912 23800 -7848
rect 23864 -7912 23884 -7848
rect 22712 -7928 23884 -7912
rect 22712 -7992 23800 -7928
rect 23864 -7992 23884 -7928
rect 22712 -8008 23884 -7992
rect 22712 -8072 23800 -8008
rect 23864 -8072 23884 -8008
rect 22712 -8088 23884 -8072
rect 22712 -8152 23800 -8088
rect 23864 -8152 23884 -8088
rect 22712 -8168 23884 -8152
rect 22712 -8232 23800 -8168
rect 23864 -8232 23884 -8168
rect 22712 -8280 23884 -8232
rect -23884 -8568 -22712 -8520
rect -23884 -8632 -22796 -8568
rect -22732 -8632 -22712 -8568
rect -23884 -8648 -22712 -8632
rect -23884 -8712 -22796 -8648
rect -22732 -8712 -22712 -8648
rect -23884 -8728 -22712 -8712
rect -23884 -8792 -22796 -8728
rect -22732 -8792 -22712 -8728
rect -23884 -8808 -22712 -8792
rect -23884 -8872 -22796 -8808
rect -22732 -8872 -22712 -8808
rect -23884 -8888 -22712 -8872
rect -23884 -8952 -22796 -8888
rect -22732 -8952 -22712 -8888
rect -23884 -8968 -22712 -8952
rect -23884 -9032 -22796 -8968
rect -22732 -9032 -22712 -8968
rect -23884 -9048 -22712 -9032
rect -23884 -9112 -22796 -9048
rect -22732 -9112 -22712 -9048
rect -23884 -9128 -22712 -9112
rect -23884 -9192 -22796 -9128
rect -22732 -9192 -22712 -9128
rect -23884 -9208 -22712 -9192
rect -23884 -9272 -22796 -9208
rect -22732 -9272 -22712 -9208
rect -23884 -9288 -22712 -9272
rect -23884 -9352 -22796 -9288
rect -22732 -9352 -22712 -9288
rect -23884 -9400 -22712 -9352
rect -22472 -8568 -21300 -8520
rect -22472 -8632 -21384 -8568
rect -21320 -8632 -21300 -8568
rect -22472 -8648 -21300 -8632
rect -22472 -8712 -21384 -8648
rect -21320 -8712 -21300 -8648
rect -22472 -8728 -21300 -8712
rect -22472 -8792 -21384 -8728
rect -21320 -8792 -21300 -8728
rect -22472 -8808 -21300 -8792
rect -22472 -8872 -21384 -8808
rect -21320 -8872 -21300 -8808
rect -22472 -8888 -21300 -8872
rect -22472 -8952 -21384 -8888
rect -21320 -8952 -21300 -8888
rect -22472 -8968 -21300 -8952
rect -22472 -9032 -21384 -8968
rect -21320 -9032 -21300 -8968
rect -22472 -9048 -21300 -9032
rect -22472 -9112 -21384 -9048
rect -21320 -9112 -21300 -9048
rect -22472 -9128 -21300 -9112
rect -22472 -9192 -21384 -9128
rect -21320 -9192 -21300 -9128
rect -22472 -9208 -21300 -9192
rect -22472 -9272 -21384 -9208
rect -21320 -9272 -21300 -9208
rect -22472 -9288 -21300 -9272
rect -22472 -9352 -21384 -9288
rect -21320 -9352 -21300 -9288
rect -22472 -9400 -21300 -9352
rect -21060 -8568 -19888 -8520
rect -21060 -8632 -19972 -8568
rect -19908 -8632 -19888 -8568
rect -21060 -8648 -19888 -8632
rect -21060 -8712 -19972 -8648
rect -19908 -8712 -19888 -8648
rect -21060 -8728 -19888 -8712
rect -21060 -8792 -19972 -8728
rect -19908 -8792 -19888 -8728
rect -21060 -8808 -19888 -8792
rect -21060 -8872 -19972 -8808
rect -19908 -8872 -19888 -8808
rect -21060 -8888 -19888 -8872
rect -21060 -8952 -19972 -8888
rect -19908 -8952 -19888 -8888
rect -21060 -8968 -19888 -8952
rect -21060 -9032 -19972 -8968
rect -19908 -9032 -19888 -8968
rect -21060 -9048 -19888 -9032
rect -21060 -9112 -19972 -9048
rect -19908 -9112 -19888 -9048
rect -21060 -9128 -19888 -9112
rect -21060 -9192 -19972 -9128
rect -19908 -9192 -19888 -9128
rect -21060 -9208 -19888 -9192
rect -21060 -9272 -19972 -9208
rect -19908 -9272 -19888 -9208
rect -21060 -9288 -19888 -9272
rect -21060 -9352 -19972 -9288
rect -19908 -9352 -19888 -9288
rect -21060 -9400 -19888 -9352
rect -19648 -8568 -18476 -8520
rect -19648 -8632 -18560 -8568
rect -18496 -8632 -18476 -8568
rect -19648 -8648 -18476 -8632
rect -19648 -8712 -18560 -8648
rect -18496 -8712 -18476 -8648
rect -19648 -8728 -18476 -8712
rect -19648 -8792 -18560 -8728
rect -18496 -8792 -18476 -8728
rect -19648 -8808 -18476 -8792
rect -19648 -8872 -18560 -8808
rect -18496 -8872 -18476 -8808
rect -19648 -8888 -18476 -8872
rect -19648 -8952 -18560 -8888
rect -18496 -8952 -18476 -8888
rect -19648 -8968 -18476 -8952
rect -19648 -9032 -18560 -8968
rect -18496 -9032 -18476 -8968
rect -19648 -9048 -18476 -9032
rect -19648 -9112 -18560 -9048
rect -18496 -9112 -18476 -9048
rect -19648 -9128 -18476 -9112
rect -19648 -9192 -18560 -9128
rect -18496 -9192 -18476 -9128
rect -19648 -9208 -18476 -9192
rect -19648 -9272 -18560 -9208
rect -18496 -9272 -18476 -9208
rect -19648 -9288 -18476 -9272
rect -19648 -9352 -18560 -9288
rect -18496 -9352 -18476 -9288
rect -19648 -9400 -18476 -9352
rect -18236 -8568 -17064 -8520
rect -18236 -8632 -17148 -8568
rect -17084 -8632 -17064 -8568
rect -18236 -8648 -17064 -8632
rect -18236 -8712 -17148 -8648
rect -17084 -8712 -17064 -8648
rect -18236 -8728 -17064 -8712
rect -18236 -8792 -17148 -8728
rect -17084 -8792 -17064 -8728
rect -18236 -8808 -17064 -8792
rect -18236 -8872 -17148 -8808
rect -17084 -8872 -17064 -8808
rect -18236 -8888 -17064 -8872
rect -18236 -8952 -17148 -8888
rect -17084 -8952 -17064 -8888
rect -18236 -8968 -17064 -8952
rect -18236 -9032 -17148 -8968
rect -17084 -9032 -17064 -8968
rect -18236 -9048 -17064 -9032
rect -18236 -9112 -17148 -9048
rect -17084 -9112 -17064 -9048
rect -18236 -9128 -17064 -9112
rect -18236 -9192 -17148 -9128
rect -17084 -9192 -17064 -9128
rect -18236 -9208 -17064 -9192
rect -18236 -9272 -17148 -9208
rect -17084 -9272 -17064 -9208
rect -18236 -9288 -17064 -9272
rect -18236 -9352 -17148 -9288
rect -17084 -9352 -17064 -9288
rect -18236 -9400 -17064 -9352
rect -16824 -8568 -15652 -8520
rect -16824 -8632 -15736 -8568
rect -15672 -8632 -15652 -8568
rect -16824 -8648 -15652 -8632
rect -16824 -8712 -15736 -8648
rect -15672 -8712 -15652 -8648
rect -16824 -8728 -15652 -8712
rect -16824 -8792 -15736 -8728
rect -15672 -8792 -15652 -8728
rect -16824 -8808 -15652 -8792
rect -16824 -8872 -15736 -8808
rect -15672 -8872 -15652 -8808
rect -16824 -8888 -15652 -8872
rect -16824 -8952 -15736 -8888
rect -15672 -8952 -15652 -8888
rect -16824 -8968 -15652 -8952
rect -16824 -9032 -15736 -8968
rect -15672 -9032 -15652 -8968
rect -16824 -9048 -15652 -9032
rect -16824 -9112 -15736 -9048
rect -15672 -9112 -15652 -9048
rect -16824 -9128 -15652 -9112
rect -16824 -9192 -15736 -9128
rect -15672 -9192 -15652 -9128
rect -16824 -9208 -15652 -9192
rect -16824 -9272 -15736 -9208
rect -15672 -9272 -15652 -9208
rect -16824 -9288 -15652 -9272
rect -16824 -9352 -15736 -9288
rect -15672 -9352 -15652 -9288
rect -16824 -9400 -15652 -9352
rect -15412 -8568 -14240 -8520
rect -15412 -8632 -14324 -8568
rect -14260 -8632 -14240 -8568
rect -15412 -8648 -14240 -8632
rect -15412 -8712 -14324 -8648
rect -14260 -8712 -14240 -8648
rect -15412 -8728 -14240 -8712
rect -15412 -8792 -14324 -8728
rect -14260 -8792 -14240 -8728
rect -15412 -8808 -14240 -8792
rect -15412 -8872 -14324 -8808
rect -14260 -8872 -14240 -8808
rect -15412 -8888 -14240 -8872
rect -15412 -8952 -14324 -8888
rect -14260 -8952 -14240 -8888
rect -15412 -8968 -14240 -8952
rect -15412 -9032 -14324 -8968
rect -14260 -9032 -14240 -8968
rect -15412 -9048 -14240 -9032
rect -15412 -9112 -14324 -9048
rect -14260 -9112 -14240 -9048
rect -15412 -9128 -14240 -9112
rect -15412 -9192 -14324 -9128
rect -14260 -9192 -14240 -9128
rect -15412 -9208 -14240 -9192
rect -15412 -9272 -14324 -9208
rect -14260 -9272 -14240 -9208
rect -15412 -9288 -14240 -9272
rect -15412 -9352 -14324 -9288
rect -14260 -9352 -14240 -9288
rect -15412 -9400 -14240 -9352
rect -14000 -8568 -12828 -8520
rect -14000 -8632 -12912 -8568
rect -12848 -8632 -12828 -8568
rect -14000 -8648 -12828 -8632
rect -14000 -8712 -12912 -8648
rect -12848 -8712 -12828 -8648
rect -14000 -8728 -12828 -8712
rect -14000 -8792 -12912 -8728
rect -12848 -8792 -12828 -8728
rect -14000 -8808 -12828 -8792
rect -14000 -8872 -12912 -8808
rect -12848 -8872 -12828 -8808
rect -14000 -8888 -12828 -8872
rect -14000 -8952 -12912 -8888
rect -12848 -8952 -12828 -8888
rect -14000 -8968 -12828 -8952
rect -14000 -9032 -12912 -8968
rect -12848 -9032 -12828 -8968
rect -14000 -9048 -12828 -9032
rect -14000 -9112 -12912 -9048
rect -12848 -9112 -12828 -9048
rect -14000 -9128 -12828 -9112
rect -14000 -9192 -12912 -9128
rect -12848 -9192 -12828 -9128
rect -14000 -9208 -12828 -9192
rect -14000 -9272 -12912 -9208
rect -12848 -9272 -12828 -9208
rect -14000 -9288 -12828 -9272
rect -14000 -9352 -12912 -9288
rect -12848 -9352 -12828 -9288
rect -14000 -9400 -12828 -9352
rect -12588 -8568 -11416 -8520
rect -12588 -8632 -11500 -8568
rect -11436 -8632 -11416 -8568
rect -12588 -8648 -11416 -8632
rect -12588 -8712 -11500 -8648
rect -11436 -8712 -11416 -8648
rect -12588 -8728 -11416 -8712
rect -12588 -8792 -11500 -8728
rect -11436 -8792 -11416 -8728
rect -12588 -8808 -11416 -8792
rect -12588 -8872 -11500 -8808
rect -11436 -8872 -11416 -8808
rect -12588 -8888 -11416 -8872
rect -12588 -8952 -11500 -8888
rect -11436 -8952 -11416 -8888
rect -12588 -8968 -11416 -8952
rect -12588 -9032 -11500 -8968
rect -11436 -9032 -11416 -8968
rect -12588 -9048 -11416 -9032
rect -12588 -9112 -11500 -9048
rect -11436 -9112 -11416 -9048
rect -12588 -9128 -11416 -9112
rect -12588 -9192 -11500 -9128
rect -11436 -9192 -11416 -9128
rect -12588 -9208 -11416 -9192
rect -12588 -9272 -11500 -9208
rect -11436 -9272 -11416 -9208
rect -12588 -9288 -11416 -9272
rect -12588 -9352 -11500 -9288
rect -11436 -9352 -11416 -9288
rect -12588 -9400 -11416 -9352
rect -11176 -8568 -10004 -8520
rect -11176 -8632 -10088 -8568
rect -10024 -8632 -10004 -8568
rect -11176 -8648 -10004 -8632
rect -11176 -8712 -10088 -8648
rect -10024 -8712 -10004 -8648
rect -11176 -8728 -10004 -8712
rect -11176 -8792 -10088 -8728
rect -10024 -8792 -10004 -8728
rect -11176 -8808 -10004 -8792
rect -11176 -8872 -10088 -8808
rect -10024 -8872 -10004 -8808
rect -11176 -8888 -10004 -8872
rect -11176 -8952 -10088 -8888
rect -10024 -8952 -10004 -8888
rect -11176 -8968 -10004 -8952
rect -11176 -9032 -10088 -8968
rect -10024 -9032 -10004 -8968
rect -11176 -9048 -10004 -9032
rect -11176 -9112 -10088 -9048
rect -10024 -9112 -10004 -9048
rect -11176 -9128 -10004 -9112
rect -11176 -9192 -10088 -9128
rect -10024 -9192 -10004 -9128
rect -11176 -9208 -10004 -9192
rect -11176 -9272 -10088 -9208
rect -10024 -9272 -10004 -9208
rect -11176 -9288 -10004 -9272
rect -11176 -9352 -10088 -9288
rect -10024 -9352 -10004 -9288
rect -11176 -9400 -10004 -9352
rect -9764 -8568 -8592 -8520
rect -9764 -8632 -8676 -8568
rect -8612 -8632 -8592 -8568
rect -9764 -8648 -8592 -8632
rect -9764 -8712 -8676 -8648
rect -8612 -8712 -8592 -8648
rect -9764 -8728 -8592 -8712
rect -9764 -8792 -8676 -8728
rect -8612 -8792 -8592 -8728
rect -9764 -8808 -8592 -8792
rect -9764 -8872 -8676 -8808
rect -8612 -8872 -8592 -8808
rect -9764 -8888 -8592 -8872
rect -9764 -8952 -8676 -8888
rect -8612 -8952 -8592 -8888
rect -9764 -8968 -8592 -8952
rect -9764 -9032 -8676 -8968
rect -8612 -9032 -8592 -8968
rect -9764 -9048 -8592 -9032
rect -9764 -9112 -8676 -9048
rect -8612 -9112 -8592 -9048
rect -9764 -9128 -8592 -9112
rect -9764 -9192 -8676 -9128
rect -8612 -9192 -8592 -9128
rect -9764 -9208 -8592 -9192
rect -9764 -9272 -8676 -9208
rect -8612 -9272 -8592 -9208
rect -9764 -9288 -8592 -9272
rect -9764 -9352 -8676 -9288
rect -8612 -9352 -8592 -9288
rect -9764 -9400 -8592 -9352
rect -8352 -8568 -7180 -8520
rect -8352 -8632 -7264 -8568
rect -7200 -8632 -7180 -8568
rect -8352 -8648 -7180 -8632
rect -8352 -8712 -7264 -8648
rect -7200 -8712 -7180 -8648
rect -8352 -8728 -7180 -8712
rect -8352 -8792 -7264 -8728
rect -7200 -8792 -7180 -8728
rect -8352 -8808 -7180 -8792
rect -8352 -8872 -7264 -8808
rect -7200 -8872 -7180 -8808
rect -8352 -8888 -7180 -8872
rect -8352 -8952 -7264 -8888
rect -7200 -8952 -7180 -8888
rect -8352 -8968 -7180 -8952
rect -8352 -9032 -7264 -8968
rect -7200 -9032 -7180 -8968
rect -8352 -9048 -7180 -9032
rect -8352 -9112 -7264 -9048
rect -7200 -9112 -7180 -9048
rect -8352 -9128 -7180 -9112
rect -8352 -9192 -7264 -9128
rect -7200 -9192 -7180 -9128
rect -8352 -9208 -7180 -9192
rect -8352 -9272 -7264 -9208
rect -7200 -9272 -7180 -9208
rect -8352 -9288 -7180 -9272
rect -8352 -9352 -7264 -9288
rect -7200 -9352 -7180 -9288
rect -8352 -9400 -7180 -9352
rect -6940 -8568 -5768 -8520
rect -6940 -8632 -5852 -8568
rect -5788 -8632 -5768 -8568
rect -6940 -8648 -5768 -8632
rect -6940 -8712 -5852 -8648
rect -5788 -8712 -5768 -8648
rect -6940 -8728 -5768 -8712
rect -6940 -8792 -5852 -8728
rect -5788 -8792 -5768 -8728
rect -6940 -8808 -5768 -8792
rect -6940 -8872 -5852 -8808
rect -5788 -8872 -5768 -8808
rect -6940 -8888 -5768 -8872
rect -6940 -8952 -5852 -8888
rect -5788 -8952 -5768 -8888
rect -6940 -8968 -5768 -8952
rect -6940 -9032 -5852 -8968
rect -5788 -9032 -5768 -8968
rect -6940 -9048 -5768 -9032
rect -6940 -9112 -5852 -9048
rect -5788 -9112 -5768 -9048
rect -6940 -9128 -5768 -9112
rect -6940 -9192 -5852 -9128
rect -5788 -9192 -5768 -9128
rect -6940 -9208 -5768 -9192
rect -6940 -9272 -5852 -9208
rect -5788 -9272 -5768 -9208
rect -6940 -9288 -5768 -9272
rect -6940 -9352 -5852 -9288
rect -5788 -9352 -5768 -9288
rect -6940 -9400 -5768 -9352
rect -5528 -8568 -4356 -8520
rect -5528 -8632 -4440 -8568
rect -4376 -8632 -4356 -8568
rect -5528 -8648 -4356 -8632
rect -5528 -8712 -4440 -8648
rect -4376 -8712 -4356 -8648
rect -5528 -8728 -4356 -8712
rect -5528 -8792 -4440 -8728
rect -4376 -8792 -4356 -8728
rect -5528 -8808 -4356 -8792
rect -5528 -8872 -4440 -8808
rect -4376 -8872 -4356 -8808
rect -5528 -8888 -4356 -8872
rect -5528 -8952 -4440 -8888
rect -4376 -8952 -4356 -8888
rect -5528 -8968 -4356 -8952
rect -5528 -9032 -4440 -8968
rect -4376 -9032 -4356 -8968
rect -5528 -9048 -4356 -9032
rect -5528 -9112 -4440 -9048
rect -4376 -9112 -4356 -9048
rect -5528 -9128 -4356 -9112
rect -5528 -9192 -4440 -9128
rect -4376 -9192 -4356 -9128
rect -5528 -9208 -4356 -9192
rect -5528 -9272 -4440 -9208
rect -4376 -9272 -4356 -9208
rect -5528 -9288 -4356 -9272
rect -5528 -9352 -4440 -9288
rect -4376 -9352 -4356 -9288
rect -5528 -9400 -4356 -9352
rect -4116 -8568 -2944 -8520
rect -4116 -8632 -3028 -8568
rect -2964 -8632 -2944 -8568
rect -4116 -8648 -2944 -8632
rect -4116 -8712 -3028 -8648
rect -2964 -8712 -2944 -8648
rect -4116 -8728 -2944 -8712
rect -4116 -8792 -3028 -8728
rect -2964 -8792 -2944 -8728
rect -4116 -8808 -2944 -8792
rect -4116 -8872 -3028 -8808
rect -2964 -8872 -2944 -8808
rect -4116 -8888 -2944 -8872
rect -4116 -8952 -3028 -8888
rect -2964 -8952 -2944 -8888
rect -4116 -8968 -2944 -8952
rect -4116 -9032 -3028 -8968
rect -2964 -9032 -2944 -8968
rect -4116 -9048 -2944 -9032
rect -4116 -9112 -3028 -9048
rect -2964 -9112 -2944 -9048
rect -4116 -9128 -2944 -9112
rect -4116 -9192 -3028 -9128
rect -2964 -9192 -2944 -9128
rect -4116 -9208 -2944 -9192
rect -4116 -9272 -3028 -9208
rect -2964 -9272 -2944 -9208
rect -4116 -9288 -2944 -9272
rect -4116 -9352 -3028 -9288
rect -2964 -9352 -2944 -9288
rect -4116 -9400 -2944 -9352
rect -2704 -8568 -1532 -8520
rect -2704 -8632 -1616 -8568
rect -1552 -8632 -1532 -8568
rect -2704 -8648 -1532 -8632
rect -2704 -8712 -1616 -8648
rect -1552 -8712 -1532 -8648
rect -2704 -8728 -1532 -8712
rect -2704 -8792 -1616 -8728
rect -1552 -8792 -1532 -8728
rect -2704 -8808 -1532 -8792
rect -2704 -8872 -1616 -8808
rect -1552 -8872 -1532 -8808
rect -2704 -8888 -1532 -8872
rect -2704 -8952 -1616 -8888
rect -1552 -8952 -1532 -8888
rect -2704 -8968 -1532 -8952
rect -2704 -9032 -1616 -8968
rect -1552 -9032 -1532 -8968
rect -2704 -9048 -1532 -9032
rect -2704 -9112 -1616 -9048
rect -1552 -9112 -1532 -9048
rect -2704 -9128 -1532 -9112
rect -2704 -9192 -1616 -9128
rect -1552 -9192 -1532 -9128
rect -2704 -9208 -1532 -9192
rect -2704 -9272 -1616 -9208
rect -1552 -9272 -1532 -9208
rect -2704 -9288 -1532 -9272
rect -2704 -9352 -1616 -9288
rect -1552 -9352 -1532 -9288
rect -2704 -9400 -1532 -9352
rect -1292 -8568 -120 -8520
rect -1292 -8632 -204 -8568
rect -140 -8632 -120 -8568
rect -1292 -8648 -120 -8632
rect -1292 -8712 -204 -8648
rect -140 -8712 -120 -8648
rect -1292 -8728 -120 -8712
rect -1292 -8792 -204 -8728
rect -140 -8792 -120 -8728
rect -1292 -8808 -120 -8792
rect -1292 -8872 -204 -8808
rect -140 -8872 -120 -8808
rect -1292 -8888 -120 -8872
rect -1292 -8952 -204 -8888
rect -140 -8952 -120 -8888
rect -1292 -8968 -120 -8952
rect -1292 -9032 -204 -8968
rect -140 -9032 -120 -8968
rect -1292 -9048 -120 -9032
rect -1292 -9112 -204 -9048
rect -140 -9112 -120 -9048
rect -1292 -9128 -120 -9112
rect -1292 -9192 -204 -9128
rect -140 -9192 -120 -9128
rect -1292 -9208 -120 -9192
rect -1292 -9272 -204 -9208
rect -140 -9272 -120 -9208
rect -1292 -9288 -120 -9272
rect -1292 -9352 -204 -9288
rect -140 -9352 -120 -9288
rect -1292 -9400 -120 -9352
rect 120 -8568 1292 -8520
rect 120 -8632 1208 -8568
rect 1272 -8632 1292 -8568
rect 120 -8648 1292 -8632
rect 120 -8712 1208 -8648
rect 1272 -8712 1292 -8648
rect 120 -8728 1292 -8712
rect 120 -8792 1208 -8728
rect 1272 -8792 1292 -8728
rect 120 -8808 1292 -8792
rect 120 -8872 1208 -8808
rect 1272 -8872 1292 -8808
rect 120 -8888 1292 -8872
rect 120 -8952 1208 -8888
rect 1272 -8952 1292 -8888
rect 120 -8968 1292 -8952
rect 120 -9032 1208 -8968
rect 1272 -9032 1292 -8968
rect 120 -9048 1292 -9032
rect 120 -9112 1208 -9048
rect 1272 -9112 1292 -9048
rect 120 -9128 1292 -9112
rect 120 -9192 1208 -9128
rect 1272 -9192 1292 -9128
rect 120 -9208 1292 -9192
rect 120 -9272 1208 -9208
rect 1272 -9272 1292 -9208
rect 120 -9288 1292 -9272
rect 120 -9352 1208 -9288
rect 1272 -9352 1292 -9288
rect 120 -9400 1292 -9352
rect 1532 -8568 2704 -8520
rect 1532 -8632 2620 -8568
rect 2684 -8632 2704 -8568
rect 1532 -8648 2704 -8632
rect 1532 -8712 2620 -8648
rect 2684 -8712 2704 -8648
rect 1532 -8728 2704 -8712
rect 1532 -8792 2620 -8728
rect 2684 -8792 2704 -8728
rect 1532 -8808 2704 -8792
rect 1532 -8872 2620 -8808
rect 2684 -8872 2704 -8808
rect 1532 -8888 2704 -8872
rect 1532 -8952 2620 -8888
rect 2684 -8952 2704 -8888
rect 1532 -8968 2704 -8952
rect 1532 -9032 2620 -8968
rect 2684 -9032 2704 -8968
rect 1532 -9048 2704 -9032
rect 1532 -9112 2620 -9048
rect 2684 -9112 2704 -9048
rect 1532 -9128 2704 -9112
rect 1532 -9192 2620 -9128
rect 2684 -9192 2704 -9128
rect 1532 -9208 2704 -9192
rect 1532 -9272 2620 -9208
rect 2684 -9272 2704 -9208
rect 1532 -9288 2704 -9272
rect 1532 -9352 2620 -9288
rect 2684 -9352 2704 -9288
rect 1532 -9400 2704 -9352
rect 2944 -8568 4116 -8520
rect 2944 -8632 4032 -8568
rect 4096 -8632 4116 -8568
rect 2944 -8648 4116 -8632
rect 2944 -8712 4032 -8648
rect 4096 -8712 4116 -8648
rect 2944 -8728 4116 -8712
rect 2944 -8792 4032 -8728
rect 4096 -8792 4116 -8728
rect 2944 -8808 4116 -8792
rect 2944 -8872 4032 -8808
rect 4096 -8872 4116 -8808
rect 2944 -8888 4116 -8872
rect 2944 -8952 4032 -8888
rect 4096 -8952 4116 -8888
rect 2944 -8968 4116 -8952
rect 2944 -9032 4032 -8968
rect 4096 -9032 4116 -8968
rect 2944 -9048 4116 -9032
rect 2944 -9112 4032 -9048
rect 4096 -9112 4116 -9048
rect 2944 -9128 4116 -9112
rect 2944 -9192 4032 -9128
rect 4096 -9192 4116 -9128
rect 2944 -9208 4116 -9192
rect 2944 -9272 4032 -9208
rect 4096 -9272 4116 -9208
rect 2944 -9288 4116 -9272
rect 2944 -9352 4032 -9288
rect 4096 -9352 4116 -9288
rect 2944 -9400 4116 -9352
rect 4356 -8568 5528 -8520
rect 4356 -8632 5444 -8568
rect 5508 -8632 5528 -8568
rect 4356 -8648 5528 -8632
rect 4356 -8712 5444 -8648
rect 5508 -8712 5528 -8648
rect 4356 -8728 5528 -8712
rect 4356 -8792 5444 -8728
rect 5508 -8792 5528 -8728
rect 4356 -8808 5528 -8792
rect 4356 -8872 5444 -8808
rect 5508 -8872 5528 -8808
rect 4356 -8888 5528 -8872
rect 4356 -8952 5444 -8888
rect 5508 -8952 5528 -8888
rect 4356 -8968 5528 -8952
rect 4356 -9032 5444 -8968
rect 5508 -9032 5528 -8968
rect 4356 -9048 5528 -9032
rect 4356 -9112 5444 -9048
rect 5508 -9112 5528 -9048
rect 4356 -9128 5528 -9112
rect 4356 -9192 5444 -9128
rect 5508 -9192 5528 -9128
rect 4356 -9208 5528 -9192
rect 4356 -9272 5444 -9208
rect 5508 -9272 5528 -9208
rect 4356 -9288 5528 -9272
rect 4356 -9352 5444 -9288
rect 5508 -9352 5528 -9288
rect 4356 -9400 5528 -9352
rect 5768 -8568 6940 -8520
rect 5768 -8632 6856 -8568
rect 6920 -8632 6940 -8568
rect 5768 -8648 6940 -8632
rect 5768 -8712 6856 -8648
rect 6920 -8712 6940 -8648
rect 5768 -8728 6940 -8712
rect 5768 -8792 6856 -8728
rect 6920 -8792 6940 -8728
rect 5768 -8808 6940 -8792
rect 5768 -8872 6856 -8808
rect 6920 -8872 6940 -8808
rect 5768 -8888 6940 -8872
rect 5768 -8952 6856 -8888
rect 6920 -8952 6940 -8888
rect 5768 -8968 6940 -8952
rect 5768 -9032 6856 -8968
rect 6920 -9032 6940 -8968
rect 5768 -9048 6940 -9032
rect 5768 -9112 6856 -9048
rect 6920 -9112 6940 -9048
rect 5768 -9128 6940 -9112
rect 5768 -9192 6856 -9128
rect 6920 -9192 6940 -9128
rect 5768 -9208 6940 -9192
rect 5768 -9272 6856 -9208
rect 6920 -9272 6940 -9208
rect 5768 -9288 6940 -9272
rect 5768 -9352 6856 -9288
rect 6920 -9352 6940 -9288
rect 5768 -9400 6940 -9352
rect 7180 -8568 8352 -8520
rect 7180 -8632 8268 -8568
rect 8332 -8632 8352 -8568
rect 7180 -8648 8352 -8632
rect 7180 -8712 8268 -8648
rect 8332 -8712 8352 -8648
rect 7180 -8728 8352 -8712
rect 7180 -8792 8268 -8728
rect 8332 -8792 8352 -8728
rect 7180 -8808 8352 -8792
rect 7180 -8872 8268 -8808
rect 8332 -8872 8352 -8808
rect 7180 -8888 8352 -8872
rect 7180 -8952 8268 -8888
rect 8332 -8952 8352 -8888
rect 7180 -8968 8352 -8952
rect 7180 -9032 8268 -8968
rect 8332 -9032 8352 -8968
rect 7180 -9048 8352 -9032
rect 7180 -9112 8268 -9048
rect 8332 -9112 8352 -9048
rect 7180 -9128 8352 -9112
rect 7180 -9192 8268 -9128
rect 8332 -9192 8352 -9128
rect 7180 -9208 8352 -9192
rect 7180 -9272 8268 -9208
rect 8332 -9272 8352 -9208
rect 7180 -9288 8352 -9272
rect 7180 -9352 8268 -9288
rect 8332 -9352 8352 -9288
rect 7180 -9400 8352 -9352
rect 8592 -8568 9764 -8520
rect 8592 -8632 9680 -8568
rect 9744 -8632 9764 -8568
rect 8592 -8648 9764 -8632
rect 8592 -8712 9680 -8648
rect 9744 -8712 9764 -8648
rect 8592 -8728 9764 -8712
rect 8592 -8792 9680 -8728
rect 9744 -8792 9764 -8728
rect 8592 -8808 9764 -8792
rect 8592 -8872 9680 -8808
rect 9744 -8872 9764 -8808
rect 8592 -8888 9764 -8872
rect 8592 -8952 9680 -8888
rect 9744 -8952 9764 -8888
rect 8592 -8968 9764 -8952
rect 8592 -9032 9680 -8968
rect 9744 -9032 9764 -8968
rect 8592 -9048 9764 -9032
rect 8592 -9112 9680 -9048
rect 9744 -9112 9764 -9048
rect 8592 -9128 9764 -9112
rect 8592 -9192 9680 -9128
rect 9744 -9192 9764 -9128
rect 8592 -9208 9764 -9192
rect 8592 -9272 9680 -9208
rect 9744 -9272 9764 -9208
rect 8592 -9288 9764 -9272
rect 8592 -9352 9680 -9288
rect 9744 -9352 9764 -9288
rect 8592 -9400 9764 -9352
rect 10004 -8568 11176 -8520
rect 10004 -8632 11092 -8568
rect 11156 -8632 11176 -8568
rect 10004 -8648 11176 -8632
rect 10004 -8712 11092 -8648
rect 11156 -8712 11176 -8648
rect 10004 -8728 11176 -8712
rect 10004 -8792 11092 -8728
rect 11156 -8792 11176 -8728
rect 10004 -8808 11176 -8792
rect 10004 -8872 11092 -8808
rect 11156 -8872 11176 -8808
rect 10004 -8888 11176 -8872
rect 10004 -8952 11092 -8888
rect 11156 -8952 11176 -8888
rect 10004 -8968 11176 -8952
rect 10004 -9032 11092 -8968
rect 11156 -9032 11176 -8968
rect 10004 -9048 11176 -9032
rect 10004 -9112 11092 -9048
rect 11156 -9112 11176 -9048
rect 10004 -9128 11176 -9112
rect 10004 -9192 11092 -9128
rect 11156 -9192 11176 -9128
rect 10004 -9208 11176 -9192
rect 10004 -9272 11092 -9208
rect 11156 -9272 11176 -9208
rect 10004 -9288 11176 -9272
rect 10004 -9352 11092 -9288
rect 11156 -9352 11176 -9288
rect 10004 -9400 11176 -9352
rect 11416 -8568 12588 -8520
rect 11416 -8632 12504 -8568
rect 12568 -8632 12588 -8568
rect 11416 -8648 12588 -8632
rect 11416 -8712 12504 -8648
rect 12568 -8712 12588 -8648
rect 11416 -8728 12588 -8712
rect 11416 -8792 12504 -8728
rect 12568 -8792 12588 -8728
rect 11416 -8808 12588 -8792
rect 11416 -8872 12504 -8808
rect 12568 -8872 12588 -8808
rect 11416 -8888 12588 -8872
rect 11416 -8952 12504 -8888
rect 12568 -8952 12588 -8888
rect 11416 -8968 12588 -8952
rect 11416 -9032 12504 -8968
rect 12568 -9032 12588 -8968
rect 11416 -9048 12588 -9032
rect 11416 -9112 12504 -9048
rect 12568 -9112 12588 -9048
rect 11416 -9128 12588 -9112
rect 11416 -9192 12504 -9128
rect 12568 -9192 12588 -9128
rect 11416 -9208 12588 -9192
rect 11416 -9272 12504 -9208
rect 12568 -9272 12588 -9208
rect 11416 -9288 12588 -9272
rect 11416 -9352 12504 -9288
rect 12568 -9352 12588 -9288
rect 11416 -9400 12588 -9352
rect 12828 -8568 14000 -8520
rect 12828 -8632 13916 -8568
rect 13980 -8632 14000 -8568
rect 12828 -8648 14000 -8632
rect 12828 -8712 13916 -8648
rect 13980 -8712 14000 -8648
rect 12828 -8728 14000 -8712
rect 12828 -8792 13916 -8728
rect 13980 -8792 14000 -8728
rect 12828 -8808 14000 -8792
rect 12828 -8872 13916 -8808
rect 13980 -8872 14000 -8808
rect 12828 -8888 14000 -8872
rect 12828 -8952 13916 -8888
rect 13980 -8952 14000 -8888
rect 12828 -8968 14000 -8952
rect 12828 -9032 13916 -8968
rect 13980 -9032 14000 -8968
rect 12828 -9048 14000 -9032
rect 12828 -9112 13916 -9048
rect 13980 -9112 14000 -9048
rect 12828 -9128 14000 -9112
rect 12828 -9192 13916 -9128
rect 13980 -9192 14000 -9128
rect 12828 -9208 14000 -9192
rect 12828 -9272 13916 -9208
rect 13980 -9272 14000 -9208
rect 12828 -9288 14000 -9272
rect 12828 -9352 13916 -9288
rect 13980 -9352 14000 -9288
rect 12828 -9400 14000 -9352
rect 14240 -8568 15412 -8520
rect 14240 -8632 15328 -8568
rect 15392 -8632 15412 -8568
rect 14240 -8648 15412 -8632
rect 14240 -8712 15328 -8648
rect 15392 -8712 15412 -8648
rect 14240 -8728 15412 -8712
rect 14240 -8792 15328 -8728
rect 15392 -8792 15412 -8728
rect 14240 -8808 15412 -8792
rect 14240 -8872 15328 -8808
rect 15392 -8872 15412 -8808
rect 14240 -8888 15412 -8872
rect 14240 -8952 15328 -8888
rect 15392 -8952 15412 -8888
rect 14240 -8968 15412 -8952
rect 14240 -9032 15328 -8968
rect 15392 -9032 15412 -8968
rect 14240 -9048 15412 -9032
rect 14240 -9112 15328 -9048
rect 15392 -9112 15412 -9048
rect 14240 -9128 15412 -9112
rect 14240 -9192 15328 -9128
rect 15392 -9192 15412 -9128
rect 14240 -9208 15412 -9192
rect 14240 -9272 15328 -9208
rect 15392 -9272 15412 -9208
rect 14240 -9288 15412 -9272
rect 14240 -9352 15328 -9288
rect 15392 -9352 15412 -9288
rect 14240 -9400 15412 -9352
rect 15652 -8568 16824 -8520
rect 15652 -8632 16740 -8568
rect 16804 -8632 16824 -8568
rect 15652 -8648 16824 -8632
rect 15652 -8712 16740 -8648
rect 16804 -8712 16824 -8648
rect 15652 -8728 16824 -8712
rect 15652 -8792 16740 -8728
rect 16804 -8792 16824 -8728
rect 15652 -8808 16824 -8792
rect 15652 -8872 16740 -8808
rect 16804 -8872 16824 -8808
rect 15652 -8888 16824 -8872
rect 15652 -8952 16740 -8888
rect 16804 -8952 16824 -8888
rect 15652 -8968 16824 -8952
rect 15652 -9032 16740 -8968
rect 16804 -9032 16824 -8968
rect 15652 -9048 16824 -9032
rect 15652 -9112 16740 -9048
rect 16804 -9112 16824 -9048
rect 15652 -9128 16824 -9112
rect 15652 -9192 16740 -9128
rect 16804 -9192 16824 -9128
rect 15652 -9208 16824 -9192
rect 15652 -9272 16740 -9208
rect 16804 -9272 16824 -9208
rect 15652 -9288 16824 -9272
rect 15652 -9352 16740 -9288
rect 16804 -9352 16824 -9288
rect 15652 -9400 16824 -9352
rect 17064 -8568 18236 -8520
rect 17064 -8632 18152 -8568
rect 18216 -8632 18236 -8568
rect 17064 -8648 18236 -8632
rect 17064 -8712 18152 -8648
rect 18216 -8712 18236 -8648
rect 17064 -8728 18236 -8712
rect 17064 -8792 18152 -8728
rect 18216 -8792 18236 -8728
rect 17064 -8808 18236 -8792
rect 17064 -8872 18152 -8808
rect 18216 -8872 18236 -8808
rect 17064 -8888 18236 -8872
rect 17064 -8952 18152 -8888
rect 18216 -8952 18236 -8888
rect 17064 -8968 18236 -8952
rect 17064 -9032 18152 -8968
rect 18216 -9032 18236 -8968
rect 17064 -9048 18236 -9032
rect 17064 -9112 18152 -9048
rect 18216 -9112 18236 -9048
rect 17064 -9128 18236 -9112
rect 17064 -9192 18152 -9128
rect 18216 -9192 18236 -9128
rect 17064 -9208 18236 -9192
rect 17064 -9272 18152 -9208
rect 18216 -9272 18236 -9208
rect 17064 -9288 18236 -9272
rect 17064 -9352 18152 -9288
rect 18216 -9352 18236 -9288
rect 17064 -9400 18236 -9352
rect 18476 -8568 19648 -8520
rect 18476 -8632 19564 -8568
rect 19628 -8632 19648 -8568
rect 18476 -8648 19648 -8632
rect 18476 -8712 19564 -8648
rect 19628 -8712 19648 -8648
rect 18476 -8728 19648 -8712
rect 18476 -8792 19564 -8728
rect 19628 -8792 19648 -8728
rect 18476 -8808 19648 -8792
rect 18476 -8872 19564 -8808
rect 19628 -8872 19648 -8808
rect 18476 -8888 19648 -8872
rect 18476 -8952 19564 -8888
rect 19628 -8952 19648 -8888
rect 18476 -8968 19648 -8952
rect 18476 -9032 19564 -8968
rect 19628 -9032 19648 -8968
rect 18476 -9048 19648 -9032
rect 18476 -9112 19564 -9048
rect 19628 -9112 19648 -9048
rect 18476 -9128 19648 -9112
rect 18476 -9192 19564 -9128
rect 19628 -9192 19648 -9128
rect 18476 -9208 19648 -9192
rect 18476 -9272 19564 -9208
rect 19628 -9272 19648 -9208
rect 18476 -9288 19648 -9272
rect 18476 -9352 19564 -9288
rect 19628 -9352 19648 -9288
rect 18476 -9400 19648 -9352
rect 19888 -8568 21060 -8520
rect 19888 -8632 20976 -8568
rect 21040 -8632 21060 -8568
rect 19888 -8648 21060 -8632
rect 19888 -8712 20976 -8648
rect 21040 -8712 21060 -8648
rect 19888 -8728 21060 -8712
rect 19888 -8792 20976 -8728
rect 21040 -8792 21060 -8728
rect 19888 -8808 21060 -8792
rect 19888 -8872 20976 -8808
rect 21040 -8872 21060 -8808
rect 19888 -8888 21060 -8872
rect 19888 -8952 20976 -8888
rect 21040 -8952 21060 -8888
rect 19888 -8968 21060 -8952
rect 19888 -9032 20976 -8968
rect 21040 -9032 21060 -8968
rect 19888 -9048 21060 -9032
rect 19888 -9112 20976 -9048
rect 21040 -9112 21060 -9048
rect 19888 -9128 21060 -9112
rect 19888 -9192 20976 -9128
rect 21040 -9192 21060 -9128
rect 19888 -9208 21060 -9192
rect 19888 -9272 20976 -9208
rect 21040 -9272 21060 -9208
rect 19888 -9288 21060 -9272
rect 19888 -9352 20976 -9288
rect 21040 -9352 21060 -9288
rect 19888 -9400 21060 -9352
rect 21300 -8568 22472 -8520
rect 21300 -8632 22388 -8568
rect 22452 -8632 22472 -8568
rect 21300 -8648 22472 -8632
rect 21300 -8712 22388 -8648
rect 22452 -8712 22472 -8648
rect 21300 -8728 22472 -8712
rect 21300 -8792 22388 -8728
rect 22452 -8792 22472 -8728
rect 21300 -8808 22472 -8792
rect 21300 -8872 22388 -8808
rect 22452 -8872 22472 -8808
rect 21300 -8888 22472 -8872
rect 21300 -8952 22388 -8888
rect 22452 -8952 22472 -8888
rect 21300 -8968 22472 -8952
rect 21300 -9032 22388 -8968
rect 22452 -9032 22472 -8968
rect 21300 -9048 22472 -9032
rect 21300 -9112 22388 -9048
rect 22452 -9112 22472 -9048
rect 21300 -9128 22472 -9112
rect 21300 -9192 22388 -9128
rect 22452 -9192 22472 -9128
rect 21300 -9208 22472 -9192
rect 21300 -9272 22388 -9208
rect 22452 -9272 22472 -9208
rect 21300 -9288 22472 -9272
rect 21300 -9352 22388 -9288
rect 22452 -9352 22472 -9288
rect 21300 -9400 22472 -9352
rect 22712 -8568 23884 -8520
rect 22712 -8632 23800 -8568
rect 23864 -8632 23884 -8568
rect 22712 -8648 23884 -8632
rect 22712 -8712 23800 -8648
rect 23864 -8712 23884 -8648
rect 22712 -8728 23884 -8712
rect 22712 -8792 23800 -8728
rect 23864 -8792 23884 -8728
rect 22712 -8808 23884 -8792
rect 22712 -8872 23800 -8808
rect 23864 -8872 23884 -8808
rect 22712 -8888 23884 -8872
rect 22712 -8952 23800 -8888
rect 23864 -8952 23884 -8888
rect 22712 -8968 23884 -8952
rect 22712 -9032 23800 -8968
rect 23864 -9032 23884 -8968
rect 22712 -9048 23884 -9032
rect 22712 -9112 23800 -9048
rect 23864 -9112 23884 -9048
rect 22712 -9128 23884 -9112
rect 22712 -9192 23800 -9128
rect 23864 -9192 23884 -9128
rect 22712 -9208 23884 -9192
rect 22712 -9272 23800 -9208
rect 23864 -9272 23884 -9208
rect 22712 -9288 23884 -9272
rect 22712 -9352 23800 -9288
rect 23864 -9352 23884 -9288
rect 22712 -9400 23884 -9352
rect -23884 -9688 -22712 -9640
rect -23884 -9752 -22796 -9688
rect -22732 -9752 -22712 -9688
rect -23884 -9768 -22712 -9752
rect -23884 -9832 -22796 -9768
rect -22732 -9832 -22712 -9768
rect -23884 -9848 -22712 -9832
rect -23884 -9912 -22796 -9848
rect -22732 -9912 -22712 -9848
rect -23884 -9928 -22712 -9912
rect -23884 -9992 -22796 -9928
rect -22732 -9992 -22712 -9928
rect -23884 -10008 -22712 -9992
rect -23884 -10072 -22796 -10008
rect -22732 -10072 -22712 -10008
rect -23884 -10088 -22712 -10072
rect -23884 -10152 -22796 -10088
rect -22732 -10152 -22712 -10088
rect -23884 -10168 -22712 -10152
rect -23884 -10232 -22796 -10168
rect -22732 -10232 -22712 -10168
rect -23884 -10248 -22712 -10232
rect -23884 -10312 -22796 -10248
rect -22732 -10312 -22712 -10248
rect -23884 -10328 -22712 -10312
rect -23884 -10392 -22796 -10328
rect -22732 -10392 -22712 -10328
rect -23884 -10408 -22712 -10392
rect -23884 -10472 -22796 -10408
rect -22732 -10472 -22712 -10408
rect -23884 -10520 -22712 -10472
rect -22472 -9688 -21300 -9640
rect -22472 -9752 -21384 -9688
rect -21320 -9752 -21300 -9688
rect -22472 -9768 -21300 -9752
rect -22472 -9832 -21384 -9768
rect -21320 -9832 -21300 -9768
rect -22472 -9848 -21300 -9832
rect -22472 -9912 -21384 -9848
rect -21320 -9912 -21300 -9848
rect -22472 -9928 -21300 -9912
rect -22472 -9992 -21384 -9928
rect -21320 -9992 -21300 -9928
rect -22472 -10008 -21300 -9992
rect -22472 -10072 -21384 -10008
rect -21320 -10072 -21300 -10008
rect -22472 -10088 -21300 -10072
rect -22472 -10152 -21384 -10088
rect -21320 -10152 -21300 -10088
rect -22472 -10168 -21300 -10152
rect -22472 -10232 -21384 -10168
rect -21320 -10232 -21300 -10168
rect -22472 -10248 -21300 -10232
rect -22472 -10312 -21384 -10248
rect -21320 -10312 -21300 -10248
rect -22472 -10328 -21300 -10312
rect -22472 -10392 -21384 -10328
rect -21320 -10392 -21300 -10328
rect -22472 -10408 -21300 -10392
rect -22472 -10472 -21384 -10408
rect -21320 -10472 -21300 -10408
rect -22472 -10520 -21300 -10472
rect -21060 -9688 -19888 -9640
rect -21060 -9752 -19972 -9688
rect -19908 -9752 -19888 -9688
rect -21060 -9768 -19888 -9752
rect -21060 -9832 -19972 -9768
rect -19908 -9832 -19888 -9768
rect -21060 -9848 -19888 -9832
rect -21060 -9912 -19972 -9848
rect -19908 -9912 -19888 -9848
rect -21060 -9928 -19888 -9912
rect -21060 -9992 -19972 -9928
rect -19908 -9992 -19888 -9928
rect -21060 -10008 -19888 -9992
rect -21060 -10072 -19972 -10008
rect -19908 -10072 -19888 -10008
rect -21060 -10088 -19888 -10072
rect -21060 -10152 -19972 -10088
rect -19908 -10152 -19888 -10088
rect -21060 -10168 -19888 -10152
rect -21060 -10232 -19972 -10168
rect -19908 -10232 -19888 -10168
rect -21060 -10248 -19888 -10232
rect -21060 -10312 -19972 -10248
rect -19908 -10312 -19888 -10248
rect -21060 -10328 -19888 -10312
rect -21060 -10392 -19972 -10328
rect -19908 -10392 -19888 -10328
rect -21060 -10408 -19888 -10392
rect -21060 -10472 -19972 -10408
rect -19908 -10472 -19888 -10408
rect -21060 -10520 -19888 -10472
rect -19648 -9688 -18476 -9640
rect -19648 -9752 -18560 -9688
rect -18496 -9752 -18476 -9688
rect -19648 -9768 -18476 -9752
rect -19648 -9832 -18560 -9768
rect -18496 -9832 -18476 -9768
rect -19648 -9848 -18476 -9832
rect -19648 -9912 -18560 -9848
rect -18496 -9912 -18476 -9848
rect -19648 -9928 -18476 -9912
rect -19648 -9992 -18560 -9928
rect -18496 -9992 -18476 -9928
rect -19648 -10008 -18476 -9992
rect -19648 -10072 -18560 -10008
rect -18496 -10072 -18476 -10008
rect -19648 -10088 -18476 -10072
rect -19648 -10152 -18560 -10088
rect -18496 -10152 -18476 -10088
rect -19648 -10168 -18476 -10152
rect -19648 -10232 -18560 -10168
rect -18496 -10232 -18476 -10168
rect -19648 -10248 -18476 -10232
rect -19648 -10312 -18560 -10248
rect -18496 -10312 -18476 -10248
rect -19648 -10328 -18476 -10312
rect -19648 -10392 -18560 -10328
rect -18496 -10392 -18476 -10328
rect -19648 -10408 -18476 -10392
rect -19648 -10472 -18560 -10408
rect -18496 -10472 -18476 -10408
rect -19648 -10520 -18476 -10472
rect -18236 -9688 -17064 -9640
rect -18236 -9752 -17148 -9688
rect -17084 -9752 -17064 -9688
rect -18236 -9768 -17064 -9752
rect -18236 -9832 -17148 -9768
rect -17084 -9832 -17064 -9768
rect -18236 -9848 -17064 -9832
rect -18236 -9912 -17148 -9848
rect -17084 -9912 -17064 -9848
rect -18236 -9928 -17064 -9912
rect -18236 -9992 -17148 -9928
rect -17084 -9992 -17064 -9928
rect -18236 -10008 -17064 -9992
rect -18236 -10072 -17148 -10008
rect -17084 -10072 -17064 -10008
rect -18236 -10088 -17064 -10072
rect -18236 -10152 -17148 -10088
rect -17084 -10152 -17064 -10088
rect -18236 -10168 -17064 -10152
rect -18236 -10232 -17148 -10168
rect -17084 -10232 -17064 -10168
rect -18236 -10248 -17064 -10232
rect -18236 -10312 -17148 -10248
rect -17084 -10312 -17064 -10248
rect -18236 -10328 -17064 -10312
rect -18236 -10392 -17148 -10328
rect -17084 -10392 -17064 -10328
rect -18236 -10408 -17064 -10392
rect -18236 -10472 -17148 -10408
rect -17084 -10472 -17064 -10408
rect -18236 -10520 -17064 -10472
rect -16824 -9688 -15652 -9640
rect -16824 -9752 -15736 -9688
rect -15672 -9752 -15652 -9688
rect -16824 -9768 -15652 -9752
rect -16824 -9832 -15736 -9768
rect -15672 -9832 -15652 -9768
rect -16824 -9848 -15652 -9832
rect -16824 -9912 -15736 -9848
rect -15672 -9912 -15652 -9848
rect -16824 -9928 -15652 -9912
rect -16824 -9992 -15736 -9928
rect -15672 -9992 -15652 -9928
rect -16824 -10008 -15652 -9992
rect -16824 -10072 -15736 -10008
rect -15672 -10072 -15652 -10008
rect -16824 -10088 -15652 -10072
rect -16824 -10152 -15736 -10088
rect -15672 -10152 -15652 -10088
rect -16824 -10168 -15652 -10152
rect -16824 -10232 -15736 -10168
rect -15672 -10232 -15652 -10168
rect -16824 -10248 -15652 -10232
rect -16824 -10312 -15736 -10248
rect -15672 -10312 -15652 -10248
rect -16824 -10328 -15652 -10312
rect -16824 -10392 -15736 -10328
rect -15672 -10392 -15652 -10328
rect -16824 -10408 -15652 -10392
rect -16824 -10472 -15736 -10408
rect -15672 -10472 -15652 -10408
rect -16824 -10520 -15652 -10472
rect -15412 -9688 -14240 -9640
rect -15412 -9752 -14324 -9688
rect -14260 -9752 -14240 -9688
rect -15412 -9768 -14240 -9752
rect -15412 -9832 -14324 -9768
rect -14260 -9832 -14240 -9768
rect -15412 -9848 -14240 -9832
rect -15412 -9912 -14324 -9848
rect -14260 -9912 -14240 -9848
rect -15412 -9928 -14240 -9912
rect -15412 -9992 -14324 -9928
rect -14260 -9992 -14240 -9928
rect -15412 -10008 -14240 -9992
rect -15412 -10072 -14324 -10008
rect -14260 -10072 -14240 -10008
rect -15412 -10088 -14240 -10072
rect -15412 -10152 -14324 -10088
rect -14260 -10152 -14240 -10088
rect -15412 -10168 -14240 -10152
rect -15412 -10232 -14324 -10168
rect -14260 -10232 -14240 -10168
rect -15412 -10248 -14240 -10232
rect -15412 -10312 -14324 -10248
rect -14260 -10312 -14240 -10248
rect -15412 -10328 -14240 -10312
rect -15412 -10392 -14324 -10328
rect -14260 -10392 -14240 -10328
rect -15412 -10408 -14240 -10392
rect -15412 -10472 -14324 -10408
rect -14260 -10472 -14240 -10408
rect -15412 -10520 -14240 -10472
rect -14000 -9688 -12828 -9640
rect -14000 -9752 -12912 -9688
rect -12848 -9752 -12828 -9688
rect -14000 -9768 -12828 -9752
rect -14000 -9832 -12912 -9768
rect -12848 -9832 -12828 -9768
rect -14000 -9848 -12828 -9832
rect -14000 -9912 -12912 -9848
rect -12848 -9912 -12828 -9848
rect -14000 -9928 -12828 -9912
rect -14000 -9992 -12912 -9928
rect -12848 -9992 -12828 -9928
rect -14000 -10008 -12828 -9992
rect -14000 -10072 -12912 -10008
rect -12848 -10072 -12828 -10008
rect -14000 -10088 -12828 -10072
rect -14000 -10152 -12912 -10088
rect -12848 -10152 -12828 -10088
rect -14000 -10168 -12828 -10152
rect -14000 -10232 -12912 -10168
rect -12848 -10232 -12828 -10168
rect -14000 -10248 -12828 -10232
rect -14000 -10312 -12912 -10248
rect -12848 -10312 -12828 -10248
rect -14000 -10328 -12828 -10312
rect -14000 -10392 -12912 -10328
rect -12848 -10392 -12828 -10328
rect -14000 -10408 -12828 -10392
rect -14000 -10472 -12912 -10408
rect -12848 -10472 -12828 -10408
rect -14000 -10520 -12828 -10472
rect -12588 -9688 -11416 -9640
rect -12588 -9752 -11500 -9688
rect -11436 -9752 -11416 -9688
rect -12588 -9768 -11416 -9752
rect -12588 -9832 -11500 -9768
rect -11436 -9832 -11416 -9768
rect -12588 -9848 -11416 -9832
rect -12588 -9912 -11500 -9848
rect -11436 -9912 -11416 -9848
rect -12588 -9928 -11416 -9912
rect -12588 -9992 -11500 -9928
rect -11436 -9992 -11416 -9928
rect -12588 -10008 -11416 -9992
rect -12588 -10072 -11500 -10008
rect -11436 -10072 -11416 -10008
rect -12588 -10088 -11416 -10072
rect -12588 -10152 -11500 -10088
rect -11436 -10152 -11416 -10088
rect -12588 -10168 -11416 -10152
rect -12588 -10232 -11500 -10168
rect -11436 -10232 -11416 -10168
rect -12588 -10248 -11416 -10232
rect -12588 -10312 -11500 -10248
rect -11436 -10312 -11416 -10248
rect -12588 -10328 -11416 -10312
rect -12588 -10392 -11500 -10328
rect -11436 -10392 -11416 -10328
rect -12588 -10408 -11416 -10392
rect -12588 -10472 -11500 -10408
rect -11436 -10472 -11416 -10408
rect -12588 -10520 -11416 -10472
rect -11176 -9688 -10004 -9640
rect -11176 -9752 -10088 -9688
rect -10024 -9752 -10004 -9688
rect -11176 -9768 -10004 -9752
rect -11176 -9832 -10088 -9768
rect -10024 -9832 -10004 -9768
rect -11176 -9848 -10004 -9832
rect -11176 -9912 -10088 -9848
rect -10024 -9912 -10004 -9848
rect -11176 -9928 -10004 -9912
rect -11176 -9992 -10088 -9928
rect -10024 -9992 -10004 -9928
rect -11176 -10008 -10004 -9992
rect -11176 -10072 -10088 -10008
rect -10024 -10072 -10004 -10008
rect -11176 -10088 -10004 -10072
rect -11176 -10152 -10088 -10088
rect -10024 -10152 -10004 -10088
rect -11176 -10168 -10004 -10152
rect -11176 -10232 -10088 -10168
rect -10024 -10232 -10004 -10168
rect -11176 -10248 -10004 -10232
rect -11176 -10312 -10088 -10248
rect -10024 -10312 -10004 -10248
rect -11176 -10328 -10004 -10312
rect -11176 -10392 -10088 -10328
rect -10024 -10392 -10004 -10328
rect -11176 -10408 -10004 -10392
rect -11176 -10472 -10088 -10408
rect -10024 -10472 -10004 -10408
rect -11176 -10520 -10004 -10472
rect -9764 -9688 -8592 -9640
rect -9764 -9752 -8676 -9688
rect -8612 -9752 -8592 -9688
rect -9764 -9768 -8592 -9752
rect -9764 -9832 -8676 -9768
rect -8612 -9832 -8592 -9768
rect -9764 -9848 -8592 -9832
rect -9764 -9912 -8676 -9848
rect -8612 -9912 -8592 -9848
rect -9764 -9928 -8592 -9912
rect -9764 -9992 -8676 -9928
rect -8612 -9992 -8592 -9928
rect -9764 -10008 -8592 -9992
rect -9764 -10072 -8676 -10008
rect -8612 -10072 -8592 -10008
rect -9764 -10088 -8592 -10072
rect -9764 -10152 -8676 -10088
rect -8612 -10152 -8592 -10088
rect -9764 -10168 -8592 -10152
rect -9764 -10232 -8676 -10168
rect -8612 -10232 -8592 -10168
rect -9764 -10248 -8592 -10232
rect -9764 -10312 -8676 -10248
rect -8612 -10312 -8592 -10248
rect -9764 -10328 -8592 -10312
rect -9764 -10392 -8676 -10328
rect -8612 -10392 -8592 -10328
rect -9764 -10408 -8592 -10392
rect -9764 -10472 -8676 -10408
rect -8612 -10472 -8592 -10408
rect -9764 -10520 -8592 -10472
rect -8352 -9688 -7180 -9640
rect -8352 -9752 -7264 -9688
rect -7200 -9752 -7180 -9688
rect -8352 -9768 -7180 -9752
rect -8352 -9832 -7264 -9768
rect -7200 -9832 -7180 -9768
rect -8352 -9848 -7180 -9832
rect -8352 -9912 -7264 -9848
rect -7200 -9912 -7180 -9848
rect -8352 -9928 -7180 -9912
rect -8352 -9992 -7264 -9928
rect -7200 -9992 -7180 -9928
rect -8352 -10008 -7180 -9992
rect -8352 -10072 -7264 -10008
rect -7200 -10072 -7180 -10008
rect -8352 -10088 -7180 -10072
rect -8352 -10152 -7264 -10088
rect -7200 -10152 -7180 -10088
rect -8352 -10168 -7180 -10152
rect -8352 -10232 -7264 -10168
rect -7200 -10232 -7180 -10168
rect -8352 -10248 -7180 -10232
rect -8352 -10312 -7264 -10248
rect -7200 -10312 -7180 -10248
rect -8352 -10328 -7180 -10312
rect -8352 -10392 -7264 -10328
rect -7200 -10392 -7180 -10328
rect -8352 -10408 -7180 -10392
rect -8352 -10472 -7264 -10408
rect -7200 -10472 -7180 -10408
rect -8352 -10520 -7180 -10472
rect -6940 -9688 -5768 -9640
rect -6940 -9752 -5852 -9688
rect -5788 -9752 -5768 -9688
rect -6940 -9768 -5768 -9752
rect -6940 -9832 -5852 -9768
rect -5788 -9832 -5768 -9768
rect -6940 -9848 -5768 -9832
rect -6940 -9912 -5852 -9848
rect -5788 -9912 -5768 -9848
rect -6940 -9928 -5768 -9912
rect -6940 -9992 -5852 -9928
rect -5788 -9992 -5768 -9928
rect -6940 -10008 -5768 -9992
rect -6940 -10072 -5852 -10008
rect -5788 -10072 -5768 -10008
rect -6940 -10088 -5768 -10072
rect -6940 -10152 -5852 -10088
rect -5788 -10152 -5768 -10088
rect -6940 -10168 -5768 -10152
rect -6940 -10232 -5852 -10168
rect -5788 -10232 -5768 -10168
rect -6940 -10248 -5768 -10232
rect -6940 -10312 -5852 -10248
rect -5788 -10312 -5768 -10248
rect -6940 -10328 -5768 -10312
rect -6940 -10392 -5852 -10328
rect -5788 -10392 -5768 -10328
rect -6940 -10408 -5768 -10392
rect -6940 -10472 -5852 -10408
rect -5788 -10472 -5768 -10408
rect -6940 -10520 -5768 -10472
rect -5528 -9688 -4356 -9640
rect -5528 -9752 -4440 -9688
rect -4376 -9752 -4356 -9688
rect -5528 -9768 -4356 -9752
rect -5528 -9832 -4440 -9768
rect -4376 -9832 -4356 -9768
rect -5528 -9848 -4356 -9832
rect -5528 -9912 -4440 -9848
rect -4376 -9912 -4356 -9848
rect -5528 -9928 -4356 -9912
rect -5528 -9992 -4440 -9928
rect -4376 -9992 -4356 -9928
rect -5528 -10008 -4356 -9992
rect -5528 -10072 -4440 -10008
rect -4376 -10072 -4356 -10008
rect -5528 -10088 -4356 -10072
rect -5528 -10152 -4440 -10088
rect -4376 -10152 -4356 -10088
rect -5528 -10168 -4356 -10152
rect -5528 -10232 -4440 -10168
rect -4376 -10232 -4356 -10168
rect -5528 -10248 -4356 -10232
rect -5528 -10312 -4440 -10248
rect -4376 -10312 -4356 -10248
rect -5528 -10328 -4356 -10312
rect -5528 -10392 -4440 -10328
rect -4376 -10392 -4356 -10328
rect -5528 -10408 -4356 -10392
rect -5528 -10472 -4440 -10408
rect -4376 -10472 -4356 -10408
rect -5528 -10520 -4356 -10472
rect -4116 -9688 -2944 -9640
rect -4116 -9752 -3028 -9688
rect -2964 -9752 -2944 -9688
rect -4116 -9768 -2944 -9752
rect -4116 -9832 -3028 -9768
rect -2964 -9832 -2944 -9768
rect -4116 -9848 -2944 -9832
rect -4116 -9912 -3028 -9848
rect -2964 -9912 -2944 -9848
rect -4116 -9928 -2944 -9912
rect -4116 -9992 -3028 -9928
rect -2964 -9992 -2944 -9928
rect -4116 -10008 -2944 -9992
rect -4116 -10072 -3028 -10008
rect -2964 -10072 -2944 -10008
rect -4116 -10088 -2944 -10072
rect -4116 -10152 -3028 -10088
rect -2964 -10152 -2944 -10088
rect -4116 -10168 -2944 -10152
rect -4116 -10232 -3028 -10168
rect -2964 -10232 -2944 -10168
rect -4116 -10248 -2944 -10232
rect -4116 -10312 -3028 -10248
rect -2964 -10312 -2944 -10248
rect -4116 -10328 -2944 -10312
rect -4116 -10392 -3028 -10328
rect -2964 -10392 -2944 -10328
rect -4116 -10408 -2944 -10392
rect -4116 -10472 -3028 -10408
rect -2964 -10472 -2944 -10408
rect -4116 -10520 -2944 -10472
rect -2704 -9688 -1532 -9640
rect -2704 -9752 -1616 -9688
rect -1552 -9752 -1532 -9688
rect -2704 -9768 -1532 -9752
rect -2704 -9832 -1616 -9768
rect -1552 -9832 -1532 -9768
rect -2704 -9848 -1532 -9832
rect -2704 -9912 -1616 -9848
rect -1552 -9912 -1532 -9848
rect -2704 -9928 -1532 -9912
rect -2704 -9992 -1616 -9928
rect -1552 -9992 -1532 -9928
rect -2704 -10008 -1532 -9992
rect -2704 -10072 -1616 -10008
rect -1552 -10072 -1532 -10008
rect -2704 -10088 -1532 -10072
rect -2704 -10152 -1616 -10088
rect -1552 -10152 -1532 -10088
rect -2704 -10168 -1532 -10152
rect -2704 -10232 -1616 -10168
rect -1552 -10232 -1532 -10168
rect -2704 -10248 -1532 -10232
rect -2704 -10312 -1616 -10248
rect -1552 -10312 -1532 -10248
rect -2704 -10328 -1532 -10312
rect -2704 -10392 -1616 -10328
rect -1552 -10392 -1532 -10328
rect -2704 -10408 -1532 -10392
rect -2704 -10472 -1616 -10408
rect -1552 -10472 -1532 -10408
rect -2704 -10520 -1532 -10472
rect -1292 -9688 -120 -9640
rect -1292 -9752 -204 -9688
rect -140 -9752 -120 -9688
rect -1292 -9768 -120 -9752
rect -1292 -9832 -204 -9768
rect -140 -9832 -120 -9768
rect -1292 -9848 -120 -9832
rect -1292 -9912 -204 -9848
rect -140 -9912 -120 -9848
rect -1292 -9928 -120 -9912
rect -1292 -9992 -204 -9928
rect -140 -9992 -120 -9928
rect -1292 -10008 -120 -9992
rect -1292 -10072 -204 -10008
rect -140 -10072 -120 -10008
rect -1292 -10088 -120 -10072
rect -1292 -10152 -204 -10088
rect -140 -10152 -120 -10088
rect -1292 -10168 -120 -10152
rect -1292 -10232 -204 -10168
rect -140 -10232 -120 -10168
rect -1292 -10248 -120 -10232
rect -1292 -10312 -204 -10248
rect -140 -10312 -120 -10248
rect -1292 -10328 -120 -10312
rect -1292 -10392 -204 -10328
rect -140 -10392 -120 -10328
rect -1292 -10408 -120 -10392
rect -1292 -10472 -204 -10408
rect -140 -10472 -120 -10408
rect -1292 -10520 -120 -10472
rect 120 -9688 1292 -9640
rect 120 -9752 1208 -9688
rect 1272 -9752 1292 -9688
rect 120 -9768 1292 -9752
rect 120 -9832 1208 -9768
rect 1272 -9832 1292 -9768
rect 120 -9848 1292 -9832
rect 120 -9912 1208 -9848
rect 1272 -9912 1292 -9848
rect 120 -9928 1292 -9912
rect 120 -9992 1208 -9928
rect 1272 -9992 1292 -9928
rect 120 -10008 1292 -9992
rect 120 -10072 1208 -10008
rect 1272 -10072 1292 -10008
rect 120 -10088 1292 -10072
rect 120 -10152 1208 -10088
rect 1272 -10152 1292 -10088
rect 120 -10168 1292 -10152
rect 120 -10232 1208 -10168
rect 1272 -10232 1292 -10168
rect 120 -10248 1292 -10232
rect 120 -10312 1208 -10248
rect 1272 -10312 1292 -10248
rect 120 -10328 1292 -10312
rect 120 -10392 1208 -10328
rect 1272 -10392 1292 -10328
rect 120 -10408 1292 -10392
rect 120 -10472 1208 -10408
rect 1272 -10472 1292 -10408
rect 120 -10520 1292 -10472
rect 1532 -9688 2704 -9640
rect 1532 -9752 2620 -9688
rect 2684 -9752 2704 -9688
rect 1532 -9768 2704 -9752
rect 1532 -9832 2620 -9768
rect 2684 -9832 2704 -9768
rect 1532 -9848 2704 -9832
rect 1532 -9912 2620 -9848
rect 2684 -9912 2704 -9848
rect 1532 -9928 2704 -9912
rect 1532 -9992 2620 -9928
rect 2684 -9992 2704 -9928
rect 1532 -10008 2704 -9992
rect 1532 -10072 2620 -10008
rect 2684 -10072 2704 -10008
rect 1532 -10088 2704 -10072
rect 1532 -10152 2620 -10088
rect 2684 -10152 2704 -10088
rect 1532 -10168 2704 -10152
rect 1532 -10232 2620 -10168
rect 2684 -10232 2704 -10168
rect 1532 -10248 2704 -10232
rect 1532 -10312 2620 -10248
rect 2684 -10312 2704 -10248
rect 1532 -10328 2704 -10312
rect 1532 -10392 2620 -10328
rect 2684 -10392 2704 -10328
rect 1532 -10408 2704 -10392
rect 1532 -10472 2620 -10408
rect 2684 -10472 2704 -10408
rect 1532 -10520 2704 -10472
rect 2944 -9688 4116 -9640
rect 2944 -9752 4032 -9688
rect 4096 -9752 4116 -9688
rect 2944 -9768 4116 -9752
rect 2944 -9832 4032 -9768
rect 4096 -9832 4116 -9768
rect 2944 -9848 4116 -9832
rect 2944 -9912 4032 -9848
rect 4096 -9912 4116 -9848
rect 2944 -9928 4116 -9912
rect 2944 -9992 4032 -9928
rect 4096 -9992 4116 -9928
rect 2944 -10008 4116 -9992
rect 2944 -10072 4032 -10008
rect 4096 -10072 4116 -10008
rect 2944 -10088 4116 -10072
rect 2944 -10152 4032 -10088
rect 4096 -10152 4116 -10088
rect 2944 -10168 4116 -10152
rect 2944 -10232 4032 -10168
rect 4096 -10232 4116 -10168
rect 2944 -10248 4116 -10232
rect 2944 -10312 4032 -10248
rect 4096 -10312 4116 -10248
rect 2944 -10328 4116 -10312
rect 2944 -10392 4032 -10328
rect 4096 -10392 4116 -10328
rect 2944 -10408 4116 -10392
rect 2944 -10472 4032 -10408
rect 4096 -10472 4116 -10408
rect 2944 -10520 4116 -10472
rect 4356 -9688 5528 -9640
rect 4356 -9752 5444 -9688
rect 5508 -9752 5528 -9688
rect 4356 -9768 5528 -9752
rect 4356 -9832 5444 -9768
rect 5508 -9832 5528 -9768
rect 4356 -9848 5528 -9832
rect 4356 -9912 5444 -9848
rect 5508 -9912 5528 -9848
rect 4356 -9928 5528 -9912
rect 4356 -9992 5444 -9928
rect 5508 -9992 5528 -9928
rect 4356 -10008 5528 -9992
rect 4356 -10072 5444 -10008
rect 5508 -10072 5528 -10008
rect 4356 -10088 5528 -10072
rect 4356 -10152 5444 -10088
rect 5508 -10152 5528 -10088
rect 4356 -10168 5528 -10152
rect 4356 -10232 5444 -10168
rect 5508 -10232 5528 -10168
rect 4356 -10248 5528 -10232
rect 4356 -10312 5444 -10248
rect 5508 -10312 5528 -10248
rect 4356 -10328 5528 -10312
rect 4356 -10392 5444 -10328
rect 5508 -10392 5528 -10328
rect 4356 -10408 5528 -10392
rect 4356 -10472 5444 -10408
rect 5508 -10472 5528 -10408
rect 4356 -10520 5528 -10472
rect 5768 -9688 6940 -9640
rect 5768 -9752 6856 -9688
rect 6920 -9752 6940 -9688
rect 5768 -9768 6940 -9752
rect 5768 -9832 6856 -9768
rect 6920 -9832 6940 -9768
rect 5768 -9848 6940 -9832
rect 5768 -9912 6856 -9848
rect 6920 -9912 6940 -9848
rect 5768 -9928 6940 -9912
rect 5768 -9992 6856 -9928
rect 6920 -9992 6940 -9928
rect 5768 -10008 6940 -9992
rect 5768 -10072 6856 -10008
rect 6920 -10072 6940 -10008
rect 5768 -10088 6940 -10072
rect 5768 -10152 6856 -10088
rect 6920 -10152 6940 -10088
rect 5768 -10168 6940 -10152
rect 5768 -10232 6856 -10168
rect 6920 -10232 6940 -10168
rect 5768 -10248 6940 -10232
rect 5768 -10312 6856 -10248
rect 6920 -10312 6940 -10248
rect 5768 -10328 6940 -10312
rect 5768 -10392 6856 -10328
rect 6920 -10392 6940 -10328
rect 5768 -10408 6940 -10392
rect 5768 -10472 6856 -10408
rect 6920 -10472 6940 -10408
rect 5768 -10520 6940 -10472
rect 7180 -9688 8352 -9640
rect 7180 -9752 8268 -9688
rect 8332 -9752 8352 -9688
rect 7180 -9768 8352 -9752
rect 7180 -9832 8268 -9768
rect 8332 -9832 8352 -9768
rect 7180 -9848 8352 -9832
rect 7180 -9912 8268 -9848
rect 8332 -9912 8352 -9848
rect 7180 -9928 8352 -9912
rect 7180 -9992 8268 -9928
rect 8332 -9992 8352 -9928
rect 7180 -10008 8352 -9992
rect 7180 -10072 8268 -10008
rect 8332 -10072 8352 -10008
rect 7180 -10088 8352 -10072
rect 7180 -10152 8268 -10088
rect 8332 -10152 8352 -10088
rect 7180 -10168 8352 -10152
rect 7180 -10232 8268 -10168
rect 8332 -10232 8352 -10168
rect 7180 -10248 8352 -10232
rect 7180 -10312 8268 -10248
rect 8332 -10312 8352 -10248
rect 7180 -10328 8352 -10312
rect 7180 -10392 8268 -10328
rect 8332 -10392 8352 -10328
rect 7180 -10408 8352 -10392
rect 7180 -10472 8268 -10408
rect 8332 -10472 8352 -10408
rect 7180 -10520 8352 -10472
rect 8592 -9688 9764 -9640
rect 8592 -9752 9680 -9688
rect 9744 -9752 9764 -9688
rect 8592 -9768 9764 -9752
rect 8592 -9832 9680 -9768
rect 9744 -9832 9764 -9768
rect 8592 -9848 9764 -9832
rect 8592 -9912 9680 -9848
rect 9744 -9912 9764 -9848
rect 8592 -9928 9764 -9912
rect 8592 -9992 9680 -9928
rect 9744 -9992 9764 -9928
rect 8592 -10008 9764 -9992
rect 8592 -10072 9680 -10008
rect 9744 -10072 9764 -10008
rect 8592 -10088 9764 -10072
rect 8592 -10152 9680 -10088
rect 9744 -10152 9764 -10088
rect 8592 -10168 9764 -10152
rect 8592 -10232 9680 -10168
rect 9744 -10232 9764 -10168
rect 8592 -10248 9764 -10232
rect 8592 -10312 9680 -10248
rect 9744 -10312 9764 -10248
rect 8592 -10328 9764 -10312
rect 8592 -10392 9680 -10328
rect 9744 -10392 9764 -10328
rect 8592 -10408 9764 -10392
rect 8592 -10472 9680 -10408
rect 9744 -10472 9764 -10408
rect 8592 -10520 9764 -10472
rect 10004 -9688 11176 -9640
rect 10004 -9752 11092 -9688
rect 11156 -9752 11176 -9688
rect 10004 -9768 11176 -9752
rect 10004 -9832 11092 -9768
rect 11156 -9832 11176 -9768
rect 10004 -9848 11176 -9832
rect 10004 -9912 11092 -9848
rect 11156 -9912 11176 -9848
rect 10004 -9928 11176 -9912
rect 10004 -9992 11092 -9928
rect 11156 -9992 11176 -9928
rect 10004 -10008 11176 -9992
rect 10004 -10072 11092 -10008
rect 11156 -10072 11176 -10008
rect 10004 -10088 11176 -10072
rect 10004 -10152 11092 -10088
rect 11156 -10152 11176 -10088
rect 10004 -10168 11176 -10152
rect 10004 -10232 11092 -10168
rect 11156 -10232 11176 -10168
rect 10004 -10248 11176 -10232
rect 10004 -10312 11092 -10248
rect 11156 -10312 11176 -10248
rect 10004 -10328 11176 -10312
rect 10004 -10392 11092 -10328
rect 11156 -10392 11176 -10328
rect 10004 -10408 11176 -10392
rect 10004 -10472 11092 -10408
rect 11156 -10472 11176 -10408
rect 10004 -10520 11176 -10472
rect 11416 -9688 12588 -9640
rect 11416 -9752 12504 -9688
rect 12568 -9752 12588 -9688
rect 11416 -9768 12588 -9752
rect 11416 -9832 12504 -9768
rect 12568 -9832 12588 -9768
rect 11416 -9848 12588 -9832
rect 11416 -9912 12504 -9848
rect 12568 -9912 12588 -9848
rect 11416 -9928 12588 -9912
rect 11416 -9992 12504 -9928
rect 12568 -9992 12588 -9928
rect 11416 -10008 12588 -9992
rect 11416 -10072 12504 -10008
rect 12568 -10072 12588 -10008
rect 11416 -10088 12588 -10072
rect 11416 -10152 12504 -10088
rect 12568 -10152 12588 -10088
rect 11416 -10168 12588 -10152
rect 11416 -10232 12504 -10168
rect 12568 -10232 12588 -10168
rect 11416 -10248 12588 -10232
rect 11416 -10312 12504 -10248
rect 12568 -10312 12588 -10248
rect 11416 -10328 12588 -10312
rect 11416 -10392 12504 -10328
rect 12568 -10392 12588 -10328
rect 11416 -10408 12588 -10392
rect 11416 -10472 12504 -10408
rect 12568 -10472 12588 -10408
rect 11416 -10520 12588 -10472
rect 12828 -9688 14000 -9640
rect 12828 -9752 13916 -9688
rect 13980 -9752 14000 -9688
rect 12828 -9768 14000 -9752
rect 12828 -9832 13916 -9768
rect 13980 -9832 14000 -9768
rect 12828 -9848 14000 -9832
rect 12828 -9912 13916 -9848
rect 13980 -9912 14000 -9848
rect 12828 -9928 14000 -9912
rect 12828 -9992 13916 -9928
rect 13980 -9992 14000 -9928
rect 12828 -10008 14000 -9992
rect 12828 -10072 13916 -10008
rect 13980 -10072 14000 -10008
rect 12828 -10088 14000 -10072
rect 12828 -10152 13916 -10088
rect 13980 -10152 14000 -10088
rect 12828 -10168 14000 -10152
rect 12828 -10232 13916 -10168
rect 13980 -10232 14000 -10168
rect 12828 -10248 14000 -10232
rect 12828 -10312 13916 -10248
rect 13980 -10312 14000 -10248
rect 12828 -10328 14000 -10312
rect 12828 -10392 13916 -10328
rect 13980 -10392 14000 -10328
rect 12828 -10408 14000 -10392
rect 12828 -10472 13916 -10408
rect 13980 -10472 14000 -10408
rect 12828 -10520 14000 -10472
rect 14240 -9688 15412 -9640
rect 14240 -9752 15328 -9688
rect 15392 -9752 15412 -9688
rect 14240 -9768 15412 -9752
rect 14240 -9832 15328 -9768
rect 15392 -9832 15412 -9768
rect 14240 -9848 15412 -9832
rect 14240 -9912 15328 -9848
rect 15392 -9912 15412 -9848
rect 14240 -9928 15412 -9912
rect 14240 -9992 15328 -9928
rect 15392 -9992 15412 -9928
rect 14240 -10008 15412 -9992
rect 14240 -10072 15328 -10008
rect 15392 -10072 15412 -10008
rect 14240 -10088 15412 -10072
rect 14240 -10152 15328 -10088
rect 15392 -10152 15412 -10088
rect 14240 -10168 15412 -10152
rect 14240 -10232 15328 -10168
rect 15392 -10232 15412 -10168
rect 14240 -10248 15412 -10232
rect 14240 -10312 15328 -10248
rect 15392 -10312 15412 -10248
rect 14240 -10328 15412 -10312
rect 14240 -10392 15328 -10328
rect 15392 -10392 15412 -10328
rect 14240 -10408 15412 -10392
rect 14240 -10472 15328 -10408
rect 15392 -10472 15412 -10408
rect 14240 -10520 15412 -10472
rect 15652 -9688 16824 -9640
rect 15652 -9752 16740 -9688
rect 16804 -9752 16824 -9688
rect 15652 -9768 16824 -9752
rect 15652 -9832 16740 -9768
rect 16804 -9832 16824 -9768
rect 15652 -9848 16824 -9832
rect 15652 -9912 16740 -9848
rect 16804 -9912 16824 -9848
rect 15652 -9928 16824 -9912
rect 15652 -9992 16740 -9928
rect 16804 -9992 16824 -9928
rect 15652 -10008 16824 -9992
rect 15652 -10072 16740 -10008
rect 16804 -10072 16824 -10008
rect 15652 -10088 16824 -10072
rect 15652 -10152 16740 -10088
rect 16804 -10152 16824 -10088
rect 15652 -10168 16824 -10152
rect 15652 -10232 16740 -10168
rect 16804 -10232 16824 -10168
rect 15652 -10248 16824 -10232
rect 15652 -10312 16740 -10248
rect 16804 -10312 16824 -10248
rect 15652 -10328 16824 -10312
rect 15652 -10392 16740 -10328
rect 16804 -10392 16824 -10328
rect 15652 -10408 16824 -10392
rect 15652 -10472 16740 -10408
rect 16804 -10472 16824 -10408
rect 15652 -10520 16824 -10472
rect 17064 -9688 18236 -9640
rect 17064 -9752 18152 -9688
rect 18216 -9752 18236 -9688
rect 17064 -9768 18236 -9752
rect 17064 -9832 18152 -9768
rect 18216 -9832 18236 -9768
rect 17064 -9848 18236 -9832
rect 17064 -9912 18152 -9848
rect 18216 -9912 18236 -9848
rect 17064 -9928 18236 -9912
rect 17064 -9992 18152 -9928
rect 18216 -9992 18236 -9928
rect 17064 -10008 18236 -9992
rect 17064 -10072 18152 -10008
rect 18216 -10072 18236 -10008
rect 17064 -10088 18236 -10072
rect 17064 -10152 18152 -10088
rect 18216 -10152 18236 -10088
rect 17064 -10168 18236 -10152
rect 17064 -10232 18152 -10168
rect 18216 -10232 18236 -10168
rect 17064 -10248 18236 -10232
rect 17064 -10312 18152 -10248
rect 18216 -10312 18236 -10248
rect 17064 -10328 18236 -10312
rect 17064 -10392 18152 -10328
rect 18216 -10392 18236 -10328
rect 17064 -10408 18236 -10392
rect 17064 -10472 18152 -10408
rect 18216 -10472 18236 -10408
rect 17064 -10520 18236 -10472
rect 18476 -9688 19648 -9640
rect 18476 -9752 19564 -9688
rect 19628 -9752 19648 -9688
rect 18476 -9768 19648 -9752
rect 18476 -9832 19564 -9768
rect 19628 -9832 19648 -9768
rect 18476 -9848 19648 -9832
rect 18476 -9912 19564 -9848
rect 19628 -9912 19648 -9848
rect 18476 -9928 19648 -9912
rect 18476 -9992 19564 -9928
rect 19628 -9992 19648 -9928
rect 18476 -10008 19648 -9992
rect 18476 -10072 19564 -10008
rect 19628 -10072 19648 -10008
rect 18476 -10088 19648 -10072
rect 18476 -10152 19564 -10088
rect 19628 -10152 19648 -10088
rect 18476 -10168 19648 -10152
rect 18476 -10232 19564 -10168
rect 19628 -10232 19648 -10168
rect 18476 -10248 19648 -10232
rect 18476 -10312 19564 -10248
rect 19628 -10312 19648 -10248
rect 18476 -10328 19648 -10312
rect 18476 -10392 19564 -10328
rect 19628 -10392 19648 -10328
rect 18476 -10408 19648 -10392
rect 18476 -10472 19564 -10408
rect 19628 -10472 19648 -10408
rect 18476 -10520 19648 -10472
rect 19888 -9688 21060 -9640
rect 19888 -9752 20976 -9688
rect 21040 -9752 21060 -9688
rect 19888 -9768 21060 -9752
rect 19888 -9832 20976 -9768
rect 21040 -9832 21060 -9768
rect 19888 -9848 21060 -9832
rect 19888 -9912 20976 -9848
rect 21040 -9912 21060 -9848
rect 19888 -9928 21060 -9912
rect 19888 -9992 20976 -9928
rect 21040 -9992 21060 -9928
rect 19888 -10008 21060 -9992
rect 19888 -10072 20976 -10008
rect 21040 -10072 21060 -10008
rect 19888 -10088 21060 -10072
rect 19888 -10152 20976 -10088
rect 21040 -10152 21060 -10088
rect 19888 -10168 21060 -10152
rect 19888 -10232 20976 -10168
rect 21040 -10232 21060 -10168
rect 19888 -10248 21060 -10232
rect 19888 -10312 20976 -10248
rect 21040 -10312 21060 -10248
rect 19888 -10328 21060 -10312
rect 19888 -10392 20976 -10328
rect 21040 -10392 21060 -10328
rect 19888 -10408 21060 -10392
rect 19888 -10472 20976 -10408
rect 21040 -10472 21060 -10408
rect 19888 -10520 21060 -10472
rect 21300 -9688 22472 -9640
rect 21300 -9752 22388 -9688
rect 22452 -9752 22472 -9688
rect 21300 -9768 22472 -9752
rect 21300 -9832 22388 -9768
rect 22452 -9832 22472 -9768
rect 21300 -9848 22472 -9832
rect 21300 -9912 22388 -9848
rect 22452 -9912 22472 -9848
rect 21300 -9928 22472 -9912
rect 21300 -9992 22388 -9928
rect 22452 -9992 22472 -9928
rect 21300 -10008 22472 -9992
rect 21300 -10072 22388 -10008
rect 22452 -10072 22472 -10008
rect 21300 -10088 22472 -10072
rect 21300 -10152 22388 -10088
rect 22452 -10152 22472 -10088
rect 21300 -10168 22472 -10152
rect 21300 -10232 22388 -10168
rect 22452 -10232 22472 -10168
rect 21300 -10248 22472 -10232
rect 21300 -10312 22388 -10248
rect 22452 -10312 22472 -10248
rect 21300 -10328 22472 -10312
rect 21300 -10392 22388 -10328
rect 22452 -10392 22472 -10328
rect 21300 -10408 22472 -10392
rect 21300 -10472 22388 -10408
rect 22452 -10472 22472 -10408
rect 21300 -10520 22472 -10472
rect 22712 -9688 23884 -9640
rect 22712 -9752 23800 -9688
rect 23864 -9752 23884 -9688
rect 22712 -9768 23884 -9752
rect 22712 -9832 23800 -9768
rect 23864 -9832 23884 -9768
rect 22712 -9848 23884 -9832
rect 22712 -9912 23800 -9848
rect 23864 -9912 23884 -9848
rect 22712 -9928 23884 -9912
rect 22712 -9992 23800 -9928
rect 23864 -9992 23884 -9928
rect 22712 -10008 23884 -9992
rect 22712 -10072 23800 -10008
rect 23864 -10072 23884 -10008
rect 22712 -10088 23884 -10072
rect 22712 -10152 23800 -10088
rect 23864 -10152 23884 -10088
rect 22712 -10168 23884 -10152
rect 22712 -10232 23800 -10168
rect 23864 -10232 23884 -10168
rect 22712 -10248 23884 -10232
rect 22712 -10312 23800 -10248
rect 23864 -10312 23884 -10248
rect 22712 -10328 23884 -10312
rect 22712 -10392 23800 -10328
rect 23864 -10392 23884 -10328
rect 22712 -10408 23884 -10392
rect 22712 -10472 23800 -10408
rect 23864 -10472 23884 -10408
rect 22712 -10520 23884 -10472
rect -23884 -10808 -22712 -10760
rect -23884 -10872 -22796 -10808
rect -22732 -10872 -22712 -10808
rect -23884 -10888 -22712 -10872
rect -23884 -10952 -22796 -10888
rect -22732 -10952 -22712 -10888
rect -23884 -10968 -22712 -10952
rect -23884 -11032 -22796 -10968
rect -22732 -11032 -22712 -10968
rect -23884 -11048 -22712 -11032
rect -23884 -11112 -22796 -11048
rect -22732 -11112 -22712 -11048
rect -23884 -11128 -22712 -11112
rect -23884 -11192 -22796 -11128
rect -22732 -11192 -22712 -11128
rect -23884 -11208 -22712 -11192
rect -23884 -11272 -22796 -11208
rect -22732 -11272 -22712 -11208
rect -23884 -11288 -22712 -11272
rect -23884 -11352 -22796 -11288
rect -22732 -11352 -22712 -11288
rect -23884 -11368 -22712 -11352
rect -23884 -11432 -22796 -11368
rect -22732 -11432 -22712 -11368
rect -23884 -11448 -22712 -11432
rect -23884 -11512 -22796 -11448
rect -22732 -11512 -22712 -11448
rect -23884 -11528 -22712 -11512
rect -23884 -11592 -22796 -11528
rect -22732 -11592 -22712 -11528
rect -23884 -11640 -22712 -11592
rect -22472 -10808 -21300 -10760
rect -22472 -10872 -21384 -10808
rect -21320 -10872 -21300 -10808
rect -22472 -10888 -21300 -10872
rect -22472 -10952 -21384 -10888
rect -21320 -10952 -21300 -10888
rect -22472 -10968 -21300 -10952
rect -22472 -11032 -21384 -10968
rect -21320 -11032 -21300 -10968
rect -22472 -11048 -21300 -11032
rect -22472 -11112 -21384 -11048
rect -21320 -11112 -21300 -11048
rect -22472 -11128 -21300 -11112
rect -22472 -11192 -21384 -11128
rect -21320 -11192 -21300 -11128
rect -22472 -11208 -21300 -11192
rect -22472 -11272 -21384 -11208
rect -21320 -11272 -21300 -11208
rect -22472 -11288 -21300 -11272
rect -22472 -11352 -21384 -11288
rect -21320 -11352 -21300 -11288
rect -22472 -11368 -21300 -11352
rect -22472 -11432 -21384 -11368
rect -21320 -11432 -21300 -11368
rect -22472 -11448 -21300 -11432
rect -22472 -11512 -21384 -11448
rect -21320 -11512 -21300 -11448
rect -22472 -11528 -21300 -11512
rect -22472 -11592 -21384 -11528
rect -21320 -11592 -21300 -11528
rect -22472 -11640 -21300 -11592
rect -21060 -10808 -19888 -10760
rect -21060 -10872 -19972 -10808
rect -19908 -10872 -19888 -10808
rect -21060 -10888 -19888 -10872
rect -21060 -10952 -19972 -10888
rect -19908 -10952 -19888 -10888
rect -21060 -10968 -19888 -10952
rect -21060 -11032 -19972 -10968
rect -19908 -11032 -19888 -10968
rect -21060 -11048 -19888 -11032
rect -21060 -11112 -19972 -11048
rect -19908 -11112 -19888 -11048
rect -21060 -11128 -19888 -11112
rect -21060 -11192 -19972 -11128
rect -19908 -11192 -19888 -11128
rect -21060 -11208 -19888 -11192
rect -21060 -11272 -19972 -11208
rect -19908 -11272 -19888 -11208
rect -21060 -11288 -19888 -11272
rect -21060 -11352 -19972 -11288
rect -19908 -11352 -19888 -11288
rect -21060 -11368 -19888 -11352
rect -21060 -11432 -19972 -11368
rect -19908 -11432 -19888 -11368
rect -21060 -11448 -19888 -11432
rect -21060 -11512 -19972 -11448
rect -19908 -11512 -19888 -11448
rect -21060 -11528 -19888 -11512
rect -21060 -11592 -19972 -11528
rect -19908 -11592 -19888 -11528
rect -21060 -11640 -19888 -11592
rect -19648 -10808 -18476 -10760
rect -19648 -10872 -18560 -10808
rect -18496 -10872 -18476 -10808
rect -19648 -10888 -18476 -10872
rect -19648 -10952 -18560 -10888
rect -18496 -10952 -18476 -10888
rect -19648 -10968 -18476 -10952
rect -19648 -11032 -18560 -10968
rect -18496 -11032 -18476 -10968
rect -19648 -11048 -18476 -11032
rect -19648 -11112 -18560 -11048
rect -18496 -11112 -18476 -11048
rect -19648 -11128 -18476 -11112
rect -19648 -11192 -18560 -11128
rect -18496 -11192 -18476 -11128
rect -19648 -11208 -18476 -11192
rect -19648 -11272 -18560 -11208
rect -18496 -11272 -18476 -11208
rect -19648 -11288 -18476 -11272
rect -19648 -11352 -18560 -11288
rect -18496 -11352 -18476 -11288
rect -19648 -11368 -18476 -11352
rect -19648 -11432 -18560 -11368
rect -18496 -11432 -18476 -11368
rect -19648 -11448 -18476 -11432
rect -19648 -11512 -18560 -11448
rect -18496 -11512 -18476 -11448
rect -19648 -11528 -18476 -11512
rect -19648 -11592 -18560 -11528
rect -18496 -11592 -18476 -11528
rect -19648 -11640 -18476 -11592
rect -18236 -10808 -17064 -10760
rect -18236 -10872 -17148 -10808
rect -17084 -10872 -17064 -10808
rect -18236 -10888 -17064 -10872
rect -18236 -10952 -17148 -10888
rect -17084 -10952 -17064 -10888
rect -18236 -10968 -17064 -10952
rect -18236 -11032 -17148 -10968
rect -17084 -11032 -17064 -10968
rect -18236 -11048 -17064 -11032
rect -18236 -11112 -17148 -11048
rect -17084 -11112 -17064 -11048
rect -18236 -11128 -17064 -11112
rect -18236 -11192 -17148 -11128
rect -17084 -11192 -17064 -11128
rect -18236 -11208 -17064 -11192
rect -18236 -11272 -17148 -11208
rect -17084 -11272 -17064 -11208
rect -18236 -11288 -17064 -11272
rect -18236 -11352 -17148 -11288
rect -17084 -11352 -17064 -11288
rect -18236 -11368 -17064 -11352
rect -18236 -11432 -17148 -11368
rect -17084 -11432 -17064 -11368
rect -18236 -11448 -17064 -11432
rect -18236 -11512 -17148 -11448
rect -17084 -11512 -17064 -11448
rect -18236 -11528 -17064 -11512
rect -18236 -11592 -17148 -11528
rect -17084 -11592 -17064 -11528
rect -18236 -11640 -17064 -11592
rect -16824 -10808 -15652 -10760
rect -16824 -10872 -15736 -10808
rect -15672 -10872 -15652 -10808
rect -16824 -10888 -15652 -10872
rect -16824 -10952 -15736 -10888
rect -15672 -10952 -15652 -10888
rect -16824 -10968 -15652 -10952
rect -16824 -11032 -15736 -10968
rect -15672 -11032 -15652 -10968
rect -16824 -11048 -15652 -11032
rect -16824 -11112 -15736 -11048
rect -15672 -11112 -15652 -11048
rect -16824 -11128 -15652 -11112
rect -16824 -11192 -15736 -11128
rect -15672 -11192 -15652 -11128
rect -16824 -11208 -15652 -11192
rect -16824 -11272 -15736 -11208
rect -15672 -11272 -15652 -11208
rect -16824 -11288 -15652 -11272
rect -16824 -11352 -15736 -11288
rect -15672 -11352 -15652 -11288
rect -16824 -11368 -15652 -11352
rect -16824 -11432 -15736 -11368
rect -15672 -11432 -15652 -11368
rect -16824 -11448 -15652 -11432
rect -16824 -11512 -15736 -11448
rect -15672 -11512 -15652 -11448
rect -16824 -11528 -15652 -11512
rect -16824 -11592 -15736 -11528
rect -15672 -11592 -15652 -11528
rect -16824 -11640 -15652 -11592
rect -15412 -10808 -14240 -10760
rect -15412 -10872 -14324 -10808
rect -14260 -10872 -14240 -10808
rect -15412 -10888 -14240 -10872
rect -15412 -10952 -14324 -10888
rect -14260 -10952 -14240 -10888
rect -15412 -10968 -14240 -10952
rect -15412 -11032 -14324 -10968
rect -14260 -11032 -14240 -10968
rect -15412 -11048 -14240 -11032
rect -15412 -11112 -14324 -11048
rect -14260 -11112 -14240 -11048
rect -15412 -11128 -14240 -11112
rect -15412 -11192 -14324 -11128
rect -14260 -11192 -14240 -11128
rect -15412 -11208 -14240 -11192
rect -15412 -11272 -14324 -11208
rect -14260 -11272 -14240 -11208
rect -15412 -11288 -14240 -11272
rect -15412 -11352 -14324 -11288
rect -14260 -11352 -14240 -11288
rect -15412 -11368 -14240 -11352
rect -15412 -11432 -14324 -11368
rect -14260 -11432 -14240 -11368
rect -15412 -11448 -14240 -11432
rect -15412 -11512 -14324 -11448
rect -14260 -11512 -14240 -11448
rect -15412 -11528 -14240 -11512
rect -15412 -11592 -14324 -11528
rect -14260 -11592 -14240 -11528
rect -15412 -11640 -14240 -11592
rect -14000 -10808 -12828 -10760
rect -14000 -10872 -12912 -10808
rect -12848 -10872 -12828 -10808
rect -14000 -10888 -12828 -10872
rect -14000 -10952 -12912 -10888
rect -12848 -10952 -12828 -10888
rect -14000 -10968 -12828 -10952
rect -14000 -11032 -12912 -10968
rect -12848 -11032 -12828 -10968
rect -14000 -11048 -12828 -11032
rect -14000 -11112 -12912 -11048
rect -12848 -11112 -12828 -11048
rect -14000 -11128 -12828 -11112
rect -14000 -11192 -12912 -11128
rect -12848 -11192 -12828 -11128
rect -14000 -11208 -12828 -11192
rect -14000 -11272 -12912 -11208
rect -12848 -11272 -12828 -11208
rect -14000 -11288 -12828 -11272
rect -14000 -11352 -12912 -11288
rect -12848 -11352 -12828 -11288
rect -14000 -11368 -12828 -11352
rect -14000 -11432 -12912 -11368
rect -12848 -11432 -12828 -11368
rect -14000 -11448 -12828 -11432
rect -14000 -11512 -12912 -11448
rect -12848 -11512 -12828 -11448
rect -14000 -11528 -12828 -11512
rect -14000 -11592 -12912 -11528
rect -12848 -11592 -12828 -11528
rect -14000 -11640 -12828 -11592
rect -12588 -10808 -11416 -10760
rect -12588 -10872 -11500 -10808
rect -11436 -10872 -11416 -10808
rect -12588 -10888 -11416 -10872
rect -12588 -10952 -11500 -10888
rect -11436 -10952 -11416 -10888
rect -12588 -10968 -11416 -10952
rect -12588 -11032 -11500 -10968
rect -11436 -11032 -11416 -10968
rect -12588 -11048 -11416 -11032
rect -12588 -11112 -11500 -11048
rect -11436 -11112 -11416 -11048
rect -12588 -11128 -11416 -11112
rect -12588 -11192 -11500 -11128
rect -11436 -11192 -11416 -11128
rect -12588 -11208 -11416 -11192
rect -12588 -11272 -11500 -11208
rect -11436 -11272 -11416 -11208
rect -12588 -11288 -11416 -11272
rect -12588 -11352 -11500 -11288
rect -11436 -11352 -11416 -11288
rect -12588 -11368 -11416 -11352
rect -12588 -11432 -11500 -11368
rect -11436 -11432 -11416 -11368
rect -12588 -11448 -11416 -11432
rect -12588 -11512 -11500 -11448
rect -11436 -11512 -11416 -11448
rect -12588 -11528 -11416 -11512
rect -12588 -11592 -11500 -11528
rect -11436 -11592 -11416 -11528
rect -12588 -11640 -11416 -11592
rect -11176 -10808 -10004 -10760
rect -11176 -10872 -10088 -10808
rect -10024 -10872 -10004 -10808
rect -11176 -10888 -10004 -10872
rect -11176 -10952 -10088 -10888
rect -10024 -10952 -10004 -10888
rect -11176 -10968 -10004 -10952
rect -11176 -11032 -10088 -10968
rect -10024 -11032 -10004 -10968
rect -11176 -11048 -10004 -11032
rect -11176 -11112 -10088 -11048
rect -10024 -11112 -10004 -11048
rect -11176 -11128 -10004 -11112
rect -11176 -11192 -10088 -11128
rect -10024 -11192 -10004 -11128
rect -11176 -11208 -10004 -11192
rect -11176 -11272 -10088 -11208
rect -10024 -11272 -10004 -11208
rect -11176 -11288 -10004 -11272
rect -11176 -11352 -10088 -11288
rect -10024 -11352 -10004 -11288
rect -11176 -11368 -10004 -11352
rect -11176 -11432 -10088 -11368
rect -10024 -11432 -10004 -11368
rect -11176 -11448 -10004 -11432
rect -11176 -11512 -10088 -11448
rect -10024 -11512 -10004 -11448
rect -11176 -11528 -10004 -11512
rect -11176 -11592 -10088 -11528
rect -10024 -11592 -10004 -11528
rect -11176 -11640 -10004 -11592
rect -9764 -10808 -8592 -10760
rect -9764 -10872 -8676 -10808
rect -8612 -10872 -8592 -10808
rect -9764 -10888 -8592 -10872
rect -9764 -10952 -8676 -10888
rect -8612 -10952 -8592 -10888
rect -9764 -10968 -8592 -10952
rect -9764 -11032 -8676 -10968
rect -8612 -11032 -8592 -10968
rect -9764 -11048 -8592 -11032
rect -9764 -11112 -8676 -11048
rect -8612 -11112 -8592 -11048
rect -9764 -11128 -8592 -11112
rect -9764 -11192 -8676 -11128
rect -8612 -11192 -8592 -11128
rect -9764 -11208 -8592 -11192
rect -9764 -11272 -8676 -11208
rect -8612 -11272 -8592 -11208
rect -9764 -11288 -8592 -11272
rect -9764 -11352 -8676 -11288
rect -8612 -11352 -8592 -11288
rect -9764 -11368 -8592 -11352
rect -9764 -11432 -8676 -11368
rect -8612 -11432 -8592 -11368
rect -9764 -11448 -8592 -11432
rect -9764 -11512 -8676 -11448
rect -8612 -11512 -8592 -11448
rect -9764 -11528 -8592 -11512
rect -9764 -11592 -8676 -11528
rect -8612 -11592 -8592 -11528
rect -9764 -11640 -8592 -11592
rect -8352 -10808 -7180 -10760
rect -8352 -10872 -7264 -10808
rect -7200 -10872 -7180 -10808
rect -8352 -10888 -7180 -10872
rect -8352 -10952 -7264 -10888
rect -7200 -10952 -7180 -10888
rect -8352 -10968 -7180 -10952
rect -8352 -11032 -7264 -10968
rect -7200 -11032 -7180 -10968
rect -8352 -11048 -7180 -11032
rect -8352 -11112 -7264 -11048
rect -7200 -11112 -7180 -11048
rect -8352 -11128 -7180 -11112
rect -8352 -11192 -7264 -11128
rect -7200 -11192 -7180 -11128
rect -8352 -11208 -7180 -11192
rect -8352 -11272 -7264 -11208
rect -7200 -11272 -7180 -11208
rect -8352 -11288 -7180 -11272
rect -8352 -11352 -7264 -11288
rect -7200 -11352 -7180 -11288
rect -8352 -11368 -7180 -11352
rect -8352 -11432 -7264 -11368
rect -7200 -11432 -7180 -11368
rect -8352 -11448 -7180 -11432
rect -8352 -11512 -7264 -11448
rect -7200 -11512 -7180 -11448
rect -8352 -11528 -7180 -11512
rect -8352 -11592 -7264 -11528
rect -7200 -11592 -7180 -11528
rect -8352 -11640 -7180 -11592
rect -6940 -10808 -5768 -10760
rect -6940 -10872 -5852 -10808
rect -5788 -10872 -5768 -10808
rect -6940 -10888 -5768 -10872
rect -6940 -10952 -5852 -10888
rect -5788 -10952 -5768 -10888
rect -6940 -10968 -5768 -10952
rect -6940 -11032 -5852 -10968
rect -5788 -11032 -5768 -10968
rect -6940 -11048 -5768 -11032
rect -6940 -11112 -5852 -11048
rect -5788 -11112 -5768 -11048
rect -6940 -11128 -5768 -11112
rect -6940 -11192 -5852 -11128
rect -5788 -11192 -5768 -11128
rect -6940 -11208 -5768 -11192
rect -6940 -11272 -5852 -11208
rect -5788 -11272 -5768 -11208
rect -6940 -11288 -5768 -11272
rect -6940 -11352 -5852 -11288
rect -5788 -11352 -5768 -11288
rect -6940 -11368 -5768 -11352
rect -6940 -11432 -5852 -11368
rect -5788 -11432 -5768 -11368
rect -6940 -11448 -5768 -11432
rect -6940 -11512 -5852 -11448
rect -5788 -11512 -5768 -11448
rect -6940 -11528 -5768 -11512
rect -6940 -11592 -5852 -11528
rect -5788 -11592 -5768 -11528
rect -6940 -11640 -5768 -11592
rect -5528 -10808 -4356 -10760
rect -5528 -10872 -4440 -10808
rect -4376 -10872 -4356 -10808
rect -5528 -10888 -4356 -10872
rect -5528 -10952 -4440 -10888
rect -4376 -10952 -4356 -10888
rect -5528 -10968 -4356 -10952
rect -5528 -11032 -4440 -10968
rect -4376 -11032 -4356 -10968
rect -5528 -11048 -4356 -11032
rect -5528 -11112 -4440 -11048
rect -4376 -11112 -4356 -11048
rect -5528 -11128 -4356 -11112
rect -5528 -11192 -4440 -11128
rect -4376 -11192 -4356 -11128
rect -5528 -11208 -4356 -11192
rect -5528 -11272 -4440 -11208
rect -4376 -11272 -4356 -11208
rect -5528 -11288 -4356 -11272
rect -5528 -11352 -4440 -11288
rect -4376 -11352 -4356 -11288
rect -5528 -11368 -4356 -11352
rect -5528 -11432 -4440 -11368
rect -4376 -11432 -4356 -11368
rect -5528 -11448 -4356 -11432
rect -5528 -11512 -4440 -11448
rect -4376 -11512 -4356 -11448
rect -5528 -11528 -4356 -11512
rect -5528 -11592 -4440 -11528
rect -4376 -11592 -4356 -11528
rect -5528 -11640 -4356 -11592
rect -4116 -10808 -2944 -10760
rect -4116 -10872 -3028 -10808
rect -2964 -10872 -2944 -10808
rect -4116 -10888 -2944 -10872
rect -4116 -10952 -3028 -10888
rect -2964 -10952 -2944 -10888
rect -4116 -10968 -2944 -10952
rect -4116 -11032 -3028 -10968
rect -2964 -11032 -2944 -10968
rect -4116 -11048 -2944 -11032
rect -4116 -11112 -3028 -11048
rect -2964 -11112 -2944 -11048
rect -4116 -11128 -2944 -11112
rect -4116 -11192 -3028 -11128
rect -2964 -11192 -2944 -11128
rect -4116 -11208 -2944 -11192
rect -4116 -11272 -3028 -11208
rect -2964 -11272 -2944 -11208
rect -4116 -11288 -2944 -11272
rect -4116 -11352 -3028 -11288
rect -2964 -11352 -2944 -11288
rect -4116 -11368 -2944 -11352
rect -4116 -11432 -3028 -11368
rect -2964 -11432 -2944 -11368
rect -4116 -11448 -2944 -11432
rect -4116 -11512 -3028 -11448
rect -2964 -11512 -2944 -11448
rect -4116 -11528 -2944 -11512
rect -4116 -11592 -3028 -11528
rect -2964 -11592 -2944 -11528
rect -4116 -11640 -2944 -11592
rect -2704 -10808 -1532 -10760
rect -2704 -10872 -1616 -10808
rect -1552 -10872 -1532 -10808
rect -2704 -10888 -1532 -10872
rect -2704 -10952 -1616 -10888
rect -1552 -10952 -1532 -10888
rect -2704 -10968 -1532 -10952
rect -2704 -11032 -1616 -10968
rect -1552 -11032 -1532 -10968
rect -2704 -11048 -1532 -11032
rect -2704 -11112 -1616 -11048
rect -1552 -11112 -1532 -11048
rect -2704 -11128 -1532 -11112
rect -2704 -11192 -1616 -11128
rect -1552 -11192 -1532 -11128
rect -2704 -11208 -1532 -11192
rect -2704 -11272 -1616 -11208
rect -1552 -11272 -1532 -11208
rect -2704 -11288 -1532 -11272
rect -2704 -11352 -1616 -11288
rect -1552 -11352 -1532 -11288
rect -2704 -11368 -1532 -11352
rect -2704 -11432 -1616 -11368
rect -1552 -11432 -1532 -11368
rect -2704 -11448 -1532 -11432
rect -2704 -11512 -1616 -11448
rect -1552 -11512 -1532 -11448
rect -2704 -11528 -1532 -11512
rect -2704 -11592 -1616 -11528
rect -1552 -11592 -1532 -11528
rect -2704 -11640 -1532 -11592
rect -1292 -10808 -120 -10760
rect -1292 -10872 -204 -10808
rect -140 -10872 -120 -10808
rect -1292 -10888 -120 -10872
rect -1292 -10952 -204 -10888
rect -140 -10952 -120 -10888
rect -1292 -10968 -120 -10952
rect -1292 -11032 -204 -10968
rect -140 -11032 -120 -10968
rect -1292 -11048 -120 -11032
rect -1292 -11112 -204 -11048
rect -140 -11112 -120 -11048
rect -1292 -11128 -120 -11112
rect -1292 -11192 -204 -11128
rect -140 -11192 -120 -11128
rect -1292 -11208 -120 -11192
rect -1292 -11272 -204 -11208
rect -140 -11272 -120 -11208
rect -1292 -11288 -120 -11272
rect -1292 -11352 -204 -11288
rect -140 -11352 -120 -11288
rect -1292 -11368 -120 -11352
rect -1292 -11432 -204 -11368
rect -140 -11432 -120 -11368
rect -1292 -11448 -120 -11432
rect -1292 -11512 -204 -11448
rect -140 -11512 -120 -11448
rect -1292 -11528 -120 -11512
rect -1292 -11592 -204 -11528
rect -140 -11592 -120 -11528
rect -1292 -11640 -120 -11592
rect 120 -10808 1292 -10760
rect 120 -10872 1208 -10808
rect 1272 -10872 1292 -10808
rect 120 -10888 1292 -10872
rect 120 -10952 1208 -10888
rect 1272 -10952 1292 -10888
rect 120 -10968 1292 -10952
rect 120 -11032 1208 -10968
rect 1272 -11032 1292 -10968
rect 120 -11048 1292 -11032
rect 120 -11112 1208 -11048
rect 1272 -11112 1292 -11048
rect 120 -11128 1292 -11112
rect 120 -11192 1208 -11128
rect 1272 -11192 1292 -11128
rect 120 -11208 1292 -11192
rect 120 -11272 1208 -11208
rect 1272 -11272 1292 -11208
rect 120 -11288 1292 -11272
rect 120 -11352 1208 -11288
rect 1272 -11352 1292 -11288
rect 120 -11368 1292 -11352
rect 120 -11432 1208 -11368
rect 1272 -11432 1292 -11368
rect 120 -11448 1292 -11432
rect 120 -11512 1208 -11448
rect 1272 -11512 1292 -11448
rect 120 -11528 1292 -11512
rect 120 -11592 1208 -11528
rect 1272 -11592 1292 -11528
rect 120 -11640 1292 -11592
rect 1532 -10808 2704 -10760
rect 1532 -10872 2620 -10808
rect 2684 -10872 2704 -10808
rect 1532 -10888 2704 -10872
rect 1532 -10952 2620 -10888
rect 2684 -10952 2704 -10888
rect 1532 -10968 2704 -10952
rect 1532 -11032 2620 -10968
rect 2684 -11032 2704 -10968
rect 1532 -11048 2704 -11032
rect 1532 -11112 2620 -11048
rect 2684 -11112 2704 -11048
rect 1532 -11128 2704 -11112
rect 1532 -11192 2620 -11128
rect 2684 -11192 2704 -11128
rect 1532 -11208 2704 -11192
rect 1532 -11272 2620 -11208
rect 2684 -11272 2704 -11208
rect 1532 -11288 2704 -11272
rect 1532 -11352 2620 -11288
rect 2684 -11352 2704 -11288
rect 1532 -11368 2704 -11352
rect 1532 -11432 2620 -11368
rect 2684 -11432 2704 -11368
rect 1532 -11448 2704 -11432
rect 1532 -11512 2620 -11448
rect 2684 -11512 2704 -11448
rect 1532 -11528 2704 -11512
rect 1532 -11592 2620 -11528
rect 2684 -11592 2704 -11528
rect 1532 -11640 2704 -11592
rect 2944 -10808 4116 -10760
rect 2944 -10872 4032 -10808
rect 4096 -10872 4116 -10808
rect 2944 -10888 4116 -10872
rect 2944 -10952 4032 -10888
rect 4096 -10952 4116 -10888
rect 2944 -10968 4116 -10952
rect 2944 -11032 4032 -10968
rect 4096 -11032 4116 -10968
rect 2944 -11048 4116 -11032
rect 2944 -11112 4032 -11048
rect 4096 -11112 4116 -11048
rect 2944 -11128 4116 -11112
rect 2944 -11192 4032 -11128
rect 4096 -11192 4116 -11128
rect 2944 -11208 4116 -11192
rect 2944 -11272 4032 -11208
rect 4096 -11272 4116 -11208
rect 2944 -11288 4116 -11272
rect 2944 -11352 4032 -11288
rect 4096 -11352 4116 -11288
rect 2944 -11368 4116 -11352
rect 2944 -11432 4032 -11368
rect 4096 -11432 4116 -11368
rect 2944 -11448 4116 -11432
rect 2944 -11512 4032 -11448
rect 4096 -11512 4116 -11448
rect 2944 -11528 4116 -11512
rect 2944 -11592 4032 -11528
rect 4096 -11592 4116 -11528
rect 2944 -11640 4116 -11592
rect 4356 -10808 5528 -10760
rect 4356 -10872 5444 -10808
rect 5508 -10872 5528 -10808
rect 4356 -10888 5528 -10872
rect 4356 -10952 5444 -10888
rect 5508 -10952 5528 -10888
rect 4356 -10968 5528 -10952
rect 4356 -11032 5444 -10968
rect 5508 -11032 5528 -10968
rect 4356 -11048 5528 -11032
rect 4356 -11112 5444 -11048
rect 5508 -11112 5528 -11048
rect 4356 -11128 5528 -11112
rect 4356 -11192 5444 -11128
rect 5508 -11192 5528 -11128
rect 4356 -11208 5528 -11192
rect 4356 -11272 5444 -11208
rect 5508 -11272 5528 -11208
rect 4356 -11288 5528 -11272
rect 4356 -11352 5444 -11288
rect 5508 -11352 5528 -11288
rect 4356 -11368 5528 -11352
rect 4356 -11432 5444 -11368
rect 5508 -11432 5528 -11368
rect 4356 -11448 5528 -11432
rect 4356 -11512 5444 -11448
rect 5508 -11512 5528 -11448
rect 4356 -11528 5528 -11512
rect 4356 -11592 5444 -11528
rect 5508 -11592 5528 -11528
rect 4356 -11640 5528 -11592
rect 5768 -10808 6940 -10760
rect 5768 -10872 6856 -10808
rect 6920 -10872 6940 -10808
rect 5768 -10888 6940 -10872
rect 5768 -10952 6856 -10888
rect 6920 -10952 6940 -10888
rect 5768 -10968 6940 -10952
rect 5768 -11032 6856 -10968
rect 6920 -11032 6940 -10968
rect 5768 -11048 6940 -11032
rect 5768 -11112 6856 -11048
rect 6920 -11112 6940 -11048
rect 5768 -11128 6940 -11112
rect 5768 -11192 6856 -11128
rect 6920 -11192 6940 -11128
rect 5768 -11208 6940 -11192
rect 5768 -11272 6856 -11208
rect 6920 -11272 6940 -11208
rect 5768 -11288 6940 -11272
rect 5768 -11352 6856 -11288
rect 6920 -11352 6940 -11288
rect 5768 -11368 6940 -11352
rect 5768 -11432 6856 -11368
rect 6920 -11432 6940 -11368
rect 5768 -11448 6940 -11432
rect 5768 -11512 6856 -11448
rect 6920 -11512 6940 -11448
rect 5768 -11528 6940 -11512
rect 5768 -11592 6856 -11528
rect 6920 -11592 6940 -11528
rect 5768 -11640 6940 -11592
rect 7180 -10808 8352 -10760
rect 7180 -10872 8268 -10808
rect 8332 -10872 8352 -10808
rect 7180 -10888 8352 -10872
rect 7180 -10952 8268 -10888
rect 8332 -10952 8352 -10888
rect 7180 -10968 8352 -10952
rect 7180 -11032 8268 -10968
rect 8332 -11032 8352 -10968
rect 7180 -11048 8352 -11032
rect 7180 -11112 8268 -11048
rect 8332 -11112 8352 -11048
rect 7180 -11128 8352 -11112
rect 7180 -11192 8268 -11128
rect 8332 -11192 8352 -11128
rect 7180 -11208 8352 -11192
rect 7180 -11272 8268 -11208
rect 8332 -11272 8352 -11208
rect 7180 -11288 8352 -11272
rect 7180 -11352 8268 -11288
rect 8332 -11352 8352 -11288
rect 7180 -11368 8352 -11352
rect 7180 -11432 8268 -11368
rect 8332 -11432 8352 -11368
rect 7180 -11448 8352 -11432
rect 7180 -11512 8268 -11448
rect 8332 -11512 8352 -11448
rect 7180 -11528 8352 -11512
rect 7180 -11592 8268 -11528
rect 8332 -11592 8352 -11528
rect 7180 -11640 8352 -11592
rect 8592 -10808 9764 -10760
rect 8592 -10872 9680 -10808
rect 9744 -10872 9764 -10808
rect 8592 -10888 9764 -10872
rect 8592 -10952 9680 -10888
rect 9744 -10952 9764 -10888
rect 8592 -10968 9764 -10952
rect 8592 -11032 9680 -10968
rect 9744 -11032 9764 -10968
rect 8592 -11048 9764 -11032
rect 8592 -11112 9680 -11048
rect 9744 -11112 9764 -11048
rect 8592 -11128 9764 -11112
rect 8592 -11192 9680 -11128
rect 9744 -11192 9764 -11128
rect 8592 -11208 9764 -11192
rect 8592 -11272 9680 -11208
rect 9744 -11272 9764 -11208
rect 8592 -11288 9764 -11272
rect 8592 -11352 9680 -11288
rect 9744 -11352 9764 -11288
rect 8592 -11368 9764 -11352
rect 8592 -11432 9680 -11368
rect 9744 -11432 9764 -11368
rect 8592 -11448 9764 -11432
rect 8592 -11512 9680 -11448
rect 9744 -11512 9764 -11448
rect 8592 -11528 9764 -11512
rect 8592 -11592 9680 -11528
rect 9744 -11592 9764 -11528
rect 8592 -11640 9764 -11592
rect 10004 -10808 11176 -10760
rect 10004 -10872 11092 -10808
rect 11156 -10872 11176 -10808
rect 10004 -10888 11176 -10872
rect 10004 -10952 11092 -10888
rect 11156 -10952 11176 -10888
rect 10004 -10968 11176 -10952
rect 10004 -11032 11092 -10968
rect 11156 -11032 11176 -10968
rect 10004 -11048 11176 -11032
rect 10004 -11112 11092 -11048
rect 11156 -11112 11176 -11048
rect 10004 -11128 11176 -11112
rect 10004 -11192 11092 -11128
rect 11156 -11192 11176 -11128
rect 10004 -11208 11176 -11192
rect 10004 -11272 11092 -11208
rect 11156 -11272 11176 -11208
rect 10004 -11288 11176 -11272
rect 10004 -11352 11092 -11288
rect 11156 -11352 11176 -11288
rect 10004 -11368 11176 -11352
rect 10004 -11432 11092 -11368
rect 11156 -11432 11176 -11368
rect 10004 -11448 11176 -11432
rect 10004 -11512 11092 -11448
rect 11156 -11512 11176 -11448
rect 10004 -11528 11176 -11512
rect 10004 -11592 11092 -11528
rect 11156 -11592 11176 -11528
rect 10004 -11640 11176 -11592
rect 11416 -10808 12588 -10760
rect 11416 -10872 12504 -10808
rect 12568 -10872 12588 -10808
rect 11416 -10888 12588 -10872
rect 11416 -10952 12504 -10888
rect 12568 -10952 12588 -10888
rect 11416 -10968 12588 -10952
rect 11416 -11032 12504 -10968
rect 12568 -11032 12588 -10968
rect 11416 -11048 12588 -11032
rect 11416 -11112 12504 -11048
rect 12568 -11112 12588 -11048
rect 11416 -11128 12588 -11112
rect 11416 -11192 12504 -11128
rect 12568 -11192 12588 -11128
rect 11416 -11208 12588 -11192
rect 11416 -11272 12504 -11208
rect 12568 -11272 12588 -11208
rect 11416 -11288 12588 -11272
rect 11416 -11352 12504 -11288
rect 12568 -11352 12588 -11288
rect 11416 -11368 12588 -11352
rect 11416 -11432 12504 -11368
rect 12568 -11432 12588 -11368
rect 11416 -11448 12588 -11432
rect 11416 -11512 12504 -11448
rect 12568 -11512 12588 -11448
rect 11416 -11528 12588 -11512
rect 11416 -11592 12504 -11528
rect 12568 -11592 12588 -11528
rect 11416 -11640 12588 -11592
rect 12828 -10808 14000 -10760
rect 12828 -10872 13916 -10808
rect 13980 -10872 14000 -10808
rect 12828 -10888 14000 -10872
rect 12828 -10952 13916 -10888
rect 13980 -10952 14000 -10888
rect 12828 -10968 14000 -10952
rect 12828 -11032 13916 -10968
rect 13980 -11032 14000 -10968
rect 12828 -11048 14000 -11032
rect 12828 -11112 13916 -11048
rect 13980 -11112 14000 -11048
rect 12828 -11128 14000 -11112
rect 12828 -11192 13916 -11128
rect 13980 -11192 14000 -11128
rect 12828 -11208 14000 -11192
rect 12828 -11272 13916 -11208
rect 13980 -11272 14000 -11208
rect 12828 -11288 14000 -11272
rect 12828 -11352 13916 -11288
rect 13980 -11352 14000 -11288
rect 12828 -11368 14000 -11352
rect 12828 -11432 13916 -11368
rect 13980 -11432 14000 -11368
rect 12828 -11448 14000 -11432
rect 12828 -11512 13916 -11448
rect 13980 -11512 14000 -11448
rect 12828 -11528 14000 -11512
rect 12828 -11592 13916 -11528
rect 13980 -11592 14000 -11528
rect 12828 -11640 14000 -11592
rect 14240 -10808 15412 -10760
rect 14240 -10872 15328 -10808
rect 15392 -10872 15412 -10808
rect 14240 -10888 15412 -10872
rect 14240 -10952 15328 -10888
rect 15392 -10952 15412 -10888
rect 14240 -10968 15412 -10952
rect 14240 -11032 15328 -10968
rect 15392 -11032 15412 -10968
rect 14240 -11048 15412 -11032
rect 14240 -11112 15328 -11048
rect 15392 -11112 15412 -11048
rect 14240 -11128 15412 -11112
rect 14240 -11192 15328 -11128
rect 15392 -11192 15412 -11128
rect 14240 -11208 15412 -11192
rect 14240 -11272 15328 -11208
rect 15392 -11272 15412 -11208
rect 14240 -11288 15412 -11272
rect 14240 -11352 15328 -11288
rect 15392 -11352 15412 -11288
rect 14240 -11368 15412 -11352
rect 14240 -11432 15328 -11368
rect 15392 -11432 15412 -11368
rect 14240 -11448 15412 -11432
rect 14240 -11512 15328 -11448
rect 15392 -11512 15412 -11448
rect 14240 -11528 15412 -11512
rect 14240 -11592 15328 -11528
rect 15392 -11592 15412 -11528
rect 14240 -11640 15412 -11592
rect 15652 -10808 16824 -10760
rect 15652 -10872 16740 -10808
rect 16804 -10872 16824 -10808
rect 15652 -10888 16824 -10872
rect 15652 -10952 16740 -10888
rect 16804 -10952 16824 -10888
rect 15652 -10968 16824 -10952
rect 15652 -11032 16740 -10968
rect 16804 -11032 16824 -10968
rect 15652 -11048 16824 -11032
rect 15652 -11112 16740 -11048
rect 16804 -11112 16824 -11048
rect 15652 -11128 16824 -11112
rect 15652 -11192 16740 -11128
rect 16804 -11192 16824 -11128
rect 15652 -11208 16824 -11192
rect 15652 -11272 16740 -11208
rect 16804 -11272 16824 -11208
rect 15652 -11288 16824 -11272
rect 15652 -11352 16740 -11288
rect 16804 -11352 16824 -11288
rect 15652 -11368 16824 -11352
rect 15652 -11432 16740 -11368
rect 16804 -11432 16824 -11368
rect 15652 -11448 16824 -11432
rect 15652 -11512 16740 -11448
rect 16804 -11512 16824 -11448
rect 15652 -11528 16824 -11512
rect 15652 -11592 16740 -11528
rect 16804 -11592 16824 -11528
rect 15652 -11640 16824 -11592
rect 17064 -10808 18236 -10760
rect 17064 -10872 18152 -10808
rect 18216 -10872 18236 -10808
rect 17064 -10888 18236 -10872
rect 17064 -10952 18152 -10888
rect 18216 -10952 18236 -10888
rect 17064 -10968 18236 -10952
rect 17064 -11032 18152 -10968
rect 18216 -11032 18236 -10968
rect 17064 -11048 18236 -11032
rect 17064 -11112 18152 -11048
rect 18216 -11112 18236 -11048
rect 17064 -11128 18236 -11112
rect 17064 -11192 18152 -11128
rect 18216 -11192 18236 -11128
rect 17064 -11208 18236 -11192
rect 17064 -11272 18152 -11208
rect 18216 -11272 18236 -11208
rect 17064 -11288 18236 -11272
rect 17064 -11352 18152 -11288
rect 18216 -11352 18236 -11288
rect 17064 -11368 18236 -11352
rect 17064 -11432 18152 -11368
rect 18216 -11432 18236 -11368
rect 17064 -11448 18236 -11432
rect 17064 -11512 18152 -11448
rect 18216 -11512 18236 -11448
rect 17064 -11528 18236 -11512
rect 17064 -11592 18152 -11528
rect 18216 -11592 18236 -11528
rect 17064 -11640 18236 -11592
rect 18476 -10808 19648 -10760
rect 18476 -10872 19564 -10808
rect 19628 -10872 19648 -10808
rect 18476 -10888 19648 -10872
rect 18476 -10952 19564 -10888
rect 19628 -10952 19648 -10888
rect 18476 -10968 19648 -10952
rect 18476 -11032 19564 -10968
rect 19628 -11032 19648 -10968
rect 18476 -11048 19648 -11032
rect 18476 -11112 19564 -11048
rect 19628 -11112 19648 -11048
rect 18476 -11128 19648 -11112
rect 18476 -11192 19564 -11128
rect 19628 -11192 19648 -11128
rect 18476 -11208 19648 -11192
rect 18476 -11272 19564 -11208
rect 19628 -11272 19648 -11208
rect 18476 -11288 19648 -11272
rect 18476 -11352 19564 -11288
rect 19628 -11352 19648 -11288
rect 18476 -11368 19648 -11352
rect 18476 -11432 19564 -11368
rect 19628 -11432 19648 -11368
rect 18476 -11448 19648 -11432
rect 18476 -11512 19564 -11448
rect 19628 -11512 19648 -11448
rect 18476 -11528 19648 -11512
rect 18476 -11592 19564 -11528
rect 19628 -11592 19648 -11528
rect 18476 -11640 19648 -11592
rect 19888 -10808 21060 -10760
rect 19888 -10872 20976 -10808
rect 21040 -10872 21060 -10808
rect 19888 -10888 21060 -10872
rect 19888 -10952 20976 -10888
rect 21040 -10952 21060 -10888
rect 19888 -10968 21060 -10952
rect 19888 -11032 20976 -10968
rect 21040 -11032 21060 -10968
rect 19888 -11048 21060 -11032
rect 19888 -11112 20976 -11048
rect 21040 -11112 21060 -11048
rect 19888 -11128 21060 -11112
rect 19888 -11192 20976 -11128
rect 21040 -11192 21060 -11128
rect 19888 -11208 21060 -11192
rect 19888 -11272 20976 -11208
rect 21040 -11272 21060 -11208
rect 19888 -11288 21060 -11272
rect 19888 -11352 20976 -11288
rect 21040 -11352 21060 -11288
rect 19888 -11368 21060 -11352
rect 19888 -11432 20976 -11368
rect 21040 -11432 21060 -11368
rect 19888 -11448 21060 -11432
rect 19888 -11512 20976 -11448
rect 21040 -11512 21060 -11448
rect 19888 -11528 21060 -11512
rect 19888 -11592 20976 -11528
rect 21040 -11592 21060 -11528
rect 19888 -11640 21060 -11592
rect 21300 -10808 22472 -10760
rect 21300 -10872 22388 -10808
rect 22452 -10872 22472 -10808
rect 21300 -10888 22472 -10872
rect 21300 -10952 22388 -10888
rect 22452 -10952 22472 -10888
rect 21300 -10968 22472 -10952
rect 21300 -11032 22388 -10968
rect 22452 -11032 22472 -10968
rect 21300 -11048 22472 -11032
rect 21300 -11112 22388 -11048
rect 22452 -11112 22472 -11048
rect 21300 -11128 22472 -11112
rect 21300 -11192 22388 -11128
rect 22452 -11192 22472 -11128
rect 21300 -11208 22472 -11192
rect 21300 -11272 22388 -11208
rect 22452 -11272 22472 -11208
rect 21300 -11288 22472 -11272
rect 21300 -11352 22388 -11288
rect 22452 -11352 22472 -11288
rect 21300 -11368 22472 -11352
rect 21300 -11432 22388 -11368
rect 22452 -11432 22472 -11368
rect 21300 -11448 22472 -11432
rect 21300 -11512 22388 -11448
rect 22452 -11512 22472 -11448
rect 21300 -11528 22472 -11512
rect 21300 -11592 22388 -11528
rect 22452 -11592 22472 -11528
rect 21300 -11640 22472 -11592
rect 22712 -10808 23884 -10760
rect 22712 -10872 23800 -10808
rect 23864 -10872 23884 -10808
rect 22712 -10888 23884 -10872
rect 22712 -10952 23800 -10888
rect 23864 -10952 23884 -10888
rect 22712 -10968 23884 -10952
rect 22712 -11032 23800 -10968
rect 23864 -11032 23884 -10968
rect 22712 -11048 23884 -11032
rect 22712 -11112 23800 -11048
rect 23864 -11112 23884 -11048
rect 22712 -11128 23884 -11112
rect 22712 -11192 23800 -11128
rect 23864 -11192 23884 -11128
rect 22712 -11208 23884 -11192
rect 22712 -11272 23800 -11208
rect 23864 -11272 23884 -11208
rect 22712 -11288 23884 -11272
rect 22712 -11352 23800 -11288
rect 23864 -11352 23884 -11288
rect 22712 -11368 23884 -11352
rect 22712 -11432 23800 -11368
rect 23864 -11432 23884 -11368
rect 22712 -11448 23884 -11432
rect 22712 -11512 23800 -11448
rect 23864 -11512 23884 -11448
rect 22712 -11528 23884 -11512
rect 22712 -11592 23800 -11528
rect 23864 -11592 23884 -11528
rect 22712 -11640 23884 -11592
rect -23884 -11928 -22712 -11880
rect -23884 -11992 -22796 -11928
rect -22732 -11992 -22712 -11928
rect -23884 -12008 -22712 -11992
rect -23884 -12072 -22796 -12008
rect -22732 -12072 -22712 -12008
rect -23884 -12088 -22712 -12072
rect -23884 -12152 -22796 -12088
rect -22732 -12152 -22712 -12088
rect -23884 -12168 -22712 -12152
rect -23884 -12232 -22796 -12168
rect -22732 -12232 -22712 -12168
rect -23884 -12248 -22712 -12232
rect -23884 -12312 -22796 -12248
rect -22732 -12312 -22712 -12248
rect -23884 -12328 -22712 -12312
rect -23884 -12392 -22796 -12328
rect -22732 -12392 -22712 -12328
rect -23884 -12408 -22712 -12392
rect -23884 -12472 -22796 -12408
rect -22732 -12472 -22712 -12408
rect -23884 -12488 -22712 -12472
rect -23884 -12552 -22796 -12488
rect -22732 -12552 -22712 -12488
rect -23884 -12568 -22712 -12552
rect -23884 -12632 -22796 -12568
rect -22732 -12632 -22712 -12568
rect -23884 -12648 -22712 -12632
rect -23884 -12712 -22796 -12648
rect -22732 -12712 -22712 -12648
rect -23884 -12760 -22712 -12712
rect -22472 -11928 -21300 -11880
rect -22472 -11992 -21384 -11928
rect -21320 -11992 -21300 -11928
rect -22472 -12008 -21300 -11992
rect -22472 -12072 -21384 -12008
rect -21320 -12072 -21300 -12008
rect -22472 -12088 -21300 -12072
rect -22472 -12152 -21384 -12088
rect -21320 -12152 -21300 -12088
rect -22472 -12168 -21300 -12152
rect -22472 -12232 -21384 -12168
rect -21320 -12232 -21300 -12168
rect -22472 -12248 -21300 -12232
rect -22472 -12312 -21384 -12248
rect -21320 -12312 -21300 -12248
rect -22472 -12328 -21300 -12312
rect -22472 -12392 -21384 -12328
rect -21320 -12392 -21300 -12328
rect -22472 -12408 -21300 -12392
rect -22472 -12472 -21384 -12408
rect -21320 -12472 -21300 -12408
rect -22472 -12488 -21300 -12472
rect -22472 -12552 -21384 -12488
rect -21320 -12552 -21300 -12488
rect -22472 -12568 -21300 -12552
rect -22472 -12632 -21384 -12568
rect -21320 -12632 -21300 -12568
rect -22472 -12648 -21300 -12632
rect -22472 -12712 -21384 -12648
rect -21320 -12712 -21300 -12648
rect -22472 -12760 -21300 -12712
rect -21060 -11928 -19888 -11880
rect -21060 -11992 -19972 -11928
rect -19908 -11992 -19888 -11928
rect -21060 -12008 -19888 -11992
rect -21060 -12072 -19972 -12008
rect -19908 -12072 -19888 -12008
rect -21060 -12088 -19888 -12072
rect -21060 -12152 -19972 -12088
rect -19908 -12152 -19888 -12088
rect -21060 -12168 -19888 -12152
rect -21060 -12232 -19972 -12168
rect -19908 -12232 -19888 -12168
rect -21060 -12248 -19888 -12232
rect -21060 -12312 -19972 -12248
rect -19908 -12312 -19888 -12248
rect -21060 -12328 -19888 -12312
rect -21060 -12392 -19972 -12328
rect -19908 -12392 -19888 -12328
rect -21060 -12408 -19888 -12392
rect -21060 -12472 -19972 -12408
rect -19908 -12472 -19888 -12408
rect -21060 -12488 -19888 -12472
rect -21060 -12552 -19972 -12488
rect -19908 -12552 -19888 -12488
rect -21060 -12568 -19888 -12552
rect -21060 -12632 -19972 -12568
rect -19908 -12632 -19888 -12568
rect -21060 -12648 -19888 -12632
rect -21060 -12712 -19972 -12648
rect -19908 -12712 -19888 -12648
rect -21060 -12760 -19888 -12712
rect -19648 -11928 -18476 -11880
rect -19648 -11992 -18560 -11928
rect -18496 -11992 -18476 -11928
rect -19648 -12008 -18476 -11992
rect -19648 -12072 -18560 -12008
rect -18496 -12072 -18476 -12008
rect -19648 -12088 -18476 -12072
rect -19648 -12152 -18560 -12088
rect -18496 -12152 -18476 -12088
rect -19648 -12168 -18476 -12152
rect -19648 -12232 -18560 -12168
rect -18496 -12232 -18476 -12168
rect -19648 -12248 -18476 -12232
rect -19648 -12312 -18560 -12248
rect -18496 -12312 -18476 -12248
rect -19648 -12328 -18476 -12312
rect -19648 -12392 -18560 -12328
rect -18496 -12392 -18476 -12328
rect -19648 -12408 -18476 -12392
rect -19648 -12472 -18560 -12408
rect -18496 -12472 -18476 -12408
rect -19648 -12488 -18476 -12472
rect -19648 -12552 -18560 -12488
rect -18496 -12552 -18476 -12488
rect -19648 -12568 -18476 -12552
rect -19648 -12632 -18560 -12568
rect -18496 -12632 -18476 -12568
rect -19648 -12648 -18476 -12632
rect -19648 -12712 -18560 -12648
rect -18496 -12712 -18476 -12648
rect -19648 -12760 -18476 -12712
rect -18236 -11928 -17064 -11880
rect -18236 -11992 -17148 -11928
rect -17084 -11992 -17064 -11928
rect -18236 -12008 -17064 -11992
rect -18236 -12072 -17148 -12008
rect -17084 -12072 -17064 -12008
rect -18236 -12088 -17064 -12072
rect -18236 -12152 -17148 -12088
rect -17084 -12152 -17064 -12088
rect -18236 -12168 -17064 -12152
rect -18236 -12232 -17148 -12168
rect -17084 -12232 -17064 -12168
rect -18236 -12248 -17064 -12232
rect -18236 -12312 -17148 -12248
rect -17084 -12312 -17064 -12248
rect -18236 -12328 -17064 -12312
rect -18236 -12392 -17148 -12328
rect -17084 -12392 -17064 -12328
rect -18236 -12408 -17064 -12392
rect -18236 -12472 -17148 -12408
rect -17084 -12472 -17064 -12408
rect -18236 -12488 -17064 -12472
rect -18236 -12552 -17148 -12488
rect -17084 -12552 -17064 -12488
rect -18236 -12568 -17064 -12552
rect -18236 -12632 -17148 -12568
rect -17084 -12632 -17064 -12568
rect -18236 -12648 -17064 -12632
rect -18236 -12712 -17148 -12648
rect -17084 -12712 -17064 -12648
rect -18236 -12760 -17064 -12712
rect -16824 -11928 -15652 -11880
rect -16824 -11992 -15736 -11928
rect -15672 -11992 -15652 -11928
rect -16824 -12008 -15652 -11992
rect -16824 -12072 -15736 -12008
rect -15672 -12072 -15652 -12008
rect -16824 -12088 -15652 -12072
rect -16824 -12152 -15736 -12088
rect -15672 -12152 -15652 -12088
rect -16824 -12168 -15652 -12152
rect -16824 -12232 -15736 -12168
rect -15672 -12232 -15652 -12168
rect -16824 -12248 -15652 -12232
rect -16824 -12312 -15736 -12248
rect -15672 -12312 -15652 -12248
rect -16824 -12328 -15652 -12312
rect -16824 -12392 -15736 -12328
rect -15672 -12392 -15652 -12328
rect -16824 -12408 -15652 -12392
rect -16824 -12472 -15736 -12408
rect -15672 -12472 -15652 -12408
rect -16824 -12488 -15652 -12472
rect -16824 -12552 -15736 -12488
rect -15672 -12552 -15652 -12488
rect -16824 -12568 -15652 -12552
rect -16824 -12632 -15736 -12568
rect -15672 -12632 -15652 -12568
rect -16824 -12648 -15652 -12632
rect -16824 -12712 -15736 -12648
rect -15672 -12712 -15652 -12648
rect -16824 -12760 -15652 -12712
rect -15412 -11928 -14240 -11880
rect -15412 -11992 -14324 -11928
rect -14260 -11992 -14240 -11928
rect -15412 -12008 -14240 -11992
rect -15412 -12072 -14324 -12008
rect -14260 -12072 -14240 -12008
rect -15412 -12088 -14240 -12072
rect -15412 -12152 -14324 -12088
rect -14260 -12152 -14240 -12088
rect -15412 -12168 -14240 -12152
rect -15412 -12232 -14324 -12168
rect -14260 -12232 -14240 -12168
rect -15412 -12248 -14240 -12232
rect -15412 -12312 -14324 -12248
rect -14260 -12312 -14240 -12248
rect -15412 -12328 -14240 -12312
rect -15412 -12392 -14324 -12328
rect -14260 -12392 -14240 -12328
rect -15412 -12408 -14240 -12392
rect -15412 -12472 -14324 -12408
rect -14260 -12472 -14240 -12408
rect -15412 -12488 -14240 -12472
rect -15412 -12552 -14324 -12488
rect -14260 -12552 -14240 -12488
rect -15412 -12568 -14240 -12552
rect -15412 -12632 -14324 -12568
rect -14260 -12632 -14240 -12568
rect -15412 -12648 -14240 -12632
rect -15412 -12712 -14324 -12648
rect -14260 -12712 -14240 -12648
rect -15412 -12760 -14240 -12712
rect -14000 -11928 -12828 -11880
rect -14000 -11992 -12912 -11928
rect -12848 -11992 -12828 -11928
rect -14000 -12008 -12828 -11992
rect -14000 -12072 -12912 -12008
rect -12848 -12072 -12828 -12008
rect -14000 -12088 -12828 -12072
rect -14000 -12152 -12912 -12088
rect -12848 -12152 -12828 -12088
rect -14000 -12168 -12828 -12152
rect -14000 -12232 -12912 -12168
rect -12848 -12232 -12828 -12168
rect -14000 -12248 -12828 -12232
rect -14000 -12312 -12912 -12248
rect -12848 -12312 -12828 -12248
rect -14000 -12328 -12828 -12312
rect -14000 -12392 -12912 -12328
rect -12848 -12392 -12828 -12328
rect -14000 -12408 -12828 -12392
rect -14000 -12472 -12912 -12408
rect -12848 -12472 -12828 -12408
rect -14000 -12488 -12828 -12472
rect -14000 -12552 -12912 -12488
rect -12848 -12552 -12828 -12488
rect -14000 -12568 -12828 -12552
rect -14000 -12632 -12912 -12568
rect -12848 -12632 -12828 -12568
rect -14000 -12648 -12828 -12632
rect -14000 -12712 -12912 -12648
rect -12848 -12712 -12828 -12648
rect -14000 -12760 -12828 -12712
rect -12588 -11928 -11416 -11880
rect -12588 -11992 -11500 -11928
rect -11436 -11992 -11416 -11928
rect -12588 -12008 -11416 -11992
rect -12588 -12072 -11500 -12008
rect -11436 -12072 -11416 -12008
rect -12588 -12088 -11416 -12072
rect -12588 -12152 -11500 -12088
rect -11436 -12152 -11416 -12088
rect -12588 -12168 -11416 -12152
rect -12588 -12232 -11500 -12168
rect -11436 -12232 -11416 -12168
rect -12588 -12248 -11416 -12232
rect -12588 -12312 -11500 -12248
rect -11436 -12312 -11416 -12248
rect -12588 -12328 -11416 -12312
rect -12588 -12392 -11500 -12328
rect -11436 -12392 -11416 -12328
rect -12588 -12408 -11416 -12392
rect -12588 -12472 -11500 -12408
rect -11436 -12472 -11416 -12408
rect -12588 -12488 -11416 -12472
rect -12588 -12552 -11500 -12488
rect -11436 -12552 -11416 -12488
rect -12588 -12568 -11416 -12552
rect -12588 -12632 -11500 -12568
rect -11436 -12632 -11416 -12568
rect -12588 -12648 -11416 -12632
rect -12588 -12712 -11500 -12648
rect -11436 -12712 -11416 -12648
rect -12588 -12760 -11416 -12712
rect -11176 -11928 -10004 -11880
rect -11176 -11992 -10088 -11928
rect -10024 -11992 -10004 -11928
rect -11176 -12008 -10004 -11992
rect -11176 -12072 -10088 -12008
rect -10024 -12072 -10004 -12008
rect -11176 -12088 -10004 -12072
rect -11176 -12152 -10088 -12088
rect -10024 -12152 -10004 -12088
rect -11176 -12168 -10004 -12152
rect -11176 -12232 -10088 -12168
rect -10024 -12232 -10004 -12168
rect -11176 -12248 -10004 -12232
rect -11176 -12312 -10088 -12248
rect -10024 -12312 -10004 -12248
rect -11176 -12328 -10004 -12312
rect -11176 -12392 -10088 -12328
rect -10024 -12392 -10004 -12328
rect -11176 -12408 -10004 -12392
rect -11176 -12472 -10088 -12408
rect -10024 -12472 -10004 -12408
rect -11176 -12488 -10004 -12472
rect -11176 -12552 -10088 -12488
rect -10024 -12552 -10004 -12488
rect -11176 -12568 -10004 -12552
rect -11176 -12632 -10088 -12568
rect -10024 -12632 -10004 -12568
rect -11176 -12648 -10004 -12632
rect -11176 -12712 -10088 -12648
rect -10024 -12712 -10004 -12648
rect -11176 -12760 -10004 -12712
rect -9764 -11928 -8592 -11880
rect -9764 -11992 -8676 -11928
rect -8612 -11992 -8592 -11928
rect -9764 -12008 -8592 -11992
rect -9764 -12072 -8676 -12008
rect -8612 -12072 -8592 -12008
rect -9764 -12088 -8592 -12072
rect -9764 -12152 -8676 -12088
rect -8612 -12152 -8592 -12088
rect -9764 -12168 -8592 -12152
rect -9764 -12232 -8676 -12168
rect -8612 -12232 -8592 -12168
rect -9764 -12248 -8592 -12232
rect -9764 -12312 -8676 -12248
rect -8612 -12312 -8592 -12248
rect -9764 -12328 -8592 -12312
rect -9764 -12392 -8676 -12328
rect -8612 -12392 -8592 -12328
rect -9764 -12408 -8592 -12392
rect -9764 -12472 -8676 -12408
rect -8612 -12472 -8592 -12408
rect -9764 -12488 -8592 -12472
rect -9764 -12552 -8676 -12488
rect -8612 -12552 -8592 -12488
rect -9764 -12568 -8592 -12552
rect -9764 -12632 -8676 -12568
rect -8612 -12632 -8592 -12568
rect -9764 -12648 -8592 -12632
rect -9764 -12712 -8676 -12648
rect -8612 -12712 -8592 -12648
rect -9764 -12760 -8592 -12712
rect -8352 -11928 -7180 -11880
rect -8352 -11992 -7264 -11928
rect -7200 -11992 -7180 -11928
rect -8352 -12008 -7180 -11992
rect -8352 -12072 -7264 -12008
rect -7200 -12072 -7180 -12008
rect -8352 -12088 -7180 -12072
rect -8352 -12152 -7264 -12088
rect -7200 -12152 -7180 -12088
rect -8352 -12168 -7180 -12152
rect -8352 -12232 -7264 -12168
rect -7200 -12232 -7180 -12168
rect -8352 -12248 -7180 -12232
rect -8352 -12312 -7264 -12248
rect -7200 -12312 -7180 -12248
rect -8352 -12328 -7180 -12312
rect -8352 -12392 -7264 -12328
rect -7200 -12392 -7180 -12328
rect -8352 -12408 -7180 -12392
rect -8352 -12472 -7264 -12408
rect -7200 -12472 -7180 -12408
rect -8352 -12488 -7180 -12472
rect -8352 -12552 -7264 -12488
rect -7200 -12552 -7180 -12488
rect -8352 -12568 -7180 -12552
rect -8352 -12632 -7264 -12568
rect -7200 -12632 -7180 -12568
rect -8352 -12648 -7180 -12632
rect -8352 -12712 -7264 -12648
rect -7200 -12712 -7180 -12648
rect -8352 -12760 -7180 -12712
rect -6940 -11928 -5768 -11880
rect -6940 -11992 -5852 -11928
rect -5788 -11992 -5768 -11928
rect -6940 -12008 -5768 -11992
rect -6940 -12072 -5852 -12008
rect -5788 -12072 -5768 -12008
rect -6940 -12088 -5768 -12072
rect -6940 -12152 -5852 -12088
rect -5788 -12152 -5768 -12088
rect -6940 -12168 -5768 -12152
rect -6940 -12232 -5852 -12168
rect -5788 -12232 -5768 -12168
rect -6940 -12248 -5768 -12232
rect -6940 -12312 -5852 -12248
rect -5788 -12312 -5768 -12248
rect -6940 -12328 -5768 -12312
rect -6940 -12392 -5852 -12328
rect -5788 -12392 -5768 -12328
rect -6940 -12408 -5768 -12392
rect -6940 -12472 -5852 -12408
rect -5788 -12472 -5768 -12408
rect -6940 -12488 -5768 -12472
rect -6940 -12552 -5852 -12488
rect -5788 -12552 -5768 -12488
rect -6940 -12568 -5768 -12552
rect -6940 -12632 -5852 -12568
rect -5788 -12632 -5768 -12568
rect -6940 -12648 -5768 -12632
rect -6940 -12712 -5852 -12648
rect -5788 -12712 -5768 -12648
rect -6940 -12760 -5768 -12712
rect -5528 -11928 -4356 -11880
rect -5528 -11992 -4440 -11928
rect -4376 -11992 -4356 -11928
rect -5528 -12008 -4356 -11992
rect -5528 -12072 -4440 -12008
rect -4376 -12072 -4356 -12008
rect -5528 -12088 -4356 -12072
rect -5528 -12152 -4440 -12088
rect -4376 -12152 -4356 -12088
rect -5528 -12168 -4356 -12152
rect -5528 -12232 -4440 -12168
rect -4376 -12232 -4356 -12168
rect -5528 -12248 -4356 -12232
rect -5528 -12312 -4440 -12248
rect -4376 -12312 -4356 -12248
rect -5528 -12328 -4356 -12312
rect -5528 -12392 -4440 -12328
rect -4376 -12392 -4356 -12328
rect -5528 -12408 -4356 -12392
rect -5528 -12472 -4440 -12408
rect -4376 -12472 -4356 -12408
rect -5528 -12488 -4356 -12472
rect -5528 -12552 -4440 -12488
rect -4376 -12552 -4356 -12488
rect -5528 -12568 -4356 -12552
rect -5528 -12632 -4440 -12568
rect -4376 -12632 -4356 -12568
rect -5528 -12648 -4356 -12632
rect -5528 -12712 -4440 -12648
rect -4376 -12712 -4356 -12648
rect -5528 -12760 -4356 -12712
rect -4116 -11928 -2944 -11880
rect -4116 -11992 -3028 -11928
rect -2964 -11992 -2944 -11928
rect -4116 -12008 -2944 -11992
rect -4116 -12072 -3028 -12008
rect -2964 -12072 -2944 -12008
rect -4116 -12088 -2944 -12072
rect -4116 -12152 -3028 -12088
rect -2964 -12152 -2944 -12088
rect -4116 -12168 -2944 -12152
rect -4116 -12232 -3028 -12168
rect -2964 -12232 -2944 -12168
rect -4116 -12248 -2944 -12232
rect -4116 -12312 -3028 -12248
rect -2964 -12312 -2944 -12248
rect -4116 -12328 -2944 -12312
rect -4116 -12392 -3028 -12328
rect -2964 -12392 -2944 -12328
rect -4116 -12408 -2944 -12392
rect -4116 -12472 -3028 -12408
rect -2964 -12472 -2944 -12408
rect -4116 -12488 -2944 -12472
rect -4116 -12552 -3028 -12488
rect -2964 -12552 -2944 -12488
rect -4116 -12568 -2944 -12552
rect -4116 -12632 -3028 -12568
rect -2964 -12632 -2944 -12568
rect -4116 -12648 -2944 -12632
rect -4116 -12712 -3028 -12648
rect -2964 -12712 -2944 -12648
rect -4116 -12760 -2944 -12712
rect -2704 -11928 -1532 -11880
rect -2704 -11992 -1616 -11928
rect -1552 -11992 -1532 -11928
rect -2704 -12008 -1532 -11992
rect -2704 -12072 -1616 -12008
rect -1552 -12072 -1532 -12008
rect -2704 -12088 -1532 -12072
rect -2704 -12152 -1616 -12088
rect -1552 -12152 -1532 -12088
rect -2704 -12168 -1532 -12152
rect -2704 -12232 -1616 -12168
rect -1552 -12232 -1532 -12168
rect -2704 -12248 -1532 -12232
rect -2704 -12312 -1616 -12248
rect -1552 -12312 -1532 -12248
rect -2704 -12328 -1532 -12312
rect -2704 -12392 -1616 -12328
rect -1552 -12392 -1532 -12328
rect -2704 -12408 -1532 -12392
rect -2704 -12472 -1616 -12408
rect -1552 -12472 -1532 -12408
rect -2704 -12488 -1532 -12472
rect -2704 -12552 -1616 -12488
rect -1552 -12552 -1532 -12488
rect -2704 -12568 -1532 -12552
rect -2704 -12632 -1616 -12568
rect -1552 -12632 -1532 -12568
rect -2704 -12648 -1532 -12632
rect -2704 -12712 -1616 -12648
rect -1552 -12712 -1532 -12648
rect -2704 -12760 -1532 -12712
rect -1292 -11928 -120 -11880
rect -1292 -11992 -204 -11928
rect -140 -11992 -120 -11928
rect -1292 -12008 -120 -11992
rect -1292 -12072 -204 -12008
rect -140 -12072 -120 -12008
rect -1292 -12088 -120 -12072
rect -1292 -12152 -204 -12088
rect -140 -12152 -120 -12088
rect -1292 -12168 -120 -12152
rect -1292 -12232 -204 -12168
rect -140 -12232 -120 -12168
rect -1292 -12248 -120 -12232
rect -1292 -12312 -204 -12248
rect -140 -12312 -120 -12248
rect -1292 -12328 -120 -12312
rect -1292 -12392 -204 -12328
rect -140 -12392 -120 -12328
rect -1292 -12408 -120 -12392
rect -1292 -12472 -204 -12408
rect -140 -12472 -120 -12408
rect -1292 -12488 -120 -12472
rect -1292 -12552 -204 -12488
rect -140 -12552 -120 -12488
rect -1292 -12568 -120 -12552
rect -1292 -12632 -204 -12568
rect -140 -12632 -120 -12568
rect -1292 -12648 -120 -12632
rect -1292 -12712 -204 -12648
rect -140 -12712 -120 -12648
rect -1292 -12760 -120 -12712
rect 120 -11928 1292 -11880
rect 120 -11992 1208 -11928
rect 1272 -11992 1292 -11928
rect 120 -12008 1292 -11992
rect 120 -12072 1208 -12008
rect 1272 -12072 1292 -12008
rect 120 -12088 1292 -12072
rect 120 -12152 1208 -12088
rect 1272 -12152 1292 -12088
rect 120 -12168 1292 -12152
rect 120 -12232 1208 -12168
rect 1272 -12232 1292 -12168
rect 120 -12248 1292 -12232
rect 120 -12312 1208 -12248
rect 1272 -12312 1292 -12248
rect 120 -12328 1292 -12312
rect 120 -12392 1208 -12328
rect 1272 -12392 1292 -12328
rect 120 -12408 1292 -12392
rect 120 -12472 1208 -12408
rect 1272 -12472 1292 -12408
rect 120 -12488 1292 -12472
rect 120 -12552 1208 -12488
rect 1272 -12552 1292 -12488
rect 120 -12568 1292 -12552
rect 120 -12632 1208 -12568
rect 1272 -12632 1292 -12568
rect 120 -12648 1292 -12632
rect 120 -12712 1208 -12648
rect 1272 -12712 1292 -12648
rect 120 -12760 1292 -12712
rect 1532 -11928 2704 -11880
rect 1532 -11992 2620 -11928
rect 2684 -11992 2704 -11928
rect 1532 -12008 2704 -11992
rect 1532 -12072 2620 -12008
rect 2684 -12072 2704 -12008
rect 1532 -12088 2704 -12072
rect 1532 -12152 2620 -12088
rect 2684 -12152 2704 -12088
rect 1532 -12168 2704 -12152
rect 1532 -12232 2620 -12168
rect 2684 -12232 2704 -12168
rect 1532 -12248 2704 -12232
rect 1532 -12312 2620 -12248
rect 2684 -12312 2704 -12248
rect 1532 -12328 2704 -12312
rect 1532 -12392 2620 -12328
rect 2684 -12392 2704 -12328
rect 1532 -12408 2704 -12392
rect 1532 -12472 2620 -12408
rect 2684 -12472 2704 -12408
rect 1532 -12488 2704 -12472
rect 1532 -12552 2620 -12488
rect 2684 -12552 2704 -12488
rect 1532 -12568 2704 -12552
rect 1532 -12632 2620 -12568
rect 2684 -12632 2704 -12568
rect 1532 -12648 2704 -12632
rect 1532 -12712 2620 -12648
rect 2684 -12712 2704 -12648
rect 1532 -12760 2704 -12712
rect 2944 -11928 4116 -11880
rect 2944 -11992 4032 -11928
rect 4096 -11992 4116 -11928
rect 2944 -12008 4116 -11992
rect 2944 -12072 4032 -12008
rect 4096 -12072 4116 -12008
rect 2944 -12088 4116 -12072
rect 2944 -12152 4032 -12088
rect 4096 -12152 4116 -12088
rect 2944 -12168 4116 -12152
rect 2944 -12232 4032 -12168
rect 4096 -12232 4116 -12168
rect 2944 -12248 4116 -12232
rect 2944 -12312 4032 -12248
rect 4096 -12312 4116 -12248
rect 2944 -12328 4116 -12312
rect 2944 -12392 4032 -12328
rect 4096 -12392 4116 -12328
rect 2944 -12408 4116 -12392
rect 2944 -12472 4032 -12408
rect 4096 -12472 4116 -12408
rect 2944 -12488 4116 -12472
rect 2944 -12552 4032 -12488
rect 4096 -12552 4116 -12488
rect 2944 -12568 4116 -12552
rect 2944 -12632 4032 -12568
rect 4096 -12632 4116 -12568
rect 2944 -12648 4116 -12632
rect 2944 -12712 4032 -12648
rect 4096 -12712 4116 -12648
rect 2944 -12760 4116 -12712
rect 4356 -11928 5528 -11880
rect 4356 -11992 5444 -11928
rect 5508 -11992 5528 -11928
rect 4356 -12008 5528 -11992
rect 4356 -12072 5444 -12008
rect 5508 -12072 5528 -12008
rect 4356 -12088 5528 -12072
rect 4356 -12152 5444 -12088
rect 5508 -12152 5528 -12088
rect 4356 -12168 5528 -12152
rect 4356 -12232 5444 -12168
rect 5508 -12232 5528 -12168
rect 4356 -12248 5528 -12232
rect 4356 -12312 5444 -12248
rect 5508 -12312 5528 -12248
rect 4356 -12328 5528 -12312
rect 4356 -12392 5444 -12328
rect 5508 -12392 5528 -12328
rect 4356 -12408 5528 -12392
rect 4356 -12472 5444 -12408
rect 5508 -12472 5528 -12408
rect 4356 -12488 5528 -12472
rect 4356 -12552 5444 -12488
rect 5508 -12552 5528 -12488
rect 4356 -12568 5528 -12552
rect 4356 -12632 5444 -12568
rect 5508 -12632 5528 -12568
rect 4356 -12648 5528 -12632
rect 4356 -12712 5444 -12648
rect 5508 -12712 5528 -12648
rect 4356 -12760 5528 -12712
rect 5768 -11928 6940 -11880
rect 5768 -11992 6856 -11928
rect 6920 -11992 6940 -11928
rect 5768 -12008 6940 -11992
rect 5768 -12072 6856 -12008
rect 6920 -12072 6940 -12008
rect 5768 -12088 6940 -12072
rect 5768 -12152 6856 -12088
rect 6920 -12152 6940 -12088
rect 5768 -12168 6940 -12152
rect 5768 -12232 6856 -12168
rect 6920 -12232 6940 -12168
rect 5768 -12248 6940 -12232
rect 5768 -12312 6856 -12248
rect 6920 -12312 6940 -12248
rect 5768 -12328 6940 -12312
rect 5768 -12392 6856 -12328
rect 6920 -12392 6940 -12328
rect 5768 -12408 6940 -12392
rect 5768 -12472 6856 -12408
rect 6920 -12472 6940 -12408
rect 5768 -12488 6940 -12472
rect 5768 -12552 6856 -12488
rect 6920 -12552 6940 -12488
rect 5768 -12568 6940 -12552
rect 5768 -12632 6856 -12568
rect 6920 -12632 6940 -12568
rect 5768 -12648 6940 -12632
rect 5768 -12712 6856 -12648
rect 6920 -12712 6940 -12648
rect 5768 -12760 6940 -12712
rect 7180 -11928 8352 -11880
rect 7180 -11992 8268 -11928
rect 8332 -11992 8352 -11928
rect 7180 -12008 8352 -11992
rect 7180 -12072 8268 -12008
rect 8332 -12072 8352 -12008
rect 7180 -12088 8352 -12072
rect 7180 -12152 8268 -12088
rect 8332 -12152 8352 -12088
rect 7180 -12168 8352 -12152
rect 7180 -12232 8268 -12168
rect 8332 -12232 8352 -12168
rect 7180 -12248 8352 -12232
rect 7180 -12312 8268 -12248
rect 8332 -12312 8352 -12248
rect 7180 -12328 8352 -12312
rect 7180 -12392 8268 -12328
rect 8332 -12392 8352 -12328
rect 7180 -12408 8352 -12392
rect 7180 -12472 8268 -12408
rect 8332 -12472 8352 -12408
rect 7180 -12488 8352 -12472
rect 7180 -12552 8268 -12488
rect 8332 -12552 8352 -12488
rect 7180 -12568 8352 -12552
rect 7180 -12632 8268 -12568
rect 8332 -12632 8352 -12568
rect 7180 -12648 8352 -12632
rect 7180 -12712 8268 -12648
rect 8332 -12712 8352 -12648
rect 7180 -12760 8352 -12712
rect 8592 -11928 9764 -11880
rect 8592 -11992 9680 -11928
rect 9744 -11992 9764 -11928
rect 8592 -12008 9764 -11992
rect 8592 -12072 9680 -12008
rect 9744 -12072 9764 -12008
rect 8592 -12088 9764 -12072
rect 8592 -12152 9680 -12088
rect 9744 -12152 9764 -12088
rect 8592 -12168 9764 -12152
rect 8592 -12232 9680 -12168
rect 9744 -12232 9764 -12168
rect 8592 -12248 9764 -12232
rect 8592 -12312 9680 -12248
rect 9744 -12312 9764 -12248
rect 8592 -12328 9764 -12312
rect 8592 -12392 9680 -12328
rect 9744 -12392 9764 -12328
rect 8592 -12408 9764 -12392
rect 8592 -12472 9680 -12408
rect 9744 -12472 9764 -12408
rect 8592 -12488 9764 -12472
rect 8592 -12552 9680 -12488
rect 9744 -12552 9764 -12488
rect 8592 -12568 9764 -12552
rect 8592 -12632 9680 -12568
rect 9744 -12632 9764 -12568
rect 8592 -12648 9764 -12632
rect 8592 -12712 9680 -12648
rect 9744 -12712 9764 -12648
rect 8592 -12760 9764 -12712
rect 10004 -11928 11176 -11880
rect 10004 -11992 11092 -11928
rect 11156 -11992 11176 -11928
rect 10004 -12008 11176 -11992
rect 10004 -12072 11092 -12008
rect 11156 -12072 11176 -12008
rect 10004 -12088 11176 -12072
rect 10004 -12152 11092 -12088
rect 11156 -12152 11176 -12088
rect 10004 -12168 11176 -12152
rect 10004 -12232 11092 -12168
rect 11156 -12232 11176 -12168
rect 10004 -12248 11176 -12232
rect 10004 -12312 11092 -12248
rect 11156 -12312 11176 -12248
rect 10004 -12328 11176 -12312
rect 10004 -12392 11092 -12328
rect 11156 -12392 11176 -12328
rect 10004 -12408 11176 -12392
rect 10004 -12472 11092 -12408
rect 11156 -12472 11176 -12408
rect 10004 -12488 11176 -12472
rect 10004 -12552 11092 -12488
rect 11156 -12552 11176 -12488
rect 10004 -12568 11176 -12552
rect 10004 -12632 11092 -12568
rect 11156 -12632 11176 -12568
rect 10004 -12648 11176 -12632
rect 10004 -12712 11092 -12648
rect 11156 -12712 11176 -12648
rect 10004 -12760 11176 -12712
rect 11416 -11928 12588 -11880
rect 11416 -11992 12504 -11928
rect 12568 -11992 12588 -11928
rect 11416 -12008 12588 -11992
rect 11416 -12072 12504 -12008
rect 12568 -12072 12588 -12008
rect 11416 -12088 12588 -12072
rect 11416 -12152 12504 -12088
rect 12568 -12152 12588 -12088
rect 11416 -12168 12588 -12152
rect 11416 -12232 12504 -12168
rect 12568 -12232 12588 -12168
rect 11416 -12248 12588 -12232
rect 11416 -12312 12504 -12248
rect 12568 -12312 12588 -12248
rect 11416 -12328 12588 -12312
rect 11416 -12392 12504 -12328
rect 12568 -12392 12588 -12328
rect 11416 -12408 12588 -12392
rect 11416 -12472 12504 -12408
rect 12568 -12472 12588 -12408
rect 11416 -12488 12588 -12472
rect 11416 -12552 12504 -12488
rect 12568 -12552 12588 -12488
rect 11416 -12568 12588 -12552
rect 11416 -12632 12504 -12568
rect 12568 -12632 12588 -12568
rect 11416 -12648 12588 -12632
rect 11416 -12712 12504 -12648
rect 12568 -12712 12588 -12648
rect 11416 -12760 12588 -12712
rect 12828 -11928 14000 -11880
rect 12828 -11992 13916 -11928
rect 13980 -11992 14000 -11928
rect 12828 -12008 14000 -11992
rect 12828 -12072 13916 -12008
rect 13980 -12072 14000 -12008
rect 12828 -12088 14000 -12072
rect 12828 -12152 13916 -12088
rect 13980 -12152 14000 -12088
rect 12828 -12168 14000 -12152
rect 12828 -12232 13916 -12168
rect 13980 -12232 14000 -12168
rect 12828 -12248 14000 -12232
rect 12828 -12312 13916 -12248
rect 13980 -12312 14000 -12248
rect 12828 -12328 14000 -12312
rect 12828 -12392 13916 -12328
rect 13980 -12392 14000 -12328
rect 12828 -12408 14000 -12392
rect 12828 -12472 13916 -12408
rect 13980 -12472 14000 -12408
rect 12828 -12488 14000 -12472
rect 12828 -12552 13916 -12488
rect 13980 -12552 14000 -12488
rect 12828 -12568 14000 -12552
rect 12828 -12632 13916 -12568
rect 13980 -12632 14000 -12568
rect 12828 -12648 14000 -12632
rect 12828 -12712 13916 -12648
rect 13980 -12712 14000 -12648
rect 12828 -12760 14000 -12712
rect 14240 -11928 15412 -11880
rect 14240 -11992 15328 -11928
rect 15392 -11992 15412 -11928
rect 14240 -12008 15412 -11992
rect 14240 -12072 15328 -12008
rect 15392 -12072 15412 -12008
rect 14240 -12088 15412 -12072
rect 14240 -12152 15328 -12088
rect 15392 -12152 15412 -12088
rect 14240 -12168 15412 -12152
rect 14240 -12232 15328 -12168
rect 15392 -12232 15412 -12168
rect 14240 -12248 15412 -12232
rect 14240 -12312 15328 -12248
rect 15392 -12312 15412 -12248
rect 14240 -12328 15412 -12312
rect 14240 -12392 15328 -12328
rect 15392 -12392 15412 -12328
rect 14240 -12408 15412 -12392
rect 14240 -12472 15328 -12408
rect 15392 -12472 15412 -12408
rect 14240 -12488 15412 -12472
rect 14240 -12552 15328 -12488
rect 15392 -12552 15412 -12488
rect 14240 -12568 15412 -12552
rect 14240 -12632 15328 -12568
rect 15392 -12632 15412 -12568
rect 14240 -12648 15412 -12632
rect 14240 -12712 15328 -12648
rect 15392 -12712 15412 -12648
rect 14240 -12760 15412 -12712
rect 15652 -11928 16824 -11880
rect 15652 -11992 16740 -11928
rect 16804 -11992 16824 -11928
rect 15652 -12008 16824 -11992
rect 15652 -12072 16740 -12008
rect 16804 -12072 16824 -12008
rect 15652 -12088 16824 -12072
rect 15652 -12152 16740 -12088
rect 16804 -12152 16824 -12088
rect 15652 -12168 16824 -12152
rect 15652 -12232 16740 -12168
rect 16804 -12232 16824 -12168
rect 15652 -12248 16824 -12232
rect 15652 -12312 16740 -12248
rect 16804 -12312 16824 -12248
rect 15652 -12328 16824 -12312
rect 15652 -12392 16740 -12328
rect 16804 -12392 16824 -12328
rect 15652 -12408 16824 -12392
rect 15652 -12472 16740 -12408
rect 16804 -12472 16824 -12408
rect 15652 -12488 16824 -12472
rect 15652 -12552 16740 -12488
rect 16804 -12552 16824 -12488
rect 15652 -12568 16824 -12552
rect 15652 -12632 16740 -12568
rect 16804 -12632 16824 -12568
rect 15652 -12648 16824 -12632
rect 15652 -12712 16740 -12648
rect 16804 -12712 16824 -12648
rect 15652 -12760 16824 -12712
rect 17064 -11928 18236 -11880
rect 17064 -11992 18152 -11928
rect 18216 -11992 18236 -11928
rect 17064 -12008 18236 -11992
rect 17064 -12072 18152 -12008
rect 18216 -12072 18236 -12008
rect 17064 -12088 18236 -12072
rect 17064 -12152 18152 -12088
rect 18216 -12152 18236 -12088
rect 17064 -12168 18236 -12152
rect 17064 -12232 18152 -12168
rect 18216 -12232 18236 -12168
rect 17064 -12248 18236 -12232
rect 17064 -12312 18152 -12248
rect 18216 -12312 18236 -12248
rect 17064 -12328 18236 -12312
rect 17064 -12392 18152 -12328
rect 18216 -12392 18236 -12328
rect 17064 -12408 18236 -12392
rect 17064 -12472 18152 -12408
rect 18216 -12472 18236 -12408
rect 17064 -12488 18236 -12472
rect 17064 -12552 18152 -12488
rect 18216 -12552 18236 -12488
rect 17064 -12568 18236 -12552
rect 17064 -12632 18152 -12568
rect 18216 -12632 18236 -12568
rect 17064 -12648 18236 -12632
rect 17064 -12712 18152 -12648
rect 18216 -12712 18236 -12648
rect 17064 -12760 18236 -12712
rect 18476 -11928 19648 -11880
rect 18476 -11992 19564 -11928
rect 19628 -11992 19648 -11928
rect 18476 -12008 19648 -11992
rect 18476 -12072 19564 -12008
rect 19628 -12072 19648 -12008
rect 18476 -12088 19648 -12072
rect 18476 -12152 19564 -12088
rect 19628 -12152 19648 -12088
rect 18476 -12168 19648 -12152
rect 18476 -12232 19564 -12168
rect 19628 -12232 19648 -12168
rect 18476 -12248 19648 -12232
rect 18476 -12312 19564 -12248
rect 19628 -12312 19648 -12248
rect 18476 -12328 19648 -12312
rect 18476 -12392 19564 -12328
rect 19628 -12392 19648 -12328
rect 18476 -12408 19648 -12392
rect 18476 -12472 19564 -12408
rect 19628 -12472 19648 -12408
rect 18476 -12488 19648 -12472
rect 18476 -12552 19564 -12488
rect 19628 -12552 19648 -12488
rect 18476 -12568 19648 -12552
rect 18476 -12632 19564 -12568
rect 19628 -12632 19648 -12568
rect 18476 -12648 19648 -12632
rect 18476 -12712 19564 -12648
rect 19628 -12712 19648 -12648
rect 18476 -12760 19648 -12712
rect 19888 -11928 21060 -11880
rect 19888 -11992 20976 -11928
rect 21040 -11992 21060 -11928
rect 19888 -12008 21060 -11992
rect 19888 -12072 20976 -12008
rect 21040 -12072 21060 -12008
rect 19888 -12088 21060 -12072
rect 19888 -12152 20976 -12088
rect 21040 -12152 21060 -12088
rect 19888 -12168 21060 -12152
rect 19888 -12232 20976 -12168
rect 21040 -12232 21060 -12168
rect 19888 -12248 21060 -12232
rect 19888 -12312 20976 -12248
rect 21040 -12312 21060 -12248
rect 19888 -12328 21060 -12312
rect 19888 -12392 20976 -12328
rect 21040 -12392 21060 -12328
rect 19888 -12408 21060 -12392
rect 19888 -12472 20976 -12408
rect 21040 -12472 21060 -12408
rect 19888 -12488 21060 -12472
rect 19888 -12552 20976 -12488
rect 21040 -12552 21060 -12488
rect 19888 -12568 21060 -12552
rect 19888 -12632 20976 -12568
rect 21040 -12632 21060 -12568
rect 19888 -12648 21060 -12632
rect 19888 -12712 20976 -12648
rect 21040 -12712 21060 -12648
rect 19888 -12760 21060 -12712
rect 21300 -11928 22472 -11880
rect 21300 -11992 22388 -11928
rect 22452 -11992 22472 -11928
rect 21300 -12008 22472 -11992
rect 21300 -12072 22388 -12008
rect 22452 -12072 22472 -12008
rect 21300 -12088 22472 -12072
rect 21300 -12152 22388 -12088
rect 22452 -12152 22472 -12088
rect 21300 -12168 22472 -12152
rect 21300 -12232 22388 -12168
rect 22452 -12232 22472 -12168
rect 21300 -12248 22472 -12232
rect 21300 -12312 22388 -12248
rect 22452 -12312 22472 -12248
rect 21300 -12328 22472 -12312
rect 21300 -12392 22388 -12328
rect 22452 -12392 22472 -12328
rect 21300 -12408 22472 -12392
rect 21300 -12472 22388 -12408
rect 22452 -12472 22472 -12408
rect 21300 -12488 22472 -12472
rect 21300 -12552 22388 -12488
rect 22452 -12552 22472 -12488
rect 21300 -12568 22472 -12552
rect 21300 -12632 22388 -12568
rect 22452 -12632 22472 -12568
rect 21300 -12648 22472 -12632
rect 21300 -12712 22388 -12648
rect 22452 -12712 22472 -12648
rect 21300 -12760 22472 -12712
rect 22712 -11928 23884 -11880
rect 22712 -11992 23800 -11928
rect 23864 -11992 23884 -11928
rect 22712 -12008 23884 -11992
rect 22712 -12072 23800 -12008
rect 23864 -12072 23884 -12008
rect 22712 -12088 23884 -12072
rect 22712 -12152 23800 -12088
rect 23864 -12152 23884 -12088
rect 22712 -12168 23884 -12152
rect 22712 -12232 23800 -12168
rect 23864 -12232 23884 -12168
rect 22712 -12248 23884 -12232
rect 22712 -12312 23800 -12248
rect 23864 -12312 23884 -12248
rect 22712 -12328 23884 -12312
rect 22712 -12392 23800 -12328
rect 23864 -12392 23884 -12328
rect 22712 -12408 23884 -12392
rect 22712 -12472 23800 -12408
rect 23864 -12472 23884 -12408
rect 22712 -12488 23884 -12472
rect 22712 -12552 23800 -12488
rect 23864 -12552 23884 -12488
rect 22712 -12568 23884 -12552
rect 22712 -12632 23800 -12568
rect 23864 -12632 23884 -12568
rect 22712 -12648 23884 -12632
rect 22712 -12712 23800 -12648
rect 23864 -12712 23884 -12648
rect 22712 -12760 23884 -12712
rect -23884 -13048 -22712 -13000
rect -23884 -13112 -22796 -13048
rect -22732 -13112 -22712 -13048
rect -23884 -13128 -22712 -13112
rect -23884 -13192 -22796 -13128
rect -22732 -13192 -22712 -13128
rect -23884 -13208 -22712 -13192
rect -23884 -13272 -22796 -13208
rect -22732 -13272 -22712 -13208
rect -23884 -13288 -22712 -13272
rect -23884 -13352 -22796 -13288
rect -22732 -13352 -22712 -13288
rect -23884 -13368 -22712 -13352
rect -23884 -13432 -22796 -13368
rect -22732 -13432 -22712 -13368
rect -23884 -13448 -22712 -13432
rect -23884 -13512 -22796 -13448
rect -22732 -13512 -22712 -13448
rect -23884 -13528 -22712 -13512
rect -23884 -13592 -22796 -13528
rect -22732 -13592 -22712 -13528
rect -23884 -13608 -22712 -13592
rect -23884 -13672 -22796 -13608
rect -22732 -13672 -22712 -13608
rect -23884 -13688 -22712 -13672
rect -23884 -13752 -22796 -13688
rect -22732 -13752 -22712 -13688
rect -23884 -13768 -22712 -13752
rect -23884 -13832 -22796 -13768
rect -22732 -13832 -22712 -13768
rect -23884 -13880 -22712 -13832
rect -22472 -13048 -21300 -13000
rect -22472 -13112 -21384 -13048
rect -21320 -13112 -21300 -13048
rect -22472 -13128 -21300 -13112
rect -22472 -13192 -21384 -13128
rect -21320 -13192 -21300 -13128
rect -22472 -13208 -21300 -13192
rect -22472 -13272 -21384 -13208
rect -21320 -13272 -21300 -13208
rect -22472 -13288 -21300 -13272
rect -22472 -13352 -21384 -13288
rect -21320 -13352 -21300 -13288
rect -22472 -13368 -21300 -13352
rect -22472 -13432 -21384 -13368
rect -21320 -13432 -21300 -13368
rect -22472 -13448 -21300 -13432
rect -22472 -13512 -21384 -13448
rect -21320 -13512 -21300 -13448
rect -22472 -13528 -21300 -13512
rect -22472 -13592 -21384 -13528
rect -21320 -13592 -21300 -13528
rect -22472 -13608 -21300 -13592
rect -22472 -13672 -21384 -13608
rect -21320 -13672 -21300 -13608
rect -22472 -13688 -21300 -13672
rect -22472 -13752 -21384 -13688
rect -21320 -13752 -21300 -13688
rect -22472 -13768 -21300 -13752
rect -22472 -13832 -21384 -13768
rect -21320 -13832 -21300 -13768
rect -22472 -13880 -21300 -13832
rect -21060 -13048 -19888 -13000
rect -21060 -13112 -19972 -13048
rect -19908 -13112 -19888 -13048
rect -21060 -13128 -19888 -13112
rect -21060 -13192 -19972 -13128
rect -19908 -13192 -19888 -13128
rect -21060 -13208 -19888 -13192
rect -21060 -13272 -19972 -13208
rect -19908 -13272 -19888 -13208
rect -21060 -13288 -19888 -13272
rect -21060 -13352 -19972 -13288
rect -19908 -13352 -19888 -13288
rect -21060 -13368 -19888 -13352
rect -21060 -13432 -19972 -13368
rect -19908 -13432 -19888 -13368
rect -21060 -13448 -19888 -13432
rect -21060 -13512 -19972 -13448
rect -19908 -13512 -19888 -13448
rect -21060 -13528 -19888 -13512
rect -21060 -13592 -19972 -13528
rect -19908 -13592 -19888 -13528
rect -21060 -13608 -19888 -13592
rect -21060 -13672 -19972 -13608
rect -19908 -13672 -19888 -13608
rect -21060 -13688 -19888 -13672
rect -21060 -13752 -19972 -13688
rect -19908 -13752 -19888 -13688
rect -21060 -13768 -19888 -13752
rect -21060 -13832 -19972 -13768
rect -19908 -13832 -19888 -13768
rect -21060 -13880 -19888 -13832
rect -19648 -13048 -18476 -13000
rect -19648 -13112 -18560 -13048
rect -18496 -13112 -18476 -13048
rect -19648 -13128 -18476 -13112
rect -19648 -13192 -18560 -13128
rect -18496 -13192 -18476 -13128
rect -19648 -13208 -18476 -13192
rect -19648 -13272 -18560 -13208
rect -18496 -13272 -18476 -13208
rect -19648 -13288 -18476 -13272
rect -19648 -13352 -18560 -13288
rect -18496 -13352 -18476 -13288
rect -19648 -13368 -18476 -13352
rect -19648 -13432 -18560 -13368
rect -18496 -13432 -18476 -13368
rect -19648 -13448 -18476 -13432
rect -19648 -13512 -18560 -13448
rect -18496 -13512 -18476 -13448
rect -19648 -13528 -18476 -13512
rect -19648 -13592 -18560 -13528
rect -18496 -13592 -18476 -13528
rect -19648 -13608 -18476 -13592
rect -19648 -13672 -18560 -13608
rect -18496 -13672 -18476 -13608
rect -19648 -13688 -18476 -13672
rect -19648 -13752 -18560 -13688
rect -18496 -13752 -18476 -13688
rect -19648 -13768 -18476 -13752
rect -19648 -13832 -18560 -13768
rect -18496 -13832 -18476 -13768
rect -19648 -13880 -18476 -13832
rect -18236 -13048 -17064 -13000
rect -18236 -13112 -17148 -13048
rect -17084 -13112 -17064 -13048
rect -18236 -13128 -17064 -13112
rect -18236 -13192 -17148 -13128
rect -17084 -13192 -17064 -13128
rect -18236 -13208 -17064 -13192
rect -18236 -13272 -17148 -13208
rect -17084 -13272 -17064 -13208
rect -18236 -13288 -17064 -13272
rect -18236 -13352 -17148 -13288
rect -17084 -13352 -17064 -13288
rect -18236 -13368 -17064 -13352
rect -18236 -13432 -17148 -13368
rect -17084 -13432 -17064 -13368
rect -18236 -13448 -17064 -13432
rect -18236 -13512 -17148 -13448
rect -17084 -13512 -17064 -13448
rect -18236 -13528 -17064 -13512
rect -18236 -13592 -17148 -13528
rect -17084 -13592 -17064 -13528
rect -18236 -13608 -17064 -13592
rect -18236 -13672 -17148 -13608
rect -17084 -13672 -17064 -13608
rect -18236 -13688 -17064 -13672
rect -18236 -13752 -17148 -13688
rect -17084 -13752 -17064 -13688
rect -18236 -13768 -17064 -13752
rect -18236 -13832 -17148 -13768
rect -17084 -13832 -17064 -13768
rect -18236 -13880 -17064 -13832
rect -16824 -13048 -15652 -13000
rect -16824 -13112 -15736 -13048
rect -15672 -13112 -15652 -13048
rect -16824 -13128 -15652 -13112
rect -16824 -13192 -15736 -13128
rect -15672 -13192 -15652 -13128
rect -16824 -13208 -15652 -13192
rect -16824 -13272 -15736 -13208
rect -15672 -13272 -15652 -13208
rect -16824 -13288 -15652 -13272
rect -16824 -13352 -15736 -13288
rect -15672 -13352 -15652 -13288
rect -16824 -13368 -15652 -13352
rect -16824 -13432 -15736 -13368
rect -15672 -13432 -15652 -13368
rect -16824 -13448 -15652 -13432
rect -16824 -13512 -15736 -13448
rect -15672 -13512 -15652 -13448
rect -16824 -13528 -15652 -13512
rect -16824 -13592 -15736 -13528
rect -15672 -13592 -15652 -13528
rect -16824 -13608 -15652 -13592
rect -16824 -13672 -15736 -13608
rect -15672 -13672 -15652 -13608
rect -16824 -13688 -15652 -13672
rect -16824 -13752 -15736 -13688
rect -15672 -13752 -15652 -13688
rect -16824 -13768 -15652 -13752
rect -16824 -13832 -15736 -13768
rect -15672 -13832 -15652 -13768
rect -16824 -13880 -15652 -13832
rect -15412 -13048 -14240 -13000
rect -15412 -13112 -14324 -13048
rect -14260 -13112 -14240 -13048
rect -15412 -13128 -14240 -13112
rect -15412 -13192 -14324 -13128
rect -14260 -13192 -14240 -13128
rect -15412 -13208 -14240 -13192
rect -15412 -13272 -14324 -13208
rect -14260 -13272 -14240 -13208
rect -15412 -13288 -14240 -13272
rect -15412 -13352 -14324 -13288
rect -14260 -13352 -14240 -13288
rect -15412 -13368 -14240 -13352
rect -15412 -13432 -14324 -13368
rect -14260 -13432 -14240 -13368
rect -15412 -13448 -14240 -13432
rect -15412 -13512 -14324 -13448
rect -14260 -13512 -14240 -13448
rect -15412 -13528 -14240 -13512
rect -15412 -13592 -14324 -13528
rect -14260 -13592 -14240 -13528
rect -15412 -13608 -14240 -13592
rect -15412 -13672 -14324 -13608
rect -14260 -13672 -14240 -13608
rect -15412 -13688 -14240 -13672
rect -15412 -13752 -14324 -13688
rect -14260 -13752 -14240 -13688
rect -15412 -13768 -14240 -13752
rect -15412 -13832 -14324 -13768
rect -14260 -13832 -14240 -13768
rect -15412 -13880 -14240 -13832
rect -14000 -13048 -12828 -13000
rect -14000 -13112 -12912 -13048
rect -12848 -13112 -12828 -13048
rect -14000 -13128 -12828 -13112
rect -14000 -13192 -12912 -13128
rect -12848 -13192 -12828 -13128
rect -14000 -13208 -12828 -13192
rect -14000 -13272 -12912 -13208
rect -12848 -13272 -12828 -13208
rect -14000 -13288 -12828 -13272
rect -14000 -13352 -12912 -13288
rect -12848 -13352 -12828 -13288
rect -14000 -13368 -12828 -13352
rect -14000 -13432 -12912 -13368
rect -12848 -13432 -12828 -13368
rect -14000 -13448 -12828 -13432
rect -14000 -13512 -12912 -13448
rect -12848 -13512 -12828 -13448
rect -14000 -13528 -12828 -13512
rect -14000 -13592 -12912 -13528
rect -12848 -13592 -12828 -13528
rect -14000 -13608 -12828 -13592
rect -14000 -13672 -12912 -13608
rect -12848 -13672 -12828 -13608
rect -14000 -13688 -12828 -13672
rect -14000 -13752 -12912 -13688
rect -12848 -13752 -12828 -13688
rect -14000 -13768 -12828 -13752
rect -14000 -13832 -12912 -13768
rect -12848 -13832 -12828 -13768
rect -14000 -13880 -12828 -13832
rect -12588 -13048 -11416 -13000
rect -12588 -13112 -11500 -13048
rect -11436 -13112 -11416 -13048
rect -12588 -13128 -11416 -13112
rect -12588 -13192 -11500 -13128
rect -11436 -13192 -11416 -13128
rect -12588 -13208 -11416 -13192
rect -12588 -13272 -11500 -13208
rect -11436 -13272 -11416 -13208
rect -12588 -13288 -11416 -13272
rect -12588 -13352 -11500 -13288
rect -11436 -13352 -11416 -13288
rect -12588 -13368 -11416 -13352
rect -12588 -13432 -11500 -13368
rect -11436 -13432 -11416 -13368
rect -12588 -13448 -11416 -13432
rect -12588 -13512 -11500 -13448
rect -11436 -13512 -11416 -13448
rect -12588 -13528 -11416 -13512
rect -12588 -13592 -11500 -13528
rect -11436 -13592 -11416 -13528
rect -12588 -13608 -11416 -13592
rect -12588 -13672 -11500 -13608
rect -11436 -13672 -11416 -13608
rect -12588 -13688 -11416 -13672
rect -12588 -13752 -11500 -13688
rect -11436 -13752 -11416 -13688
rect -12588 -13768 -11416 -13752
rect -12588 -13832 -11500 -13768
rect -11436 -13832 -11416 -13768
rect -12588 -13880 -11416 -13832
rect -11176 -13048 -10004 -13000
rect -11176 -13112 -10088 -13048
rect -10024 -13112 -10004 -13048
rect -11176 -13128 -10004 -13112
rect -11176 -13192 -10088 -13128
rect -10024 -13192 -10004 -13128
rect -11176 -13208 -10004 -13192
rect -11176 -13272 -10088 -13208
rect -10024 -13272 -10004 -13208
rect -11176 -13288 -10004 -13272
rect -11176 -13352 -10088 -13288
rect -10024 -13352 -10004 -13288
rect -11176 -13368 -10004 -13352
rect -11176 -13432 -10088 -13368
rect -10024 -13432 -10004 -13368
rect -11176 -13448 -10004 -13432
rect -11176 -13512 -10088 -13448
rect -10024 -13512 -10004 -13448
rect -11176 -13528 -10004 -13512
rect -11176 -13592 -10088 -13528
rect -10024 -13592 -10004 -13528
rect -11176 -13608 -10004 -13592
rect -11176 -13672 -10088 -13608
rect -10024 -13672 -10004 -13608
rect -11176 -13688 -10004 -13672
rect -11176 -13752 -10088 -13688
rect -10024 -13752 -10004 -13688
rect -11176 -13768 -10004 -13752
rect -11176 -13832 -10088 -13768
rect -10024 -13832 -10004 -13768
rect -11176 -13880 -10004 -13832
rect -9764 -13048 -8592 -13000
rect -9764 -13112 -8676 -13048
rect -8612 -13112 -8592 -13048
rect -9764 -13128 -8592 -13112
rect -9764 -13192 -8676 -13128
rect -8612 -13192 -8592 -13128
rect -9764 -13208 -8592 -13192
rect -9764 -13272 -8676 -13208
rect -8612 -13272 -8592 -13208
rect -9764 -13288 -8592 -13272
rect -9764 -13352 -8676 -13288
rect -8612 -13352 -8592 -13288
rect -9764 -13368 -8592 -13352
rect -9764 -13432 -8676 -13368
rect -8612 -13432 -8592 -13368
rect -9764 -13448 -8592 -13432
rect -9764 -13512 -8676 -13448
rect -8612 -13512 -8592 -13448
rect -9764 -13528 -8592 -13512
rect -9764 -13592 -8676 -13528
rect -8612 -13592 -8592 -13528
rect -9764 -13608 -8592 -13592
rect -9764 -13672 -8676 -13608
rect -8612 -13672 -8592 -13608
rect -9764 -13688 -8592 -13672
rect -9764 -13752 -8676 -13688
rect -8612 -13752 -8592 -13688
rect -9764 -13768 -8592 -13752
rect -9764 -13832 -8676 -13768
rect -8612 -13832 -8592 -13768
rect -9764 -13880 -8592 -13832
rect -8352 -13048 -7180 -13000
rect -8352 -13112 -7264 -13048
rect -7200 -13112 -7180 -13048
rect -8352 -13128 -7180 -13112
rect -8352 -13192 -7264 -13128
rect -7200 -13192 -7180 -13128
rect -8352 -13208 -7180 -13192
rect -8352 -13272 -7264 -13208
rect -7200 -13272 -7180 -13208
rect -8352 -13288 -7180 -13272
rect -8352 -13352 -7264 -13288
rect -7200 -13352 -7180 -13288
rect -8352 -13368 -7180 -13352
rect -8352 -13432 -7264 -13368
rect -7200 -13432 -7180 -13368
rect -8352 -13448 -7180 -13432
rect -8352 -13512 -7264 -13448
rect -7200 -13512 -7180 -13448
rect -8352 -13528 -7180 -13512
rect -8352 -13592 -7264 -13528
rect -7200 -13592 -7180 -13528
rect -8352 -13608 -7180 -13592
rect -8352 -13672 -7264 -13608
rect -7200 -13672 -7180 -13608
rect -8352 -13688 -7180 -13672
rect -8352 -13752 -7264 -13688
rect -7200 -13752 -7180 -13688
rect -8352 -13768 -7180 -13752
rect -8352 -13832 -7264 -13768
rect -7200 -13832 -7180 -13768
rect -8352 -13880 -7180 -13832
rect -6940 -13048 -5768 -13000
rect -6940 -13112 -5852 -13048
rect -5788 -13112 -5768 -13048
rect -6940 -13128 -5768 -13112
rect -6940 -13192 -5852 -13128
rect -5788 -13192 -5768 -13128
rect -6940 -13208 -5768 -13192
rect -6940 -13272 -5852 -13208
rect -5788 -13272 -5768 -13208
rect -6940 -13288 -5768 -13272
rect -6940 -13352 -5852 -13288
rect -5788 -13352 -5768 -13288
rect -6940 -13368 -5768 -13352
rect -6940 -13432 -5852 -13368
rect -5788 -13432 -5768 -13368
rect -6940 -13448 -5768 -13432
rect -6940 -13512 -5852 -13448
rect -5788 -13512 -5768 -13448
rect -6940 -13528 -5768 -13512
rect -6940 -13592 -5852 -13528
rect -5788 -13592 -5768 -13528
rect -6940 -13608 -5768 -13592
rect -6940 -13672 -5852 -13608
rect -5788 -13672 -5768 -13608
rect -6940 -13688 -5768 -13672
rect -6940 -13752 -5852 -13688
rect -5788 -13752 -5768 -13688
rect -6940 -13768 -5768 -13752
rect -6940 -13832 -5852 -13768
rect -5788 -13832 -5768 -13768
rect -6940 -13880 -5768 -13832
rect -5528 -13048 -4356 -13000
rect -5528 -13112 -4440 -13048
rect -4376 -13112 -4356 -13048
rect -5528 -13128 -4356 -13112
rect -5528 -13192 -4440 -13128
rect -4376 -13192 -4356 -13128
rect -5528 -13208 -4356 -13192
rect -5528 -13272 -4440 -13208
rect -4376 -13272 -4356 -13208
rect -5528 -13288 -4356 -13272
rect -5528 -13352 -4440 -13288
rect -4376 -13352 -4356 -13288
rect -5528 -13368 -4356 -13352
rect -5528 -13432 -4440 -13368
rect -4376 -13432 -4356 -13368
rect -5528 -13448 -4356 -13432
rect -5528 -13512 -4440 -13448
rect -4376 -13512 -4356 -13448
rect -5528 -13528 -4356 -13512
rect -5528 -13592 -4440 -13528
rect -4376 -13592 -4356 -13528
rect -5528 -13608 -4356 -13592
rect -5528 -13672 -4440 -13608
rect -4376 -13672 -4356 -13608
rect -5528 -13688 -4356 -13672
rect -5528 -13752 -4440 -13688
rect -4376 -13752 -4356 -13688
rect -5528 -13768 -4356 -13752
rect -5528 -13832 -4440 -13768
rect -4376 -13832 -4356 -13768
rect -5528 -13880 -4356 -13832
rect -4116 -13048 -2944 -13000
rect -4116 -13112 -3028 -13048
rect -2964 -13112 -2944 -13048
rect -4116 -13128 -2944 -13112
rect -4116 -13192 -3028 -13128
rect -2964 -13192 -2944 -13128
rect -4116 -13208 -2944 -13192
rect -4116 -13272 -3028 -13208
rect -2964 -13272 -2944 -13208
rect -4116 -13288 -2944 -13272
rect -4116 -13352 -3028 -13288
rect -2964 -13352 -2944 -13288
rect -4116 -13368 -2944 -13352
rect -4116 -13432 -3028 -13368
rect -2964 -13432 -2944 -13368
rect -4116 -13448 -2944 -13432
rect -4116 -13512 -3028 -13448
rect -2964 -13512 -2944 -13448
rect -4116 -13528 -2944 -13512
rect -4116 -13592 -3028 -13528
rect -2964 -13592 -2944 -13528
rect -4116 -13608 -2944 -13592
rect -4116 -13672 -3028 -13608
rect -2964 -13672 -2944 -13608
rect -4116 -13688 -2944 -13672
rect -4116 -13752 -3028 -13688
rect -2964 -13752 -2944 -13688
rect -4116 -13768 -2944 -13752
rect -4116 -13832 -3028 -13768
rect -2964 -13832 -2944 -13768
rect -4116 -13880 -2944 -13832
rect -2704 -13048 -1532 -13000
rect -2704 -13112 -1616 -13048
rect -1552 -13112 -1532 -13048
rect -2704 -13128 -1532 -13112
rect -2704 -13192 -1616 -13128
rect -1552 -13192 -1532 -13128
rect -2704 -13208 -1532 -13192
rect -2704 -13272 -1616 -13208
rect -1552 -13272 -1532 -13208
rect -2704 -13288 -1532 -13272
rect -2704 -13352 -1616 -13288
rect -1552 -13352 -1532 -13288
rect -2704 -13368 -1532 -13352
rect -2704 -13432 -1616 -13368
rect -1552 -13432 -1532 -13368
rect -2704 -13448 -1532 -13432
rect -2704 -13512 -1616 -13448
rect -1552 -13512 -1532 -13448
rect -2704 -13528 -1532 -13512
rect -2704 -13592 -1616 -13528
rect -1552 -13592 -1532 -13528
rect -2704 -13608 -1532 -13592
rect -2704 -13672 -1616 -13608
rect -1552 -13672 -1532 -13608
rect -2704 -13688 -1532 -13672
rect -2704 -13752 -1616 -13688
rect -1552 -13752 -1532 -13688
rect -2704 -13768 -1532 -13752
rect -2704 -13832 -1616 -13768
rect -1552 -13832 -1532 -13768
rect -2704 -13880 -1532 -13832
rect -1292 -13048 -120 -13000
rect -1292 -13112 -204 -13048
rect -140 -13112 -120 -13048
rect -1292 -13128 -120 -13112
rect -1292 -13192 -204 -13128
rect -140 -13192 -120 -13128
rect -1292 -13208 -120 -13192
rect -1292 -13272 -204 -13208
rect -140 -13272 -120 -13208
rect -1292 -13288 -120 -13272
rect -1292 -13352 -204 -13288
rect -140 -13352 -120 -13288
rect -1292 -13368 -120 -13352
rect -1292 -13432 -204 -13368
rect -140 -13432 -120 -13368
rect -1292 -13448 -120 -13432
rect -1292 -13512 -204 -13448
rect -140 -13512 -120 -13448
rect -1292 -13528 -120 -13512
rect -1292 -13592 -204 -13528
rect -140 -13592 -120 -13528
rect -1292 -13608 -120 -13592
rect -1292 -13672 -204 -13608
rect -140 -13672 -120 -13608
rect -1292 -13688 -120 -13672
rect -1292 -13752 -204 -13688
rect -140 -13752 -120 -13688
rect -1292 -13768 -120 -13752
rect -1292 -13832 -204 -13768
rect -140 -13832 -120 -13768
rect -1292 -13880 -120 -13832
rect 120 -13048 1292 -13000
rect 120 -13112 1208 -13048
rect 1272 -13112 1292 -13048
rect 120 -13128 1292 -13112
rect 120 -13192 1208 -13128
rect 1272 -13192 1292 -13128
rect 120 -13208 1292 -13192
rect 120 -13272 1208 -13208
rect 1272 -13272 1292 -13208
rect 120 -13288 1292 -13272
rect 120 -13352 1208 -13288
rect 1272 -13352 1292 -13288
rect 120 -13368 1292 -13352
rect 120 -13432 1208 -13368
rect 1272 -13432 1292 -13368
rect 120 -13448 1292 -13432
rect 120 -13512 1208 -13448
rect 1272 -13512 1292 -13448
rect 120 -13528 1292 -13512
rect 120 -13592 1208 -13528
rect 1272 -13592 1292 -13528
rect 120 -13608 1292 -13592
rect 120 -13672 1208 -13608
rect 1272 -13672 1292 -13608
rect 120 -13688 1292 -13672
rect 120 -13752 1208 -13688
rect 1272 -13752 1292 -13688
rect 120 -13768 1292 -13752
rect 120 -13832 1208 -13768
rect 1272 -13832 1292 -13768
rect 120 -13880 1292 -13832
rect 1532 -13048 2704 -13000
rect 1532 -13112 2620 -13048
rect 2684 -13112 2704 -13048
rect 1532 -13128 2704 -13112
rect 1532 -13192 2620 -13128
rect 2684 -13192 2704 -13128
rect 1532 -13208 2704 -13192
rect 1532 -13272 2620 -13208
rect 2684 -13272 2704 -13208
rect 1532 -13288 2704 -13272
rect 1532 -13352 2620 -13288
rect 2684 -13352 2704 -13288
rect 1532 -13368 2704 -13352
rect 1532 -13432 2620 -13368
rect 2684 -13432 2704 -13368
rect 1532 -13448 2704 -13432
rect 1532 -13512 2620 -13448
rect 2684 -13512 2704 -13448
rect 1532 -13528 2704 -13512
rect 1532 -13592 2620 -13528
rect 2684 -13592 2704 -13528
rect 1532 -13608 2704 -13592
rect 1532 -13672 2620 -13608
rect 2684 -13672 2704 -13608
rect 1532 -13688 2704 -13672
rect 1532 -13752 2620 -13688
rect 2684 -13752 2704 -13688
rect 1532 -13768 2704 -13752
rect 1532 -13832 2620 -13768
rect 2684 -13832 2704 -13768
rect 1532 -13880 2704 -13832
rect 2944 -13048 4116 -13000
rect 2944 -13112 4032 -13048
rect 4096 -13112 4116 -13048
rect 2944 -13128 4116 -13112
rect 2944 -13192 4032 -13128
rect 4096 -13192 4116 -13128
rect 2944 -13208 4116 -13192
rect 2944 -13272 4032 -13208
rect 4096 -13272 4116 -13208
rect 2944 -13288 4116 -13272
rect 2944 -13352 4032 -13288
rect 4096 -13352 4116 -13288
rect 2944 -13368 4116 -13352
rect 2944 -13432 4032 -13368
rect 4096 -13432 4116 -13368
rect 2944 -13448 4116 -13432
rect 2944 -13512 4032 -13448
rect 4096 -13512 4116 -13448
rect 2944 -13528 4116 -13512
rect 2944 -13592 4032 -13528
rect 4096 -13592 4116 -13528
rect 2944 -13608 4116 -13592
rect 2944 -13672 4032 -13608
rect 4096 -13672 4116 -13608
rect 2944 -13688 4116 -13672
rect 2944 -13752 4032 -13688
rect 4096 -13752 4116 -13688
rect 2944 -13768 4116 -13752
rect 2944 -13832 4032 -13768
rect 4096 -13832 4116 -13768
rect 2944 -13880 4116 -13832
rect 4356 -13048 5528 -13000
rect 4356 -13112 5444 -13048
rect 5508 -13112 5528 -13048
rect 4356 -13128 5528 -13112
rect 4356 -13192 5444 -13128
rect 5508 -13192 5528 -13128
rect 4356 -13208 5528 -13192
rect 4356 -13272 5444 -13208
rect 5508 -13272 5528 -13208
rect 4356 -13288 5528 -13272
rect 4356 -13352 5444 -13288
rect 5508 -13352 5528 -13288
rect 4356 -13368 5528 -13352
rect 4356 -13432 5444 -13368
rect 5508 -13432 5528 -13368
rect 4356 -13448 5528 -13432
rect 4356 -13512 5444 -13448
rect 5508 -13512 5528 -13448
rect 4356 -13528 5528 -13512
rect 4356 -13592 5444 -13528
rect 5508 -13592 5528 -13528
rect 4356 -13608 5528 -13592
rect 4356 -13672 5444 -13608
rect 5508 -13672 5528 -13608
rect 4356 -13688 5528 -13672
rect 4356 -13752 5444 -13688
rect 5508 -13752 5528 -13688
rect 4356 -13768 5528 -13752
rect 4356 -13832 5444 -13768
rect 5508 -13832 5528 -13768
rect 4356 -13880 5528 -13832
rect 5768 -13048 6940 -13000
rect 5768 -13112 6856 -13048
rect 6920 -13112 6940 -13048
rect 5768 -13128 6940 -13112
rect 5768 -13192 6856 -13128
rect 6920 -13192 6940 -13128
rect 5768 -13208 6940 -13192
rect 5768 -13272 6856 -13208
rect 6920 -13272 6940 -13208
rect 5768 -13288 6940 -13272
rect 5768 -13352 6856 -13288
rect 6920 -13352 6940 -13288
rect 5768 -13368 6940 -13352
rect 5768 -13432 6856 -13368
rect 6920 -13432 6940 -13368
rect 5768 -13448 6940 -13432
rect 5768 -13512 6856 -13448
rect 6920 -13512 6940 -13448
rect 5768 -13528 6940 -13512
rect 5768 -13592 6856 -13528
rect 6920 -13592 6940 -13528
rect 5768 -13608 6940 -13592
rect 5768 -13672 6856 -13608
rect 6920 -13672 6940 -13608
rect 5768 -13688 6940 -13672
rect 5768 -13752 6856 -13688
rect 6920 -13752 6940 -13688
rect 5768 -13768 6940 -13752
rect 5768 -13832 6856 -13768
rect 6920 -13832 6940 -13768
rect 5768 -13880 6940 -13832
rect 7180 -13048 8352 -13000
rect 7180 -13112 8268 -13048
rect 8332 -13112 8352 -13048
rect 7180 -13128 8352 -13112
rect 7180 -13192 8268 -13128
rect 8332 -13192 8352 -13128
rect 7180 -13208 8352 -13192
rect 7180 -13272 8268 -13208
rect 8332 -13272 8352 -13208
rect 7180 -13288 8352 -13272
rect 7180 -13352 8268 -13288
rect 8332 -13352 8352 -13288
rect 7180 -13368 8352 -13352
rect 7180 -13432 8268 -13368
rect 8332 -13432 8352 -13368
rect 7180 -13448 8352 -13432
rect 7180 -13512 8268 -13448
rect 8332 -13512 8352 -13448
rect 7180 -13528 8352 -13512
rect 7180 -13592 8268 -13528
rect 8332 -13592 8352 -13528
rect 7180 -13608 8352 -13592
rect 7180 -13672 8268 -13608
rect 8332 -13672 8352 -13608
rect 7180 -13688 8352 -13672
rect 7180 -13752 8268 -13688
rect 8332 -13752 8352 -13688
rect 7180 -13768 8352 -13752
rect 7180 -13832 8268 -13768
rect 8332 -13832 8352 -13768
rect 7180 -13880 8352 -13832
rect 8592 -13048 9764 -13000
rect 8592 -13112 9680 -13048
rect 9744 -13112 9764 -13048
rect 8592 -13128 9764 -13112
rect 8592 -13192 9680 -13128
rect 9744 -13192 9764 -13128
rect 8592 -13208 9764 -13192
rect 8592 -13272 9680 -13208
rect 9744 -13272 9764 -13208
rect 8592 -13288 9764 -13272
rect 8592 -13352 9680 -13288
rect 9744 -13352 9764 -13288
rect 8592 -13368 9764 -13352
rect 8592 -13432 9680 -13368
rect 9744 -13432 9764 -13368
rect 8592 -13448 9764 -13432
rect 8592 -13512 9680 -13448
rect 9744 -13512 9764 -13448
rect 8592 -13528 9764 -13512
rect 8592 -13592 9680 -13528
rect 9744 -13592 9764 -13528
rect 8592 -13608 9764 -13592
rect 8592 -13672 9680 -13608
rect 9744 -13672 9764 -13608
rect 8592 -13688 9764 -13672
rect 8592 -13752 9680 -13688
rect 9744 -13752 9764 -13688
rect 8592 -13768 9764 -13752
rect 8592 -13832 9680 -13768
rect 9744 -13832 9764 -13768
rect 8592 -13880 9764 -13832
rect 10004 -13048 11176 -13000
rect 10004 -13112 11092 -13048
rect 11156 -13112 11176 -13048
rect 10004 -13128 11176 -13112
rect 10004 -13192 11092 -13128
rect 11156 -13192 11176 -13128
rect 10004 -13208 11176 -13192
rect 10004 -13272 11092 -13208
rect 11156 -13272 11176 -13208
rect 10004 -13288 11176 -13272
rect 10004 -13352 11092 -13288
rect 11156 -13352 11176 -13288
rect 10004 -13368 11176 -13352
rect 10004 -13432 11092 -13368
rect 11156 -13432 11176 -13368
rect 10004 -13448 11176 -13432
rect 10004 -13512 11092 -13448
rect 11156 -13512 11176 -13448
rect 10004 -13528 11176 -13512
rect 10004 -13592 11092 -13528
rect 11156 -13592 11176 -13528
rect 10004 -13608 11176 -13592
rect 10004 -13672 11092 -13608
rect 11156 -13672 11176 -13608
rect 10004 -13688 11176 -13672
rect 10004 -13752 11092 -13688
rect 11156 -13752 11176 -13688
rect 10004 -13768 11176 -13752
rect 10004 -13832 11092 -13768
rect 11156 -13832 11176 -13768
rect 10004 -13880 11176 -13832
rect 11416 -13048 12588 -13000
rect 11416 -13112 12504 -13048
rect 12568 -13112 12588 -13048
rect 11416 -13128 12588 -13112
rect 11416 -13192 12504 -13128
rect 12568 -13192 12588 -13128
rect 11416 -13208 12588 -13192
rect 11416 -13272 12504 -13208
rect 12568 -13272 12588 -13208
rect 11416 -13288 12588 -13272
rect 11416 -13352 12504 -13288
rect 12568 -13352 12588 -13288
rect 11416 -13368 12588 -13352
rect 11416 -13432 12504 -13368
rect 12568 -13432 12588 -13368
rect 11416 -13448 12588 -13432
rect 11416 -13512 12504 -13448
rect 12568 -13512 12588 -13448
rect 11416 -13528 12588 -13512
rect 11416 -13592 12504 -13528
rect 12568 -13592 12588 -13528
rect 11416 -13608 12588 -13592
rect 11416 -13672 12504 -13608
rect 12568 -13672 12588 -13608
rect 11416 -13688 12588 -13672
rect 11416 -13752 12504 -13688
rect 12568 -13752 12588 -13688
rect 11416 -13768 12588 -13752
rect 11416 -13832 12504 -13768
rect 12568 -13832 12588 -13768
rect 11416 -13880 12588 -13832
rect 12828 -13048 14000 -13000
rect 12828 -13112 13916 -13048
rect 13980 -13112 14000 -13048
rect 12828 -13128 14000 -13112
rect 12828 -13192 13916 -13128
rect 13980 -13192 14000 -13128
rect 12828 -13208 14000 -13192
rect 12828 -13272 13916 -13208
rect 13980 -13272 14000 -13208
rect 12828 -13288 14000 -13272
rect 12828 -13352 13916 -13288
rect 13980 -13352 14000 -13288
rect 12828 -13368 14000 -13352
rect 12828 -13432 13916 -13368
rect 13980 -13432 14000 -13368
rect 12828 -13448 14000 -13432
rect 12828 -13512 13916 -13448
rect 13980 -13512 14000 -13448
rect 12828 -13528 14000 -13512
rect 12828 -13592 13916 -13528
rect 13980 -13592 14000 -13528
rect 12828 -13608 14000 -13592
rect 12828 -13672 13916 -13608
rect 13980 -13672 14000 -13608
rect 12828 -13688 14000 -13672
rect 12828 -13752 13916 -13688
rect 13980 -13752 14000 -13688
rect 12828 -13768 14000 -13752
rect 12828 -13832 13916 -13768
rect 13980 -13832 14000 -13768
rect 12828 -13880 14000 -13832
rect 14240 -13048 15412 -13000
rect 14240 -13112 15328 -13048
rect 15392 -13112 15412 -13048
rect 14240 -13128 15412 -13112
rect 14240 -13192 15328 -13128
rect 15392 -13192 15412 -13128
rect 14240 -13208 15412 -13192
rect 14240 -13272 15328 -13208
rect 15392 -13272 15412 -13208
rect 14240 -13288 15412 -13272
rect 14240 -13352 15328 -13288
rect 15392 -13352 15412 -13288
rect 14240 -13368 15412 -13352
rect 14240 -13432 15328 -13368
rect 15392 -13432 15412 -13368
rect 14240 -13448 15412 -13432
rect 14240 -13512 15328 -13448
rect 15392 -13512 15412 -13448
rect 14240 -13528 15412 -13512
rect 14240 -13592 15328 -13528
rect 15392 -13592 15412 -13528
rect 14240 -13608 15412 -13592
rect 14240 -13672 15328 -13608
rect 15392 -13672 15412 -13608
rect 14240 -13688 15412 -13672
rect 14240 -13752 15328 -13688
rect 15392 -13752 15412 -13688
rect 14240 -13768 15412 -13752
rect 14240 -13832 15328 -13768
rect 15392 -13832 15412 -13768
rect 14240 -13880 15412 -13832
rect 15652 -13048 16824 -13000
rect 15652 -13112 16740 -13048
rect 16804 -13112 16824 -13048
rect 15652 -13128 16824 -13112
rect 15652 -13192 16740 -13128
rect 16804 -13192 16824 -13128
rect 15652 -13208 16824 -13192
rect 15652 -13272 16740 -13208
rect 16804 -13272 16824 -13208
rect 15652 -13288 16824 -13272
rect 15652 -13352 16740 -13288
rect 16804 -13352 16824 -13288
rect 15652 -13368 16824 -13352
rect 15652 -13432 16740 -13368
rect 16804 -13432 16824 -13368
rect 15652 -13448 16824 -13432
rect 15652 -13512 16740 -13448
rect 16804 -13512 16824 -13448
rect 15652 -13528 16824 -13512
rect 15652 -13592 16740 -13528
rect 16804 -13592 16824 -13528
rect 15652 -13608 16824 -13592
rect 15652 -13672 16740 -13608
rect 16804 -13672 16824 -13608
rect 15652 -13688 16824 -13672
rect 15652 -13752 16740 -13688
rect 16804 -13752 16824 -13688
rect 15652 -13768 16824 -13752
rect 15652 -13832 16740 -13768
rect 16804 -13832 16824 -13768
rect 15652 -13880 16824 -13832
rect 17064 -13048 18236 -13000
rect 17064 -13112 18152 -13048
rect 18216 -13112 18236 -13048
rect 17064 -13128 18236 -13112
rect 17064 -13192 18152 -13128
rect 18216 -13192 18236 -13128
rect 17064 -13208 18236 -13192
rect 17064 -13272 18152 -13208
rect 18216 -13272 18236 -13208
rect 17064 -13288 18236 -13272
rect 17064 -13352 18152 -13288
rect 18216 -13352 18236 -13288
rect 17064 -13368 18236 -13352
rect 17064 -13432 18152 -13368
rect 18216 -13432 18236 -13368
rect 17064 -13448 18236 -13432
rect 17064 -13512 18152 -13448
rect 18216 -13512 18236 -13448
rect 17064 -13528 18236 -13512
rect 17064 -13592 18152 -13528
rect 18216 -13592 18236 -13528
rect 17064 -13608 18236 -13592
rect 17064 -13672 18152 -13608
rect 18216 -13672 18236 -13608
rect 17064 -13688 18236 -13672
rect 17064 -13752 18152 -13688
rect 18216 -13752 18236 -13688
rect 17064 -13768 18236 -13752
rect 17064 -13832 18152 -13768
rect 18216 -13832 18236 -13768
rect 17064 -13880 18236 -13832
rect 18476 -13048 19648 -13000
rect 18476 -13112 19564 -13048
rect 19628 -13112 19648 -13048
rect 18476 -13128 19648 -13112
rect 18476 -13192 19564 -13128
rect 19628 -13192 19648 -13128
rect 18476 -13208 19648 -13192
rect 18476 -13272 19564 -13208
rect 19628 -13272 19648 -13208
rect 18476 -13288 19648 -13272
rect 18476 -13352 19564 -13288
rect 19628 -13352 19648 -13288
rect 18476 -13368 19648 -13352
rect 18476 -13432 19564 -13368
rect 19628 -13432 19648 -13368
rect 18476 -13448 19648 -13432
rect 18476 -13512 19564 -13448
rect 19628 -13512 19648 -13448
rect 18476 -13528 19648 -13512
rect 18476 -13592 19564 -13528
rect 19628 -13592 19648 -13528
rect 18476 -13608 19648 -13592
rect 18476 -13672 19564 -13608
rect 19628 -13672 19648 -13608
rect 18476 -13688 19648 -13672
rect 18476 -13752 19564 -13688
rect 19628 -13752 19648 -13688
rect 18476 -13768 19648 -13752
rect 18476 -13832 19564 -13768
rect 19628 -13832 19648 -13768
rect 18476 -13880 19648 -13832
rect 19888 -13048 21060 -13000
rect 19888 -13112 20976 -13048
rect 21040 -13112 21060 -13048
rect 19888 -13128 21060 -13112
rect 19888 -13192 20976 -13128
rect 21040 -13192 21060 -13128
rect 19888 -13208 21060 -13192
rect 19888 -13272 20976 -13208
rect 21040 -13272 21060 -13208
rect 19888 -13288 21060 -13272
rect 19888 -13352 20976 -13288
rect 21040 -13352 21060 -13288
rect 19888 -13368 21060 -13352
rect 19888 -13432 20976 -13368
rect 21040 -13432 21060 -13368
rect 19888 -13448 21060 -13432
rect 19888 -13512 20976 -13448
rect 21040 -13512 21060 -13448
rect 19888 -13528 21060 -13512
rect 19888 -13592 20976 -13528
rect 21040 -13592 21060 -13528
rect 19888 -13608 21060 -13592
rect 19888 -13672 20976 -13608
rect 21040 -13672 21060 -13608
rect 19888 -13688 21060 -13672
rect 19888 -13752 20976 -13688
rect 21040 -13752 21060 -13688
rect 19888 -13768 21060 -13752
rect 19888 -13832 20976 -13768
rect 21040 -13832 21060 -13768
rect 19888 -13880 21060 -13832
rect 21300 -13048 22472 -13000
rect 21300 -13112 22388 -13048
rect 22452 -13112 22472 -13048
rect 21300 -13128 22472 -13112
rect 21300 -13192 22388 -13128
rect 22452 -13192 22472 -13128
rect 21300 -13208 22472 -13192
rect 21300 -13272 22388 -13208
rect 22452 -13272 22472 -13208
rect 21300 -13288 22472 -13272
rect 21300 -13352 22388 -13288
rect 22452 -13352 22472 -13288
rect 21300 -13368 22472 -13352
rect 21300 -13432 22388 -13368
rect 22452 -13432 22472 -13368
rect 21300 -13448 22472 -13432
rect 21300 -13512 22388 -13448
rect 22452 -13512 22472 -13448
rect 21300 -13528 22472 -13512
rect 21300 -13592 22388 -13528
rect 22452 -13592 22472 -13528
rect 21300 -13608 22472 -13592
rect 21300 -13672 22388 -13608
rect 22452 -13672 22472 -13608
rect 21300 -13688 22472 -13672
rect 21300 -13752 22388 -13688
rect 22452 -13752 22472 -13688
rect 21300 -13768 22472 -13752
rect 21300 -13832 22388 -13768
rect 22452 -13832 22472 -13768
rect 21300 -13880 22472 -13832
rect 22712 -13048 23884 -13000
rect 22712 -13112 23800 -13048
rect 23864 -13112 23884 -13048
rect 22712 -13128 23884 -13112
rect 22712 -13192 23800 -13128
rect 23864 -13192 23884 -13128
rect 22712 -13208 23884 -13192
rect 22712 -13272 23800 -13208
rect 23864 -13272 23884 -13208
rect 22712 -13288 23884 -13272
rect 22712 -13352 23800 -13288
rect 23864 -13352 23884 -13288
rect 22712 -13368 23884 -13352
rect 22712 -13432 23800 -13368
rect 23864 -13432 23884 -13368
rect 22712 -13448 23884 -13432
rect 22712 -13512 23800 -13448
rect 23864 -13512 23884 -13448
rect 22712 -13528 23884 -13512
rect 22712 -13592 23800 -13528
rect 23864 -13592 23884 -13528
rect 22712 -13608 23884 -13592
rect 22712 -13672 23800 -13608
rect 23864 -13672 23884 -13608
rect 22712 -13688 23884 -13672
rect 22712 -13752 23800 -13688
rect 23864 -13752 23884 -13688
rect 22712 -13768 23884 -13752
rect 22712 -13832 23800 -13768
rect 23864 -13832 23884 -13768
rect 22712 -13880 23884 -13832
rect -23884 -14168 -22712 -14120
rect -23884 -14232 -22796 -14168
rect -22732 -14232 -22712 -14168
rect -23884 -14248 -22712 -14232
rect -23884 -14312 -22796 -14248
rect -22732 -14312 -22712 -14248
rect -23884 -14328 -22712 -14312
rect -23884 -14392 -22796 -14328
rect -22732 -14392 -22712 -14328
rect -23884 -14408 -22712 -14392
rect -23884 -14472 -22796 -14408
rect -22732 -14472 -22712 -14408
rect -23884 -14488 -22712 -14472
rect -23884 -14552 -22796 -14488
rect -22732 -14552 -22712 -14488
rect -23884 -14568 -22712 -14552
rect -23884 -14632 -22796 -14568
rect -22732 -14632 -22712 -14568
rect -23884 -14648 -22712 -14632
rect -23884 -14712 -22796 -14648
rect -22732 -14712 -22712 -14648
rect -23884 -14728 -22712 -14712
rect -23884 -14792 -22796 -14728
rect -22732 -14792 -22712 -14728
rect -23884 -14808 -22712 -14792
rect -23884 -14872 -22796 -14808
rect -22732 -14872 -22712 -14808
rect -23884 -14888 -22712 -14872
rect -23884 -14952 -22796 -14888
rect -22732 -14952 -22712 -14888
rect -23884 -15000 -22712 -14952
rect -22472 -14168 -21300 -14120
rect -22472 -14232 -21384 -14168
rect -21320 -14232 -21300 -14168
rect -22472 -14248 -21300 -14232
rect -22472 -14312 -21384 -14248
rect -21320 -14312 -21300 -14248
rect -22472 -14328 -21300 -14312
rect -22472 -14392 -21384 -14328
rect -21320 -14392 -21300 -14328
rect -22472 -14408 -21300 -14392
rect -22472 -14472 -21384 -14408
rect -21320 -14472 -21300 -14408
rect -22472 -14488 -21300 -14472
rect -22472 -14552 -21384 -14488
rect -21320 -14552 -21300 -14488
rect -22472 -14568 -21300 -14552
rect -22472 -14632 -21384 -14568
rect -21320 -14632 -21300 -14568
rect -22472 -14648 -21300 -14632
rect -22472 -14712 -21384 -14648
rect -21320 -14712 -21300 -14648
rect -22472 -14728 -21300 -14712
rect -22472 -14792 -21384 -14728
rect -21320 -14792 -21300 -14728
rect -22472 -14808 -21300 -14792
rect -22472 -14872 -21384 -14808
rect -21320 -14872 -21300 -14808
rect -22472 -14888 -21300 -14872
rect -22472 -14952 -21384 -14888
rect -21320 -14952 -21300 -14888
rect -22472 -15000 -21300 -14952
rect -21060 -14168 -19888 -14120
rect -21060 -14232 -19972 -14168
rect -19908 -14232 -19888 -14168
rect -21060 -14248 -19888 -14232
rect -21060 -14312 -19972 -14248
rect -19908 -14312 -19888 -14248
rect -21060 -14328 -19888 -14312
rect -21060 -14392 -19972 -14328
rect -19908 -14392 -19888 -14328
rect -21060 -14408 -19888 -14392
rect -21060 -14472 -19972 -14408
rect -19908 -14472 -19888 -14408
rect -21060 -14488 -19888 -14472
rect -21060 -14552 -19972 -14488
rect -19908 -14552 -19888 -14488
rect -21060 -14568 -19888 -14552
rect -21060 -14632 -19972 -14568
rect -19908 -14632 -19888 -14568
rect -21060 -14648 -19888 -14632
rect -21060 -14712 -19972 -14648
rect -19908 -14712 -19888 -14648
rect -21060 -14728 -19888 -14712
rect -21060 -14792 -19972 -14728
rect -19908 -14792 -19888 -14728
rect -21060 -14808 -19888 -14792
rect -21060 -14872 -19972 -14808
rect -19908 -14872 -19888 -14808
rect -21060 -14888 -19888 -14872
rect -21060 -14952 -19972 -14888
rect -19908 -14952 -19888 -14888
rect -21060 -15000 -19888 -14952
rect -19648 -14168 -18476 -14120
rect -19648 -14232 -18560 -14168
rect -18496 -14232 -18476 -14168
rect -19648 -14248 -18476 -14232
rect -19648 -14312 -18560 -14248
rect -18496 -14312 -18476 -14248
rect -19648 -14328 -18476 -14312
rect -19648 -14392 -18560 -14328
rect -18496 -14392 -18476 -14328
rect -19648 -14408 -18476 -14392
rect -19648 -14472 -18560 -14408
rect -18496 -14472 -18476 -14408
rect -19648 -14488 -18476 -14472
rect -19648 -14552 -18560 -14488
rect -18496 -14552 -18476 -14488
rect -19648 -14568 -18476 -14552
rect -19648 -14632 -18560 -14568
rect -18496 -14632 -18476 -14568
rect -19648 -14648 -18476 -14632
rect -19648 -14712 -18560 -14648
rect -18496 -14712 -18476 -14648
rect -19648 -14728 -18476 -14712
rect -19648 -14792 -18560 -14728
rect -18496 -14792 -18476 -14728
rect -19648 -14808 -18476 -14792
rect -19648 -14872 -18560 -14808
rect -18496 -14872 -18476 -14808
rect -19648 -14888 -18476 -14872
rect -19648 -14952 -18560 -14888
rect -18496 -14952 -18476 -14888
rect -19648 -15000 -18476 -14952
rect -18236 -14168 -17064 -14120
rect -18236 -14232 -17148 -14168
rect -17084 -14232 -17064 -14168
rect -18236 -14248 -17064 -14232
rect -18236 -14312 -17148 -14248
rect -17084 -14312 -17064 -14248
rect -18236 -14328 -17064 -14312
rect -18236 -14392 -17148 -14328
rect -17084 -14392 -17064 -14328
rect -18236 -14408 -17064 -14392
rect -18236 -14472 -17148 -14408
rect -17084 -14472 -17064 -14408
rect -18236 -14488 -17064 -14472
rect -18236 -14552 -17148 -14488
rect -17084 -14552 -17064 -14488
rect -18236 -14568 -17064 -14552
rect -18236 -14632 -17148 -14568
rect -17084 -14632 -17064 -14568
rect -18236 -14648 -17064 -14632
rect -18236 -14712 -17148 -14648
rect -17084 -14712 -17064 -14648
rect -18236 -14728 -17064 -14712
rect -18236 -14792 -17148 -14728
rect -17084 -14792 -17064 -14728
rect -18236 -14808 -17064 -14792
rect -18236 -14872 -17148 -14808
rect -17084 -14872 -17064 -14808
rect -18236 -14888 -17064 -14872
rect -18236 -14952 -17148 -14888
rect -17084 -14952 -17064 -14888
rect -18236 -15000 -17064 -14952
rect -16824 -14168 -15652 -14120
rect -16824 -14232 -15736 -14168
rect -15672 -14232 -15652 -14168
rect -16824 -14248 -15652 -14232
rect -16824 -14312 -15736 -14248
rect -15672 -14312 -15652 -14248
rect -16824 -14328 -15652 -14312
rect -16824 -14392 -15736 -14328
rect -15672 -14392 -15652 -14328
rect -16824 -14408 -15652 -14392
rect -16824 -14472 -15736 -14408
rect -15672 -14472 -15652 -14408
rect -16824 -14488 -15652 -14472
rect -16824 -14552 -15736 -14488
rect -15672 -14552 -15652 -14488
rect -16824 -14568 -15652 -14552
rect -16824 -14632 -15736 -14568
rect -15672 -14632 -15652 -14568
rect -16824 -14648 -15652 -14632
rect -16824 -14712 -15736 -14648
rect -15672 -14712 -15652 -14648
rect -16824 -14728 -15652 -14712
rect -16824 -14792 -15736 -14728
rect -15672 -14792 -15652 -14728
rect -16824 -14808 -15652 -14792
rect -16824 -14872 -15736 -14808
rect -15672 -14872 -15652 -14808
rect -16824 -14888 -15652 -14872
rect -16824 -14952 -15736 -14888
rect -15672 -14952 -15652 -14888
rect -16824 -15000 -15652 -14952
rect -15412 -14168 -14240 -14120
rect -15412 -14232 -14324 -14168
rect -14260 -14232 -14240 -14168
rect -15412 -14248 -14240 -14232
rect -15412 -14312 -14324 -14248
rect -14260 -14312 -14240 -14248
rect -15412 -14328 -14240 -14312
rect -15412 -14392 -14324 -14328
rect -14260 -14392 -14240 -14328
rect -15412 -14408 -14240 -14392
rect -15412 -14472 -14324 -14408
rect -14260 -14472 -14240 -14408
rect -15412 -14488 -14240 -14472
rect -15412 -14552 -14324 -14488
rect -14260 -14552 -14240 -14488
rect -15412 -14568 -14240 -14552
rect -15412 -14632 -14324 -14568
rect -14260 -14632 -14240 -14568
rect -15412 -14648 -14240 -14632
rect -15412 -14712 -14324 -14648
rect -14260 -14712 -14240 -14648
rect -15412 -14728 -14240 -14712
rect -15412 -14792 -14324 -14728
rect -14260 -14792 -14240 -14728
rect -15412 -14808 -14240 -14792
rect -15412 -14872 -14324 -14808
rect -14260 -14872 -14240 -14808
rect -15412 -14888 -14240 -14872
rect -15412 -14952 -14324 -14888
rect -14260 -14952 -14240 -14888
rect -15412 -15000 -14240 -14952
rect -14000 -14168 -12828 -14120
rect -14000 -14232 -12912 -14168
rect -12848 -14232 -12828 -14168
rect -14000 -14248 -12828 -14232
rect -14000 -14312 -12912 -14248
rect -12848 -14312 -12828 -14248
rect -14000 -14328 -12828 -14312
rect -14000 -14392 -12912 -14328
rect -12848 -14392 -12828 -14328
rect -14000 -14408 -12828 -14392
rect -14000 -14472 -12912 -14408
rect -12848 -14472 -12828 -14408
rect -14000 -14488 -12828 -14472
rect -14000 -14552 -12912 -14488
rect -12848 -14552 -12828 -14488
rect -14000 -14568 -12828 -14552
rect -14000 -14632 -12912 -14568
rect -12848 -14632 -12828 -14568
rect -14000 -14648 -12828 -14632
rect -14000 -14712 -12912 -14648
rect -12848 -14712 -12828 -14648
rect -14000 -14728 -12828 -14712
rect -14000 -14792 -12912 -14728
rect -12848 -14792 -12828 -14728
rect -14000 -14808 -12828 -14792
rect -14000 -14872 -12912 -14808
rect -12848 -14872 -12828 -14808
rect -14000 -14888 -12828 -14872
rect -14000 -14952 -12912 -14888
rect -12848 -14952 -12828 -14888
rect -14000 -15000 -12828 -14952
rect -12588 -14168 -11416 -14120
rect -12588 -14232 -11500 -14168
rect -11436 -14232 -11416 -14168
rect -12588 -14248 -11416 -14232
rect -12588 -14312 -11500 -14248
rect -11436 -14312 -11416 -14248
rect -12588 -14328 -11416 -14312
rect -12588 -14392 -11500 -14328
rect -11436 -14392 -11416 -14328
rect -12588 -14408 -11416 -14392
rect -12588 -14472 -11500 -14408
rect -11436 -14472 -11416 -14408
rect -12588 -14488 -11416 -14472
rect -12588 -14552 -11500 -14488
rect -11436 -14552 -11416 -14488
rect -12588 -14568 -11416 -14552
rect -12588 -14632 -11500 -14568
rect -11436 -14632 -11416 -14568
rect -12588 -14648 -11416 -14632
rect -12588 -14712 -11500 -14648
rect -11436 -14712 -11416 -14648
rect -12588 -14728 -11416 -14712
rect -12588 -14792 -11500 -14728
rect -11436 -14792 -11416 -14728
rect -12588 -14808 -11416 -14792
rect -12588 -14872 -11500 -14808
rect -11436 -14872 -11416 -14808
rect -12588 -14888 -11416 -14872
rect -12588 -14952 -11500 -14888
rect -11436 -14952 -11416 -14888
rect -12588 -15000 -11416 -14952
rect -11176 -14168 -10004 -14120
rect -11176 -14232 -10088 -14168
rect -10024 -14232 -10004 -14168
rect -11176 -14248 -10004 -14232
rect -11176 -14312 -10088 -14248
rect -10024 -14312 -10004 -14248
rect -11176 -14328 -10004 -14312
rect -11176 -14392 -10088 -14328
rect -10024 -14392 -10004 -14328
rect -11176 -14408 -10004 -14392
rect -11176 -14472 -10088 -14408
rect -10024 -14472 -10004 -14408
rect -11176 -14488 -10004 -14472
rect -11176 -14552 -10088 -14488
rect -10024 -14552 -10004 -14488
rect -11176 -14568 -10004 -14552
rect -11176 -14632 -10088 -14568
rect -10024 -14632 -10004 -14568
rect -11176 -14648 -10004 -14632
rect -11176 -14712 -10088 -14648
rect -10024 -14712 -10004 -14648
rect -11176 -14728 -10004 -14712
rect -11176 -14792 -10088 -14728
rect -10024 -14792 -10004 -14728
rect -11176 -14808 -10004 -14792
rect -11176 -14872 -10088 -14808
rect -10024 -14872 -10004 -14808
rect -11176 -14888 -10004 -14872
rect -11176 -14952 -10088 -14888
rect -10024 -14952 -10004 -14888
rect -11176 -15000 -10004 -14952
rect -9764 -14168 -8592 -14120
rect -9764 -14232 -8676 -14168
rect -8612 -14232 -8592 -14168
rect -9764 -14248 -8592 -14232
rect -9764 -14312 -8676 -14248
rect -8612 -14312 -8592 -14248
rect -9764 -14328 -8592 -14312
rect -9764 -14392 -8676 -14328
rect -8612 -14392 -8592 -14328
rect -9764 -14408 -8592 -14392
rect -9764 -14472 -8676 -14408
rect -8612 -14472 -8592 -14408
rect -9764 -14488 -8592 -14472
rect -9764 -14552 -8676 -14488
rect -8612 -14552 -8592 -14488
rect -9764 -14568 -8592 -14552
rect -9764 -14632 -8676 -14568
rect -8612 -14632 -8592 -14568
rect -9764 -14648 -8592 -14632
rect -9764 -14712 -8676 -14648
rect -8612 -14712 -8592 -14648
rect -9764 -14728 -8592 -14712
rect -9764 -14792 -8676 -14728
rect -8612 -14792 -8592 -14728
rect -9764 -14808 -8592 -14792
rect -9764 -14872 -8676 -14808
rect -8612 -14872 -8592 -14808
rect -9764 -14888 -8592 -14872
rect -9764 -14952 -8676 -14888
rect -8612 -14952 -8592 -14888
rect -9764 -15000 -8592 -14952
rect -8352 -14168 -7180 -14120
rect -8352 -14232 -7264 -14168
rect -7200 -14232 -7180 -14168
rect -8352 -14248 -7180 -14232
rect -8352 -14312 -7264 -14248
rect -7200 -14312 -7180 -14248
rect -8352 -14328 -7180 -14312
rect -8352 -14392 -7264 -14328
rect -7200 -14392 -7180 -14328
rect -8352 -14408 -7180 -14392
rect -8352 -14472 -7264 -14408
rect -7200 -14472 -7180 -14408
rect -8352 -14488 -7180 -14472
rect -8352 -14552 -7264 -14488
rect -7200 -14552 -7180 -14488
rect -8352 -14568 -7180 -14552
rect -8352 -14632 -7264 -14568
rect -7200 -14632 -7180 -14568
rect -8352 -14648 -7180 -14632
rect -8352 -14712 -7264 -14648
rect -7200 -14712 -7180 -14648
rect -8352 -14728 -7180 -14712
rect -8352 -14792 -7264 -14728
rect -7200 -14792 -7180 -14728
rect -8352 -14808 -7180 -14792
rect -8352 -14872 -7264 -14808
rect -7200 -14872 -7180 -14808
rect -8352 -14888 -7180 -14872
rect -8352 -14952 -7264 -14888
rect -7200 -14952 -7180 -14888
rect -8352 -15000 -7180 -14952
rect -6940 -14168 -5768 -14120
rect -6940 -14232 -5852 -14168
rect -5788 -14232 -5768 -14168
rect -6940 -14248 -5768 -14232
rect -6940 -14312 -5852 -14248
rect -5788 -14312 -5768 -14248
rect -6940 -14328 -5768 -14312
rect -6940 -14392 -5852 -14328
rect -5788 -14392 -5768 -14328
rect -6940 -14408 -5768 -14392
rect -6940 -14472 -5852 -14408
rect -5788 -14472 -5768 -14408
rect -6940 -14488 -5768 -14472
rect -6940 -14552 -5852 -14488
rect -5788 -14552 -5768 -14488
rect -6940 -14568 -5768 -14552
rect -6940 -14632 -5852 -14568
rect -5788 -14632 -5768 -14568
rect -6940 -14648 -5768 -14632
rect -6940 -14712 -5852 -14648
rect -5788 -14712 -5768 -14648
rect -6940 -14728 -5768 -14712
rect -6940 -14792 -5852 -14728
rect -5788 -14792 -5768 -14728
rect -6940 -14808 -5768 -14792
rect -6940 -14872 -5852 -14808
rect -5788 -14872 -5768 -14808
rect -6940 -14888 -5768 -14872
rect -6940 -14952 -5852 -14888
rect -5788 -14952 -5768 -14888
rect -6940 -15000 -5768 -14952
rect -5528 -14168 -4356 -14120
rect -5528 -14232 -4440 -14168
rect -4376 -14232 -4356 -14168
rect -5528 -14248 -4356 -14232
rect -5528 -14312 -4440 -14248
rect -4376 -14312 -4356 -14248
rect -5528 -14328 -4356 -14312
rect -5528 -14392 -4440 -14328
rect -4376 -14392 -4356 -14328
rect -5528 -14408 -4356 -14392
rect -5528 -14472 -4440 -14408
rect -4376 -14472 -4356 -14408
rect -5528 -14488 -4356 -14472
rect -5528 -14552 -4440 -14488
rect -4376 -14552 -4356 -14488
rect -5528 -14568 -4356 -14552
rect -5528 -14632 -4440 -14568
rect -4376 -14632 -4356 -14568
rect -5528 -14648 -4356 -14632
rect -5528 -14712 -4440 -14648
rect -4376 -14712 -4356 -14648
rect -5528 -14728 -4356 -14712
rect -5528 -14792 -4440 -14728
rect -4376 -14792 -4356 -14728
rect -5528 -14808 -4356 -14792
rect -5528 -14872 -4440 -14808
rect -4376 -14872 -4356 -14808
rect -5528 -14888 -4356 -14872
rect -5528 -14952 -4440 -14888
rect -4376 -14952 -4356 -14888
rect -5528 -15000 -4356 -14952
rect -4116 -14168 -2944 -14120
rect -4116 -14232 -3028 -14168
rect -2964 -14232 -2944 -14168
rect -4116 -14248 -2944 -14232
rect -4116 -14312 -3028 -14248
rect -2964 -14312 -2944 -14248
rect -4116 -14328 -2944 -14312
rect -4116 -14392 -3028 -14328
rect -2964 -14392 -2944 -14328
rect -4116 -14408 -2944 -14392
rect -4116 -14472 -3028 -14408
rect -2964 -14472 -2944 -14408
rect -4116 -14488 -2944 -14472
rect -4116 -14552 -3028 -14488
rect -2964 -14552 -2944 -14488
rect -4116 -14568 -2944 -14552
rect -4116 -14632 -3028 -14568
rect -2964 -14632 -2944 -14568
rect -4116 -14648 -2944 -14632
rect -4116 -14712 -3028 -14648
rect -2964 -14712 -2944 -14648
rect -4116 -14728 -2944 -14712
rect -4116 -14792 -3028 -14728
rect -2964 -14792 -2944 -14728
rect -4116 -14808 -2944 -14792
rect -4116 -14872 -3028 -14808
rect -2964 -14872 -2944 -14808
rect -4116 -14888 -2944 -14872
rect -4116 -14952 -3028 -14888
rect -2964 -14952 -2944 -14888
rect -4116 -15000 -2944 -14952
rect -2704 -14168 -1532 -14120
rect -2704 -14232 -1616 -14168
rect -1552 -14232 -1532 -14168
rect -2704 -14248 -1532 -14232
rect -2704 -14312 -1616 -14248
rect -1552 -14312 -1532 -14248
rect -2704 -14328 -1532 -14312
rect -2704 -14392 -1616 -14328
rect -1552 -14392 -1532 -14328
rect -2704 -14408 -1532 -14392
rect -2704 -14472 -1616 -14408
rect -1552 -14472 -1532 -14408
rect -2704 -14488 -1532 -14472
rect -2704 -14552 -1616 -14488
rect -1552 -14552 -1532 -14488
rect -2704 -14568 -1532 -14552
rect -2704 -14632 -1616 -14568
rect -1552 -14632 -1532 -14568
rect -2704 -14648 -1532 -14632
rect -2704 -14712 -1616 -14648
rect -1552 -14712 -1532 -14648
rect -2704 -14728 -1532 -14712
rect -2704 -14792 -1616 -14728
rect -1552 -14792 -1532 -14728
rect -2704 -14808 -1532 -14792
rect -2704 -14872 -1616 -14808
rect -1552 -14872 -1532 -14808
rect -2704 -14888 -1532 -14872
rect -2704 -14952 -1616 -14888
rect -1552 -14952 -1532 -14888
rect -2704 -15000 -1532 -14952
rect -1292 -14168 -120 -14120
rect -1292 -14232 -204 -14168
rect -140 -14232 -120 -14168
rect -1292 -14248 -120 -14232
rect -1292 -14312 -204 -14248
rect -140 -14312 -120 -14248
rect -1292 -14328 -120 -14312
rect -1292 -14392 -204 -14328
rect -140 -14392 -120 -14328
rect -1292 -14408 -120 -14392
rect -1292 -14472 -204 -14408
rect -140 -14472 -120 -14408
rect -1292 -14488 -120 -14472
rect -1292 -14552 -204 -14488
rect -140 -14552 -120 -14488
rect -1292 -14568 -120 -14552
rect -1292 -14632 -204 -14568
rect -140 -14632 -120 -14568
rect -1292 -14648 -120 -14632
rect -1292 -14712 -204 -14648
rect -140 -14712 -120 -14648
rect -1292 -14728 -120 -14712
rect -1292 -14792 -204 -14728
rect -140 -14792 -120 -14728
rect -1292 -14808 -120 -14792
rect -1292 -14872 -204 -14808
rect -140 -14872 -120 -14808
rect -1292 -14888 -120 -14872
rect -1292 -14952 -204 -14888
rect -140 -14952 -120 -14888
rect -1292 -15000 -120 -14952
rect 120 -14168 1292 -14120
rect 120 -14232 1208 -14168
rect 1272 -14232 1292 -14168
rect 120 -14248 1292 -14232
rect 120 -14312 1208 -14248
rect 1272 -14312 1292 -14248
rect 120 -14328 1292 -14312
rect 120 -14392 1208 -14328
rect 1272 -14392 1292 -14328
rect 120 -14408 1292 -14392
rect 120 -14472 1208 -14408
rect 1272 -14472 1292 -14408
rect 120 -14488 1292 -14472
rect 120 -14552 1208 -14488
rect 1272 -14552 1292 -14488
rect 120 -14568 1292 -14552
rect 120 -14632 1208 -14568
rect 1272 -14632 1292 -14568
rect 120 -14648 1292 -14632
rect 120 -14712 1208 -14648
rect 1272 -14712 1292 -14648
rect 120 -14728 1292 -14712
rect 120 -14792 1208 -14728
rect 1272 -14792 1292 -14728
rect 120 -14808 1292 -14792
rect 120 -14872 1208 -14808
rect 1272 -14872 1292 -14808
rect 120 -14888 1292 -14872
rect 120 -14952 1208 -14888
rect 1272 -14952 1292 -14888
rect 120 -15000 1292 -14952
rect 1532 -14168 2704 -14120
rect 1532 -14232 2620 -14168
rect 2684 -14232 2704 -14168
rect 1532 -14248 2704 -14232
rect 1532 -14312 2620 -14248
rect 2684 -14312 2704 -14248
rect 1532 -14328 2704 -14312
rect 1532 -14392 2620 -14328
rect 2684 -14392 2704 -14328
rect 1532 -14408 2704 -14392
rect 1532 -14472 2620 -14408
rect 2684 -14472 2704 -14408
rect 1532 -14488 2704 -14472
rect 1532 -14552 2620 -14488
rect 2684 -14552 2704 -14488
rect 1532 -14568 2704 -14552
rect 1532 -14632 2620 -14568
rect 2684 -14632 2704 -14568
rect 1532 -14648 2704 -14632
rect 1532 -14712 2620 -14648
rect 2684 -14712 2704 -14648
rect 1532 -14728 2704 -14712
rect 1532 -14792 2620 -14728
rect 2684 -14792 2704 -14728
rect 1532 -14808 2704 -14792
rect 1532 -14872 2620 -14808
rect 2684 -14872 2704 -14808
rect 1532 -14888 2704 -14872
rect 1532 -14952 2620 -14888
rect 2684 -14952 2704 -14888
rect 1532 -15000 2704 -14952
rect 2944 -14168 4116 -14120
rect 2944 -14232 4032 -14168
rect 4096 -14232 4116 -14168
rect 2944 -14248 4116 -14232
rect 2944 -14312 4032 -14248
rect 4096 -14312 4116 -14248
rect 2944 -14328 4116 -14312
rect 2944 -14392 4032 -14328
rect 4096 -14392 4116 -14328
rect 2944 -14408 4116 -14392
rect 2944 -14472 4032 -14408
rect 4096 -14472 4116 -14408
rect 2944 -14488 4116 -14472
rect 2944 -14552 4032 -14488
rect 4096 -14552 4116 -14488
rect 2944 -14568 4116 -14552
rect 2944 -14632 4032 -14568
rect 4096 -14632 4116 -14568
rect 2944 -14648 4116 -14632
rect 2944 -14712 4032 -14648
rect 4096 -14712 4116 -14648
rect 2944 -14728 4116 -14712
rect 2944 -14792 4032 -14728
rect 4096 -14792 4116 -14728
rect 2944 -14808 4116 -14792
rect 2944 -14872 4032 -14808
rect 4096 -14872 4116 -14808
rect 2944 -14888 4116 -14872
rect 2944 -14952 4032 -14888
rect 4096 -14952 4116 -14888
rect 2944 -15000 4116 -14952
rect 4356 -14168 5528 -14120
rect 4356 -14232 5444 -14168
rect 5508 -14232 5528 -14168
rect 4356 -14248 5528 -14232
rect 4356 -14312 5444 -14248
rect 5508 -14312 5528 -14248
rect 4356 -14328 5528 -14312
rect 4356 -14392 5444 -14328
rect 5508 -14392 5528 -14328
rect 4356 -14408 5528 -14392
rect 4356 -14472 5444 -14408
rect 5508 -14472 5528 -14408
rect 4356 -14488 5528 -14472
rect 4356 -14552 5444 -14488
rect 5508 -14552 5528 -14488
rect 4356 -14568 5528 -14552
rect 4356 -14632 5444 -14568
rect 5508 -14632 5528 -14568
rect 4356 -14648 5528 -14632
rect 4356 -14712 5444 -14648
rect 5508 -14712 5528 -14648
rect 4356 -14728 5528 -14712
rect 4356 -14792 5444 -14728
rect 5508 -14792 5528 -14728
rect 4356 -14808 5528 -14792
rect 4356 -14872 5444 -14808
rect 5508 -14872 5528 -14808
rect 4356 -14888 5528 -14872
rect 4356 -14952 5444 -14888
rect 5508 -14952 5528 -14888
rect 4356 -15000 5528 -14952
rect 5768 -14168 6940 -14120
rect 5768 -14232 6856 -14168
rect 6920 -14232 6940 -14168
rect 5768 -14248 6940 -14232
rect 5768 -14312 6856 -14248
rect 6920 -14312 6940 -14248
rect 5768 -14328 6940 -14312
rect 5768 -14392 6856 -14328
rect 6920 -14392 6940 -14328
rect 5768 -14408 6940 -14392
rect 5768 -14472 6856 -14408
rect 6920 -14472 6940 -14408
rect 5768 -14488 6940 -14472
rect 5768 -14552 6856 -14488
rect 6920 -14552 6940 -14488
rect 5768 -14568 6940 -14552
rect 5768 -14632 6856 -14568
rect 6920 -14632 6940 -14568
rect 5768 -14648 6940 -14632
rect 5768 -14712 6856 -14648
rect 6920 -14712 6940 -14648
rect 5768 -14728 6940 -14712
rect 5768 -14792 6856 -14728
rect 6920 -14792 6940 -14728
rect 5768 -14808 6940 -14792
rect 5768 -14872 6856 -14808
rect 6920 -14872 6940 -14808
rect 5768 -14888 6940 -14872
rect 5768 -14952 6856 -14888
rect 6920 -14952 6940 -14888
rect 5768 -15000 6940 -14952
rect 7180 -14168 8352 -14120
rect 7180 -14232 8268 -14168
rect 8332 -14232 8352 -14168
rect 7180 -14248 8352 -14232
rect 7180 -14312 8268 -14248
rect 8332 -14312 8352 -14248
rect 7180 -14328 8352 -14312
rect 7180 -14392 8268 -14328
rect 8332 -14392 8352 -14328
rect 7180 -14408 8352 -14392
rect 7180 -14472 8268 -14408
rect 8332 -14472 8352 -14408
rect 7180 -14488 8352 -14472
rect 7180 -14552 8268 -14488
rect 8332 -14552 8352 -14488
rect 7180 -14568 8352 -14552
rect 7180 -14632 8268 -14568
rect 8332 -14632 8352 -14568
rect 7180 -14648 8352 -14632
rect 7180 -14712 8268 -14648
rect 8332 -14712 8352 -14648
rect 7180 -14728 8352 -14712
rect 7180 -14792 8268 -14728
rect 8332 -14792 8352 -14728
rect 7180 -14808 8352 -14792
rect 7180 -14872 8268 -14808
rect 8332 -14872 8352 -14808
rect 7180 -14888 8352 -14872
rect 7180 -14952 8268 -14888
rect 8332 -14952 8352 -14888
rect 7180 -15000 8352 -14952
rect 8592 -14168 9764 -14120
rect 8592 -14232 9680 -14168
rect 9744 -14232 9764 -14168
rect 8592 -14248 9764 -14232
rect 8592 -14312 9680 -14248
rect 9744 -14312 9764 -14248
rect 8592 -14328 9764 -14312
rect 8592 -14392 9680 -14328
rect 9744 -14392 9764 -14328
rect 8592 -14408 9764 -14392
rect 8592 -14472 9680 -14408
rect 9744 -14472 9764 -14408
rect 8592 -14488 9764 -14472
rect 8592 -14552 9680 -14488
rect 9744 -14552 9764 -14488
rect 8592 -14568 9764 -14552
rect 8592 -14632 9680 -14568
rect 9744 -14632 9764 -14568
rect 8592 -14648 9764 -14632
rect 8592 -14712 9680 -14648
rect 9744 -14712 9764 -14648
rect 8592 -14728 9764 -14712
rect 8592 -14792 9680 -14728
rect 9744 -14792 9764 -14728
rect 8592 -14808 9764 -14792
rect 8592 -14872 9680 -14808
rect 9744 -14872 9764 -14808
rect 8592 -14888 9764 -14872
rect 8592 -14952 9680 -14888
rect 9744 -14952 9764 -14888
rect 8592 -15000 9764 -14952
rect 10004 -14168 11176 -14120
rect 10004 -14232 11092 -14168
rect 11156 -14232 11176 -14168
rect 10004 -14248 11176 -14232
rect 10004 -14312 11092 -14248
rect 11156 -14312 11176 -14248
rect 10004 -14328 11176 -14312
rect 10004 -14392 11092 -14328
rect 11156 -14392 11176 -14328
rect 10004 -14408 11176 -14392
rect 10004 -14472 11092 -14408
rect 11156 -14472 11176 -14408
rect 10004 -14488 11176 -14472
rect 10004 -14552 11092 -14488
rect 11156 -14552 11176 -14488
rect 10004 -14568 11176 -14552
rect 10004 -14632 11092 -14568
rect 11156 -14632 11176 -14568
rect 10004 -14648 11176 -14632
rect 10004 -14712 11092 -14648
rect 11156 -14712 11176 -14648
rect 10004 -14728 11176 -14712
rect 10004 -14792 11092 -14728
rect 11156 -14792 11176 -14728
rect 10004 -14808 11176 -14792
rect 10004 -14872 11092 -14808
rect 11156 -14872 11176 -14808
rect 10004 -14888 11176 -14872
rect 10004 -14952 11092 -14888
rect 11156 -14952 11176 -14888
rect 10004 -15000 11176 -14952
rect 11416 -14168 12588 -14120
rect 11416 -14232 12504 -14168
rect 12568 -14232 12588 -14168
rect 11416 -14248 12588 -14232
rect 11416 -14312 12504 -14248
rect 12568 -14312 12588 -14248
rect 11416 -14328 12588 -14312
rect 11416 -14392 12504 -14328
rect 12568 -14392 12588 -14328
rect 11416 -14408 12588 -14392
rect 11416 -14472 12504 -14408
rect 12568 -14472 12588 -14408
rect 11416 -14488 12588 -14472
rect 11416 -14552 12504 -14488
rect 12568 -14552 12588 -14488
rect 11416 -14568 12588 -14552
rect 11416 -14632 12504 -14568
rect 12568 -14632 12588 -14568
rect 11416 -14648 12588 -14632
rect 11416 -14712 12504 -14648
rect 12568 -14712 12588 -14648
rect 11416 -14728 12588 -14712
rect 11416 -14792 12504 -14728
rect 12568 -14792 12588 -14728
rect 11416 -14808 12588 -14792
rect 11416 -14872 12504 -14808
rect 12568 -14872 12588 -14808
rect 11416 -14888 12588 -14872
rect 11416 -14952 12504 -14888
rect 12568 -14952 12588 -14888
rect 11416 -15000 12588 -14952
rect 12828 -14168 14000 -14120
rect 12828 -14232 13916 -14168
rect 13980 -14232 14000 -14168
rect 12828 -14248 14000 -14232
rect 12828 -14312 13916 -14248
rect 13980 -14312 14000 -14248
rect 12828 -14328 14000 -14312
rect 12828 -14392 13916 -14328
rect 13980 -14392 14000 -14328
rect 12828 -14408 14000 -14392
rect 12828 -14472 13916 -14408
rect 13980 -14472 14000 -14408
rect 12828 -14488 14000 -14472
rect 12828 -14552 13916 -14488
rect 13980 -14552 14000 -14488
rect 12828 -14568 14000 -14552
rect 12828 -14632 13916 -14568
rect 13980 -14632 14000 -14568
rect 12828 -14648 14000 -14632
rect 12828 -14712 13916 -14648
rect 13980 -14712 14000 -14648
rect 12828 -14728 14000 -14712
rect 12828 -14792 13916 -14728
rect 13980 -14792 14000 -14728
rect 12828 -14808 14000 -14792
rect 12828 -14872 13916 -14808
rect 13980 -14872 14000 -14808
rect 12828 -14888 14000 -14872
rect 12828 -14952 13916 -14888
rect 13980 -14952 14000 -14888
rect 12828 -15000 14000 -14952
rect 14240 -14168 15412 -14120
rect 14240 -14232 15328 -14168
rect 15392 -14232 15412 -14168
rect 14240 -14248 15412 -14232
rect 14240 -14312 15328 -14248
rect 15392 -14312 15412 -14248
rect 14240 -14328 15412 -14312
rect 14240 -14392 15328 -14328
rect 15392 -14392 15412 -14328
rect 14240 -14408 15412 -14392
rect 14240 -14472 15328 -14408
rect 15392 -14472 15412 -14408
rect 14240 -14488 15412 -14472
rect 14240 -14552 15328 -14488
rect 15392 -14552 15412 -14488
rect 14240 -14568 15412 -14552
rect 14240 -14632 15328 -14568
rect 15392 -14632 15412 -14568
rect 14240 -14648 15412 -14632
rect 14240 -14712 15328 -14648
rect 15392 -14712 15412 -14648
rect 14240 -14728 15412 -14712
rect 14240 -14792 15328 -14728
rect 15392 -14792 15412 -14728
rect 14240 -14808 15412 -14792
rect 14240 -14872 15328 -14808
rect 15392 -14872 15412 -14808
rect 14240 -14888 15412 -14872
rect 14240 -14952 15328 -14888
rect 15392 -14952 15412 -14888
rect 14240 -15000 15412 -14952
rect 15652 -14168 16824 -14120
rect 15652 -14232 16740 -14168
rect 16804 -14232 16824 -14168
rect 15652 -14248 16824 -14232
rect 15652 -14312 16740 -14248
rect 16804 -14312 16824 -14248
rect 15652 -14328 16824 -14312
rect 15652 -14392 16740 -14328
rect 16804 -14392 16824 -14328
rect 15652 -14408 16824 -14392
rect 15652 -14472 16740 -14408
rect 16804 -14472 16824 -14408
rect 15652 -14488 16824 -14472
rect 15652 -14552 16740 -14488
rect 16804 -14552 16824 -14488
rect 15652 -14568 16824 -14552
rect 15652 -14632 16740 -14568
rect 16804 -14632 16824 -14568
rect 15652 -14648 16824 -14632
rect 15652 -14712 16740 -14648
rect 16804 -14712 16824 -14648
rect 15652 -14728 16824 -14712
rect 15652 -14792 16740 -14728
rect 16804 -14792 16824 -14728
rect 15652 -14808 16824 -14792
rect 15652 -14872 16740 -14808
rect 16804 -14872 16824 -14808
rect 15652 -14888 16824 -14872
rect 15652 -14952 16740 -14888
rect 16804 -14952 16824 -14888
rect 15652 -15000 16824 -14952
rect 17064 -14168 18236 -14120
rect 17064 -14232 18152 -14168
rect 18216 -14232 18236 -14168
rect 17064 -14248 18236 -14232
rect 17064 -14312 18152 -14248
rect 18216 -14312 18236 -14248
rect 17064 -14328 18236 -14312
rect 17064 -14392 18152 -14328
rect 18216 -14392 18236 -14328
rect 17064 -14408 18236 -14392
rect 17064 -14472 18152 -14408
rect 18216 -14472 18236 -14408
rect 17064 -14488 18236 -14472
rect 17064 -14552 18152 -14488
rect 18216 -14552 18236 -14488
rect 17064 -14568 18236 -14552
rect 17064 -14632 18152 -14568
rect 18216 -14632 18236 -14568
rect 17064 -14648 18236 -14632
rect 17064 -14712 18152 -14648
rect 18216 -14712 18236 -14648
rect 17064 -14728 18236 -14712
rect 17064 -14792 18152 -14728
rect 18216 -14792 18236 -14728
rect 17064 -14808 18236 -14792
rect 17064 -14872 18152 -14808
rect 18216 -14872 18236 -14808
rect 17064 -14888 18236 -14872
rect 17064 -14952 18152 -14888
rect 18216 -14952 18236 -14888
rect 17064 -15000 18236 -14952
rect 18476 -14168 19648 -14120
rect 18476 -14232 19564 -14168
rect 19628 -14232 19648 -14168
rect 18476 -14248 19648 -14232
rect 18476 -14312 19564 -14248
rect 19628 -14312 19648 -14248
rect 18476 -14328 19648 -14312
rect 18476 -14392 19564 -14328
rect 19628 -14392 19648 -14328
rect 18476 -14408 19648 -14392
rect 18476 -14472 19564 -14408
rect 19628 -14472 19648 -14408
rect 18476 -14488 19648 -14472
rect 18476 -14552 19564 -14488
rect 19628 -14552 19648 -14488
rect 18476 -14568 19648 -14552
rect 18476 -14632 19564 -14568
rect 19628 -14632 19648 -14568
rect 18476 -14648 19648 -14632
rect 18476 -14712 19564 -14648
rect 19628 -14712 19648 -14648
rect 18476 -14728 19648 -14712
rect 18476 -14792 19564 -14728
rect 19628 -14792 19648 -14728
rect 18476 -14808 19648 -14792
rect 18476 -14872 19564 -14808
rect 19628 -14872 19648 -14808
rect 18476 -14888 19648 -14872
rect 18476 -14952 19564 -14888
rect 19628 -14952 19648 -14888
rect 18476 -15000 19648 -14952
rect 19888 -14168 21060 -14120
rect 19888 -14232 20976 -14168
rect 21040 -14232 21060 -14168
rect 19888 -14248 21060 -14232
rect 19888 -14312 20976 -14248
rect 21040 -14312 21060 -14248
rect 19888 -14328 21060 -14312
rect 19888 -14392 20976 -14328
rect 21040 -14392 21060 -14328
rect 19888 -14408 21060 -14392
rect 19888 -14472 20976 -14408
rect 21040 -14472 21060 -14408
rect 19888 -14488 21060 -14472
rect 19888 -14552 20976 -14488
rect 21040 -14552 21060 -14488
rect 19888 -14568 21060 -14552
rect 19888 -14632 20976 -14568
rect 21040 -14632 21060 -14568
rect 19888 -14648 21060 -14632
rect 19888 -14712 20976 -14648
rect 21040 -14712 21060 -14648
rect 19888 -14728 21060 -14712
rect 19888 -14792 20976 -14728
rect 21040 -14792 21060 -14728
rect 19888 -14808 21060 -14792
rect 19888 -14872 20976 -14808
rect 21040 -14872 21060 -14808
rect 19888 -14888 21060 -14872
rect 19888 -14952 20976 -14888
rect 21040 -14952 21060 -14888
rect 19888 -15000 21060 -14952
rect 21300 -14168 22472 -14120
rect 21300 -14232 22388 -14168
rect 22452 -14232 22472 -14168
rect 21300 -14248 22472 -14232
rect 21300 -14312 22388 -14248
rect 22452 -14312 22472 -14248
rect 21300 -14328 22472 -14312
rect 21300 -14392 22388 -14328
rect 22452 -14392 22472 -14328
rect 21300 -14408 22472 -14392
rect 21300 -14472 22388 -14408
rect 22452 -14472 22472 -14408
rect 21300 -14488 22472 -14472
rect 21300 -14552 22388 -14488
rect 22452 -14552 22472 -14488
rect 21300 -14568 22472 -14552
rect 21300 -14632 22388 -14568
rect 22452 -14632 22472 -14568
rect 21300 -14648 22472 -14632
rect 21300 -14712 22388 -14648
rect 22452 -14712 22472 -14648
rect 21300 -14728 22472 -14712
rect 21300 -14792 22388 -14728
rect 22452 -14792 22472 -14728
rect 21300 -14808 22472 -14792
rect 21300 -14872 22388 -14808
rect 22452 -14872 22472 -14808
rect 21300 -14888 22472 -14872
rect 21300 -14952 22388 -14888
rect 22452 -14952 22472 -14888
rect 21300 -15000 22472 -14952
rect 22712 -14168 23884 -14120
rect 22712 -14232 23800 -14168
rect 23864 -14232 23884 -14168
rect 22712 -14248 23884 -14232
rect 22712 -14312 23800 -14248
rect 23864 -14312 23884 -14248
rect 22712 -14328 23884 -14312
rect 22712 -14392 23800 -14328
rect 23864 -14392 23884 -14328
rect 22712 -14408 23884 -14392
rect 22712 -14472 23800 -14408
rect 23864 -14472 23884 -14408
rect 22712 -14488 23884 -14472
rect 22712 -14552 23800 -14488
rect 23864 -14552 23884 -14488
rect 22712 -14568 23884 -14552
rect 22712 -14632 23800 -14568
rect 23864 -14632 23884 -14568
rect 22712 -14648 23884 -14632
rect 22712 -14712 23800 -14648
rect 23864 -14712 23884 -14648
rect 22712 -14728 23884 -14712
rect 22712 -14792 23800 -14728
rect 23864 -14792 23884 -14728
rect 22712 -14808 23884 -14792
rect 22712 -14872 23800 -14808
rect 23864 -14872 23884 -14808
rect 22712 -14888 23884 -14872
rect 22712 -14952 23800 -14888
rect 23864 -14952 23884 -14888
rect 22712 -15000 23884 -14952
rect -23884 -15288 -22712 -15240
rect -23884 -15352 -22796 -15288
rect -22732 -15352 -22712 -15288
rect -23884 -15368 -22712 -15352
rect -23884 -15432 -22796 -15368
rect -22732 -15432 -22712 -15368
rect -23884 -15448 -22712 -15432
rect -23884 -15512 -22796 -15448
rect -22732 -15512 -22712 -15448
rect -23884 -15528 -22712 -15512
rect -23884 -15592 -22796 -15528
rect -22732 -15592 -22712 -15528
rect -23884 -15608 -22712 -15592
rect -23884 -15672 -22796 -15608
rect -22732 -15672 -22712 -15608
rect -23884 -15688 -22712 -15672
rect -23884 -15752 -22796 -15688
rect -22732 -15752 -22712 -15688
rect -23884 -15768 -22712 -15752
rect -23884 -15832 -22796 -15768
rect -22732 -15832 -22712 -15768
rect -23884 -15848 -22712 -15832
rect -23884 -15912 -22796 -15848
rect -22732 -15912 -22712 -15848
rect -23884 -15928 -22712 -15912
rect -23884 -15992 -22796 -15928
rect -22732 -15992 -22712 -15928
rect -23884 -16008 -22712 -15992
rect -23884 -16072 -22796 -16008
rect -22732 -16072 -22712 -16008
rect -23884 -16120 -22712 -16072
rect -22472 -15288 -21300 -15240
rect -22472 -15352 -21384 -15288
rect -21320 -15352 -21300 -15288
rect -22472 -15368 -21300 -15352
rect -22472 -15432 -21384 -15368
rect -21320 -15432 -21300 -15368
rect -22472 -15448 -21300 -15432
rect -22472 -15512 -21384 -15448
rect -21320 -15512 -21300 -15448
rect -22472 -15528 -21300 -15512
rect -22472 -15592 -21384 -15528
rect -21320 -15592 -21300 -15528
rect -22472 -15608 -21300 -15592
rect -22472 -15672 -21384 -15608
rect -21320 -15672 -21300 -15608
rect -22472 -15688 -21300 -15672
rect -22472 -15752 -21384 -15688
rect -21320 -15752 -21300 -15688
rect -22472 -15768 -21300 -15752
rect -22472 -15832 -21384 -15768
rect -21320 -15832 -21300 -15768
rect -22472 -15848 -21300 -15832
rect -22472 -15912 -21384 -15848
rect -21320 -15912 -21300 -15848
rect -22472 -15928 -21300 -15912
rect -22472 -15992 -21384 -15928
rect -21320 -15992 -21300 -15928
rect -22472 -16008 -21300 -15992
rect -22472 -16072 -21384 -16008
rect -21320 -16072 -21300 -16008
rect -22472 -16120 -21300 -16072
rect -21060 -15288 -19888 -15240
rect -21060 -15352 -19972 -15288
rect -19908 -15352 -19888 -15288
rect -21060 -15368 -19888 -15352
rect -21060 -15432 -19972 -15368
rect -19908 -15432 -19888 -15368
rect -21060 -15448 -19888 -15432
rect -21060 -15512 -19972 -15448
rect -19908 -15512 -19888 -15448
rect -21060 -15528 -19888 -15512
rect -21060 -15592 -19972 -15528
rect -19908 -15592 -19888 -15528
rect -21060 -15608 -19888 -15592
rect -21060 -15672 -19972 -15608
rect -19908 -15672 -19888 -15608
rect -21060 -15688 -19888 -15672
rect -21060 -15752 -19972 -15688
rect -19908 -15752 -19888 -15688
rect -21060 -15768 -19888 -15752
rect -21060 -15832 -19972 -15768
rect -19908 -15832 -19888 -15768
rect -21060 -15848 -19888 -15832
rect -21060 -15912 -19972 -15848
rect -19908 -15912 -19888 -15848
rect -21060 -15928 -19888 -15912
rect -21060 -15992 -19972 -15928
rect -19908 -15992 -19888 -15928
rect -21060 -16008 -19888 -15992
rect -21060 -16072 -19972 -16008
rect -19908 -16072 -19888 -16008
rect -21060 -16120 -19888 -16072
rect -19648 -15288 -18476 -15240
rect -19648 -15352 -18560 -15288
rect -18496 -15352 -18476 -15288
rect -19648 -15368 -18476 -15352
rect -19648 -15432 -18560 -15368
rect -18496 -15432 -18476 -15368
rect -19648 -15448 -18476 -15432
rect -19648 -15512 -18560 -15448
rect -18496 -15512 -18476 -15448
rect -19648 -15528 -18476 -15512
rect -19648 -15592 -18560 -15528
rect -18496 -15592 -18476 -15528
rect -19648 -15608 -18476 -15592
rect -19648 -15672 -18560 -15608
rect -18496 -15672 -18476 -15608
rect -19648 -15688 -18476 -15672
rect -19648 -15752 -18560 -15688
rect -18496 -15752 -18476 -15688
rect -19648 -15768 -18476 -15752
rect -19648 -15832 -18560 -15768
rect -18496 -15832 -18476 -15768
rect -19648 -15848 -18476 -15832
rect -19648 -15912 -18560 -15848
rect -18496 -15912 -18476 -15848
rect -19648 -15928 -18476 -15912
rect -19648 -15992 -18560 -15928
rect -18496 -15992 -18476 -15928
rect -19648 -16008 -18476 -15992
rect -19648 -16072 -18560 -16008
rect -18496 -16072 -18476 -16008
rect -19648 -16120 -18476 -16072
rect -18236 -15288 -17064 -15240
rect -18236 -15352 -17148 -15288
rect -17084 -15352 -17064 -15288
rect -18236 -15368 -17064 -15352
rect -18236 -15432 -17148 -15368
rect -17084 -15432 -17064 -15368
rect -18236 -15448 -17064 -15432
rect -18236 -15512 -17148 -15448
rect -17084 -15512 -17064 -15448
rect -18236 -15528 -17064 -15512
rect -18236 -15592 -17148 -15528
rect -17084 -15592 -17064 -15528
rect -18236 -15608 -17064 -15592
rect -18236 -15672 -17148 -15608
rect -17084 -15672 -17064 -15608
rect -18236 -15688 -17064 -15672
rect -18236 -15752 -17148 -15688
rect -17084 -15752 -17064 -15688
rect -18236 -15768 -17064 -15752
rect -18236 -15832 -17148 -15768
rect -17084 -15832 -17064 -15768
rect -18236 -15848 -17064 -15832
rect -18236 -15912 -17148 -15848
rect -17084 -15912 -17064 -15848
rect -18236 -15928 -17064 -15912
rect -18236 -15992 -17148 -15928
rect -17084 -15992 -17064 -15928
rect -18236 -16008 -17064 -15992
rect -18236 -16072 -17148 -16008
rect -17084 -16072 -17064 -16008
rect -18236 -16120 -17064 -16072
rect -16824 -15288 -15652 -15240
rect -16824 -15352 -15736 -15288
rect -15672 -15352 -15652 -15288
rect -16824 -15368 -15652 -15352
rect -16824 -15432 -15736 -15368
rect -15672 -15432 -15652 -15368
rect -16824 -15448 -15652 -15432
rect -16824 -15512 -15736 -15448
rect -15672 -15512 -15652 -15448
rect -16824 -15528 -15652 -15512
rect -16824 -15592 -15736 -15528
rect -15672 -15592 -15652 -15528
rect -16824 -15608 -15652 -15592
rect -16824 -15672 -15736 -15608
rect -15672 -15672 -15652 -15608
rect -16824 -15688 -15652 -15672
rect -16824 -15752 -15736 -15688
rect -15672 -15752 -15652 -15688
rect -16824 -15768 -15652 -15752
rect -16824 -15832 -15736 -15768
rect -15672 -15832 -15652 -15768
rect -16824 -15848 -15652 -15832
rect -16824 -15912 -15736 -15848
rect -15672 -15912 -15652 -15848
rect -16824 -15928 -15652 -15912
rect -16824 -15992 -15736 -15928
rect -15672 -15992 -15652 -15928
rect -16824 -16008 -15652 -15992
rect -16824 -16072 -15736 -16008
rect -15672 -16072 -15652 -16008
rect -16824 -16120 -15652 -16072
rect -15412 -15288 -14240 -15240
rect -15412 -15352 -14324 -15288
rect -14260 -15352 -14240 -15288
rect -15412 -15368 -14240 -15352
rect -15412 -15432 -14324 -15368
rect -14260 -15432 -14240 -15368
rect -15412 -15448 -14240 -15432
rect -15412 -15512 -14324 -15448
rect -14260 -15512 -14240 -15448
rect -15412 -15528 -14240 -15512
rect -15412 -15592 -14324 -15528
rect -14260 -15592 -14240 -15528
rect -15412 -15608 -14240 -15592
rect -15412 -15672 -14324 -15608
rect -14260 -15672 -14240 -15608
rect -15412 -15688 -14240 -15672
rect -15412 -15752 -14324 -15688
rect -14260 -15752 -14240 -15688
rect -15412 -15768 -14240 -15752
rect -15412 -15832 -14324 -15768
rect -14260 -15832 -14240 -15768
rect -15412 -15848 -14240 -15832
rect -15412 -15912 -14324 -15848
rect -14260 -15912 -14240 -15848
rect -15412 -15928 -14240 -15912
rect -15412 -15992 -14324 -15928
rect -14260 -15992 -14240 -15928
rect -15412 -16008 -14240 -15992
rect -15412 -16072 -14324 -16008
rect -14260 -16072 -14240 -16008
rect -15412 -16120 -14240 -16072
rect -14000 -15288 -12828 -15240
rect -14000 -15352 -12912 -15288
rect -12848 -15352 -12828 -15288
rect -14000 -15368 -12828 -15352
rect -14000 -15432 -12912 -15368
rect -12848 -15432 -12828 -15368
rect -14000 -15448 -12828 -15432
rect -14000 -15512 -12912 -15448
rect -12848 -15512 -12828 -15448
rect -14000 -15528 -12828 -15512
rect -14000 -15592 -12912 -15528
rect -12848 -15592 -12828 -15528
rect -14000 -15608 -12828 -15592
rect -14000 -15672 -12912 -15608
rect -12848 -15672 -12828 -15608
rect -14000 -15688 -12828 -15672
rect -14000 -15752 -12912 -15688
rect -12848 -15752 -12828 -15688
rect -14000 -15768 -12828 -15752
rect -14000 -15832 -12912 -15768
rect -12848 -15832 -12828 -15768
rect -14000 -15848 -12828 -15832
rect -14000 -15912 -12912 -15848
rect -12848 -15912 -12828 -15848
rect -14000 -15928 -12828 -15912
rect -14000 -15992 -12912 -15928
rect -12848 -15992 -12828 -15928
rect -14000 -16008 -12828 -15992
rect -14000 -16072 -12912 -16008
rect -12848 -16072 -12828 -16008
rect -14000 -16120 -12828 -16072
rect -12588 -15288 -11416 -15240
rect -12588 -15352 -11500 -15288
rect -11436 -15352 -11416 -15288
rect -12588 -15368 -11416 -15352
rect -12588 -15432 -11500 -15368
rect -11436 -15432 -11416 -15368
rect -12588 -15448 -11416 -15432
rect -12588 -15512 -11500 -15448
rect -11436 -15512 -11416 -15448
rect -12588 -15528 -11416 -15512
rect -12588 -15592 -11500 -15528
rect -11436 -15592 -11416 -15528
rect -12588 -15608 -11416 -15592
rect -12588 -15672 -11500 -15608
rect -11436 -15672 -11416 -15608
rect -12588 -15688 -11416 -15672
rect -12588 -15752 -11500 -15688
rect -11436 -15752 -11416 -15688
rect -12588 -15768 -11416 -15752
rect -12588 -15832 -11500 -15768
rect -11436 -15832 -11416 -15768
rect -12588 -15848 -11416 -15832
rect -12588 -15912 -11500 -15848
rect -11436 -15912 -11416 -15848
rect -12588 -15928 -11416 -15912
rect -12588 -15992 -11500 -15928
rect -11436 -15992 -11416 -15928
rect -12588 -16008 -11416 -15992
rect -12588 -16072 -11500 -16008
rect -11436 -16072 -11416 -16008
rect -12588 -16120 -11416 -16072
rect -11176 -15288 -10004 -15240
rect -11176 -15352 -10088 -15288
rect -10024 -15352 -10004 -15288
rect -11176 -15368 -10004 -15352
rect -11176 -15432 -10088 -15368
rect -10024 -15432 -10004 -15368
rect -11176 -15448 -10004 -15432
rect -11176 -15512 -10088 -15448
rect -10024 -15512 -10004 -15448
rect -11176 -15528 -10004 -15512
rect -11176 -15592 -10088 -15528
rect -10024 -15592 -10004 -15528
rect -11176 -15608 -10004 -15592
rect -11176 -15672 -10088 -15608
rect -10024 -15672 -10004 -15608
rect -11176 -15688 -10004 -15672
rect -11176 -15752 -10088 -15688
rect -10024 -15752 -10004 -15688
rect -11176 -15768 -10004 -15752
rect -11176 -15832 -10088 -15768
rect -10024 -15832 -10004 -15768
rect -11176 -15848 -10004 -15832
rect -11176 -15912 -10088 -15848
rect -10024 -15912 -10004 -15848
rect -11176 -15928 -10004 -15912
rect -11176 -15992 -10088 -15928
rect -10024 -15992 -10004 -15928
rect -11176 -16008 -10004 -15992
rect -11176 -16072 -10088 -16008
rect -10024 -16072 -10004 -16008
rect -11176 -16120 -10004 -16072
rect -9764 -15288 -8592 -15240
rect -9764 -15352 -8676 -15288
rect -8612 -15352 -8592 -15288
rect -9764 -15368 -8592 -15352
rect -9764 -15432 -8676 -15368
rect -8612 -15432 -8592 -15368
rect -9764 -15448 -8592 -15432
rect -9764 -15512 -8676 -15448
rect -8612 -15512 -8592 -15448
rect -9764 -15528 -8592 -15512
rect -9764 -15592 -8676 -15528
rect -8612 -15592 -8592 -15528
rect -9764 -15608 -8592 -15592
rect -9764 -15672 -8676 -15608
rect -8612 -15672 -8592 -15608
rect -9764 -15688 -8592 -15672
rect -9764 -15752 -8676 -15688
rect -8612 -15752 -8592 -15688
rect -9764 -15768 -8592 -15752
rect -9764 -15832 -8676 -15768
rect -8612 -15832 -8592 -15768
rect -9764 -15848 -8592 -15832
rect -9764 -15912 -8676 -15848
rect -8612 -15912 -8592 -15848
rect -9764 -15928 -8592 -15912
rect -9764 -15992 -8676 -15928
rect -8612 -15992 -8592 -15928
rect -9764 -16008 -8592 -15992
rect -9764 -16072 -8676 -16008
rect -8612 -16072 -8592 -16008
rect -9764 -16120 -8592 -16072
rect -8352 -15288 -7180 -15240
rect -8352 -15352 -7264 -15288
rect -7200 -15352 -7180 -15288
rect -8352 -15368 -7180 -15352
rect -8352 -15432 -7264 -15368
rect -7200 -15432 -7180 -15368
rect -8352 -15448 -7180 -15432
rect -8352 -15512 -7264 -15448
rect -7200 -15512 -7180 -15448
rect -8352 -15528 -7180 -15512
rect -8352 -15592 -7264 -15528
rect -7200 -15592 -7180 -15528
rect -8352 -15608 -7180 -15592
rect -8352 -15672 -7264 -15608
rect -7200 -15672 -7180 -15608
rect -8352 -15688 -7180 -15672
rect -8352 -15752 -7264 -15688
rect -7200 -15752 -7180 -15688
rect -8352 -15768 -7180 -15752
rect -8352 -15832 -7264 -15768
rect -7200 -15832 -7180 -15768
rect -8352 -15848 -7180 -15832
rect -8352 -15912 -7264 -15848
rect -7200 -15912 -7180 -15848
rect -8352 -15928 -7180 -15912
rect -8352 -15992 -7264 -15928
rect -7200 -15992 -7180 -15928
rect -8352 -16008 -7180 -15992
rect -8352 -16072 -7264 -16008
rect -7200 -16072 -7180 -16008
rect -8352 -16120 -7180 -16072
rect -6940 -15288 -5768 -15240
rect -6940 -15352 -5852 -15288
rect -5788 -15352 -5768 -15288
rect -6940 -15368 -5768 -15352
rect -6940 -15432 -5852 -15368
rect -5788 -15432 -5768 -15368
rect -6940 -15448 -5768 -15432
rect -6940 -15512 -5852 -15448
rect -5788 -15512 -5768 -15448
rect -6940 -15528 -5768 -15512
rect -6940 -15592 -5852 -15528
rect -5788 -15592 -5768 -15528
rect -6940 -15608 -5768 -15592
rect -6940 -15672 -5852 -15608
rect -5788 -15672 -5768 -15608
rect -6940 -15688 -5768 -15672
rect -6940 -15752 -5852 -15688
rect -5788 -15752 -5768 -15688
rect -6940 -15768 -5768 -15752
rect -6940 -15832 -5852 -15768
rect -5788 -15832 -5768 -15768
rect -6940 -15848 -5768 -15832
rect -6940 -15912 -5852 -15848
rect -5788 -15912 -5768 -15848
rect -6940 -15928 -5768 -15912
rect -6940 -15992 -5852 -15928
rect -5788 -15992 -5768 -15928
rect -6940 -16008 -5768 -15992
rect -6940 -16072 -5852 -16008
rect -5788 -16072 -5768 -16008
rect -6940 -16120 -5768 -16072
rect -5528 -15288 -4356 -15240
rect -5528 -15352 -4440 -15288
rect -4376 -15352 -4356 -15288
rect -5528 -15368 -4356 -15352
rect -5528 -15432 -4440 -15368
rect -4376 -15432 -4356 -15368
rect -5528 -15448 -4356 -15432
rect -5528 -15512 -4440 -15448
rect -4376 -15512 -4356 -15448
rect -5528 -15528 -4356 -15512
rect -5528 -15592 -4440 -15528
rect -4376 -15592 -4356 -15528
rect -5528 -15608 -4356 -15592
rect -5528 -15672 -4440 -15608
rect -4376 -15672 -4356 -15608
rect -5528 -15688 -4356 -15672
rect -5528 -15752 -4440 -15688
rect -4376 -15752 -4356 -15688
rect -5528 -15768 -4356 -15752
rect -5528 -15832 -4440 -15768
rect -4376 -15832 -4356 -15768
rect -5528 -15848 -4356 -15832
rect -5528 -15912 -4440 -15848
rect -4376 -15912 -4356 -15848
rect -5528 -15928 -4356 -15912
rect -5528 -15992 -4440 -15928
rect -4376 -15992 -4356 -15928
rect -5528 -16008 -4356 -15992
rect -5528 -16072 -4440 -16008
rect -4376 -16072 -4356 -16008
rect -5528 -16120 -4356 -16072
rect -4116 -15288 -2944 -15240
rect -4116 -15352 -3028 -15288
rect -2964 -15352 -2944 -15288
rect -4116 -15368 -2944 -15352
rect -4116 -15432 -3028 -15368
rect -2964 -15432 -2944 -15368
rect -4116 -15448 -2944 -15432
rect -4116 -15512 -3028 -15448
rect -2964 -15512 -2944 -15448
rect -4116 -15528 -2944 -15512
rect -4116 -15592 -3028 -15528
rect -2964 -15592 -2944 -15528
rect -4116 -15608 -2944 -15592
rect -4116 -15672 -3028 -15608
rect -2964 -15672 -2944 -15608
rect -4116 -15688 -2944 -15672
rect -4116 -15752 -3028 -15688
rect -2964 -15752 -2944 -15688
rect -4116 -15768 -2944 -15752
rect -4116 -15832 -3028 -15768
rect -2964 -15832 -2944 -15768
rect -4116 -15848 -2944 -15832
rect -4116 -15912 -3028 -15848
rect -2964 -15912 -2944 -15848
rect -4116 -15928 -2944 -15912
rect -4116 -15992 -3028 -15928
rect -2964 -15992 -2944 -15928
rect -4116 -16008 -2944 -15992
rect -4116 -16072 -3028 -16008
rect -2964 -16072 -2944 -16008
rect -4116 -16120 -2944 -16072
rect -2704 -15288 -1532 -15240
rect -2704 -15352 -1616 -15288
rect -1552 -15352 -1532 -15288
rect -2704 -15368 -1532 -15352
rect -2704 -15432 -1616 -15368
rect -1552 -15432 -1532 -15368
rect -2704 -15448 -1532 -15432
rect -2704 -15512 -1616 -15448
rect -1552 -15512 -1532 -15448
rect -2704 -15528 -1532 -15512
rect -2704 -15592 -1616 -15528
rect -1552 -15592 -1532 -15528
rect -2704 -15608 -1532 -15592
rect -2704 -15672 -1616 -15608
rect -1552 -15672 -1532 -15608
rect -2704 -15688 -1532 -15672
rect -2704 -15752 -1616 -15688
rect -1552 -15752 -1532 -15688
rect -2704 -15768 -1532 -15752
rect -2704 -15832 -1616 -15768
rect -1552 -15832 -1532 -15768
rect -2704 -15848 -1532 -15832
rect -2704 -15912 -1616 -15848
rect -1552 -15912 -1532 -15848
rect -2704 -15928 -1532 -15912
rect -2704 -15992 -1616 -15928
rect -1552 -15992 -1532 -15928
rect -2704 -16008 -1532 -15992
rect -2704 -16072 -1616 -16008
rect -1552 -16072 -1532 -16008
rect -2704 -16120 -1532 -16072
rect -1292 -15288 -120 -15240
rect -1292 -15352 -204 -15288
rect -140 -15352 -120 -15288
rect -1292 -15368 -120 -15352
rect -1292 -15432 -204 -15368
rect -140 -15432 -120 -15368
rect -1292 -15448 -120 -15432
rect -1292 -15512 -204 -15448
rect -140 -15512 -120 -15448
rect -1292 -15528 -120 -15512
rect -1292 -15592 -204 -15528
rect -140 -15592 -120 -15528
rect -1292 -15608 -120 -15592
rect -1292 -15672 -204 -15608
rect -140 -15672 -120 -15608
rect -1292 -15688 -120 -15672
rect -1292 -15752 -204 -15688
rect -140 -15752 -120 -15688
rect -1292 -15768 -120 -15752
rect -1292 -15832 -204 -15768
rect -140 -15832 -120 -15768
rect -1292 -15848 -120 -15832
rect -1292 -15912 -204 -15848
rect -140 -15912 -120 -15848
rect -1292 -15928 -120 -15912
rect -1292 -15992 -204 -15928
rect -140 -15992 -120 -15928
rect -1292 -16008 -120 -15992
rect -1292 -16072 -204 -16008
rect -140 -16072 -120 -16008
rect -1292 -16120 -120 -16072
rect 120 -15288 1292 -15240
rect 120 -15352 1208 -15288
rect 1272 -15352 1292 -15288
rect 120 -15368 1292 -15352
rect 120 -15432 1208 -15368
rect 1272 -15432 1292 -15368
rect 120 -15448 1292 -15432
rect 120 -15512 1208 -15448
rect 1272 -15512 1292 -15448
rect 120 -15528 1292 -15512
rect 120 -15592 1208 -15528
rect 1272 -15592 1292 -15528
rect 120 -15608 1292 -15592
rect 120 -15672 1208 -15608
rect 1272 -15672 1292 -15608
rect 120 -15688 1292 -15672
rect 120 -15752 1208 -15688
rect 1272 -15752 1292 -15688
rect 120 -15768 1292 -15752
rect 120 -15832 1208 -15768
rect 1272 -15832 1292 -15768
rect 120 -15848 1292 -15832
rect 120 -15912 1208 -15848
rect 1272 -15912 1292 -15848
rect 120 -15928 1292 -15912
rect 120 -15992 1208 -15928
rect 1272 -15992 1292 -15928
rect 120 -16008 1292 -15992
rect 120 -16072 1208 -16008
rect 1272 -16072 1292 -16008
rect 120 -16120 1292 -16072
rect 1532 -15288 2704 -15240
rect 1532 -15352 2620 -15288
rect 2684 -15352 2704 -15288
rect 1532 -15368 2704 -15352
rect 1532 -15432 2620 -15368
rect 2684 -15432 2704 -15368
rect 1532 -15448 2704 -15432
rect 1532 -15512 2620 -15448
rect 2684 -15512 2704 -15448
rect 1532 -15528 2704 -15512
rect 1532 -15592 2620 -15528
rect 2684 -15592 2704 -15528
rect 1532 -15608 2704 -15592
rect 1532 -15672 2620 -15608
rect 2684 -15672 2704 -15608
rect 1532 -15688 2704 -15672
rect 1532 -15752 2620 -15688
rect 2684 -15752 2704 -15688
rect 1532 -15768 2704 -15752
rect 1532 -15832 2620 -15768
rect 2684 -15832 2704 -15768
rect 1532 -15848 2704 -15832
rect 1532 -15912 2620 -15848
rect 2684 -15912 2704 -15848
rect 1532 -15928 2704 -15912
rect 1532 -15992 2620 -15928
rect 2684 -15992 2704 -15928
rect 1532 -16008 2704 -15992
rect 1532 -16072 2620 -16008
rect 2684 -16072 2704 -16008
rect 1532 -16120 2704 -16072
rect 2944 -15288 4116 -15240
rect 2944 -15352 4032 -15288
rect 4096 -15352 4116 -15288
rect 2944 -15368 4116 -15352
rect 2944 -15432 4032 -15368
rect 4096 -15432 4116 -15368
rect 2944 -15448 4116 -15432
rect 2944 -15512 4032 -15448
rect 4096 -15512 4116 -15448
rect 2944 -15528 4116 -15512
rect 2944 -15592 4032 -15528
rect 4096 -15592 4116 -15528
rect 2944 -15608 4116 -15592
rect 2944 -15672 4032 -15608
rect 4096 -15672 4116 -15608
rect 2944 -15688 4116 -15672
rect 2944 -15752 4032 -15688
rect 4096 -15752 4116 -15688
rect 2944 -15768 4116 -15752
rect 2944 -15832 4032 -15768
rect 4096 -15832 4116 -15768
rect 2944 -15848 4116 -15832
rect 2944 -15912 4032 -15848
rect 4096 -15912 4116 -15848
rect 2944 -15928 4116 -15912
rect 2944 -15992 4032 -15928
rect 4096 -15992 4116 -15928
rect 2944 -16008 4116 -15992
rect 2944 -16072 4032 -16008
rect 4096 -16072 4116 -16008
rect 2944 -16120 4116 -16072
rect 4356 -15288 5528 -15240
rect 4356 -15352 5444 -15288
rect 5508 -15352 5528 -15288
rect 4356 -15368 5528 -15352
rect 4356 -15432 5444 -15368
rect 5508 -15432 5528 -15368
rect 4356 -15448 5528 -15432
rect 4356 -15512 5444 -15448
rect 5508 -15512 5528 -15448
rect 4356 -15528 5528 -15512
rect 4356 -15592 5444 -15528
rect 5508 -15592 5528 -15528
rect 4356 -15608 5528 -15592
rect 4356 -15672 5444 -15608
rect 5508 -15672 5528 -15608
rect 4356 -15688 5528 -15672
rect 4356 -15752 5444 -15688
rect 5508 -15752 5528 -15688
rect 4356 -15768 5528 -15752
rect 4356 -15832 5444 -15768
rect 5508 -15832 5528 -15768
rect 4356 -15848 5528 -15832
rect 4356 -15912 5444 -15848
rect 5508 -15912 5528 -15848
rect 4356 -15928 5528 -15912
rect 4356 -15992 5444 -15928
rect 5508 -15992 5528 -15928
rect 4356 -16008 5528 -15992
rect 4356 -16072 5444 -16008
rect 5508 -16072 5528 -16008
rect 4356 -16120 5528 -16072
rect 5768 -15288 6940 -15240
rect 5768 -15352 6856 -15288
rect 6920 -15352 6940 -15288
rect 5768 -15368 6940 -15352
rect 5768 -15432 6856 -15368
rect 6920 -15432 6940 -15368
rect 5768 -15448 6940 -15432
rect 5768 -15512 6856 -15448
rect 6920 -15512 6940 -15448
rect 5768 -15528 6940 -15512
rect 5768 -15592 6856 -15528
rect 6920 -15592 6940 -15528
rect 5768 -15608 6940 -15592
rect 5768 -15672 6856 -15608
rect 6920 -15672 6940 -15608
rect 5768 -15688 6940 -15672
rect 5768 -15752 6856 -15688
rect 6920 -15752 6940 -15688
rect 5768 -15768 6940 -15752
rect 5768 -15832 6856 -15768
rect 6920 -15832 6940 -15768
rect 5768 -15848 6940 -15832
rect 5768 -15912 6856 -15848
rect 6920 -15912 6940 -15848
rect 5768 -15928 6940 -15912
rect 5768 -15992 6856 -15928
rect 6920 -15992 6940 -15928
rect 5768 -16008 6940 -15992
rect 5768 -16072 6856 -16008
rect 6920 -16072 6940 -16008
rect 5768 -16120 6940 -16072
rect 7180 -15288 8352 -15240
rect 7180 -15352 8268 -15288
rect 8332 -15352 8352 -15288
rect 7180 -15368 8352 -15352
rect 7180 -15432 8268 -15368
rect 8332 -15432 8352 -15368
rect 7180 -15448 8352 -15432
rect 7180 -15512 8268 -15448
rect 8332 -15512 8352 -15448
rect 7180 -15528 8352 -15512
rect 7180 -15592 8268 -15528
rect 8332 -15592 8352 -15528
rect 7180 -15608 8352 -15592
rect 7180 -15672 8268 -15608
rect 8332 -15672 8352 -15608
rect 7180 -15688 8352 -15672
rect 7180 -15752 8268 -15688
rect 8332 -15752 8352 -15688
rect 7180 -15768 8352 -15752
rect 7180 -15832 8268 -15768
rect 8332 -15832 8352 -15768
rect 7180 -15848 8352 -15832
rect 7180 -15912 8268 -15848
rect 8332 -15912 8352 -15848
rect 7180 -15928 8352 -15912
rect 7180 -15992 8268 -15928
rect 8332 -15992 8352 -15928
rect 7180 -16008 8352 -15992
rect 7180 -16072 8268 -16008
rect 8332 -16072 8352 -16008
rect 7180 -16120 8352 -16072
rect 8592 -15288 9764 -15240
rect 8592 -15352 9680 -15288
rect 9744 -15352 9764 -15288
rect 8592 -15368 9764 -15352
rect 8592 -15432 9680 -15368
rect 9744 -15432 9764 -15368
rect 8592 -15448 9764 -15432
rect 8592 -15512 9680 -15448
rect 9744 -15512 9764 -15448
rect 8592 -15528 9764 -15512
rect 8592 -15592 9680 -15528
rect 9744 -15592 9764 -15528
rect 8592 -15608 9764 -15592
rect 8592 -15672 9680 -15608
rect 9744 -15672 9764 -15608
rect 8592 -15688 9764 -15672
rect 8592 -15752 9680 -15688
rect 9744 -15752 9764 -15688
rect 8592 -15768 9764 -15752
rect 8592 -15832 9680 -15768
rect 9744 -15832 9764 -15768
rect 8592 -15848 9764 -15832
rect 8592 -15912 9680 -15848
rect 9744 -15912 9764 -15848
rect 8592 -15928 9764 -15912
rect 8592 -15992 9680 -15928
rect 9744 -15992 9764 -15928
rect 8592 -16008 9764 -15992
rect 8592 -16072 9680 -16008
rect 9744 -16072 9764 -16008
rect 8592 -16120 9764 -16072
rect 10004 -15288 11176 -15240
rect 10004 -15352 11092 -15288
rect 11156 -15352 11176 -15288
rect 10004 -15368 11176 -15352
rect 10004 -15432 11092 -15368
rect 11156 -15432 11176 -15368
rect 10004 -15448 11176 -15432
rect 10004 -15512 11092 -15448
rect 11156 -15512 11176 -15448
rect 10004 -15528 11176 -15512
rect 10004 -15592 11092 -15528
rect 11156 -15592 11176 -15528
rect 10004 -15608 11176 -15592
rect 10004 -15672 11092 -15608
rect 11156 -15672 11176 -15608
rect 10004 -15688 11176 -15672
rect 10004 -15752 11092 -15688
rect 11156 -15752 11176 -15688
rect 10004 -15768 11176 -15752
rect 10004 -15832 11092 -15768
rect 11156 -15832 11176 -15768
rect 10004 -15848 11176 -15832
rect 10004 -15912 11092 -15848
rect 11156 -15912 11176 -15848
rect 10004 -15928 11176 -15912
rect 10004 -15992 11092 -15928
rect 11156 -15992 11176 -15928
rect 10004 -16008 11176 -15992
rect 10004 -16072 11092 -16008
rect 11156 -16072 11176 -16008
rect 10004 -16120 11176 -16072
rect 11416 -15288 12588 -15240
rect 11416 -15352 12504 -15288
rect 12568 -15352 12588 -15288
rect 11416 -15368 12588 -15352
rect 11416 -15432 12504 -15368
rect 12568 -15432 12588 -15368
rect 11416 -15448 12588 -15432
rect 11416 -15512 12504 -15448
rect 12568 -15512 12588 -15448
rect 11416 -15528 12588 -15512
rect 11416 -15592 12504 -15528
rect 12568 -15592 12588 -15528
rect 11416 -15608 12588 -15592
rect 11416 -15672 12504 -15608
rect 12568 -15672 12588 -15608
rect 11416 -15688 12588 -15672
rect 11416 -15752 12504 -15688
rect 12568 -15752 12588 -15688
rect 11416 -15768 12588 -15752
rect 11416 -15832 12504 -15768
rect 12568 -15832 12588 -15768
rect 11416 -15848 12588 -15832
rect 11416 -15912 12504 -15848
rect 12568 -15912 12588 -15848
rect 11416 -15928 12588 -15912
rect 11416 -15992 12504 -15928
rect 12568 -15992 12588 -15928
rect 11416 -16008 12588 -15992
rect 11416 -16072 12504 -16008
rect 12568 -16072 12588 -16008
rect 11416 -16120 12588 -16072
rect 12828 -15288 14000 -15240
rect 12828 -15352 13916 -15288
rect 13980 -15352 14000 -15288
rect 12828 -15368 14000 -15352
rect 12828 -15432 13916 -15368
rect 13980 -15432 14000 -15368
rect 12828 -15448 14000 -15432
rect 12828 -15512 13916 -15448
rect 13980 -15512 14000 -15448
rect 12828 -15528 14000 -15512
rect 12828 -15592 13916 -15528
rect 13980 -15592 14000 -15528
rect 12828 -15608 14000 -15592
rect 12828 -15672 13916 -15608
rect 13980 -15672 14000 -15608
rect 12828 -15688 14000 -15672
rect 12828 -15752 13916 -15688
rect 13980 -15752 14000 -15688
rect 12828 -15768 14000 -15752
rect 12828 -15832 13916 -15768
rect 13980 -15832 14000 -15768
rect 12828 -15848 14000 -15832
rect 12828 -15912 13916 -15848
rect 13980 -15912 14000 -15848
rect 12828 -15928 14000 -15912
rect 12828 -15992 13916 -15928
rect 13980 -15992 14000 -15928
rect 12828 -16008 14000 -15992
rect 12828 -16072 13916 -16008
rect 13980 -16072 14000 -16008
rect 12828 -16120 14000 -16072
rect 14240 -15288 15412 -15240
rect 14240 -15352 15328 -15288
rect 15392 -15352 15412 -15288
rect 14240 -15368 15412 -15352
rect 14240 -15432 15328 -15368
rect 15392 -15432 15412 -15368
rect 14240 -15448 15412 -15432
rect 14240 -15512 15328 -15448
rect 15392 -15512 15412 -15448
rect 14240 -15528 15412 -15512
rect 14240 -15592 15328 -15528
rect 15392 -15592 15412 -15528
rect 14240 -15608 15412 -15592
rect 14240 -15672 15328 -15608
rect 15392 -15672 15412 -15608
rect 14240 -15688 15412 -15672
rect 14240 -15752 15328 -15688
rect 15392 -15752 15412 -15688
rect 14240 -15768 15412 -15752
rect 14240 -15832 15328 -15768
rect 15392 -15832 15412 -15768
rect 14240 -15848 15412 -15832
rect 14240 -15912 15328 -15848
rect 15392 -15912 15412 -15848
rect 14240 -15928 15412 -15912
rect 14240 -15992 15328 -15928
rect 15392 -15992 15412 -15928
rect 14240 -16008 15412 -15992
rect 14240 -16072 15328 -16008
rect 15392 -16072 15412 -16008
rect 14240 -16120 15412 -16072
rect 15652 -15288 16824 -15240
rect 15652 -15352 16740 -15288
rect 16804 -15352 16824 -15288
rect 15652 -15368 16824 -15352
rect 15652 -15432 16740 -15368
rect 16804 -15432 16824 -15368
rect 15652 -15448 16824 -15432
rect 15652 -15512 16740 -15448
rect 16804 -15512 16824 -15448
rect 15652 -15528 16824 -15512
rect 15652 -15592 16740 -15528
rect 16804 -15592 16824 -15528
rect 15652 -15608 16824 -15592
rect 15652 -15672 16740 -15608
rect 16804 -15672 16824 -15608
rect 15652 -15688 16824 -15672
rect 15652 -15752 16740 -15688
rect 16804 -15752 16824 -15688
rect 15652 -15768 16824 -15752
rect 15652 -15832 16740 -15768
rect 16804 -15832 16824 -15768
rect 15652 -15848 16824 -15832
rect 15652 -15912 16740 -15848
rect 16804 -15912 16824 -15848
rect 15652 -15928 16824 -15912
rect 15652 -15992 16740 -15928
rect 16804 -15992 16824 -15928
rect 15652 -16008 16824 -15992
rect 15652 -16072 16740 -16008
rect 16804 -16072 16824 -16008
rect 15652 -16120 16824 -16072
rect 17064 -15288 18236 -15240
rect 17064 -15352 18152 -15288
rect 18216 -15352 18236 -15288
rect 17064 -15368 18236 -15352
rect 17064 -15432 18152 -15368
rect 18216 -15432 18236 -15368
rect 17064 -15448 18236 -15432
rect 17064 -15512 18152 -15448
rect 18216 -15512 18236 -15448
rect 17064 -15528 18236 -15512
rect 17064 -15592 18152 -15528
rect 18216 -15592 18236 -15528
rect 17064 -15608 18236 -15592
rect 17064 -15672 18152 -15608
rect 18216 -15672 18236 -15608
rect 17064 -15688 18236 -15672
rect 17064 -15752 18152 -15688
rect 18216 -15752 18236 -15688
rect 17064 -15768 18236 -15752
rect 17064 -15832 18152 -15768
rect 18216 -15832 18236 -15768
rect 17064 -15848 18236 -15832
rect 17064 -15912 18152 -15848
rect 18216 -15912 18236 -15848
rect 17064 -15928 18236 -15912
rect 17064 -15992 18152 -15928
rect 18216 -15992 18236 -15928
rect 17064 -16008 18236 -15992
rect 17064 -16072 18152 -16008
rect 18216 -16072 18236 -16008
rect 17064 -16120 18236 -16072
rect 18476 -15288 19648 -15240
rect 18476 -15352 19564 -15288
rect 19628 -15352 19648 -15288
rect 18476 -15368 19648 -15352
rect 18476 -15432 19564 -15368
rect 19628 -15432 19648 -15368
rect 18476 -15448 19648 -15432
rect 18476 -15512 19564 -15448
rect 19628 -15512 19648 -15448
rect 18476 -15528 19648 -15512
rect 18476 -15592 19564 -15528
rect 19628 -15592 19648 -15528
rect 18476 -15608 19648 -15592
rect 18476 -15672 19564 -15608
rect 19628 -15672 19648 -15608
rect 18476 -15688 19648 -15672
rect 18476 -15752 19564 -15688
rect 19628 -15752 19648 -15688
rect 18476 -15768 19648 -15752
rect 18476 -15832 19564 -15768
rect 19628 -15832 19648 -15768
rect 18476 -15848 19648 -15832
rect 18476 -15912 19564 -15848
rect 19628 -15912 19648 -15848
rect 18476 -15928 19648 -15912
rect 18476 -15992 19564 -15928
rect 19628 -15992 19648 -15928
rect 18476 -16008 19648 -15992
rect 18476 -16072 19564 -16008
rect 19628 -16072 19648 -16008
rect 18476 -16120 19648 -16072
rect 19888 -15288 21060 -15240
rect 19888 -15352 20976 -15288
rect 21040 -15352 21060 -15288
rect 19888 -15368 21060 -15352
rect 19888 -15432 20976 -15368
rect 21040 -15432 21060 -15368
rect 19888 -15448 21060 -15432
rect 19888 -15512 20976 -15448
rect 21040 -15512 21060 -15448
rect 19888 -15528 21060 -15512
rect 19888 -15592 20976 -15528
rect 21040 -15592 21060 -15528
rect 19888 -15608 21060 -15592
rect 19888 -15672 20976 -15608
rect 21040 -15672 21060 -15608
rect 19888 -15688 21060 -15672
rect 19888 -15752 20976 -15688
rect 21040 -15752 21060 -15688
rect 19888 -15768 21060 -15752
rect 19888 -15832 20976 -15768
rect 21040 -15832 21060 -15768
rect 19888 -15848 21060 -15832
rect 19888 -15912 20976 -15848
rect 21040 -15912 21060 -15848
rect 19888 -15928 21060 -15912
rect 19888 -15992 20976 -15928
rect 21040 -15992 21060 -15928
rect 19888 -16008 21060 -15992
rect 19888 -16072 20976 -16008
rect 21040 -16072 21060 -16008
rect 19888 -16120 21060 -16072
rect 21300 -15288 22472 -15240
rect 21300 -15352 22388 -15288
rect 22452 -15352 22472 -15288
rect 21300 -15368 22472 -15352
rect 21300 -15432 22388 -15368
rect 22452 -15432 22472 -15368
rect 21300 -15448 22472 -15432
rect 21300 -15512 22388 -15448
rect 22452 -15512 22472 -15448
rect 21300 -15528 22472 -15512
rect 21300 -15592 22388 -15528
rect 22452 -15592 22472 -15528
rect 21300 -15608 22472 -15592
rect 21300 -15672 22388 -15608
rect 22452 -15672 22472 -15608
rect 21300 -15688 22472 -15672
rect 21300 -15752 22388 -15688
rect 22452 -15752 22472 -15688
rect 21300 -15768 22472 -15752
rect 21300 -15832 22388 -15768
rect 22452 -15832 22472 -15768
rect 21300 -15848 22472 -15832
rect 21300 -15912 22388 -15848
rect 22452 -15912 22472 -15848
rect 21300 -15928 22472 -15912
rect 21300 -15992 22388 -15928
rect 22452 -15992 22472 -15928
rect 21300 -16008 22472 -15992
rect 21300 -16072 22388 -16008
rect 22452 -16072 22472 -16008
rect 21300 -16120 22472 -16072
rect 22712 -15288 23884 -15240
rect 22712 -15352 23800 -15288
rect 23864 -15352 23884 -15288
rect 22712 -15368 23884 -15352
rect 22712 -15432 23800 -15368
rect 23864 -15432 23884 -15368
rect 22712 -15448 23884 -15432
rect 22712 -15512 23800 -15448
rect 23864 -15512 23884 -15448
rect 22712 -15528 23884 -15512
rect 22712 -15592 23800 -15528
rect 23864 -15592 23884 -15528
rect 22712 -15608 23884 -15592
rect 22712 -15672 23800 -15608
rect 23864 -15672 23884 -15608
rect 22712 -15688 23884 -15672
rect 22712 -15752 23800 -15688
rect 23864 -15752 23884 -15688
rect 22712 -15768 23884 -15752
rect 22712 -15832 23800 -15768
rect 23864 -15832 23884 -15768
rect 22712 -15848 23884 -15832
rect 22712 -15912 23800 -15848
rect 23864 -15912 23884 -15848
rect 22712 -15928 23884 -15912
rect 22712 -15992 23800 -15928
rect 23864 -15992 23884 -15928
rect 22712 -16008 23884 -15992
rect 22712 -16072 23800 -16008
rect 23864 -16072 23884 -16008
rect 22712 -16120 23884 -16072
rect -23884 -16408 -22712 -16360
rect -23884 -16472 -22796 -16408
rect -22732 -16472 -22712 -16408
rect -23884 -16488 -22712 -16472
rect -23884 -16552 -22796 -16488
rect -22732 -16552 -22712 -16488
rect -23884 -16568 -22712 -16552
rect -23884 -16632 -22796 -16568
rect -22732 -16632 -22712 -16568
rect -23884 -16648 -22712 -16632
rect -23884 -16712 -22796 -16648
rect -22732 -16712 -22712 -16648
rect -23884 -16728 -22712 -16712
rect -23884 -16792 -22796 -16728
rect -22732 -16792 -22712 -16728
rect -23884 -16808 -22712 -16792
rect -23884 -16872 -22796 -16808
rect -22732 -16872 -22712 -16808
rect -23884 -16888 -22712 -16872
rect -23884 -16952 -22796 -16888
rect -22732 -16952 -22712 -16888
rect -23884 -16968 -22712 -16952
rect -23884 -17032 -22796 -16968
rect -22732 -17032 -22712 -16968
rect -23884 -17048 -22712 -17032
rect -23884 -17112 -22796 -17048
rect -22732 -17112 -22712 -17048
rect -23884 -17128 -22712 -17112
rect -23884 -17192 -22796 -17128
rect -22732 -17192 -22712 -17128
rect -23884 -17240 -22712 -17192
rect -22472 -16408 -21300 -16360
rect -22472 -16472 -21384 -16408
rect -21320 -16472 -21300 -16408
rect -22472 -16488 -21300 -16472
rect -22472 -16552 -21384 -16488
rect -21320 -16552 -21300 -16488
rect -22472 -16568 -21300 -16552
rect -22472 -16632 -21384 -16568
rect -21320 -16632 -21300 -16568
rect -22472 -16648 -21300 -16632
rect -22472 -16712 -21384 -16648
rect -21320 -16712 -21300 -16648
rect -22472 -16728 -21300 -16712
rect -22472 -16792 -21384 -16728
rect -21320 -16792 -21300 -16728
rect -22472 -16808 -21300 -16792
rect -22472 -16872 -21384 -16808
rect -21320 -16872 -21300 -16808
rect -22472 -16888 -21300 -16872
rect -22472 -16952 -21384 -16888
rect -21320 -16952 -21300 -16888
rect -22472 -16968 -21300 -16952
rect -22472 -17032 -21384 -16968
rect -21320 -17032 -21300 -16968
rect -22472 -17048 -21300 -17032
rect -22472 -17112 -21384 -17048
rect -21320 -17112 -21300 -17048
rect -22472 -17128 -21300 -17112
rect -22472 -17192 -21384 -17128
rect -21320 -17192 -21300 -17128
rect -22472 -17240 -21300 -17192
rect -21060 -16408 -19888 -16360
rect -21060 -16472 -19972 -16408
rect -19908 -16472 -19888 -16408
rect -21060 -16488 -19888 -16472
rect -21060 -16552 -19972 -16488
rect -19908 -16552 -19888 -16488
rect -21060 -16568 -19888 -16552
rect -21060 -16632 -19972 -16568
rect -19908 -16632 -19888 -16568
rect -21060 -16648 -19888 -16632
rect -21060 -16712 -19972 -16648
rect -19908 -16712 -19888 -16648
rect -21060 -16728 -19888 -16712
rect -21060 -16792 -19972 -16728
rect -19908 -16792 -19888 -16728
rect -21060 -16808 -19888 -16792
rect -21060 -16872 -19972 -16808
rect -19908 -16872 -19888 -16808
rect -21060 -16888 -19888 -16872
rect -21060 -16952 -19972 -16888
rect -19908 -16952 -19888 -16888
rect -21060 -16968 -19888 -16952
rect -21060 -17032 -19972 -16968
rect -19908 -17032 -19888 -16968
rect -21060 -17048 -19888 -17032
rect -21060 -17112 -19972 -17048
rect -19908 -17112 -19888 -17048
rect -21060 -17128 -19888 -17112
rect -21060 -17192 -19972 -17128
rect -19908 -17192 -19888 -17128
rect -21060 -17240 -19888 -17192
rect -19648 -16408 -18476 -16360
rect -19648 -16472 -18560 -16408
rect -18496 -16472 -18476 -16408
rect -19648 -16488 -18476 -16472
rect -19648 -16552 -18560 -16488
rect -18496 -16552 -18476 -16488
rect -19648 -16568 -18476 -16552
rect -19648 -16632 -18560 -16568
rect -18496 -16632 -18476 -16568
rect -19648 -16648 -18476 -16632
rect -19648 -16712 -18560 -16648
rect -18496 -16712 -18476 -16648
rect -19648 -16728 -18476 -16712
rect -19648 -16792 -18560 -16728
rect -18496 -16792 -18476 -16728
rect -19648 -16808 -18476 -16792
rect -19648 -16872 -18560 -16808
rect -18496 -16872 -18476 -16808
rect -19648 -16888 -18476 -16872
rect -19648 -16952 -18560 -16888
rect -18496 -16952 -18476 -16888
rect -19648 -16968 -18476 -16952
rect -19648 -17032 -18560 -16968
rect -18496 -17032 -18476 -16968
rect -19648 -17048 -18476 -17032
rect -19648 -17112 -18560 -17048
rect -18496 -17112 -18476 -17048
rect -19648 -17128 -18476 -17112
rect -19648 -17192 -18560 -17128
rect -18496 -17192 -18476 -17128
rect -19648 -17240 -18476 -17192
rect -18236 -16408 -17064 -16360
rect -18236 -16472 -17148 -16408
rect -17084 -16472 -17064 -16408
rect -18236 -16488 -17064 -16472
rect -18236 -16552 -17148 -16488
rect -17084 -16552 -17064 -16488
rect -18236 -16568 -17064 -16552
rect -18236 -16632 -17148 -16568
rect -17084 -16632 -17064 -16568
rect -18236 -16648 -17064 -16632
rect -18236 -16712 -17148 -16648
rect -17084 -16712 -17064 -16648
rect -18236 -16728 -17064 -16712
rect -18236 -16792 -17148 -16728
rect -17084 -16792 -17064 -16728
rect -18236 -16808 -17064 -16792
rect -18236 -16872 -17148 -16808
rect -17084 -16872 -17064 -16808
rect -18236 -16888 -17064 -16872
rect -18236 -16952 -17148 -16888
rect -17084 -16952 -17064 -16888
rect -18236 -16968 -17064 -16952
rect -18236 -17032 -17148 -16968
rect -17084 -17032 -17064 -16968
rect -18236 -17048 -17064 -17032
rect -18236 -17112 -17148 -17048
rect -17084 -17112 -17064 -17048
rect -18236 -17128 -17064 -17112
rect -18236 -17192 -17148 -17128
rect -17084 -17192 -17064 -17128
rect -18236 -17240 -17064 -17192
rect -16824 -16408 -15652 -16360
rect -16824 -16472 -15736 -16408
rect -15672 -16472 -15652 -16408
rect -16824 -16488 -15652 -16472
rect -16824 -16552 -15736 -16488
rect -15672 -16552 -15652 -16488
rect -16824 -16568 -15652 -16552
rect -16824 -16632 -15736 -16568
rect -15672 -16632 -15652 -16568
rect -16824 -16648 -15652 -16632
rect -16824 -16712 -15736 -16648
rect -15672 -16712 -15652 -16648
rect -16824 -16728 -15652 -16712
rect -16824 -16792 -15736 -16728
rect -15672 -16792 -15652 -16728
rect -16824 -16808 -15652 -16792
rect -16824 -16872 -15736 -16808
rect -15672 -16872 -15652 -16808
rect -16824 -16888 -15652 -16872
rect -16824 -16952 -15736 -16888
rect -15672 -16952 -15652 -16888
rect -16824 -16968 -15652 -16952
rect -16824 -17032 -15736 -16968
rect -15672 -17032 -15652 -16968
rect -16824 -17048 -15652 -17032
rect -16824 -17112 -15736 -17048
rect -15672 -17112 -15652 -17048
rect -16824 -17128 -15652 -17112
rect -16824 -17192 -15736 -17128
rect -15672 -17192 -15652 -17128
rect -16824 -17240 -15652 -17192
rect -15412 -16408 -14240 -16360
rect -15412 -16472 -14324 -16408
rect -14260 -16472 -14240 -16408
rect -15412 -16488 -14240 -16472
rect -15412 -16552 -14324 -16488
rect -14260 -16552 -14240 -16488
rect -15412 -16568 -14240 -16552
rect -15412 -16632 -14324 -16568
rect -14260 -16632 -14240 -16568
rect -15412 -16648 -14240 -16632
rect -15412 -16712 -14324 -16648
rect -14260 -16712 -14240 -16648
rect -15412 -16728 -14240 -16712
rect -15412 -16792 -14324 -16728
rect -14260 -16792 -14240 -16728
rect -15412 -16808 -14240 -16792
rect -15412 -16872 -14324 -16808
rect -14260 -16872 -14240 -16808
rect -15412 -16888 -14240 -16872
rect -15412 -16952 -14324 -16888
rect -14260 -16952 -14240 -16888
rect -15412 -16968 -14240 -16952
rect -15412 -17032 -14324 -16968
rect -14260 -17032 -14240 -16968
rect -15412 -17048 -14240 -17032
rect -15412 -17112 -14324 -17048
rect -14260 -17112 -14240 -17048
rect -15412 -17128 -14240 -17112
rect -15412 -17192 -14324 -17128
rect -14260 -17192 -14240 -17128
rect -15412 -17240 -14240 -17192
rect -14000 -16408 -12828 -16360
rect -14000 -16472 -12912 -16408
rect -12848 -16472 -12828 -16408
rect -14000 -16488 -12828 -16472
rect -14000 -16552 -12912 -16488
rect -12848 -16552 -12828 -16488
rect -14000 -16568 -12828 -16552
rect -14000 -16632 -12912 -16568
rect -12848 -16632 -12828 -16568
rect -14000 -16648 -12828 -16632
rect -14000 -16712 -12912 -16648
rect -12848 -16712 -12828 -16648
rect -14000 -16728 -12828 -16712
rect -14000 -16792 -12912 -16728
rect -12848 -16792 -12828 -16728
rect -14000 -16808 -12828 -16792
rect -14000 -16872 -12912 -16808
rect -12848 -16872 -12828 -16808
rect -14000 -16888 -12828 -16872
rect -14000 -16952 -12912 -16888
rect -12848 -16952 -12828 -16888
rect -14000 -16968 -12828 -16952
rect -14000 -17032 -12912 -16968
rect -12848 -17032 -12828 -16968
rect -14000 -17048 -12828 -17032
rect -14000 -17112 -12912 -17048
rect -12848 -17112 -12828 -17048
rect -14000 -17128 -12828 -17112
rect -14000 -17192 -12912 -17128
rect -12848 -17192 -12828 -17128
rect -14000 -17240 -12828 -17192
rect -12588 -16408 -11416 -16360
rect -12588 -16472 -11500 -16408
rect -11436 -16472 -11416 -16408
rect -12588 -16488 -11416 -16472
rect -12588 -16552 -11500 -16488
rect -11436 -16552 -11416 -16488
rect -12588 -16568 -11416 -16552
rect -12588 -16632 -11500 -16568
rect -11436 -16632 -11416 -16568
rect -12588 -16648 -11416 -16632
rect -12588 -16712 -11500 -16648
rect -11436 -16712 -11416 -16648
rect -12588 -16728 -11416 -16712
rect -12588 -16792 -11500 -16728
rect -11436 -16792 -11416 -16728
rect -12588 -16808 -11416 -16792
rect -12588 -16872 -11500 -16808
rect -11436 -16872 -11416 -16808
rect -12588 -16888 -11416 -16872
rect -12588 -16952 -11500 -16888
rect -11436 -16952 -11416 -16888
rect -12588 -16968 -11416 -16952
rect -12588 -17032 -11500 -16968
rect -11436 -17032 -11416 -16968
rect -12588 -17048 -11416 -17032
rect -12588 -17112 -11500 -17048
rect -11436 -17112 -11416 -17048
rect -12588 -17128 -11416 -17112
rect -12588 -17192 -11500 -17128
rect -11436 -17192 -11416 -17128
rect -12588 -17240 -11416 -17192
rect -11176 -16408 -10004 -16360
rect -11176 -16472 -10088 -16408
rect -10024 -16472 -10004 -16408
rect -11176 -16488 -10004 -16472
rect -11176 -16552 -10088 -16488
rect -10024 -16552 -10004 -16488
rect -11176 -16568 -10004 -16552
rect -11176 -16632 -10088 -16568
rect -10024 -16632 -10004 -16568
rect -11176 -16648 -10004 -16632
rect -11176 -16712 -10088 -16648
rect -10024 -16712 -10004 -16648
rect -11176 -16728 -10004 -16712
rect -11176 -16792 -10088 -16728
rect -10024 -16792 -10004 -16728
rect -11176 -16808 -10004 -16792
rect -11176 -16872 -10088 -16808
rect -10024 -16872 -10004 -16808
rect -11176 -16888 -10004 -16872
rect -11176 -16952 -10088 -16888
rect -10024 -16952 -10004 -16888
rect -11176 -16968 -10004 -16952
rect -11176 -17032 -10088 -16968
rect -10024 -17032 -10004 -16968
rect -11176 -17048 -10004 -17032
rect -11176 -17112 -10088 -17048
rect -10024 -17112 -10004 -17048
rect -11176 -17128 -10004 -17112
rect -11176 -17192 -10088 -17128
rect -10024 -17192 -10004 -17128
rect -11176 -17240 -10004 -17192
rect -9764 -16408 -8592 -16360
rect -9764 -16472 -8676 -16408
rect -8612 -16472 -8592 -16408
rect -9764 -16488 -8592 -16472
rect -9764 -16552 -8676 -16488
rect -8612 -16552 -8592 -16488
rect -9764 -16568 -8592 -16552
rect -9764 -16632 -8676 -16568
rect -8612 -16632 -8592 -16568
rect -9764 -16648 -8592 -16632
rect -9764 -16712 -8676 -16648
rect -8612 -16712 -8592 -16648
rect -9764 -16728 -8592 -16712
rect -9764 -16792 -8676 -16728
rect -8612 -16792 -8592 -16728
rect -9764 -16808 -8592 -16792
rect -9764 -16872 -8676 -16808
rect -8612 -16872 -8592 -16808
rect -9764 -16888 -8592 -16872
rect -9764 -16952 -8676 -16888
rect -8612 -16952 -8592 -16888
rect -9764 -16968 -8592 -16952
rect -9764 -17032 -8676 -16968
rect -8612 -17032 -8592 -16968
rect -9764 -17048 -8592 -17032
rect -9764 -17112 -8676 -17048
rect -8612 -17112 -8592 -17048
rect -9764 -17128 -8592 -17112
rect -9764 -17192 -8676 -17128
rect -8612 -17192 -8592 -17128
rect -9764 -17240 -8592 -17192
rect -8352 -16408 -7180 -16360
rect -8352 -16472 -7264 -16408
rect -7200 -16472 -7180 -16408
rect -8352 -16488 -7180 -16472
rect -8352 -16552 -7264 -16488
rect -7200 -16552 -7180 -16488
rect -8352 -16568 -7180 -16552
rect -8352 -16632 -7264 -16568
rect -7200 -16632 -7180 -16568
rect -8352 -16648 -7180 -16632
rect -8352 -16712 -7264 -16648
rect -7200 -16712 -7180 -16648
rect -8352 -16728 -7180 -16712
rect -8352 -16792 -7264 -16728
rect -7200 -16792 -7180 -16728
rect -8352 -16808 -7180 -16792
rect -8352 -16872 -7264 -16808
rect -7200 -16872 -7180 -16808
rect -8352 -16888 -7180 -16872
rect -8352 -16952 -7264 -16888
rect -7200 -16952 -7180 -16888
rect -8352 -16968 -7180 -16952
rect -8352 -17032 -7264 -16968
rect -7200 -17032 -7180 -16968
rect -8352 -17048 -7180 -17032
rect -8352 -17112 -7264 -17048
rect -7200 -17112 -7180 -17048
rect -8352 -17128 -7180 -17112
rect -8352 -17192 -7264 -17128
rect -7200 -17192 -7180 -17128
rect -8352 -17240 -7180 -17192
rect -6940 -16408 -5768 -16360
rect -6940 -16472 -5852 -16408
rect -5788 -16472 -5768 -16408
rect -6940 -16488 -5768 -16472
rect -6940 -16552 -5852 -16488
rect -5788 -16552 -5768 -16488
rect -6940 -16568 -5768 -16552
rect -6940 -16632 -5852 -16568
rect -5788 -16632 -5768 -16568
rect -6940 -16648 -5768 -16632
rect -6940 -16712 -5852 -16648
rect -5788 -16712 -5768 -16648
rect -6940 -16728 -5768 -16712
rect -6940 -16792 -5852 -16728
rect -5788 -16792 -5768 -16728
rect -6940 -16808 -5768 -16792
rect -6940 -16872 -5852 -16808
rect -5788 -16872 -5768 -16808
rect -6940 -16888 -5768 -16872
rect -6940 -16952 -5852 -16888
rect -5788 -16952 -5768 -16888
rect -6940 -16968 -5768 -16952
rect -6940 -17032 -5852 -16968
rect -5788 -17032 -5768 -16968
rect -6940 -17048 -5768 -17032
rect -6940 -17112 -5852 -17048
rect -5788 -17112 -5768 -17048
rect -6940 -17128 -5768 -17112
rect -6940 -17192 -5852 -17128
rect -5788 -17192 -5768 -17128
rect -6940 -17240 -5768 -17192
rect -5528 -16408 -4356 -16360
rect -5528 -16472 -4440 -16408
rect -4376 -16472 -4356 -16408
rect -5528 -16488 -4356 -16472
rect -5528 -16552 -4440 -16488
rect -4376 -16552 -4356 -16488
rect -5528 -16568 -4356 -16552
rect -5528 -16632 -4440 -16568
rect -4376 -16632 -4356 -16568
rect -5528 -16648 -4356 -16632
rect -5528 -16712 -4440 -16648
rect -4376 -16712 -4356 -16648
rect -5528 -16728 -4356 -16712
rect -5528 -16792 -4440 -16728
rect -4376 -16792 -4356 -16728
rect -5528 -16808 -4356 -16792
rect -5528 -16872 -4440 -16808
rect -4376 -16872 -4356 -16808
rect -5528 -16888 -4356 -16872
rect -5528 -16952 -4440 -16888
rect -4376 -16952 -4356 -16888
rect -5528 -16968 -4356 -16952
rect -5528 -17032 -4440 -16968
rect -4376 -17032 -4356 -16968
rect -5528 -17048 -4356 -17032
rect -5528 -17112 -4440 -17048
rect -4376 -17112 -4356 -17048
rect -5528 -17128 -4356 -17112
rect -5528 -17192 -4440 -17128
rect -4376 -17192 -4356 -17128
rect -5528 -17240 -4356 -17192
rect -4116 -16408 -2944 -16360
rect -4116 -16472 -3028 -16408
rect -2964 -16472 -2944 -16408
rect -4116 -16488 -2944 -16472
rect -4116 -16552 -3028 -16488
rect -2964 -16552 -2944 -16488
rect -4116 -16568 -2944 -16552
rect -4116 -16632 -3028 -16568
rect -2964 -16632 -2944 -16568
rect -4116 -16648 -2944 -16632
rect -4116 -16712 -3028 -16648
rect -2964 -16712 -2944 -16648
rect -4116 -16728 -2944 -16712
rect -4116 -16792 -3028 -16728
rect -2964 -16792 -2944 -16728
rect -4116 -16808 -2944 -16792
rect -4116 -16872 -3028 -16808
rect -2964 -16872 -2944 -16808
rect -4116 -16888 -2944 -16872
rect -4116 -16952 -3028 -16888
rect -2964 -16952 -2944 -16888
rect -4116 -16968 -2944 -16952
rect -4116 -17032 -3028 -16968
rect -2964 -17032 -2944 -16968
rect -4116 -17048 -2944 -17032
rect -4116 -17112 -3028 -17048
rect -2964 -17112 -2944 -17048
rect -4116 -17128 -2944 -17112
rect -4116 -17192 -3028 -17128
rect -2964 -17192 -2944 -17128
rect -4116 -17240 -2944 -17192
rect -2704 -16408 -1532 -16360
rect -2704 -16472 -1616 -16408
rect -1552 -16472 -1532 -16408
rect -2704 -16488 -1532 -16472
rect -2704 -16552 -1616 -16488
rect -1552 -16552 -1532 -16488
rect -2704 -16568 -1532 -16552
rect -2704 -16632 -1616 -16568
rect -1552 -16632 -1532 -16568
rect -2704 -16648 -1532 -16632
rect -2704 -16712 -1616 -16648
rect -1552 -16712 -1532 -16648
rect -2704 -16728 -1532 -16712
rect -2704 -16792 -1616 -16728
rect -1552 -16792 -1532 -16728
rect -2704 -16808 -1532 -16792
rect -2704 -16872 -1616 -16808
rect -1552 -16872 -1532 -16808
rect -2704 -16888 -1532 -16872
rect -2704 -16952 -1616 -16888
rect -1552 -16952 -1532 -16888
rect -2704 -16968 -1532 -16952
rect -2704 -17032 -1616 -16968
rect -1552 -17032 -1532 -16968
rect -2704 -17048 -1532 -17032
rect -2704 -17112 -1616 -17048
rect -1552 -17112 -1532 -17048
rect -2704 -17128 -1532 -17112
rect -2704 -17192 -1616 -17128
rect -1552 -17192 -1532 -17128
rect -2704 -17240 -1532 -17192
rect -1292 -16408 -120 -16360
rect -1292 -16472 -204 -16408
rect -140 -16472 -120 -16408
rect -1292 -16488 -120 -16472
rect -1292 -16552 -204 -16488
rect -140 -16552 -120 -16488
rect -1292 -16568 -120 -16552
rect -1292 -16632 -204 -16568
rect -140 -16632 -120 -16568
rect -1292 -16648 -120 -16632
rect -1292 -16712 -204 -16648
rect -140 -16712 -120 -16648
rect -1292 -16728 -120 -16712
rect -1292 -16792 -204 -16728
rect -140 -16792 -120 -16728
rect -1292 -16808 -120 -16792
rect -1292 -16872 -204 -16808
rect -140 -16872 -120 -16808
rect -1292 -16888 -120 -16872
rect -1292 -16952 -204 -16888
rect -140 -16952 -120 -16888
rect -1292 -16968 -120 -16952
rect -1292 -17032 -204 -16968
rect -140 -17032 -120 -16968
rect -1292 -17048 -120 -17032
rect -1292 -17112 -204 -17048
rect -140 -17112 -120 -17048
rect -1292 -17128 -120 -17112
rect -1292 -17192 -204 -17128
rect -140 -17192 -120 -17128
rect -1292 -17240 -120 -17192
rect 120 -16408 1292 -16360
rect 120 -16472 1208 -16408
rect 1272 -16472 1292 -16408
rect 120 -16488 1292 -16472
rect 120 -16552 1208 -16488
rect 1272 -16552 1292 -16488
rect 120 -16568 1292 -16552
rect 120 -16632 1208 -16568
rect 1272 -16632 1292 -16568
rect 120 -16648 1292 -16632
rect 120 -16712 1208 -16648
rect 1272 -16712 1292 -16648
rect 120 -16728 1292 -16712
rect 120 -16792 1208 -16728
rect 1272 -16792 1292 -16728
rect 120 -16808 1292 -16792
rect 120 -16872 1208 -16808
rect 1272 -16872 1292 -16808
rect 120 -16888 1292 -16872
rect 120 -16952 1208 -16888
rect 1272 -16952 1292 -16888
rect 120 -16968 1292 -16952
rect 120 -17032 1208 -16968
rect 1272 -17032 1292 -16968
rect 120 -17048 1292 -17032
rect 120 -17112 1208 -17048
rect 1272 -17112 1292 -17048
rect 120 -17128 1292 -17112
rect 120 -17192 1208 -17128
rect 1272 -17192 1292 -17128
rect 120 -17240 1292 -17192
rect 1532 -16408 2704 -16360
rect 1532 -16472 2620 -16408
rect 2684 -16472 2704 -16408
rect 1532 -16488 2704 -16472
rect 1532 -16552 2620 -16488
rect 2684 -16552 2704 -16488
rect 1532 -16568 2704 -16552
rect 1532 -16632 2620 -16568
rect 2684 -16632 2704 -16568
rect 1532 -16648 2704 -16632
rect 1532 -16712 2620 -16648
rect 2684 -16712 2704 -16648
rect 1532 -16728 2704 -16712
rect 1532 -16792 2620 -16728
rect 2684 -16792 2704 -16728
rect 1532 -16808 2704 -16792
rect 1532 -16872 2620 -16808
rect 2684 -16872 2704 -16808
rect 1532 -16888 2704 -16872
rect 1532 -16952 2620 -16888
rect 2684 -16952 2704 -16888
rect 1532 -16968 2704 -16952
rect 1532 -17032 2620 -16968
rect 2684 -17032 2704 -16968
rect 1532 -17048 2704 -17032
rect 1532 -17112 2620 -17048
rect 2684 -17112 2704 -17048
rect 1532 -17128 2704 -17112
rect 1532 -17192 2620 -17128
rect 2684 -17192 2704 -17128
rect 1532 -17240 2704 -17192
rect 2944 -16408 4116 -16360
rect 2944 -16472 4032 -16408
rect 4096 -16472 4116 -16408
rect 2944 -16488 4116 -16472
rect 2944 -16552 4032 -16488
rect 4096 -16552 4116 -16488
rect 2944 -16568 4116 -16552
rect 2944 -16632 4032 -16568
rect 4096 -16632 4116 -16568
rect 2944 -16648 4116 -16632
rect 2944 -16712 4032 -16648
rect 4096 -16712 4116 -16648
rect 2944 -16728 4116 -16712
rect 2944 -16792 4032 -16728
rect 4096 -16792 4116 -16728
rect 2944 -16808 4116 -16792
rect 2944 -16872 4032 -16808
rect 4096 -16872 4116 -16808
rect 2944 -16888 4116 -16872
rect 2944 -16952 4032 -16888
rect 4096 -16952 4116 -16888
rect 2944 -16968 4116 -16952
rect 2944 -17032 4032 -16968
rect 4096 -17032 4116 -16968
rect 2944 -17048 4116 -17032
rect 2944 -17112 4032 -17048
rect 4096 -17112 4116 -17048
rect 2944 -17128 4116 -17112
rect 2944 -17192 4032 -17128
rect 4096 -17192 4116 -17128
rect 2944 -17240 4116 -17192
rect 4356 -16408 5528 -16360
rect 4356 -16472 5444 -16408
rect 5508 -16472 5528 -16408
rect 4356 -16488 5528 -16472
rect 4356 -16552 5444 -16488
rect 5508 -16552 5528 -16488
rect 4356 -16568 5528 -16552
rect 4356 -16632 5444 -16568
rect 5508 -16632 5528 -16568
rect 4356 -16648 5528 -16632
rect 4356 -16712 5444 -16648
rect 5508 -16712 5528 -16648
rect 4356 -16728 5528 -16712
rect 4356 -16792 5444 -16728
rect 5508 -16792 5528 -16728
rect 4356 -16808 5528 -16792
rect 4356 -16872 5444 -16808
rect 5508 -16872 5528 -16808
rect 4356 -16888 5528 -16872
rect 4356 -16952 5444 -16888
rect 5508 -16952 5528 -16888
rect 4356 -16968 5528 -16952
rect 4356 -17032 5444 -16968
rect 5508 -17032 5528 -16968
rect 4356 -17048 5528 -17032
rect 4356 -17112 5444 -17048
rect 5508 -17112 5528 -17048
rect 4356 -17128 5528 -17112
rect 4356 -17192 5444 -17128
rect 5508 -17192 5528 -17128
rect 4356 -17240 5528 -17192
rect 5768 -16408 6940 -16360
rect 5768 -16472 6856 -16408
rect 6920 -16472 6940 -16408
rect 5768 -16488 6940 -16472
rect 5768 -16552 6856 -16488
rect 6920 -16552 6940 -16488
rect 5768 -16568 6940 -16552
rect 5768 -16632 6856 -16568
rect 6920 -16632 6940 -16568
rect 5768 -16648 6940 -16632
rect 5768 -16712 6856 -16648
rect 6920 -16712 6940 -16648
rect 5768 -16728 6940 -16712
rect 5768 -16792 6856 -16728
rect 6920 -16792 6940 -16728
rect 5768 -16808 6940 -16792
rect 5768 -16872 6856 -16808
rect 6920 -16872 6940 -16808
rect 5768 -16888 6940 -16872
rect 5768 -16952 6856 -16888
rect 6920 -16952 6940 -16888
rect 5768 -16968 6940 -16952
rect 5768 -17032 6856 -16968
rect 6920 -17032 6940 -16968
rect 5768 -17048 6940 -17032
rect 5768 -17112 6856 -17048
rect 6920 -17112 6940 -17048
rect 5768 -17128 6940 -17112
rect 5768 -17192 6856 -17128
rect 6920 -17192 6940 -17128
rect 5768 -17240 6940 -17192
rect 7180 -16408 8352 -16360
rect 7180 -16472 8268 -16408
rect 8332 -16472 8352 -16408
rect 7180 -16488 8352 -16472
rect 7180 -16552 8268 -16488
rect 8332 -16552 8352 -16488
rect 7180 -16568 8352 -16552
rect 7180 -16632 8268 -16568
rect 8332 -16632 8352 -16568
rect 7180 -16648 8352 -16632
rect 7180 -16712 8268 -16648
rect 8332 -16712 8352 -16648
rect 7180 -16728 8352 -16712
rect 7180 -16792 8268 -16728
rect 8332 -16792 8352 -16728
rect 7180 -16808 8352 -16792
rect 7180 -16872 8268 -16808
rect 8332 -16872 8352 -16808
rect 7180 -16888 8352 -16872
rect 7180 -16952 8268 -16888
rect 8332 -16952 8352 -16888
rect 7180 -16968 8352 -16952
rect 7180 -17032 8268 -16968
rect 8332 -17032 8352 -16968
rect 7180 -17048 8352 -17032
rect 7180 -17112 8268 -17048
rect 8332 -17112 8352 -17048
rect 7180 -17128 8352 -17112
rect 7180 -17192 8268 -17128
rect 8332 -17192 8352 -17128
rect 7180 -17240 8352 -17192
rect 8592 -16408 9764 -16360
rect 8592 -16472 9680 -16408
rect 9744 -16472 9764 -16408
rect 8592 -16488 9764 -16472
rect 8592 -16552 9680 -16488
rect 9744 -16552 9764 -16488
rect 8592 -16568 9764 -16552
rect 8592 -16632 9680 -16568
rect 9744 -16632 9764 -16568
rect 8592 -16648 9764 -16632
rect 8592 -16712 9680 -16648
rect 9744 -16712 9764 -16648
rect 8592 -16728 9764 -16712
rect 8592 -16792 9680 -16728
rect 9744 -16792 9764 -16728
rect 8592 -16808 9764 -16792
rect 8592 -16872 9680 -16808
rect 9744 -16872 9764 -16808
rect 8592 -16888 9764 -16872
rect 8592 -16952 9680 -16888
rect 9744 -16952 9764 -16888
rect 8592 -16968 9764 -16952
rect 8592 -17032 9680 -16968
rect 9744 -17032 9764 -16968
rect 8592 -17048 9764 -17032
rect 8592 -17112 9680 -17048
rect 9744 -17112 9764 -17048
rect 8592 -17128 9764 -17112
rect 8592 -17192 9680 -17128
rect 9744 -17192 9764 -17128
rect 8592 -17240 9764 -17192
rect 10004 -16408 11176 -16360
rect 10004 -16472 11092 -16408
rect 11156 -16472 11176 -16408
rect 10004 -16488 11176 -16472
rect 10004 -16552 11092 -16488
rect 11156 -16552 11176 -16488
rect 10004 -16568 11176 -16552
rect 10004 -16632 11092 -16568
rect 11156 -16632 11176 -16568
rect 10004 -16648 11176 -16632
rect 10004 -16712 11092 -16648
rect 11156 -16712 11176 -16648
rect 10004 -16728 11176 -16712
rect 10004 -16792 11092 -16728
rect 11156 -16792 11176 -16728
rect 10004 -16808 11176 -16792
rect 10004 -16872 11092 -16808
rect 11156 -16872 11176 -16808
rect 10004 -16888 11176 -16872
rect 10004 -16952 11092 -16888
rect 11156 -16952 11176 -16888
rect 10004 -16968 11176 -16952
rect 10004 -17032 11092 -16968
rect 11156 -17032 11176 -16968
rect 10004 -17048 11176 -17032
rect 10004 -17112 11092 -17048
rect 11156 -17112 11176 -17048
rect 10004 -17128 11176 -17112
rect 10004 -17192 11092 -17128
rect 11156 -17192 11176 -17128
rect 10004 -17240 11176 -17192
rect 11416 -16408 12588 -16360
rect 11416 -16472 12504 -16408
rect 12568 -16472 12588 -16408
rect 11416 -16488 12588 -16472
rect 11416 -16552 12504 -16488
rect 12568 -16552 12588 -16488
rect 11416 -16568 12588 -16552
rect 11416 -16632 12504 -16568
rect 12568 -16632 12588 -16568
rect 11416 -16648 12588 -16632
rect 11416 -16712 12504 -16648
rect 12568 -16712 12588 -16648
rect 11416 -16728 12588 -16712
rect 11416 -16792 12504 -16728
rect 12568 -16792 12588 -16728
rect 11416 -16808 12588 -16792
rect 11416 -16872 12504 -16808
rect 12568 -16872 12588 -16808
rect 11416 -16888 12588 -16872
rect 11416 -16952 12504 -16888
rect 12568 -16952 12588 -16888
rect 11416 -16968 12588 -16952
rect 11416 -17032 12504 -16968
rect 12568 -17032 12588 -16968
rect 11416 -17048 12588 -17032
rect 11416 -17112 12504 -17048
rect 12568 -17112 12588 -17048
rect 11416 -17128 12588 -17112
rect 11416 -17192 12504 -17128
rect 12568 -17192 12588 -17128
rect 11416 -17240 12588 -17192
rect 12828 -16408 14000 -16360
rect 12828 -16472 13916 -16408
rect 13980 -16472 14000 -16408
rect 12828 -16488 14000 -16472
rect 12828 -16552 13916 -16488
rect 13980 -16552 14000 -16488
rect 12828 -16568 14000 -16552
rect 12828 -16632 13916 -16568
rect 13980 -16632 14000 -16568
rect 12828 -16648 14000 -16632
rect 12828 -16712 13916 -16648
rect 13980 -16712 14000 -16648
rect 12828 -16728 14000 -16712
rect 12828 -16792 13916 -16728
rect 13980 -16792 14000 -16728
rect 12828 -16808 14000 -16792
rect 12828 -16872 13916 -16808
rect 13980 -16872 14000 -16808
rect 12828 -16888 14000 -16872
rect 12828 -16952 13916 -16888
rect 13980 -16952 14000 -16888
rect 12828 -16968 14000 -16952
rect 12828 -17032 13916 -16968
rect 13980 -17032 14000 -16968
rect 12828 -17048 14000 -17032
rect 12828 -17112 13916 -17048
rect 13980 -17112 14000 -17048
rect 12828 -17128 14000 -17112
rect 12828 -17192 13916 -17128
rect 13980 -17192 14000 -17128
rect 12828 -17240 14000 -17192
rect 14240 -16408 15412 -16360
rect 14240 -16472 15328 -16408
rect 15392 -16472 15412 -16408
rect 14240 -16488 15412 -16472
rect 14240 -16552 15328 -16488
rect 15392 -16552 15412 -16488
rect 14240 -16568 15412 -16552
rect 14240 -16632 15328 -16568
rect 15392 -16632 15412 -16568
rect 14240 -16648 15412 -16632
rect 14240 -16712 15328 -16648
rect 15392 -16712 15412 -16648
rect 14240 -16728 15412 -16712
rect 14240 -16792 15328 -16728
rect 15392 -16792 15412 -16728
rect 14240 -16808 15412 -16792
rect 14240 -16872 15328 -16808
rect 15392 -16872 15412 -16808
rect 14240 -16888 15412 -16872
rect 14240 -16952 15328 -16888
rect 15392 -16952 15412 -16888
rect 14240 -16968 15412 -16952
rect 14240 -17032 15328 -16968
rect 15392 -17032 15412 -16968
rect 14240 -17048 15412 -17032
rect 14240 -17112 15328 -17048
rect 15392 -17112 15412 -17048
rect 14240 -17128 15412 -17112
rect 14240 -17192 15328 -17128
rect 15392 -17192 15412 -17128
rect 14240 -17240 15412 -17192
rect 15652 -16408 16824 -16360
rect 15652 -16472 16740 -16408
rect 16804 -16472 16824 -16408
rect 15652 -16488 16824 -16472
rect 15652 -16552 16740 -16488
rect 16804 -16552 16824 -16488
rect 15652 -16568 16824 -16552
rect 15652 -16632 16740 -16568
rect 16804 -16632 16824 -16568
rect 15652 -16648 16824 -16632
rect 15652 -16712 16740 -16648
rect 16804 -16712 16824 -16648
rect 15652 -16728 16824 -16712
rect 15652 -16792 16740 -16728
rect 16804 -16792 16824 -16728
rect 15652 -16808 16824 -16792
rect 15652 -16872 16740 -16808
rect 16804 -16872 16824 -16808
rect 15652 -16888 16824 -16872
rect 15652 -16952 16740 -16888
rect 16804 -16952 16824 -16888
rect 15652 -16968 16824 -16952
rect 15652 -17032 16740 -16968
rect 16804 -17032 16824 -16968
rect 15652 -17048 16824 -17032
rect 15652 -17112 16740 -17048
rect 16804 -17112 16824 -17048
rect 15652 -17128 16824 -17112
rect 15652 -17192 16740 -17128
rect 16804 -17192 16824 -17128
rect 15652 -17240 16824 -17192
rect 17064 -16408 18236 -16360
rect 17064 -16472 18152 -16408
rect 18216 -16472 18236 -16408
rect 17064 -16488 18236 -16472
rect 17064 -16552 18152 -16488
rect 18216 -16552 18236 -16488
rect 17064 -16568 18236 -16552
rect 17064 -16632 18152 -16568
rect 18216 -16632 18236 -16568
rect 17064 -16648 18236 -16632
rect 17064 -16712 18152 -16648
rect 18216 -16712 18236 -16648
rect 17064 -16728 18236 -16712
rect 17064 -16792 18152 -16728
rect 18216 -16792 18236 -16728
rect 17064 -16808 18236 -16792
rect 17064 -16872 18152 -16808
rect 18216 -16872 18236 -16808
rect 17064 -16888 18236 -16872
rect 17064 -16952 18152 -16888
rect 18216 -16952 18236 -16888
rect 17064 -16968 18236 -16952
rect 17064 -17032 18152 -16968
rect 18216 -17032 18236 -16968
rect 17064 -17048 18236 -17032
rect 17064 -17112 18152 -17048
rect 18216 -17112 18236 -17048
rect 17064 -17128 18236 -17112
rect 17064 -17192 18152 -17128
rect 18216 -17192 18236 -17128
rect 17064 -17240 18236 -17192
rect 18476 -16408 19648 -16360
rect 18476 -16472 19564 -16408
rect 19628 -16472 19648 -16408
rect 18476 -16488 19648 -16472
rect 18476 -16552 19564 -16488
rect 19628 -16552 19648 -16488
rect 18476 -16568 19648 -16552
rect 18476 -16632 19564 -16568
rect 19628 -16632 19648 -16568
rect 18476 -16648 19648 -16632
rect 18476 -16712 19564 -16648
rect 19628 -16712 19648 -16648
rect 18476 -16728 19648 -16712
rect 18476 -16792 19564 -16728
rect 19628 -16792 19648 -16728
rect 18476 -16808 19648 -16792
rect 18476 -16872 19564 -16808
rect 19628 -16872 19648 -16808
rect 18476 -16888 19648 -16872
rect 18476 -16952 19564 -16888
rect 19628 -16952 19648 -16888
rect 18476 -16968 19648 -16952
rect 18476 -17032 19564 -16968
rect 19628 -17032 19648 -16968
rect 18476 -17048 19648 -17032
rect 18476 -17112 19564 -17048
rect 19628 -17112 19648 -17048
rect 18476 -17128 19648 -17112
rect 18476 -17192 19564 -17128
rect 19628 -17192 19648 -17128
rect 18476 -17240 19648 -17192
rect 19888 -16408 21060 -16360
rect 19888 -16472 20976 -16408
rect 21040 -16472 21060 -16408
rect 19888 -16488 21060 -16472
rect 19888 -16552 20976 -16488
rect 21040 -16552 21060 -16488
rect 19888 -16568 21060 -16552
rect 19888 -16632 20976 -16568
rect 21040 -16632 21060 -16568
rect 19888 -16648 21060 -16632
rect 19888 -16712 20976 -16648
rect 21040 -16712 21060 -16648
rect 19888 -16728 21060 -16712
rect 19888 -16792 20976 -16728
rect 21040 -16792 21060 -16728
rect 19888 -16808 21060 -16792
rect 19888 -16872 20976 -16808
rect 21040 -16872 21060 -16808
rect 19888 -16888 21060 -16872
rect 19888 -16952 20976 -16888
rect 21040 -16952 21060 -16888
rect 19888 -16968 21060 -16952
rect 19888 -17032 20976 -16968
rect 21040 -17032 21060 -16968
rect 19888 -17048 21060 -17032
rect 19888 -17112 20976 -17048
rect 21040 -17112 21060 -17048
rect 19888 -17128 21060 -17112
rect 19888 -17192 20976 -17128
rect 21040 -17192 21060 -17128
rect 19888 -17240 21060 -17192
rect 21300 -16408 22472 -16360
rect 21300 -16472 22388 -16408
rect 22452 -16472 22472 -16408
rect 21300 -16488 22472 -16472
rect 21300 -16552 22388 -16488
rect 22452 -16552 22472 -16488
rect 21300 -16568 22472 -16552
rect 21300 -16632 22388 -16568
rect 22452 -16632 22472 -16568
rect 21300 -16648 22472 -16632
rect 21300 -16712 22388 -16648
rect 22452 -16712 22472 -16648
rect 21300 -16728 22472 -16712
rect 21300 -16792 22388 -16728
rect 22452 -16792 22472 -16728
rect 21300 -16808 22472 -16792
rect 21300 -16872 22388 -16808
rect 22452 -16872 22472 -16808
rect 21300 -16888 22472 -16872
rect 21300 -16952 22388 -16888
rect 22452 -16952 22472 -16888
rect 21300 -16968 22472 -16952
rect 21300 -17032 22388 -16968
rect 22452 -17032 22472 -16968
rect 21300 -17048 22472 -17032
rect 21300 -17112 22388 -17048
rect 22452 -17112 22472 -17048
rect 21300 -17128 22472 -17112
rect 21300 -17192 22388 -17128
rect 22452 -17192 22472 -17128
rect 21300 -17240 22472 -17192
rect 22712 -16408 23884 -16360
rect 22712 -16472 23800 -16408
rect 23864 -16472 23884 -16408
rect 22712 -16488 23884 -16472
rect 22712 -16552 23800 -16488
rect 23864 -16552 23884 -16488
rect 22712 -16568 23884 -16552
rect 22712 -16632 23800 -16568
rect 23864 -16632 23884 -16568
rect 22712 -16648 23884 -16632
rect 22712 -16712 23800 -16648
rect 23864 -16712 23884 -16648
rect 22712 -16728 23884 -16712
rect 22712 -16792 23800 -16728
rect 23864 -16792 23884 -16728
rect 22712 -16808 23884 -16792
rect 22712 -16872 23800 -16808
rect 23864 -16872 23884 -16808
rect 22712 -16888 23884 -16872
rect 22712 -16952 23800 -16888
rect 23864 -16952 23884 -16888
rect 22712 -16968 23884 -16952
rect 22712 -17032 23800 -16968
rect 23864 -17032 23884 -16968
rect 22712 -17048 23884 -17032
rect 22712 -17112 23800 -17048
rect 23864 -17112 23884 -17048
rect 22712 -17128 23884 -17112
rect 22712 -17192 23800 -17128
rect 23864 -17192 23884 -17128
rect 22712 -17240 23884 -17192
rect -23884 -17528 -22712 -17480
rect -23884 -17592 -22796 -17528
rect -22732 -17592 -22712 -17528
rect -23884 -17608 -22712 -17592
rect -23884 -17672 -22796 -17608
rect -22732 -17672 -22712 -17608
rect -23884 -17688 -22712 -17672
rect -23884 -17752 -22796 -17688
rect -22732 -17752 -22712 -17688
rect -23884 -17768 -22712 -17752
rect -23884 -17832 -22796 -17768
rect -22732 -17832 -22712 -17768
rect -23884 -17848 -22712 -17832
rect -23884 -17912 -22796 -17848
rect -22732 -17912 -22712 -17848
rect -23884 -17928 -22712 -17912
rect -23884 -17992 -22796 -17928
rect -22732 -17992 -22712 -17928
rect -23884 -18008 -22712 -17992
rect -23884 -18072 -22796 -18008
rect -22732 -18072 -22712 -18008
rect -23884 -18088 -22712 -18072
rect -23884 -18152 -22796 -18088
rect -22732 -18152 -22712 -18088
rect -23884 -18168 -22712 -18152
rect -23884 -18232 -22796 -18168
rect -22732 -18232 -22712 -18168
rect -23884 -18248 -22712 -18232
rect -23884 -18312 -22796 -18248
rect -22732 -18312 -22712 -18248
rect -23884 -18360 -22712 -18312
rect -22472 -17528 -21300 -17480
rect -22472 -17592 -21384 -17528
rect -21320 -17592 -21300 -17528
rect -22472 -17608 -21300 -17592
rect -22472 -17672 -21384 -17608
rect -21320 -17672 -21300 -17608
rect -22472 -17688 -21300 -17672
rect -22472 -17752 -21384 -17688
rect -21320 -17752 -21300 -17688
rect -22472 -17768 -21300 -17752
rect -22472 -17832 -21384 -17768
rect -21320 -17832 -21300 -17768
rect -22472 -17848 -21300 -17832
rect -22472 -17912 -21384 -17848
rect -21320 -17912 -21300 -17848
rect -22472 -17928 -21300 -17912
rect -22472 -17992 -21384 -17928
rect -21320 -17992 -21300 -17928
rect -22472 -18008 -21300 -17992
rect -22472 -18072 -21384 -18008
rect -21320 -18072 -21300 -18008
rect -22472 -18088 -21300 -18072
rect -22472 -18152 -21384 -18088
rect -21320 -18152 -21300 -18088
rect -22472 -18168 -21300 -18152
rect -22472 -18232 -21384 -18168
rect -21320 -18232 -21300 -18168
rect -22472 -18248 -21300 -18232
rect -22472 -18312 -21384 -18248
rect -21320 -18312 -21300 -18248
rect -22472 -18360 -21300 -18312
rect -21060 -17528 -19888 -17480
rect -21060 -17592 -19972 -17528
rect -19908 -17592 -19888 -17528
rect -21060 -17608 -19888 -17592
rect -21060 -17672 -19972 -17608
rect -19908 -17672 -19888 -17608
rect -21060 -17688 -19888 -17672
rect -21060 -17752 -19972 -17688
rect -19908 -17752 -19888 -17688
rect -21060 -17768 -19888 -17752
rect -21060 -17832 -19972 -17768
rect -19908 -17832 -19888 -17768
rect -21060 -17848 -19888 -17832
rect -21060 -17912 -19972 -17848
rect -19908 -17912 -19888 -17848
rect -21060 -17928 -19888 -17912
rect -21060 -17992 -19972 -17928
rect -19908 -17992 -19888 -17928
rect -21060 -18008 -19888 -17992
rect -21060 -18072 -19972 -18008
rect -19908 -18072 -19888 -18008
rect -21060 -18088 -19888 -18072
rect -21060 -18152 -19972 -18088
rect -19908 -18152 -19888 -18088
rect -21060 -18168 -19888 -18152
rect -21060 -18232 -19972 -18168
rect -19908 -18232 -19888 -18168
rect -21060 -18248 -19888 -18232
rect -21060 -18312 -19972 -18248
rect -19908 -18312 -19888 -18248
rect -21060 -18360 -19888 -18312
rect -19648 -17528 -18476 -17480
rect -19648 -17592 -18560 -17528
rect -18496 -17592 -18476 -17528
rect -19648 -17608 -18476 -17592
rect -19648 -17672 -18560 -17608
rect -18496 -17672 -18476 -17608
rect -19648 -17688 -18476 -17672
rect -19648 -17752 -18560 -17688
rect -18496 -17752 -18476 -17688
rect -19648 -17768 -18476 -17752
rect -19648 -17832 -18560 -17768
rect -18496 -17832 -18476 -17768
rect -19648 -17848 -18476 -17832
rect -19648 -17912 -18560 -17848
rect -18496 -17912 -18476 -17848
rect -19648 -17928 -18476 -17912
rect -19648 -17992 -18560 -17928
rect -18496 -17992 -18476 -17928
rect -19648 -18008 -18476 -17992
rect -19648 -18072 -18560 -18008
rect -18496 -18072 -18476 -18008
rect -19648 -18088 -18476 -18072
rect -19648 -18152 -18560 -18088
rect -18496 -18152 -18476 -18088
rect -19648 -18168 -18476 -18152
rect -19648 -18232 -18560 -18168
rect -18496 -18232 -18476 -18168
rect -19648 -18248 -18476 -18232
rect -19648 -18312 -18560 -18248
rect -18496 -18312 -18476 -18248
rect -19648 -18360 -18476 -18312
rect -18236 -17528 -17064 -17480
rect -18236 -17592 -17148 -17528
rect -17084 -17592 -17064 -17528
rect -18236 -17608 -17064 -17592
rect -18236 -17672 -17148 -17608
rect -17084 -17672 -17064 -17608
rect -18236 -17688 -17064 -17672
rect -18236 -17752 -17148 -17688
rect -17084 -17752 -17064 -17688
rect -18236 -17768 -17064 -17752
rect -18236 -17832 -17148 -17768
rect -17084 -17832 -17064 -17768
rect -18236 -17848 -17064 -17832
rect -18236 -17912 -17148 -17848
rect -17084 -17912 -17064 -17848
rect -18236 -17928 -17064 -17912
rect -18236 -17992 -17148 -17928
rect -17084 -17992 -17064 -17928
rect -18236 -18008 -17064 -17992
rect -18236 -18072 -17148 -18008
rect -17084 -18072 -17064 -18008
rect -18236 -18088 -17064 -18072
rect -18236 -18152 -17148 -18088
rect -17084 -18152 -17064 -18088
rect -18236 -18168 -17064 -18152
rect -18236 -18232 -17148 -18168
rect -17084 -18232 -17064 -18168
rect -18236 -18248 -17064 -18232
rect -18236 -18312 -17148 -18248
rect -17084 -18312 -17064 -18248
rect -18236 -18360 -17064 -18312
rect -16824 -17528 -15652 -17480
rect -16824 -17592 -15736 -17528
rect -15672 -17592 -15652 -17528
rect -16824 -17608 -15652 -17592
rect -16824 -17672 -15736 -17608
rect -15672 -17672 -15652 -17608
rect -16824 -17688 -15652 -17672
rect -16824 -17752 -15736 -17688
rect -15672 -17752 -15652 -17688
rect -16824 -17768 -15652 -17752
rect -16824 -17832 -15736 -17768
rect -15672 -17832 -15652 -17768
rect -16824 -17848 -15652 -17832
rect -16824 -17912 -15736 -17848
rect -15672 -17912 -15652 -17848
rect -16824 -17928 -15652 -17912
rect -16824 -17992 -15736 -17928
rect -15672 -17992 -15652 -17928
rect -16824 -18008 -15652 -17992
rect -16824 -18072 -15736 -18008
rect -15672 -18072 -15652 -18008
rect -16824 -18088 -15652 -18072
rect -16824 -18152 -15736 -18088
rect -15672 -18152 -15652 -18088
rect -16824 -18168 -15652 -18152
rect -16824 -18232 -15736 -18168
rect -15672 -18232 -15652 -18168
rect -16824 -18248 -15652 -18232
rect -16824 -18312 -15736 -18248
rect -15672 -18312 -15652 -18248
rect -16824 -18360 -15652 -18312
rect -15412 -17528 -14240 -17480
rect -15412 -17592 -14324 -17528
rect -14260 -17592 -14240 -17528
rect -15412 -17608 -14240 -17592
rect -15412 -17672 -14324 -17608
rect -14260 -17672 -14240 -17608
rect -15412 -17688 -14240 -17672
rect -15412 -17752 -14324 -17688
rect -14260 -17752 -14240 -17688
rect -15412 -17768 -14240 -17752
rect -15412 -17832 -14324 -17768
rect -14260 -17832 -14240 -17768
rect -15412 -17848 -14240 -17832
rect -15412 -17912 -14324 -17848
rect -14260 -17912 -14240 -17848
rect -15412 -17928 -14240 -17912
rect -15412 -17992 -14324 -17928
rect -14260 -17992 -14240 -17928
rect -15412 -18008 -14240 -17992
rect -15412 -18072 -14324 -18008
rect -14260 -18072 -14240 -18008
rect -15412 -18088 -14240 -18072
rect -15412 -18152 -14324 -18088
rect -14260 -18152 -14240 -18088
rect -15412 -18168 -14240 -18152
rect -15412 -18232 -14324 -18168
rect -14260 -18232 -14240 -18168
rect -15412 -18248 -14240 -18232
rect -15412 -18312 -14324 -18248
rect -14260 -18312 -14240 -18248
rect -15412 -18360 -14240 -18312
rect -14000 -17528 -12828 -17480
rect -14000 -17592 -12912 -17528
rect -12848 -17592 -12828 -17528
rect -14000 -17608 -12828 -17592
rect -14000 -17672 -12912 -17608
rect -12848 -17672 -12828 -17608
rect -14000 -17688 -12828 -17672
rect -14000 -17752 -12912 -17688
rect -12848 -17752 -12828 -17688
rect -14000 -17768 -12828 -17752
rect -14000 -17832 -12912 -17768
rect -12848 -17832 -12828 -17768
rect -14000 -17848 -12828 -17832
rect -14000 -17912 -12912 -17848
rect -12848 -17912 -12828 -17848
rect -14000 -17928 -12828 -17912
rect -14000 -17992 -12912 -17928
rect -12848 -17992 -12828 -17928
rect -14000 -18008 -12828 -17992
rect -14000 -18072 -12912 -18008
rect -12848 -18072 -12828 -18008
rect -14000 -18088 -12828 -18072
rect -14000 -18152 -12912 -18088
rect -12848 -18152 -12828 -18088
rect -14000 -18168 -12828 -18152
rect -14000 -18232 -12912 -18168
rect -12848 -18232 -12828 -18168
rect -14000 -18248 -12828 -18232
rect -14000 -18312 -12912 -18248
rect -12848 -18312 -12828 -18248
rect -14000 -18360 -12828 -18312
rect -12588 -17528 -11416 -17480
rect -12588 -17592 -11500 -17528
rect -11436 -17592 -11416 -17528
rect -12588 -17608 -11416 -17592
rect -12588 -17672 -11500 -17608
rect -11436 -17672 -11416 -17608
rect -12588 -17688 -11416 -17672
rect -12588 -17752 -11500 -17688
rect -11436 -17752 -11416 -17688
rect -12588 -17768 -11416 -17752
rect -12588 -17832 -11500 -17768
rect -11436 -17832 -11416 -17768
rect -12588 -17848 -11416 -17832
rect -12588 -17912 -11500 -17848
rect -11436 -17912 -11416 -17848
rect -12588 -17928 -11416 -17912
rect -12588 -17992 -11500 -17928
rect -11436 -17992 -11416 -17928
rect -12588 -18008 -11416 -17992
rect -12588 -18072 -11500 -18008
rect -11436 -18072 -11416 -18008
rect -12588 -18088 -11416 -18072
rect -12588 -18152 -11500 -18088
rect -11436 -18152 -11416 -18088
rect -12588 -18168 -11416 -18152
rect -12588 -18232 -11500 -18168
rect -11436 -18232 -11416 -18168
rect -12588 -18248 -11416 -18232
rect -12588 -18312 -11500 -18248
rect -11436 -18312 -11416 -18248
rect -12588 -18360 -11416 -18312
rect -11176 -17528 -10004 -17480
rect -11176 -17592 -10088 -17528
rect -10024 -17592 -10004 -17528
rect -11176 -17608 -10004 -17592
rect -11176 -17672 -10088 -17608
rect -10024 -17672 -10004 -17608
rect -11176 -17688 -10004 -17672
rect -11176 -17752 -10088 -17688
rect -10024 -17752 -10004 -17688
rect -11176 -17768 -10004 -17752
rect -11176 -17832 -10088 -17768
rect -10024 -17832 -10004 -17768
rect -11176 -17848 -10004 -17832
rect -11176 -17912 -10088 -17848
rect -10024 -17912 -10004 -17848
rect -11176 -17928 -10004 -17912
rect -11176 -17992 -10088 -17928
rect -10024 -17992 -10004 -17928
rect -11176 -18008 -10004 -17992
rect -11176 -18072 -10088 -18008
rect -10024 -18072 -10004 -18008
rect -11176 -18088 -10004 -18072
rect -11176 -18152 -10088 -18088
rect -10024 -18152 -10004 -18088
rect -11176 -18168 -10004 -18152
rect -11176 -18232 -10088 -18168
rect -10024 -18232 -10004 -18168
rect -11176 -18248 -10004 -18232
rect -11176 -18312 -10088 -18248
rect -10024 -18312 -10004 -18248
rect -11176 -18360 -10004 -18312
rect -9764 -17528 -8592 -17480
rect -9764 -17592 -8676 -17528
rect -8612 -17592 -8592 -17528
rect -9764 -17608 -8592 -17592
rect -9764 -17672 -8676 -17608
rect -8612 -17672 -8592 -17608
rect -9764 -17688 -8592 -17672
rect -9764 -17752 -8676 -17688
rect -8612 -17752 -8592 -17688
rect -9764 -17768 -8592 -17752
rect -9764 -17832 -8676 -17768
rect -8612 -17832 -8592 -17768
rect -9764 -17848 -8592 -17832
rect -9764 -17912 -8676 -17848
rect -8612 -17912 -8592 -17848
rect -9764 -17928 -8592 -17912
rect -9764 -17992 -8676 -17928
rect -8612 -17992 -8592 -17928
rect -9764 -18008 -8592 -17992
rect -9764 -18072 -8676 -18008
rect -8612 -18072 -8592 -18008
rect -9764 -18088 -8592 -18072
rect -9764 -18152 -8676 -18088
rect -8612 -18152 -8592 -18088
rect -9764 -18168 -8592 -18152
rect -9764 -18232 -8676 -18168
rect -8612 -18232 -8592 -18168
rect -9764 -18248 -8592 -18232
rect -9764 -18312 -8676 -18248
rect -8612 -18312 -8592 -18248
rect -9764 -18360 -8592 -18312
rect -8352 -17528 -7180 -17480
rect -8352 -17592 -7264 -17528
rect -7200 -17592 -7180 -17528
rect -8352 -17608 -7180 -17592
rect -8352 -17672 -7264 -17608
rect -7200 -17672 -7180 -17608
rect -8352 -17688 -7180 -17672
rect -8352 -17752 -7264 -17688
rect -7200 -17752 -7180 -17688
rect -8352 -17768 -7180 -17752
rect -8352 -17832 -7264 -17768
rect -7200 -17832 -7180 -17768
rect -8352 -17848 -7180 -17832
rect -8352 -17912 -7264 -17848
rect -7200 -17912 -7180 -17848
rect -8352 -17928 -7180 -17912
rect -8352 -17992 -7264 -17928
rect -7200 -17992 -7180 -17928
rect -8352 -18008 -7180 -17992
rect -8352 -18072 -7264 -18008
rect -7200 -18072 -7180 -18008
rect -8352 -18088 -7180 -18072
rect -8352 -18152 -7264 -18088
rect -7200 -18152 -7180 -18088
rect -8352 -18168 -7180 -18152
rect -8352 -18232 -7264 -18168
rect -7200 -18232 -7180 -18168
rect -8352 -18248 -7180 -18232
rect -8352 -18312 -7264 -18248
rect -7200 -18312 -7180 -18248
rect -8352 -18360 -7180 -18312
rect -6940 -17528 -5768 -17480
rect -6940 -17592 -5852 -17528
rect -5788 -17592 -5768 -17528
rect -6940 -17608 -5768 -17592
rect -6940 -17672 -5852 -17608
rect -5788 -17672 -5768 -17608
rect -6940 -17688 -5768 -17672
rect -6940 -17752 -5852 -17688
rect -5788 -17752 -5768 -17688
rect -6940 -17768 -5768 -17752
rect -6940 -17832 -5852 -17768
rect -5788 -17832 -5768 -17768
rect -6940 -17848 -5768 -17832
rect -6940 -17912 -5852 -17848
rect -5788 -17912 -5768 -17848
rect -6940 -17928 -5768 -17912
rect -6940 -17992 -5852 -17928
rect -5788 -17992 -5768 -17928
rect -6940 -18008 -5768 -17992
rect -6940 -18072 -5852 -18008
rect -5788 -18072 -5768 -18008
rect -6940 -18088 -5768 -18072
rect -6940 -18152 -5852 -18088
rect -5788 -18152 -5768 -18088
rect -6940 -18168 -5768 -18152
rect -6940 -18232 -5852 -18168
rect -5788 -18232 -5768 -18168
rect -6940 -18248 -5768 -18232
rect -6940 -18312 -5852 -18248
rect -5788 -18312 -5768 -18248
rect -6940 -18360 -5768 -18312
rect -5528 -17528 -4356 -17480
rect -5528 -17592 -4440 -17528
rect -4376 -17592 -4356 -17528
rect -5528 -17608 -4356 -17592
rect -5528 -17672 -4440 -17608
rect -4376 -17672 -4356 -17608
rect -5528 -17688 -4356 -17672
rect -5528 -17752 -4440 -17688
rect -4376 -17752 -4356 -17688
rect -5528 -17768 -4356 -17752
rect -5528 -17832 -4440 -17768
rect -4376 -17832 -4356 -17768
rect -5528 -17848 -4356 -17832
rect -5528 -17912 -4440 -17848
rect -4376 -17912 -4356 -17848
rect -5528 -17928 -4356 -17912
rect -5528 -17992 -4440 -17928
rect -4376 -17992 -4356 -17928
rect -5528 -18008 -4356 -17992
rect -5528 -18072 -4440 -18008
rect -4376 -18072 -4356 -18008
rect -5528 -18088 -4356 -18072
rect -5528 -18152 -4440 -18088
rect -4376 -18152 -4356 -18088
rect -5528 -18168 -4356 -18152
rect -5528 -18232 -4440 -18168
rect -4376 -18232 -4356 -18168
rect -5528 -18248 -4356 -18232
rect -5528 -18312 -4440 -18248
rect -4376 -18312 -4356 -18248
rect -5528 -18360 -4356 -18312
rect -4116 -17528 -2944 -17480
rect -4116 -17592 -3028 -17528
rect -2964 -17592 -2944 -17528
rect -4116 -17608 -2944 -17592
rect -4116 -17672 -3028 -17608
rect -2964 -17672 -2944 -17608
rect -4116 -17688 -2944 -17672
rect -4116 -17752 -3028 -17688
rect -2964 -17752 -2944 -17688
rect -4116 -17768 -2944 -17752
rect -4116 -17832 -3028 -17768
rect -2964 -17832 -2944 -17768
rect -4116 -17848 -2944 -17832
rect -4116 -17912 -3028 -17848
rect -2964 -17912 -2944 -17848
rect -4116 -17928 -2944 -17912
rect -4116 -17992 -3028 -17928
rect -2964 -17992 -2944 -17928
rect -4116 -18008 -2944 -17992
rect -4116 -18072 -3028 -18008
rect -2964 -18072 -2944 -18008
rect -4116 -18088 -2944 -18072
rect -4116 -18152 -3028 -18088
rect -2964 -18152 -2944 -18088
rect -4116 -18168 -2944 -18152
rect -4116 -18232 -3028 -18168
rect -2964 -18232 -2944 -18168
rect -4116 -18248 -2944 -18232
rect -4116 -18312 -3028 -18248
rect -2964 -18312 -2944 -18248
rect -4116 -18360 -2944 -18312
rect -2704 -17528 -1532 -17480
rect -2704 -17592 -1616 -17528
rect -1552 -17592 -1532 -17528
rect -2704 -17608 -1532 -17592
rect -2704 -17672 -1616 -17608
rect -1552 -17672 -1532 -17608
rect -2704 -17688 -1532 -17672
rect -2704 -17752 -1616 -17688
rect -1552 -17752 -1532 -17688
rect -2704 -17768 -1532 -17752
rect -2704 -17832 -1616 -17768
rect -1552 -17832 -1532 -17768
rect -2704 -17848 -1532 -17832
rect -2704 -17912 -1616 -17848
rect -1552 -17912 -1532 -17848
rect -2704 -17928 -1532 -17912
rect -2704 -17992 -1616 -17928
rect -1552 -17992 -1532 -17928
rect -2704 -18008 -1532 -17992
rect -2704 -18072 -1616 -18008
rect -1552 -18072 -1532 -18008
rect -2704 -18088 -1532 -18072
rect -2704 -18152 -1616 -18088
rect -1552 -18152 -1532 -18088
rect -2704 -18168 -1532 -18152
rect -2704 -18232 -1616 -18168
rect -1552 -18232 -1532 -18168
rect -2704 -18248 -1532 -18232
rect -2704 -18312 -1616 -18248
rect -1552 -18312 -1532 -18248
rect -2704 -18360 -1532 -18312
rect -1292 -17528 -120 -17480
rect -1292 -17592 -204 -17528
rect -140 -17592 -120 -17528
rect -1292 -17608 -120 -17592
rect -1292 -17672 -204 -17608
rect -140 -17672 -120 -17608
rect -1292 -17688 -120 -17672
rect -1292 -17752 -204 -17688
rect -140 -17752 -120 -17688
rect -1292 -17768 -120 -17752
rect -1292 -17832 -204 -17768
rect -140 -17832 -120 -17768
rect -1292 -17848 -120 -17832
rect -1292 -17912 -204 -17848
rect -140 -17912 -120 -17848
rect -1292 -17928 -120 -17912
rect -1292 -17992 -204 -17928
rect -140 -17992 -120 -17928
rect -1292 -18008 -120 -17992
rect -1292 -18072 -204 -18008
rect -140 -18072 -120 -18008
rect -1292 -18088 -120 -18072
rect -1292 -18152 -204 -18088
rect -140 -18152 -120 -18088
rect -1292 -18168 -120 -18152
rect -1292 -18232 -204 -18168
rect -140 -18232 -120 -18168
rect -1292 -18248 -120 -18232
rect -1292 -18312 -204 -18248
rect -140 -18312 -120 -18248
rect -1292 -18360 -120 -18312
rect 120 -17528 1292 -17480
rect 120 -17592 1208 -17528
rect 1272 -17592 1292 -17528
rect 120 -17608 1292 -17592
rect 120 -17672 1208 -17608
rect 1272 -17672 1292 -17608
rect 120 -17688 1292 -17672
rect 120 -17752 1208 -17688
rect 1272 -17752 1292 -17688
rect 120 -17768 1292 -17752
rect 120 -17832 1208 -17768
rect 1272 -17832 1292 -17768
rect 120 -17848 1292 -17832
rect 120 -17912 1208 -17848
rect 1272 -17912 1292 -17848
rect 120 -17928 1292 -17912
rect 120 -17992 1208 -17928
rect 1272 -17992 1292 -17928
rect 120 -18008 1292 -17992
rect 120 -18072 1208 -18008
rect 1272 -18072 1292 -18008
rect 120 -18088 1292 -18072
rect 120 -18152 1208 -18088
rect 1272 -18152 1292 -18088
rect 120 -18168 1292 -18152
rect 120 -18232 1208 -18168
rect 1272 -18232 1292 -18168
rect 120 -18248 1292 -18232
rect 120 -18312 1208 -18248
rect 1272 -18312 1292 -18248
rect 120 -18360 1292 -18312
rect 1532 -17528 2704 -17480
rect 1532 -17592 2620 -17528
rect 2684 -17592 2704 -17528
rect 1532 -17608 2704 -17592
rect 1532 -17672 2620 -17608
rect 2684 -17672 2704 -17608
rect 1532 -17688 2704 -17672
rect 1532 -17752 2620 -17688
rect 2684 -17752 2704 -17688
rect 1532 -17768 2704 -17752
rect 1532 -17832 2620 -17768
rect 2684 -17832 2704 -17768
rect 1532 -17848 2704 -17832
rect 1532 -17912 2620 -17848
rect 2684 -17912 2704 -17848
rect 1532 -17928 2704 -17912
rect 1532 -17992 2620 -17928
rect 2684 -17992 2704 -17928
rect 1532 -18008 2704 -17992
rect 1532 -18072 2620 -18008
rect 2684 -18072 2704 -18008
rect 1532 -18088 2704 -18072
rect 1532 -18152 2620 -18088
rect 2684 -18152 2704 -18088
rect 1532 -18168 2704 -18152
rect 1532 -18232 2620 -18168
rect 2684 -18232 2704 -18168
rect 1532 -18248 2704 -18232
rect 1532 -18312 2620 -18248
rect 2684 -18312 2704 -18248
rect 1532 -18360 2704 -18312
rect 2944 -17528 4116 -17480
rect 2944 -17592 4032 -17528
rect 4096 -17592 4116 -17528
rect 2944 -17608 4116 -17592
rect 2944 -17672 4032 -17608
rect 4096 -17672 4116 -17608
rect 2944 -17688 4116 -17672
rect 2944 -17752 4032 -17688
rect 4096 -17752 4116 -17688
rect 2944 -17768 4116 -17752
rect 2944 -17832 4032 -17768
rect 4096 -17832 4116 -17768
rect 2944 -17848 4116 -17832
rect 2944 -17912 4032 -17848
rect 4096 -17912 4116 -17848
rect 2944 -17928 4116 -17912
rect 2944 -17992 4032 -17928
rect 4096 -17992 4116 -17928
rect 2944 -18008 4116 -17992
rect 2944 -18072 4032 -18008
rect 4096 -18072 4116 -18008
rect 2944 -18088 4116 -18072
rect 2944 -18152 4032 -18088
rect 4096 -18152 4116 -18088
rect 2944 -18168 4116 -18152
rect 2944 -18232 4032 -18168
rect 4096 -18232 4116 -18168
rect 2944 -18248 4116 -18232
rect 2944 -18312 4032 -18248
rect 4096 -18312 4116 -18248
rect 2944 -18360 4116 -18312
rect 4356 -17528 5528 -17480
rect 4356 -17592 5444 -17528
rect 5508 -17592 5528 -17528
rect 4356 -17608 5528 -17592
rect 4356 -17672 5444 -17608
rect 5508 -17672 5528 -17608
rect 4356 -17688 5528 -17672
rect 4356 -17752 5444 -17688
rect 5508 -17752 5528 -17688
rect 4356 -17768 5528 -17752
rect 4356 -17832 5444 -17768
rect 5508 -17832 5528 -17768
rect 4356 -17848 5528 -17832
rect 4356 -17912 5444 -17848
rect 5508 -17912 5528 -17848
rect 4356 -17928 5528 -17912
rect 4356 -17992 5444 -17928
rect 5508 -17992 5528 -17928
rect 4356 -18008 5528 -17992
rect 4356 -18072 5444 -18008
rect 5508 -18072 5528 -18008
rect 4356 -18088 5528 -18072
rect 4356 -18152 5444 -18088
rect 5508 -18152 5528 -18088
rect 4356 -18168 5528 -18152
rect 4356 -18232 5444 -18168
rect 5508 -18232 5528 -18168
rect 4356 -18248 5528 -18232
rect 4356 -18312 5444 -18248
rect 5508 -18312 5528 -18248
rect 4356 -18360 5528 -18312
rect 5768 -17528 6940 -17480
rect 5768 -17592 6856 -17528
rect 6920 -17592 6940 -17528
rect 5768 -17608 6940 -17592
rect 5768 -17672 6856 -17608
rect 6920 -17672 6940 -17608
rect 5768 -17688 6940 -17672
rect 5768 -17752 6856 -17688
rect 6920 -17752 6940 -17688
rect 5768 -17768 6940 -17752
rect 5768 -17832 6856 -17768
rect 6920 -17832 6940 -17768
rect 5768 -17848 6940 -17832
rect 5768 -17912 6856 -17848
rect 6920 -17912 6940 -17848
rect 5768 -17928 6940 -17912
rect 5768 -17992 6856 -17928
rect 6920 -17992 6940 -17928
rect 5768 -18008 6940 -17992
rect 5768 -18072 6856 -18008
rect 6920 -18072 6940 -18008
rect 5768 -18088 6940 -18072
rect 5768 -18152 6856 -18088
rect 6920 -18152 6940 -18088
rect 5768 -18168 6940 -18152
rect 5768 -18232 6856 -18168
rect 6920 -18232 6940 -18168
rect 5768 -18248 6940 -18232
rect 5768 -18312 6856 -18248
rect 6920 -18312 6940 -18248
rect 5768 -18360 6940 -18312
rect 7180 -17528 8352 -17480
rect 7180 -17592 8268 -17528
rect 8332 -17592 8352 -17528
rect 7180 -17608 8352 -17592
rect 7180 -17672 8268 -17608
rect 8332 -17672 8352 -17608
rect 7180 -17688 8352 -17672
rect 7180 -17752 8268 -17688
rect 8332 -17752 8352 -17688
rect 7180 -17768 8352 -17752
rect 7180 -17832 8268 -17768
rect 8332 -17832 8352 -17768
rect 7180 -17848 8352 -17832
rect 7180 -17912 8268 -17848
rect 8332 -17912 8352 -17848
rect 7180 -17928 8352 -17912
rect 7180 -17992 8268 -17928
rect 8332 -17992 8352 -17928
rect 7180 -18008 8352 -17992
rect 7180 -18072 8268 -18008
rect 8332 -18072 8352 -18008
rect 7180 -18088 8352 -18072
rect 7180 -18152 8268 -18088
rect 8332 -18152 8352 -18088
rect 7180 -18168 8352 -18152
rect 7180 -18232 8268 -18168
rect 8332 -18232 8352 -18168
rect 7180 -18248 8352 -18232
rect 7180 -18312 8268 -18248
rect 8332 -18312 8352 -18248
rect 7180 -18360 8352 -18312
rect 8592 -17528 9764 -17480
rect 8592 -17592 9680 -17528
rect 9744 -17592 9764 -17528
rect 8592 -17608 9764 -17592
rect 8592 -17672 9680 -17608
rect 9744 -17672 9764 -17608
rect 8592 -17688 9764 -17672
rect 8592 -17752 9680 -17688
rect 9744 -17752 9764 -17688
rect 8592 -17768 9764 -17752
rect 8592 -17832 9680 -17768
rect 9744 -17832 9764 -17768
rect 8592 -17848 9764 -17832
rect 8592 -17912 9680 -17848
rect 9744 -17912 9764 -17848
rect 8592 -17928 9764 -17912
rect 8592 -17992 9680 -17928
rect 9744 -17992 9764 -17928
rect 8592 -18008 9764 -17992
rect 8592 -18072 9680 -18008
rect 9744 -18072 9764 -18008
rect 8592 -18088 9764 -18072
rect 8592 -18152 9680 -18088
rect 9744 -18152 9764 -18088
rect 8592 -18168 9764 -18152
rect 8592 -18232 9680 -18168
rect 9744 -18232 9764 -18168
rect 8592 -18248 9764 -18232
rect 8592 -18312 9680 -18248
rect 9744 -18312 9764 -18248
rect 8592 -18360 9764 -18312
rect 10004 -17528 11176 -17480
rect 10004 -17592 11092 -17528
rect 11156 -17592 11176 -17528
rect 10004 -17608 11176 -17592
rect 10004 -17672 11092 -17608
rect 11156 -17672 11176 -17608
rect 10004 -17688 11176 -17672
rect 10004 -17752 11092 -17688
rect 11156 -17752 11176 -17688
rect 10004 -17768 11176 -17752
rect 10004 -17832 11092 -17768
rect 11156 -17832 11176 -17768
rect 10004 -17848 11176 -17832
rect 10004 -17912 11092 -17848
rect 11156 -17912 11176 -17848
rect 10004 -17928 11176 -17912
rect 10004 -17992 11092 -17928
rect 11156 -17992 11176 -17928
rect 10004 -18008 11176 -17992
rect 10004 -18072 11092 -18008
rect 11156 -18072 11176 -18008
rect 10004 -18088 11176 -18072
rect 10004 -18152 11092 -18088
rect 11156 -18152 11176 -18088
rect 10004 -18168 11176 -18152
rect 10004 -18232 11092 -18168
rect 11156 -18232 11176 -18168
rect 10004 -18248 11176 -18232
rect 10004 -18312 11092 -18248
rect 11156 -18312 11176 -18248
rect 10004 -18360 11176 -18312
rect 11416 -17528 12588 -17480
rect 11416 -17592 12504 -17528
rect 12568 -17592 12588 -17528
rect 11416 -17608 12588 -17592
rect 11416 -17672 12504 -17608
rect 12568 -17672 12588 -17608
rect 11416 -17688 12588 -17672
rect 11416 -17752 12504 -17688
rect 12568 -17752 12588 -17688
rect 11416 -17768 12588 -17752
rect 11416 -17832 12504 -17768
rect 12568 -17832 12588 -17768
rect 11416 -17848 12588 -17832
rect 11416 -17912 12504 -17848
rect 12568 -17912 12588 -17848
rect 11416 -17928 12588 -17912
rect 11416 -17992 12504 -17928
rect 12568 -17992 12588 -17928
rect 11416 -18008 12588 -17992
rect 11416 -18072 12504 -18008
rect 12568 -18072 12588 -18008
rect 11416 -18088 12588 -18072
rect 11416 -18152 12504 -18088
rect 12568 -18152 12588 -18088
rect 11416 -18168 12588 -18152
rect 11416 -18232 12504 -18168
rect 12568 -18232 12588 -18168
rect 11416 -18248 12588 -18232
rect 11416 -18312 12504 -18248
rect 12568 -18312 12588 -18248
rect 11416 -18360 12588 -18312
rect 12828 -17528 14000 -17480
rect 12828 -17592 13916 -17528
rect 13980 -17592 14000 -17528
rect 12828 -17608 14000 -17592
rect 12828 -17672 13916 -17608
rect 13980 -17672 14000 -17608
rect 12828 -17688 14000 -17672
rect 12828 -17752 13916 -17688
rect 13980 -17752 14000 -17688
rect 12828 -17768 14000 -17752
rect 12828 -17832 13916 -17768
rect 13980 -17832 14000 -17768
rect 12828 -17848 14000 -17832
rect 12828 -17912 13916 -17848
rect 13980 -17912 14000 -17848
rect 12828 -17928 14000 -17912
rect 12828 -17992 13916 -17928
rect 13980 -17992 14000 -17928
rect 12828 -18008 14000 -17992
rect 12828 -18072 13916 -18008
rect 13980 -18072 14000 -18008
rect 12828 -18088 14000 -18072
rect 12828 -18152 13916 -18088
rect 13980 -18152 14000 -18088
rect 12828 -18168 14000 -18152
rect 12828 -18232 13916 -18168
rect 13980 -18232 14000 -18168
rect 12828 -18248 14000 -18232
rect 12828 -18312 13916 -18248
rect 13980 -18312 14000 -18248
rect 12828 -18360 14000 -18312
rect 14240 -17528 15412 -17480
rect 14240 -17592 15328 -17528
rect 15392 -17592 15412 -17528
rect 14240 -17608 15412 -17592
rect 14240 -17672 15328 -17608
rect 15392 -17672 15412 -17608
rect 14240 -17688 15412 -17672
rect 14240 -17752 15328 -17688
rect 15392 -17752 15412 -17688
rect 14240 -17768 15412 -17752
rect 14240 -17832 15328 -17768
rect 15392 -17832 15412 -17768
rect 14240 -17848 15412 -17832
rect 14240 -17912 15328 -17848
rect 15392 -17912 15412 -17848
rect 14240 -17928 15412 -17912
rect 14240 -17992 15328 -17928
rect 15392 -17992 15412 -17928
rect 14240 -18008 15412 -17992
rect 14240 -18072 15328 -18008
rect 15392 -18072 15412 -18008
rect 14240 -18088 15412 -18072
rect 14240 -18152 15328 -18088
rect 15392 -18152 15412 -18088
rect 14240 -18168 15412 -18152
rect 14240 -18232 15328 -18168
rect 15392 -18232 15412 -18168
rect 14240 -18248 15412 -18232
rect 14240 -18312 15328 -18248
rect 15392 -18312 15412 -18248
rect 14240 -18360 15412 -18312
rect 15652 -17528 16824 -17480
rect 15652 -17592 16740 -17528
rect 16804 -17592 16824 -17528
rect 15652 -17608 16824 -17592
rect 15652 -17672 16740 -17608
rect 16804 -17672 16824 -17608
rect 15652 -17688 16824 -17672
rect 15652 -17752 16740 -17688
rect 16804 -17752 16824 -17688
rect 15652 -17768 16824 -17752
rect 15652 -17832 16740 -17768
rect 16804 -17832 16824 -17768
rect 15652 -17848 16824 -17832
rect 15652 -17912 16740 -17848
rect 16804 -17912 16824 -17848
rect 15652 -17928 16824 -17912
rect 15652 -17992 16740 -17928
rect 16804 -17992 16824 -17928
rect 15652 -18008 16824 -17992
rect 15652 -18072 16740 -18008
rect 16804 -18072 16824 -18008
rect 15652 -18088 16824 -18072
rect 15652 -18152 16740 -18088
rect 16804 -18152 16824 -18088
rect 15652 -18168 16824 -18152
rect 15652 -18232 16740 -18168
rect 16804 -18232 16824 -18168
rect 15652 -18248 16824 -18232
rect 15652 -18312 16740 -18248
rect 16804 -18312 16824 -18248
rect 15652 -18360 16824 -18312
rect 17064 -17528 18236 -17480
rect 17064 -17592 18152 -17528
rect 18216 -17592 18236 -17528
rect 17064 -17608 18236 -17592
rect 17064 -17672 18152 -17608
rect 18216 -17672 18236 -17608
rect 17064 -17688 18236 -17672
rect 17064 -17752 18152 -17688
rect 18216 -17752 18236 -17688
rect 17064 -17768 18236 -17752
rect 17064 -17832 18152 -17768
rect 18216 -17832 18236 -17768
rect 17064 -17848 18236 -17832
rect 17064 -17912 18152 -17848
rect 18216 -17912 18236 -17848
rect 17064 -17928 18236 -17912
rect 17064 -17992 18152 -17928
rect 18216 -17992 18236 -17928
rect 17064 -18008 18236 -17992
rect 17064 -18072 18152 -18008
rect 18216 -18072 18236 -18008
rect 17064 -18088 18236 -18072
rect 17064 -18152 18152 -18088
rect 18216 -18152 18236 -18088
rect 17064 -18168 18236 -18152
rect 17064 -18232 18152 -18168
rect 18216 -18232 18236 -18168
rect 17064 -18248 18236 -18232
rect 17064 -18312 18152 -18248
rect 18216 -18312 18236 -18248
rect 17064 -18360 18236 -18312
rect 18476 -17528 19648 -17480
rect 18476 -17592 19564 -17528
rect 19628 -17592 19648 -17528
rect 18476 -17608 19648 -17592
rect 18476 -17672 19564 -17608
rect 19628 -17672 19648 -17608
rect 18476 -17688 19648 -17672
rect 18476 -17752 19564 -17688
rect 19628 -17752 19648 -17688
rect 18476 -17768 19648 -17752
rect 18476 -17832 19564 -17768
rect 19628 -17832 19648 -17768
rect 18476 -17848 19648 -17832
rect 18476 -17912 19564 -17848
rect 19628 -17912 19648 -17848
rect 18476 -17928 19648 -17912
rect 18476 -17992 19564 -17928
rect 19628 -17992 19648 -17928
rect 18476 -18008 19648 -17992
rect 18476 -18072 19564 -18008
rect 19628 -18072 19648 -18008
rect 18476 -18088 19648 -18072
rect 18476 -18152 19564 -18088
rect 19628 -18152 19648 -18088
rect 18476 -18168 19648 -18152
rect 18476 -18232 19564 -18168
rect 19628 -18232 19648 -18168
rect 18476 -18248 19648 -18232
rect 18476 -18312 19564 -18248
rect 19628 -18312 19648 -18248
rect 18476 -18360 19648 -18312
rect 19888 -17528 21060 -17480
rect 19888 -17592 20976 -17528
rect 21040 -17592 21060 -17528
rect 19888 -17608 21060 -17592
rect 19888 -17672 20976 -17608
rect 21040 -17672 21060 -17608
rect 19888 -17688 21060 -17672
rect 19888 -17752 20976 -17688
rect 21040 -17752 21060 -17688
rect 19888 -17768 21060 -17752
rect 19888 -17832 20976 -17768
rect 21040 -17832 21060 -17768
rect 19888 -17848 21060 -17832
rect 19888 -17912 20976 -17848
rect 21040 -17912 21060 -17848
rect 19888 -17928 21060 -17912
rect 19888 -17992 20976 -17928
rect 21040 -17992 21060 -17928
rect 19888 -18008 21060 -17992
rect 19888 -18072 20976 -18008
rect 21040 -18072 21060 -18008
rect 19888 -18088 21060 -18072
rect 19888 -18152 20976 -18088
rect 21040 -18152 21060 -18088
rect 19888 -18168 21060 -18152
rect 19888 -18232 20976 -18168
rect 21040 -18232 21060 -18168
rect 19888 -18248 21060 -18232
rect 19888 -18312 20976 -18248
rect 21040 -18312 21060 -18248
rect 19888 -18360 21060 -18312
rect 21300 -17528 22472 -17480
rect 21300 -17592 22388 -17528
rect 22452 -17592 22472 -17528
rect 21300 -17608 22472 -17592
rect 21300 -17672 22388 -17608
rect 22452 -17672 22472 -17608
rect 21300 -17688 22472 -17672
rect 21300 -17752 22388 -17688
rect 22452 -17752 22472 -17688
rect 21300 -17768 22472 -17752
rect 21300 -17832 22388 -17768
rect 22452 -17832 22472 -17768
rect 21300 -17848 22472 -17832
rect 21300 -17912 22388 -17848
rect 22452 -17912 22472 -17848
rect 21300 -17928 22472 -17912
rect 21300 -17992 22388 -17928
rect 22452 -17992 22472 -17928
rect 21300 -18008 22472 -17992
rect 21300 -18072 22388 -18008
rect 22452 -18072 22472 -18008
rect 21300 -18088 22472 -18072
rect 21300 -18152 22388 -18088
rect 22452 -18152 22472 -18088
rect 21300 -18168 22472 -18152
rect 21300 -18232 22388 -18168
rect 22452 -18232 22472 -18168
rect 21300 -18248 22472 -18232
rect 21300 -18312 22388 -18248
rect 22452 -18312 22472 -18248
rect 21300 -18360 22472 -18312
rect 22712 -17528 23884 -17480
rect 22712 -17592 23800 -17528
rect 23864 -17592 23884 -17528
rect 22712 -17608 23884 -17592
rect 22712 -17672 23800 -17608
rect 23864 -17672 23884 -17608
rect 22712 -17688 23884 -17672
rect 22712 -17752 23800 -17688
rect 23864 -17752 23884 -17688
rect 22712 -17768 23884 -17752
rect 22712 -17832 23800 -17768
rect 23864 -17832 23884 -17768
rect 22712 -17848 23884 -17832
rect 22712 -17912 23800 -17848
rect 23864 -17912 23884 -17848
rect 22712 -17928 23884 -17912
rect 22712 -17992 23800 -17928
rect 23864 -17992 23884 -17928
rect 22712 -18008 23884 -17992
rect 22712 -18072 23800 -18008
rect 23864 -18072 23884 -18008
rect 22712 -18088 23884 -18072
rect 22712 -18152 23800 -18088
rect 23864 -18152 23884 -18088
rect 22712 -18168 23884 -18152
rect 22712 -18232 23800 -18168
rect 23864 -18232 23884 -18168
rect 22712 -18248 23884 -18232
rect 22712 -18312 23800 -18248
rect 23864 -18312 23884 -18248
rect 22712 -18360 23884 -18312
<< via3 >>
rect -22796 18248 -22732 18312
rect -22796 18168 -22732 18232
rect -22796 18088 -22732 18152
rect -22796 18008 -22732 18072
rect -22796 17928 -22732 17992
rect -22796 17848 -22732 17912
rect -22796 17768 -22732 17832
rect -22796 17688 -22732 17752
rect -22796 17608 -22732 17672
rect -22796 17528 -22732 17592
rect -21384 18248 -21320 18312
rect -21384 18168 -21320 18232
rect -21384 18088 -21320 18152
rect -21384 18008 -21320 18072
rect -21384 17928 -21320 17992
rect -21384 17848 -21320 17912
rect -21384 17768 -21320 17832
rect -21384 17688 -21320 17752
rect -21384 17608 -21320 17672
rect -21384 17528 -21320 17592
rect -19972 18248 -19908 18312
rect -19972 18168 -19908 18232
rect -19972 18088 -19908 18152
rect -19972 18008 -19908 18072
rect -19972 17928 -19908 17992
rect -19972 17848 -19908 17912
rect -19972 17768 -19908 17832
rect -19972 17688 -19908 17752
rect -19972 17608 -19908 17672
rect -19972 17528 -19908 17592
rect -18560 18248 -18496 18312
rect -18560 18168 -18496 18232
rect -18560 18088 -18496 18152
rect -18560 18008 -18496 18072
rect -18560 17928 -18496 17992
rect -18560 17848 -18496 17912
rect -18560 17768 -18496 17832
rect -18560 17688 -18496 17752
rect -18560 17608 -18496 17672
rect -18560 17528 -18496 17592
rect -17148 18248 -17084 18312
rect -17148 18168 -17084 18232
rect -17148 18088 -17084 18152
rect -17148 18008 -17084 18072
rect -17148 17928 -17084 17992
rect -17148 17848 -17084 17912
rect -17148 17768 -17084 17832
rect -17148 17688 -17084 17752
rect -17148 17608 -17084 17672
rect -17148 17528 -17084 17592
rect -15736 18248 -15672 18312
rect -15736 18168 -15672 18232
rect -15736 18088 -15672 18152
rect -15736 18008 -15672 18072
rect -15736 17928 -15672 17992
rect -15736 17848 -15672 17912
rect -15736 17768 -15672 17832
rect -15736 17688 -15672 17752
rect -15736 17608 -15672 17672
rect -15736 17528 -15672 17592
rect -14324 18248 -14260 18312
rect -14324 18168 -14260 18232
rect -14324 18088 -14260 18152
rect -14324 18008 -14260 18072
rect -14324 17928 -14260 17992
rect -14324 17848 -14260 17912
rect -14324 17768 -14260 17832
rect -14324 17688 -14260 17752
rect -14324 17608 -14260 17672
rect -14324 17528 -14260 17592
rect -12912 18248 -12848 18312
rect -12912 18168 -12848 18232
rect -12912 18088 -12848 18152
rect -12912 18008 -12848 18072
rect -12912 17928 -12848 17992
rect -12912 17848 -12848 17912
rect -12912 17768 -12848 17832
rect -12912 17688 -12848 17752
rect -12912 17608 -12848 17672
rect -12912 17528 -12848 17592
rect -11500 18248 -11436 18312
rect -11500 18168 -11436 18232
rect -11500 18088 -11436 18152
rect -11500 18008 -11436 18072
rect -11500 17928 -11436 17992
rect -11500 17848 -11436 17912
rect -11500 17768 -11436 17832
rect -11500 17688 -11436 17752
rect -11500 17608 -11436 17672
rect -11500 17528 -11436 17592
rect -10088 18248 -10024 18312
rect -10088 18168 -10024 18232
rect -10088 18088 -10024 18152
rect -10088 18008 -10024 18072
rect -10088 17928 -10024 17992
rect -10088 17848 -10024 17912
rect -10088 17768 -10024 17832
rect -10088 17688 -10024 17752
rect -10088 17608 -10024 17672
rect -10088 17528 -10024 17592
rect -8676 18248 -8612 18312
rect -8676 18168 -8612 18232
rect -8676 18088 -8612 18152
rect -8676 18008 -8612 18072
rect -8676 17928 -8612 17992
rect -8676 17848 -8612 17912
rect -8676 17768 -8612 17832
rect -8676 17688 -8612 17752
rect -8676 17608 -8612 17672
rect -8676 17528 -8612 17592
rect -7264 18248 -7200 18312
rect -7264 18168 -7200 18232
rect -7264 18088 -7200 18152
rect -7264 18008 -7200 18072
rect -7264 17928 -7200 17992
rect -7264 17848 -7200 17912
rect -7264 17768 -7200 17832
rect -7264 17688 -7200 17752
rect -7264 17608 -7200 17672
rect -7264 17528 -7200 17592
rect -5852 18248 -5788 18312
rect -5852 18168 -5788 18232
rect -5852 18088 -5788 18152
rect -5852 18008 -5788 18072
rect -5852 17928 -5788 17992
rect -5852 17848 -5788 17912
rect -5852 17768 -5788 17832
rect -5852 17688 -5788 17752
rect -5852 17608 -5788 17672
rect -5852 17528 -5788 17592
rect -4440 18248 -4376 18312
rect -4440 18168 -4376 18232
rect -4440 18088 -4376 18152
rect -4440 18008 -4376 18072
rect -4440 17928 -4376 17992
rect -4440 17848 -4376 17912
rect -4440 17768 -4376 17832
rect -4440 17688 -4376 17752
rect -4440 17608 -4376 17672
rect -4440 17528 -4376 17592
rect -3028 18248 -2964 18312
rect -3028 18168 -2964 18232
rect -3028 18088 -2964 18152
rect -3028 18008 -2964 18072
rect -3028 17928 -2964 17992
rect -3028 17848 -2964 17912
rect -3028 17768 -2964 17832
rect -3028 17688 -2964 17752
rect -3028 17608 -2964 17672
rect -3028 17528 -2964 17592
rect -1616 18248 -1552 18312
rect -1616 18168 -1552 18232
rect -1616 18088 -1552 18152
rect -1616 18008 -1552 18072
rect -1616 17928 -1552 17992
rect -1616 17848 -1552 17912
rect -1616 17768 -1552 17832
rect -1616 17688 -1552 17752
rect -1616 17608 -1552 17672
rect -1616 17528 -1552 17592
rect -204 18248 -140 18312
rect -204 18168 -140 18232
rect -204 18088 -140 18152
rect -204 18008 -140 18072
rect -204 17928 -140 17992
rect -204 17848 -140 17912
rect -204 17768 -140 17832
rect -204 17688 -140 17752
rect -204 17608 -140 17672
rect -204 17528 -140 17592
rect 1208 18248 1272 18312
rect 1208 18168 1272 18232
rect 1208 18088 1272 18152
rect 1208 18008 1272 18072
rect 1208 17928 1272 17992
rect 1208 17848 1272 17912
rect 1208 17768 1272 17832
rect 1208 17688 1272 17752
rect 1208 17608 1272 17672
rect 1208 17528 1272 17592
rect 2620 18248 2684 18312
rect 2620 18168 2684 18232
rect 2620 18088 2684 18152
rect 2620 18008 2684 18072
rect 2620 17928 2684 17992
rect 2620 17848 2684 17912
rect 2620 17768 2684 17832
rect 2620 17688 2684 17752
rect 2620 17608 2684 17672
rect 2620 17528 2684 17592
rect 4032 18248 4096 18312
rect 4032 18168 4096 18232
rect 4032 18088 4096 18152
rect 4032 18008 4096 18072
rect 4032 17928 4096 17992
rect 4032 17848 4096 17912
rect 4032 17768 4096 17832
rect 4032 17688 4096 17752
rect 4032 17608 4096 17672
rect 4032 17528 4096 17592
rect 5444 18248 5508 18312
rect 5444 18168 5508 18232
rect 5444 18088 5508 18152
rect 5444 18008 5508 18072
rect 5444 17928 5508 17992
rect 5444 17848 5508 17912
rect 5444 17768 5508 17832
rect 5444 17688 5508 17752
rect 5444 17608 5508 17672
rect 5444 17528 5508 17592
rect 6856 18248 6920 18312
rect 6856 18168 6920 18232
rect 6856 18088 6920 18152
rect 6856 18008 6920 18072
rect 6856 17928 6920 17992
rect 6856 17848 6920 17912
rect 6856 17768 6920 17832
rect 6856 17688 6920 17752
rect 6856 17608 6920 17672
rect 6856 17528 6920 17592
rect 8268 18248 8332 18312
rect 8268 18168 8332 18232
rect 8268 18088 8332 18152
rect 8268 18008 8332 18072
rect 8268 17928 8332 17992
rect 8268 17848 8332 17912
rect 8268 17768 8332 17832
rect 8268 17688 8332 17752
rect 8268 17608 8332 17672
rect 8268 17528 8332 17592
rect 9680 18248 9744 18312
rect 9680 18168 9744 18232
rect 9680 18088 9744 18152
rect 9680 18008 9744 18072
rect 9680 17928 9744 17992
rect 9680 17848 9744 17912
rect 9680 17768 9744 17832
rect 9680 17688 9744 17752
rect 9680 17608 9744 17672
rect 9680 17528 9744 17592
rect 11092 18248 11156 18312
rect 11092 18168 11156 18232
rect 11092 18088 11156 18152
rect 11092 18008 11156 18072
rect 11092 17928 11156 17992
rect 11092 17848 11156 17912
rect 11092 17768 11156 17832
rect 11092 17688 11156 17752
rect 11092 17608 11156 17672
rect 11092 17528 11156 17592
rect 12504 18248 12568 18312
rect 12504 18168 12568 18232
rect 12504 18088 12568 18152
rect 12504 18008 12568 18072
rect 12504 17928 12568 17992
rect 12504 17848 12568 17912
rect 12504 17768 12568 17832
rect 12504 17688 12568 17752
rect 12504 17608 12568 17672
rect 12504 17528 12568 17592
rect 13916 18248 13980 18312
rect 13916 18168 13980 18232
rect 13916 18088 13980 18152
rect 13916 18008 13980 18072
rect 13916 17928 13980 17992
rect 13916 17848 13980 17912
rect 13916 17768 13980 17832
rect 13916 17688 13980 17752
rect 13916 17608 13980 17672
rect 13916 17528 13980 17592
rect 15328 18248 15392 18312
rect 15328 18168 15392 18232
rect 15328 18088 15392 18152
rect 15328 18008 15392 18072
rect 15328 17928 15392 17992
rect 15328 17848 15392 17912
rect 15328 17768 15392 17832
rect 15328 17688 15392 17752
rect 15328 17608 15392 17672
rect 15328 17528 15392 17592
rect 16740 18248 16804 18312
rect 16740 18168 16804 18232
rect 16740 18088 16804 18152
rect 16740 18008 16804 18072
rect 16740 17928 16804 17992
rect 16740 17848 16804 17912
rect 16740 17768 16804 17832
rect 16740 17688 16804 17752
rect 16740 17608 16804 17672
rect 16740 17528 16804 17592
rect 18152 18248 18216 18312
rect 18152 18168 18216 18232
rect 18152 18088 18216 18152
rect 18152 18008 18216 18072
rect 18152 17928 18216 17992
rect 18152 17848 18216 17912
rect 18152 17768 18216 17832
rect 18152 17688 18216 17752
rect 18152 17608 18216 17672
rect 18152 17528 18216 17592
rect 19564 18248 19628 18312
rect 19564 18168 19628 18232
rect 19564 18088 19628 18152
rect 19564 18008 19628 18072
rect 19564 17928 19628 17992
rect 19564 17848 19628 17912
rect 19564 17768 19628 17832
rect 19564 17688 19628 17752
rect 19564 17608 19628 17672
rect 19564 17528 19628 17592
rect 20976 18248 21040 18312
rect 20976 18168 21040 18232
rect 20976 18088 21040 18152
rect 20976 18008 21040 18072
rect 20976 17928 21040 17992
rect 20976 17848 21040 17912
rect 20976 17768 21040 17832
rect 20976 17688 21040 17752
rect 20976 17608 21040 17672
rect 20976 17528 21040 17592
rect 22388 18248 22452 18312
rect 22388 18168 22452 18232
rect 22388 18088 22452 18152
rect 22388 18008 22452 18072
rect 22388 17928 22452 17992
rect 22388 17848 22452 17912
rect 22388 17768 22452 17832
rect 22388 17688 22452 17752
rect 22388 17608 22452 17672
rect 22388 17528 22452 17592
rect 23800 18248 23864 18312
rect 23800 18168 23864 18232
rect 23800 18088 23864 18152
rect 23800 18008 23864 18072
rect 23800 17928 23864 17992
rect 23800 17848 23864 17912
rect 23800 17768 23864 17832
rect 23800 17688 23864 17752
rect 23800 17608 23864 17672
rect 23800 17528 23864 17592
rect -22796 17128 -22732 17192
rect -22796 17048 -22732 17112
rect -22796 16968 -22732 17032
rect -22796 16888 -22732 16952
rect -22796 16808 -22732 16872
rect -22796 16728 -22732 16792
rect -22796 16648 -22732 16712
rect -22796 16568 -22732 16632
rect -22796 16488 -22732 16552
rect -22796 16408 -22732 16472
rect -21384 17128 -21320 17192
rect -21384 17048 -21320 17112
rect -21384 16968 -21320 17032
rect -21384 16888 -21320 16952
rect -21384 16808 -21320 16872
rect -21384 16728 -21320 16792
rect -21384 16648 -21320 16712
rect -21384 16568 -21320 16632
rect -21384 16488 -21320 16552
rect -21384 16408 -21320 16472
rect -19972 17128 -19908 17192
rect -19972 17048 -19908 17112
rect -19972 16968 -19908 17032
rect -19972 16888 -19908 16952
rect -19972 16808 -19908 16872
rect -19972 16728 -19908 16792
rect -19972 16648 -19908 16712
rect -19972 16568 -19908 16632
rect -19972 16488 -19908 16552
rect -19972 16408 -19908 16472
rect -18560 17128 -18496 17192
rect -18560 17048 -18496 17112
rect -18560 16968 -18496 17032
rect -18560 16888 -18496 16952
rect -18560 16808 -18496 16872
rect -18560 16728 -18496 16792
rect -18560 16648 -18496 16712
rect -18560 16568 -18496 16632
rect -18560 16488 -18496 16552
rect -18560 16408 -18496 16472
rect -17148 17128 -17084 17192
rect -17148 17048 -17084 17112
rect -17148 16968 -17084 17032
rect -17148 16888 -17084 16952
rect -17148 16808 -17084 16872
rect -17148 16728 -17084 16792
rect -17148 16648 -17084 16712
rect -17148 16568 -17084 16632
rect -17148 16488 -17084 16552
rect -17148 16408 -17084 16472
rect -15736 17128 -15672 17192
rect -15736 17048 -15672 17112
rect -15736 16968 -15672 17032
rect -15736 16888 -15672 16952
rect -15736 16808 -15672 16872
rect -15736 16728 -15672 16792
rect -15736 16648 -15672 16712
rect -15736 16568 -15672 16632
rect -15736 16488 -15672 16552
rect -15736 16408 -15672 16472
rect -14324 17128 -14260 17192
rect -14324 17048 -14260 17112
rect -14324 16968 -14260 17032
rect -14324 16888 -14260 16952
rect -14324 16808 -14260 16872
rect -14324 16728 -14260 16792
rect -14324 16648 -14260 16712
rect -14324 16568 -14260 16632
rect -14324 16488 -14260 16552
rect -14324 16408 -14260 16472
rect -12912 17128 -12848 17192
rect -12912 17048 -12848 17112
rect -12912 16968 -12848 17032
rect -12912 16888 -12848 16952
rect -12912 16808 -12848 16872
rect -12912 16728 -12848 16792
rect -12912 16648 -12848 16712
rect -12912 16568 -12848 16632
rect -12912 16488 -12848 16552
rect -12912 16408 -12848 16472
rect -11500 17128 -11436 17192
rect -11500 17048 -11436 17112
rect -11500 16968 -11436 17032
rect -11500 16888 -11436 16952
rect -11500 16808 -11436 16872
rect -11500 16728 -11436 16792
rect -11500 16648 -11436 16712
rect -11500 16568 -11436 16632
rect -11500 16488 -11436 16552
rect -11500 16408 -11436 16472
rect -10088 17128 -10024 17192
rect -10088 17048 -10024 17112
rect -10088 16968 -10024 17032
rect -10088 16888 -10024 16952
rect -10088 16808 -10024 16872
rect -10088 16728 -10024 16792
rect -10088 16648 -10024 16712
rect -10088 16568 -10024 16632
rect -10088 16488 -10024 16552
rect -10088 16408 -10024 16472
rect -8676 17128 -8612 17192
rect -8676 17048 -8612 17112
rect -8676 16968 -8612 17032
rect -8676 16888 -8612 16952
rect -8676 16808 -8612 16872
rect -8676 16728 -8612 16792
rect -8676 16648 -8612 16712
rect -8676 16568 -8612 16632
rect -8676 16488 -8612 16552
rect -8676 16408 -8612 16472
rect -7264 17128 -7200 17192
rect -7264 17048 -7200 17112
rect -7264 16968 -7200 17032
rect -7264 16888 -7200 16952
rect -7264 16808 -7200 16872
rect -7264 16728 -7200 16792
rect -7264 16648 -7200 16712
rect -7264 16568 -7200 16632
rect -7264 16488 -7200 16552
rect -7264 16408 -7200 16472
rect -5852 17128 -5788 17192
rect -5852 17048 -5788 17112
rect -5852 16968 -5788 17032
rect -5852 16888 -5788 16952
rect -5852 16808 -5788 16872
rect -5852 16728 -5788 16792
rect -5852 16648 -5788 16712
rect -5852 16568 -5788 16632
rect -5852 16488 -5788 16552
rect -5852 16408 -5788 16472
rect -4440 17128 -4376 17192
rect -4440 17048 -4376 17112
rect -4440 16968 -4376 17032
rect -4440 16888 -4376 16952
rect -4440 16808 -4376 16872
rect -4440 16728 -4376 16792
rect -4440 16648 -4376 16712
rect -4440 16568 -4376 16632
rect -4440 16488 -4376 16552
rect -4440 16408 -4376 16472
rect -3028 17128 -2964 17192
rect -3028 17048 -2964 17112
rect -3028 16968 -2964 17032
rect -3028 16888 -2964 16952
rect -3028 16808 -2964 16872
rect -3028 16728 -2964 16792
rect -3028 16648 -2964 16712
rect -3028 16568 -2964 16632
rect -3028 16488 -2964 16552
rect -3028 16408 -2964 16472
rect -1616 17128 -1552 17192
rect -1616 17048 -1552 17112
rect -1616 16968 -1552 17032
rect -1616 16888 -1552 16952
rect -1616 16808 -1552 16872
rect -1616 16728 -1552 16792
rect -1616 16648 -1552 16712
rect -1616 16568 -1552 16632
rect -1616 16488 -1552 16552
rect -1616 16408 -1552 16472
rect -204 17128 -140 17192
rect -204 17048 -140 17112
rect -204 16968 -140 17032
rect -204 16888 -140 16952
rect -204 16808 -140 16872
rect -204 16728 -140 16792
rect -204 16648 -140 16712
rect -204 16568 -140 16632
rect -204 16488 -140 16552
rect -204 16408 -140 16472
rect 1208 17128 1272 17192
rect 1208 17048 1272 17112
rect 1208 16968 1272 17032
rect 1208 16888 1272 16952
rect 1208 16808 1272 16872
rect 1208 16728 1272 16792
rect 1208 16648 1272 16712
rect 1208 16568 1272 16632
rect 1208 16488 1272 16552
rect 1208 16408 1272 16472
rect 2620 17128 2684 17192
rect 2620 17048 2684 17112
rect 2620 16968 2684 17032
rect 2620 16888 2684 16952
rect 2620 16808 2684 16872
rect 2620 16728 2684 16792
rect 2620 16648 2684 16712
rect 2620 16568 2684 16632
rect 2620 16488 2684 16552
rect 2620 16408 2684 16472
rect 4032 17128 4096 17192
rect 4032 17048 4096 17112
rect 4032 16968 4096 17032
rect 4032 16888 4096 16952
rect 4032 16808 4096 16872
rect 4032 16728 4096 16792
rect 4032 16648 4096 16712
rect 4032 16568 4096 16632
rect 4032 16488 4096 16552
rect 4032 16408 4096 16472
rect 5444 17128 5508 17192
rect 5444 17048 5508 17112
rect 5444 16968 5508 17032
rect 5444 16888 5508 16952
rect 5444 16808 5508 16872
rect 5444 16728 5508 16792
rect 5444 16648 5508 16712
rect 5444 16568 5508 16632
rect 5444 16488 5508 16552
rect 5444 16408 5508 16472
rect 6856 17128 6920 17192
rect 6856 17048 6920 17112
rect 6856 16968 6920 17032
rect 6856 16888 6920 16952
rect 6856 16808 6920 16872
rect 6856 16728 6920 16792
rect 6856 16648 6920 16712
rect 6856 16568 6920 16632
rect 6856 16488 6920 16552
rect 6856 16408 6920 16472
rect 8268 17128 8332 17192
rect 8268 17048 8332 17112
rect 8268 16968 8332 17032
rect 8268 16888 8332 16952
rect 8268 16808 8332 16872
rect 8268 16728 8332 16792
rect 8268 16648 8332 16712
rect 8268 16568 8332 16632
rect 8268 16488 8332 16552
rect 8268 16408 8332 16472
rect 9680 17128 9744 17192
rect 9680 17048 9744 17112
rect 9680 16968 9744 17032
rect 9680 16888 9744 16952
rect 9680 16808 9744 16872
rect 9680 16728 9744 16792
rect 9680 16648 9744 16712
rect 9680 16568 9744 16632
rect 9680 16488 9744 16552
rect 9680 16408 9744 16472
rect 11092 17128 11156 17192
rect 11092 17048 11156 17112
rect 11092 16968 11156 17032
rect 11092 16888 11156 16952
rect 11092 16808 11156 16872
rect 11092 16728 11156 16792
rect 11092 16648 11156 16712
rect 11092 16568 11156 16632
rect 11092 16488 11156 16552
rect 11092 16408 11156 16472
rect 12504 17128 12568 17192
rect 12504 17048 12568 17112
rect 12504 16968 12568 17032
rect 12504 16888 12568 16952
rect 12504 16808 12568 16872
rect 12504 16728 12568 16792
rect 12504 16648 12568 16712
rect 12504 16568 12568 16632
rect 12504 16488 12568 16552
rect 12504 16408 12568 16472
rect 13916 17128 13980 17192
rect 13916 17048 13980 17112
rect 13916 16968 13980 17032
rect 13916 16888 13980 16952
rect 13916 16808 13980 16872
rect 13916 16728 13980 16792
rect 13916 16648 13980 16712
rect 13916 16568 13980 16632
rect 13916 16488 13980 16552
rect 13916 16408 13980 16472
rect 15328 17128 15392 17192
rect 15328 17048 15392 17112
rect 15328 16968 15392 17032
rect 15328 16888 15392 16952
rect 15328 16808 15392 16872
rect 15328 16728 15392 16792
rect 15328 16648 15392 16712
rect 15328 16568 15392 16632
rect 15328 16488 15392 16552
rect 15328 16408 15392 16472
rect 16740 17128 16804 17192
rect 16740 17048 16804 17112
rect 16740 16968 16804 17032
rect 16740 16888 16804 16952
rect 16740 16808 16804 16872
rect 16740 16728 16804 16792
rect 16740 16648 16804 16712
rect 16740 16568 16804 16632
rect 16740 16488 16804 16552
rect 16740 16408 16804 16472
rect 18152 17128 18216 17192
rect 18152 17048 18216 17112
rect 18152 16968 18216 17032
rect 18152 16888 18216 16952
rect 18152 16808 18216 16872
rect 18152 16728 18216 16792
rect 18152 16648 18216 16712
rect 18152 16568 18216 16632
rect 18152 16488 18216 16552
rect 18152 16408 18216 16472
rect 19564 17128 19628 17192
rect 19564 17048 19628 17112
rect 19564 16968 19628 17032
rect 19564 16888 19628 16952
rect 19564 16808 19628 16872
rect 19564 16728 19628 16792
rect 19564 16648 19628 16712
rect 19564 16568 19628 16632
rect 19564 16488 19628 16552
rect 19564 16408 19628 16472
rect 20976 17128 21040 17192
rect 20976 17048 21040 17112
rect 20976 16968 21040 17032
rect 20976 16888 21040 16952
rect 20976 16808 21040 16872
rect 20976 16728 21040 16792
rect 20976 16648 21040 16712
rect 20976 16568 21040 16632
rect 20976 16488 21040 16552
rect 20976 16408 21040 16472
rect 22388 17128 22452 17192
rect 22388 17048 22452 17112
rect 22388 16968 22452 17032
rect 22388 16888 22452 16952
rect 22388 16808 22452 16872
rect 22388 16728 22452 16792
rect 22388 16648 22452 16712
rect 22388 16568 22452 16632
rect 22388 16488 22452 16552
rect 22388 16408 22452 16472
rect 23800 17128 23864 17192
rect 23800 17048 23864 17112
rect 23800 16968 23864 17032
rect 23800 16888 23864 16952
rect 23800 16808 23864 16872
rect 23800 16728 23864 16792
rect 23800 16648 23864 16712
rect 23800 16568 23864 16632
rect 23800 16488 23864 16552
rect 23800 16408 23864 16472
rect -22796 16008 -22732 16072
rect -22796 15928 -22732 15992
rect -22796 15848 -22732 15912
rect -22796 15768 -22732 15832
rect -22796 15688 -22732 15752
rect -22796 15608 -22732 15672
rect -22796 15528 -22732 15592
rect -22796 15448 -22732 15512
rect -22796 15368 -22732 15432
rect -22796 15288 -22732 15352
rect -21384 16008 -21320 16072
rect -21384 15928 -21320 15992
rect -21384 15848 -21320 15912
rect -21384 15768 -21320 15832
rect -21384 15688 -21320 15752
rect -21384 15608 -21320 15672
rect -21384 15528 -21320 15592
rect -21384 15448 -21320 15512
rect -21384 15368 -21320 15432
rect -21384 15288 -21320 15352
rect -19972 16008 -19908 16072
rect -19972 15928 -19908 15992
rect -19972 15848 -19908 15912
rect -19972 15768 -19908 15832
rect -19972 15688 -19908 15752
rect -19972 15608 -19908 15672
rect -19972 15528 -19908 15592
rect -19972 15448 -19908 15512
rect -19972 15368 -19908 15432
rect -19972 15288 -19908 15352
rect -18560 16008 -18496 16072
rect -18560 15928 -18496 15992
rect -18560 15848 -18496 15912
rect -18560 15768 -18496 15832
rect -18560 15688 -18496 15752
rect -18560 15608 -18496 15672
rect -18560 15528 -18496 15592
rect -18560 15448 -18496 15512
rect -18560 15368 -18496 15432
rect -18560 15288 -18496 15352
rect -17148 16008 -17084 16072
rect -17148 15928 -17084 15992
rect -17148 15848 -17084 15912
rect -17148 15768 -17084 15832
rect -17148 15688 -17084 15752
rect -17148 15608 -17084 15672
rect -17148 15528 -17084 15592
rect -17148 15448 -17084 15512
rect -17148 15368 -17084 15432
rect -17148 15288 -17084 15352
rect -15736 16008 -15672 16072
rect -15736 15928 -15672 15992
rect -15736 15848 -15672 15912
rect -15736 15768 -15672 15832
rect -15736 15688 -15672 15752
rect -15736 15608 -15672 15672
rect -15736 15528 -15672 15592
rect -15736 15448 -15672 15512
rect -15736 15368 -15672 15432
rect -15736 15288 -15672 15352
rect -14324 16008 -14260 16072
rect -14324 15928 -14260 15992
rect -14324 15848 -14260 15912
rect -14324 15768 -14260 15832
rect -14324 15688 -14260 15752
rect -14324 15608 -14260 15672
rect -14324 15528 -14260 15592
rect -14324 15448 -14260 15512
rect -14324 15368 -14260 15432
rect -14324 15288 -14260 15352
rect -12912 16008 -12848 16072
rect -12912 15928 -12848 15992
rect -12912 15848 -12848 15912
rect -12912 15768 -12848 15832
rect -12912 15688 -12848 15752
rect -12912 15608 -12848 15672
rect -12912 15528 -12848 15592
rect -12912 15448 -12848 15512
rect -12912 15368 -12848 15432
rect -12912 15288 -12848 15352
rect -11500 16008 -11436 16072
rect -11500 15928 -11436 15992
rect -11500 15848 -11436 15912
rect -11500 15768 -11436 15832
rect -11500 15688 -11436 15752
rect -11500 15608 -11436 15672
rect -11500 15528 -11436 15592
rect -11500 15448 -11436 15512
rect -11500 15368 -11436 15432
rect -11500 15288 -11436 15352
rect -10088 16008 -10024 16072
rect -10088 15928 -10024 15992
rect -10088 15848 -10024 15912
rect -10088 15768 -10024 15832
rect -10088 15688 -10024 15752
rect -10088 15608 -10024 15672
rect -10088 15528 -10024 15592
rect -10088 15448 -10024 15512
rect -10088 15368 -10024 15432
rect -10088 15288 -10024 15352
rect -8676 16008 -8612 16072
rect -8676 15928 -8612 15992
rect -8676 15848 -8612 15912
rect -8676 15768 -8612 15832
rect -8676 15688 -8612 15752
rect -8676 15608 -8612 15672
rect -8676 15528 -8612 15592
rect -8676 15448 -8612 15512
rect -8676 15368 -8612 15432
rect -8676 15288 -8612 15352
rect -7264 16008 -7200 16072
rect -7264 15928 -7200 15992
rect -7264 15848 -7200 15912
rect -7264 15768 -7200 15832
rect -7264 15688 -7200 15752
rect -7264 15608 -7200 15672
rect -7264 15528 -7200 15592
rect -7264 15448 -7200 15512
rect -7264 15368 -7200 15432
rect -7264 15288 -7200 15352
rect -5852 16008 -5788 16072
rect -5852 15928 -5788 15992
rect -5852 15848 -5788 15912
rect -5852 15768 -5788 15832
rect -5852 15688 -5788 15752
rect -5852 15608 -5788 15672
rect -5852 15528 -5788 15592
rect -5852 15448 -5788 15512
rect -5852 15368 -5788 15432
rect -5852 15288 -5788 15352
rect -4440 16008 -4376 16072
rect -4440 15928 -4376 15992
rect -4440 15848 -4376 15912
rect -4440 15768 -4376 15832
rect -4440 15688 -4376 15752
rect -4440 15608 -4376 15672
rect -4440 15528 -4376 15592
rect -4440 15448 -4376 15512
rect -4440 15368 -4376 15432
rect -4440 15288 -4376 15352
rect -3028 16008 -2964 16072
rect -3028 15928 -2964 15992
rect -3028 15848 -2964 15912
rect -3028 15768 -2964 15832
rect -3028 15688 -2964 15752
rect -3028 15608 -2964 15672
rect -3028 15528 -2964 15592
rect -3028 15448 -2964 15512
rect -3028 15368 -2964 15432
rect -3028 15288 -2964 15352
rect -1616 16008 -1552 16072
rect -1616 15928 -1552 15992
rect -1616 15848 -1552 15912
rect -1616 15768 -1552 15832
rect -1616 15688 -1552 15752
rect -1616 15608 -1552 15672
rect -1616 15528 -1552 15592
rect -1616 15448 -1552 15512
rect -1616 15368 -1552 15432
rect -1616 15288 -1552 15352
rect -204 16008 -140 16072
rect -204 15928 -140 15992
rect -204 15848 -140 15912
rect -204 15768 -140 15832
rect -204 15688 -140 15752
rect -204 15608 -140 15672
rect -204 15528 -140 15592
rect -204 15448 -140 15512
rect -204 15368 -140 15432
rect -204 15288 -140 15352
rect 1208 16008 1272 16072
rect 1208 15928 1272 15992
rect 1208 15848 1272 15912
rect 1208 15768 1272 15832
rect 1208 15688 1272 15752
rect 1208 15608 1272 15672
rect 1208 15528 1272 15592
rect 1208 15448 1272 15512
rect 1208 15368 1272 15432
rect 1208 15288 1272 15352
rect 2620 16008 2684 16072
rect 2620 15928 2684 15992
rect 2620 15848 2684 15912
rect 2620 15768 2684 15832
rect 2620 15688 2684 15752
rect 2620 15608 2684 15672
rect 2620 15528 2684 15592
rect 2620 15448 2684 15512
rect 2620 15368 2684 15432
rect 2620 15288 2684 15352
rect 4032 16008 4096 16072
rect 4032 15928 4096 15992
rect 4032 15848 4096 15912
rect 4032 15768 4096 15832
rect 4032 15688 4096 15752
rect 4032 15608 4096 15672
rect 4032 15528 4096 15592
rect 4032 15448 4096 15512
rect 4032 15368 4096 15432
rect 4032 15288 4096 15352
rect 5444 16008 5508 16072
rect 5444 15928 5508 15992
rect 5444 15848 5508 15912
rect 5444 15768 5508 15832
rect 5444 15688 5508 15752
rect 5444 15608 5508 15672
rect 5444 15528 5508 15592
rect 5444 15448 5508 15512
rect 5444 15368 5508 15432
rect 5444 15288 5508 15352
rect 6856 16008 6920 16072
rect 6856 15928 6920 15992
rect 6856 15848 6920 15912
rect 6856 15768 6920 15832
rect 6856 15688 6920 15752
rect 6856 15608 6920 15672
rect 6856 15528 6920 15592
rect 6856 15448 6920 15512
rect 6856 15368 6920 15432
rect 6856 15288 6920 15352
rect 8268 16008 8332 16072
rect 8268 15928 8332 15992
rect 8268 15848 8332 15912
rect 8268 15768 8332 15832
rect 8268 15688 8332 15752
rect 8268 15608 8332 15672
rect 8268 15528 8332 15592
rect 8268 15448 8332 15512
rect 8268 15368 8332 15432
rect 8268 15288 8332 15352
rect 9680 16008 9744 16072
rect 9680 15928 9744 15992
rect 9680 15848 9744 15912
rect 9680 15768 9744 15832
rect 9680 15688 9744 15752
rect 9680 15608 9744 15672
rect 9680 15528 9744 15592
rect 9680 15448 9744 15512
rect 9680 15368 9744 15432
rect 9680 15288 9744 15352
rect 11092 16008 11156 16072
rect 11092 15928 11156 15992
rect 11092 15848 11156 15912
rect 11092 15768 11156 15832
rect 11092 15688 11156 15752
rect 11092 15608 11156 15672
rect 11092 15528 11156 15592
rect 11092 15448 11156 15512
rect 11092 15368 11156 15432
rect 11092 15288 11156 15352
rect 12504 16008 12568 16072
rect 12504 15928 12568 15992
rect 12504 15848 12568 15912
rect 12504 15768 12568 15832
rect 12504 15688 12568 15752
rect 12504 15608 12568 15672
rect 12504 15528 12568 15592
rect 12504 15448 12568 15512
rect 12504 15368 12568 15432
rect 12504 15288 12568 15352
rect 13916 16008 13980 16072
rect 13916 15928 13980 15992
rect 13916 15848 13980 15912
rect 13916 15768 13980 15832
rect 13916 15688 13980 15752
rect 13916 15608 13980 15672
rect 13916 15528 13980 15592
rect 13916 15448 13980 15512
rect 13916 15368 13980 15432
rect 13916 15288 13980 15352
rect 15328 16008 15392 16072
rect 15328 15928 15392 15992
rect 15328 15848 15392 15912
rect 15328 15768 15392 15832
rect 15328 15688 15392 15752
rect 15328 15608 15392 15672
rect 15328 15528 15392 15592
rect 15328 15448 15392 15512
rect 15328 15368 15392 15432
rect 15328 15288 15392 15352
rect 16740 16008 16804 16072
rect 16740 15928 16804 15992
rect 16740 15848 16804 15912
rect 16740 15768 16804 15832
rect 16740 15688 16804 15752
rect 16740 15608 16804 15672
rect 16740 15528 16804 15592
rect 16740 15448 16804 15512
rect 16740 15368 16804 15432
rect 16740 15288 16804 15352
rect 18152 16008 18216 16072
rect 18152 15928 18216 15992
rect 18152 15848 18216 15912
rect 18152 15768 18216 15832
rect 18152 15688 18216 15752
rect 18152 15608 18216 15672
rect 18152 15528 18216 15592
rect 18152 15448 18216 15512
rect 18152 15368 18216 15432
rect 18152 15288 18216 15352
rect 19564 16008 19628 16072
rect 19564 15928 19628 15992
rect 19564 15848 19628 15912
rect 19564 15768 19628 15832
rect 19564 15688 19628 15752
rect 19564 15608 19628 15672
rect 19564 15528 19628 15592
rect 19564 15448 19628 15512
rect 19564 15368 19628 15432
rect 19564 15288 19628 15352
rect 20976 16008 21040 16072
rect 20976 15928 21040 15992
rect 20976 15848 21040 15912
rect 20976 15768 21040 15832
rect 20976 15688 21040 15752
rect 20976 15608 21040 15672
rect 20976 15528 21040 15592
rect 20976 15448 21040 15512
rect 20976 15368 21040 15432
rect 20976 15288 21040 15352
rect 22388 16008 22452 16072
rect 22388 15928 22452 15992
rect 22388 15848 22452 15912
rect 22388 15768 22452 15832
rect 22388 15688 22452 15752
rect 22388 15608 22452 15672
rect 22388 15528 22452 15592
rect 22388 15448 22452 15512
rect 22388 15368 22452 15432
rect 22388 15288 22452 15352
rect 23800 16008 23864 16072
rect 23800 15928 23864 15992
rect 23800 15848 23864 15912
rect 23800 15768 23864 15832
rect 23800 15688 23864 15752
rect 23800 15608 23864 15672
rect 23800 15528 23864 15592
rect 23800 15448 23864 15512
rect 23800 15368 23864 15432
rect 23800 15288 23864 15352
rect -22796 14888 -22732 14952
rect -22796 14808 -22732 14872
rect -22796 14728 -22732 14792
rect -22796 14648 -22732 14712
rect -22796 14568 -22732 14632
rect -22796 14488 -22732 14552
rect -22796 14408 -22732 14472
rect -22796 14328 -22732 14392
rect -22796 14248 -22732 14312
rect -22796 14168 -22732 14232
rect -21384 14888 -21320 14952
rect -21384 14808 -21320 14872
rect -21384 14728 -21320 14792
rect -21384 14648 -21320 14712
rect -21384 14568 -21320 14632
rect -21384 14488 -21320 14552
rect -21384 14408 -21320 14472
rect -21384 14328 -21320 14392
rect -21384 14248 -21320 14312
rect -21384 14168 -21320 14232
rect -19972 14888 -19908 14952
rect -19972 14808 -19908 14872
rect -19972 14728 -19908 14792
rect -19972 14648 -19908 14712
rect -19972 14568 -19908 14632
rect -19972 14488 -19908 14552
rect -19972 14408 -19908 14472
rect -19972 14328 -19908 14392
rect -19972 14248 -19908 14312
rect -19972 14168 -19908 14232
rect -18560 14888 -18496 14952
rect -18560 14808 -18496 14872
rect -18560 14728 -18496 14792
rect -18560 14648 -18496 14712
rect -18560 14568 -18496 14632
rect -18560 14488 -18496 14552
rect -18560 14408 -18496 14472
rect -18560 14328 -18496 14392
rect -18560 14248 -18496 14312
rect -18560 14168 -18496 14232
rect -17148 14888 -17084 14952
rect -17148 14808 -17084 14872
rect -17148 14728 -17084 14792
rect -17148 14648 -17084 14712
rect -17148 14568 -17084 14632
rect -17148 14488 -17084 14552
rect -17148 14408 -17084 14472
rect -17148 14328 -17084 14392
rect -17148 14248 -17084 14312
rect -17148 14168 -17084 14232
rect -15736 14888 -15672 14952
rect -15736 14808 -15672 14872
rect -15736 14728 -15672 14792
rect -15736 14648 -15672 14712
rect -15736 14568 -15672 14632
rect -15736 14488 -15672 14552
rect -15736 14408 -15672 14472
rect -15736 14328 -15672 14392
rect -15736 14248 -15672 14312
rect -15736 14168 -15672 14232
rect -14324 14888 -14260 14952
rect -14324 14808 -14260 14872
rect -14324 14728 -14260 14792
rect -14324 14648 -14260 14712
rect -14324 14568 -14260 14632
rect -14324 14488 -14260 14552
rect -14324 14408 -14260 14472
rect -14324 14328 -14260 14392
rect -14324 14248 -14260 14312
rect -14324 14168 -14260 14232
rect -12912 14888 -12848 14952
rect -12912 14808 -12848 14872
rect -12912 14728 -12848 14792
rect -12912 14648 -12848 14712
rect -12912 14568 -12848 14632
rect -12912 14488 -12848 14552
rect -12912 14408 -12848 14472
rect -12912 14328 -12848 14392
rect -12912 14248 -12848 14312
rect -12912 14168 -12848 14232
rect -11500 14888 -11436 14952
rect -11500 14808 -11436 14872
rect -11500 14728 -11436 14792
rect -11500 14648 -11436 14712
rect -11500 14568 -11436 14632
rect -11500 14488 -11436 14552
rect -11500 14408 -11436 14472
rect -11500 14328 -11436 14392
rect -11500 14248 -11436 14312
rect -11500 14168 -11436 14232
rect -10088 14888 -10024 14952
rect -10088 14808 -10024 14872
rect -10088 14728 -10024 14792
rect -10088 14648 -10024 14712
rect -10088 14568 -10024 14632
rect -10088 14488 -10024 14552
rect -10088 14408 -10024 14472
rect -10088 14328 -10024 14392
rect -10088 14248 -10024 14312
rect -10088 14168 -10024 14232
rect -8676 14888 -8612 14952
rect -8676 14808 -8612 14872
rect -8676 14728 -8612 14792
rect -8676 14648 -8612 14712
rect -8676 14568 -8612 14632
rect -8676 14488 -8612 14552
rect -8676 14408 -8612 14472
rect -8676 14328 -8612 14392
rect -8676 14248 -8612 14312
rect -8676 14168 -8612 14232
rect -7264 14888 -7200 14952
rect -7264 14808 -7200 14872
rect -7264 14728 -7200 14792
rect -7264 14648 -7200 14712
rect -7264 14568 -7200 14632
rect -7264 14488 -7200 14552
rect -7264 14408 -7200 14472
rect -7264 14328 -7200 14392
rect -7264 14248 -7200 14312
rect -7264 14168 -7200 14232
rect -5852 14888 -5788 14952
rect -5852 14808 -5788 14872
rect -5852 14728 -5788 14792
rect -5852 14648 -5788 14712
rect -5852 14568 -5788 14632
rect -5852 14488 -5788 14552
rect -5852 14408 -5788 14472
rect -5852 14328 -5788 14392
rect -5852 14248 -5788 14312
rect -5852 14168 -5788 14232
rect -4440 14888 -4376 14952
rect -4440 14808 -4376 14872
rect -4440 14728 -4376 14792
rect -4440 14648 -4376 14712
rect -4440 14568 -4376 14632
rect -4440 14488 -4376 14552
rect -4440 14408 -4376 14472
rect -4440 14328 -4376 14392
rect -4440 14248 -4376 14312
rect -4440 14168 -4376 14232
rect -3028 14888 -2964 14952
rect -3028 14808 -2964 14872
rect -3028 14728 -2964 14792
rect -3028 14648 -2964 14712
rect -3028 14568 -2964 14632
rect -3028 14488 -2964 14552
rect -3028 14408 -2964 14472
rect -3028 14328 -2964 14392
rect -3028 14248 -2964 14312
rect -3028 14168 -2964 14232
rect -1616 14888 -1552 14952
rect -1616 14808 -1552 14872
rect -1616 14728 -1552 14792
rect -1616 14648 -1552 14712
rect -1616 14568 -1552 14632
rect -1616 14488 -1552 14552
rect -1616 14408 -1552 14472
rect -1616 14328 -1552 14392
rect -1616 14248 -1552 14312
rect -1616 14168 -1552 14232
rect -204 14888 -140 14952
rect -204 14808 -140 14872
rect -204 14728 -140 14792
rect -204 14648 -140 14712
rect -204 14568 -140 14632
rect -204 14488 -140 14552
rect -204 14408 -140 14472
rect -204 14328 -140 14392
rect -204 14248 -140 14312
rect -204 14168 -140 14232
rect 1208 14888 1272 14952
rect 1208 14808 1272 14872
rect 1208 14728 1272 14792
rect 1208 14648 1272 14712
rect 1208 14568 1272 14632
rect 1208 14488 1272 14552
rect 1208 14408 1272 14472
rect 1208 14328 1272 14392
rect 1208 14248 1272 14312
rect 1208 14168 1272 14232
rect 2620 14888 2684 14952
rect 2620 14808 2684 14872
rect 2620 14728 2684 14792
rect 2620 14648 2684 14712
rect 2620 14568 2684 14632
rect 2620 14488 2684 14552
rect 2620 14408 2684 14472
rect 2620 14328 2684 14392
rect 2620 14248 2684 14312
rect 2620 14168 2684 14232
rect 4032 14888 4096 14952
rect 4032 14808 4096 14872
rect 4032 14728 4096 14792
rect 4032 14648 4096 14712
rect 4032 14568 4096 14632
rect 4032 14488 4096 14552
rect 4032 14408 4096 14472
rect 4032 14328 4096 14392
rect 4032 14248 4096 14312
rect 4032 14168 4096 14232
rect 5444 14888 5508 14952
rect 5444 14808 5508 14872
rect 5444 14728 5508 14792
rect 5444 14648 5508 14712
rect 5444 14568 5508 14632
rect 5444 14488 5508 14552
rect 5444 14408 5508 14472
rect 5444 14328 5508 14392
rect 5444 14248 5508 14312
rect 5444 14168 5508 14232
rect 6856 14888 6920 14952
rect 6856 14808 6920 14872
rect 6856 14728 6920 14792
rect 6856 14648 6920 14712
rect 6856 14568 6920 14632
rect 6856 14488 6920 14552
rect 6856 14408 6920 14472
rect 6856 14328 6920 14392
rect 6856 14248 6920 14312
rect 6856 14168 6920 14232
rect 8268 14888 8332 14952
rect 8268 14808 8332 14872
rect 8268 14728 8332 14792
rect 8268 14648 8332 14712
rect 8268 14568 8332 14632
rect 8268 14488 8332 14552
rect 8268 14408 8332 14472
rect 8268 14328 8332 14392
rect 8268 14248 8332 14312
rect 8268 14168 8332 14232
rect 9680 14888 9744 14952
rect 9680 14808 9744 14872
rect 9680 14728 9744 14792
rect 9680 14648 9744 14712
rect 9680 14568 9744 14632
rect 9680 14488 9744 14552
rect 9680 14408 9744 14472
rect 9680 14328 9744 14392
rect 9680 14248 9744 14312
rect 9680 14168 9744 14232
rect 11092 14888 11156 14952
rect 11092 14808 11156 14872
rect 11092 14728 11156 14792
rect 11092 14648 11156 14712
rect 11092 14568 11156 14632
rect 11092 14488 11156 14552
rect 11092 14408 11156 14472
rect 11092 14328 11156 14392
rect 11092 14248 11156 14312
rect 11092 14168 11156 14232
rect 12504 14888 12568 14952
rect 12504 14808 12568 14872
rect 12504 14728 12568 14792
rect 12504 14648 12568 14712
rect 12504 14568 12568 14632
rect 12504 14488 12568 14552
rect 12504 14408 12568 14472
rect 12504 14328 12568 14392
rect 12504 14248 12568 14312
rect 12504 14168 12568 14232
rect 13916 14888 13980 14952
rect 13916 14808 13980 14872
rect 13916 14728 13980 14792
rect 13916 14648 13980 14712
rect 13916 14568 13980 14632
rect 13916 14488 13980 14552
rect 13916 14408 13980 14472
rect 13916 14328 13980 14392
rect 13916 14248 13980 14312
rect 13916 14168 13980 14232
rect 15328 14888 15392 14952
rect 15328 14808 15392 14872
rect 15328 14728 15392 14792
rect 15328 14648 15392 14712
rect 15328 14568 15392 14632
rect 15328 14488 15392 14552
rect 15328 14408 15392 14472
rect 15328 14328 15392 14392
rect 15328 14248 15392 14312
rect 15328 14168 15392 14232
rect 16740 14888 16804 14952
rect 16740 14808 16804 14872
rect 16740 14728 16804 14792
rect 16740 14648 16804 14712
rect 16740 14568 16804 14632
rect 16740 14488 16804 14552
rect 16740 14408 16804 14472
rect 16740 14328 16804 14392
rect 16740 14248 16804 14312
rect 16740 14168 16804 14232
rect 18152 14888 18216 14952
rect 18152 14808 18216 14872
rect 18152 14728 18216 14792
rect 18152 14648 18216 14712
rect 18152 14568 18216 14632
rect 18152 14488 18216 14552
rect 18152 14408 18216 14472
rect 18152 14328 18216 14392
rect 18152 14248 18216 14312
rect 18152 14168 18216 14232
rect 19564 14888 19628 14952
rect 19564 14808 19628 14872
rect 19564 14728 19628 14792
rect 19564 14648 19628 14712
rect 19564 14568 19628 14632
rect 19564 14488 19628 14552
rect 19564 14408 19628 14472
rect 19564 14328 19628 14392
rect 19564 14248 19628 14312
rect 19564 14168 19628 14232
rect 20976 14888 21040 14952
rect 20976 14808 21040 14872
rect 20976 14728 21040 14792
rect 20976 14648 21040 14712
rect 20976 14568 21040 14632
rect 20976 14488 21040 14552
rect 20976 14408 21040 14472
rect 20976 14328 21040 14392
rect 20976 14248 21040 14312
rect 20976 14168 21040 14232
rect 22388 14888 22452 14952
rect 22388 14808 22452 14872
rect 22388 14728 22452 14792
rect 22388 14648 22452 14712
rect 22388 14568 22452 14632
rect 22388 14488 22452 14552
rect 22388 14408 22452 14472
rect 22388 14328 22452 14392
rect 22388 14248 22452 14312
rect 22388 14168 22452 14232
rect 23800 14888 23864 14952
rect 23800 14808 23864 14872
rect 23800 14728 23864 14792
rect 23800 14648 23864 14712
rect 23800 14568 23864 14632
rect 23800 14488 23864 14552
rect 23800 14408 23864 14472
rect 23800 14328 23864 14392
rect 23800 14248 23864 14312
rect 23800 14168 23864 14232
rect -22796 13768 -22732 13832
rect -22796 13688 -22732 13752
rect -22796 13608 -22732 13672
rect -22796 13528 -22732 13592
rect -22796 13448 -22732 13512
rect -22796 13368 -22732 13432
rect -22796 13288 -22732 13352
rect -22796 13208 -22732 13272
rect -22796 13128 -22732 13192
rect -22796 13048 -22732 13112
rect -21384 13768 -21320 13832
rect -21384 13688 -21320 13752
rect -21384 13608 -21320 13672
rect -21384 13528 -21320 13592
rect -21384 13448 -21320 13512
rect -21384 13368 -21320 13432
rect -21384 13288 -21320 13352
rect -21384 13208 -21320 13272
rect -21384 13128 -21320 13192
rect -21384 13048 -21320 13112
rect -19972 13768 -19908 13832
rect -19972 13688 -19908 13752
rect -19972 13608 -19908 13672
rect -19972 13528 -19908 13592
rect -19972 13448 -19908 13512
rect -19972 13368 -19908 13432
rect -19972 13288 -19908 13352
rect -19972 13208 -19908 13272
rect -19972 13128 -19908 13192
rect -19972 13048 -19908 13112
rect -18560 13768 -18496 13832
rect -18560 13688 -18496 13752
rect -18560 13608 -18496 13672
rect -18560 13528 -18496 13592
rect -18560 13448 -18496 13512
rect -18560 13368 -18496 13432
rect -18560 13288 -18496 13352
rect -18560 13208 -18496 13272
rect -18560 13128 -18496 13192
rect -18560 13048 -18496 13112
rect -17148 13768 -17084 13832
rect -17148 13688 -17084 13752
rect -17148 13608 -17084 13672
rect -17148 13528 -17084 13592
rect -17148 13448 -17084 13512
rect -17148 13368 -17084 13432
rect -17148 13288 -17084 13352
rect -17148 13208 -17084 13272
rect -17148 13128 -17084 13192
rect -17148 13048 -17084 13112
rect -15736 13768 -15672 13832
rect -15736 13688 -15672 13752
rect -15736 13608 -15672 13672
rect -15736 13528 -15672 13592
rect -15736 13448 -15672 13512
rect -15736 13368 -15672 13432
rect -15736 13288 -15672 13352
rect -15736 13208 -15672 13272
rect -15736 13128 -15672 13192
rect -15736 13048 -15672 13112
rect -14324 13768 -14260 13832
rect -14324 13688 -14260 13752
rect -14324 13608 -14260 13672
rect -14324 13528 -14260 13592
rect -14324 13448 -14260 13512
rect -14324 13368 -14260 13432
rect -14324 13288 -14260 13352
rect -14324 13208 -14260 13272
rect -14324 13128 -14260 13192
rect -14324 13048 -14260 13112
rect -12912 13768 -12848 13832
rect -12912 13688 -12848 13752
rect -12912 13608 -12848 13672
rect -12912 13528 -12848 13592
rect -12912 13448 -12848 13512
rect -12912 13368 -12848 13432
rect -12912 13288 -12848 13352
rect -12912 13208 -12848 13272
rect -12912 13128 -12848 13192
rect -12912 13048 -12848 13112
rect -11500 13768 -11436 13832
rect -11500 13688 -11436 13752
rect -11500 13608 -11436 13672
rect -11500 13528 -11436 13592
rect -11500 13448 -11436 13512
rect -11500 13368 -11436 13432
rect -11500 13288 -11436 13352
rect -11500 13208 -11436 13272
rect -11500 13128 -11436 13192
rect -11500 13048 -11436 13112
rect -10088 13768 -10024 13832
rect -10088 13688 -10024 13752
rect -10088 13608 -10024 13672
rect -10088 13528 -10024 13592
rect -10088 13448 -10024 13512
rect -10088 13368 -10024 13432
rect -10088 13288 -10024 13352
rect -10088 13208 -10024 13272
rect -10088 13128 -10024 13192
rect -10088 13048 -10024 13112
rect -8676 13768 -8612 13832
rect -8676 13688 -8612 13752
rect -8676 13608 -8612 13672
rect -8676 13528 -8612 13592
rect -8676 13448 -8612 13512
rect -8676 13368 -8612 13432
rect -8676 13288 -8612 13352
rect -8676 13208 -8612 13272
rect -8676 13128 -8612 13192
rect -8676 13048 -8612 13112
rect -7264 13768 -7200 13832
rect -7264 13688 -7200 13752
rect -7264 13608 -7200 13672
rect -7264 13528 -7200 13592
rect -7264 13448 -7200 13512
rect -7264 13368 -7200 13432
rect -7264 13288 -7200 13352
rect -7264 13208 -7200 13272
rect -7264 13128 -7200 13192
rect -7264 13048 -7200 13112
rect -5852 13768 -5788 13832
rect -5852 13688 -5788 13752
rect -5852 13608 -5788 13672
rect -5852 13528 -5788 13592
rect -5852 13448 -5788 13512
rect -5852 13368 -5788 13432
rect -5852 13288 -5788 13352
rect -5852 13208 -5788 13272
rect -5852 13128 -5788 13192
rect -5852 13048 -5788 13112
rect -4440 13768 -4376 13832
rect -4440 13688 -4376 13752
rect -4440 13608 -4376 13672
rect -4440 13528 -4376 13592
rect -4440 13448 -4376 13512
rect -4440 13368 -4376 13432
rect -4440 13288 -4376 13352
rect -4440 13208 -4376 13272
rect -4440 13128 -4376 13192
rect -4440 13048 -4376 13112
rect -3028 13768 -2964 13832
rect -3028 13688 -2964 13752
rect -3028 13608 -2964 13672
rect -3028 13528 -2964 13592
rect -3028 13448 -2964 13512
rect -3028 13368 -2964 13432
rect -3028 13288 -2964 13352
rect -3028 13208 -2964 13272
rect -3028 13128 -2964 13192
rect -3028 13048 -2964 13112
rect -1616 13768 -1552 13832
rect -1616 13688 -1552 13752
rect -1616 13608 -1552 13672
rect -1616 13528 -1552 13592
rect -1616 13448 -1552 13512
rect -1616 13368 -1552 13432
rect -1616 13288 -1552 13352
rect -1616 13208 -1552 13272
rect -1616 13128 -1552 13192
rect -1616 13048 -1552 13112
rect -204 13768 -140 13832
rect -204 13688 -140 13752
rect -204 13608 -140 13672
rect -204 13528 -140 13592
rect -204 13448 -140 13512
rect -204 13368 -140 13432
rect -204 13288 -140 13352
rect -204 13208 -140 13272
rect -204 13128 -140 13192
rect -204 13048 -140 13112
rect 1208 13768 1272 13832
rect 1208 13688 1272 13752
rect 1208 13608 1272 13672
rect 1208 13528 1272 13592
rect 1208 13448 1272 13512
rect 1208 13368 1272 13432
rect 1208 13288 1272 13352
rect 1208 13208 1272 13272
rect 1208 13128 1272 13192
rect 1208 13048 1272 13112
rect 2620 13768 2684 13832
rect 2620 13688 2684 13752
rect 2620 13608 2684 13672
rect 2620 13528 2684 13592
rect 2620 13448 2684 13512
rect 2620 13368 2684 13432
rect 2620 13288 2684 13352
rect 2620 13208 2684 13272
rect 2620 13128 2684 13192
rect 2620 13048 2684 13112
rect 4032 13768 4096 13832
rect 4032 13688 4096 13752
rect 4032 13608 4096 13672
rect 4032 13528 4096 13592
rect 4032 13448 4096 13512
rect 4032 13368 4096 13432
rect 4032 13288 4096 13352
rect 4032 13208 4096 13272
rect 4032 13128 4096 13192
rect 4032 13048 4096 13112
rect 5444 13768 5508 13832
rect 5444 13688 5508 13752
rect 5444 13608 5508 13672
rect 5444 13528 5508 13592
rect 5444 13448 5508 13512
rect 5444 13368 5508 13432
rect 5444 13288 5508 13352
rect 5444 13208 5508 13272
rect 5444 13128 5508 13192
rect 5444 13048 5508 13112
rect 6856 13768 6920 13832
rect 6856 13688 6920 13752
rect 6856 13608 6920 13672
rect 6856 13528 6920 13592
rect 6856 13448 6920 13512
rect 6856 13368 6920 13432
rect 6856 13288 6920 13352
rect 6856 13208 6920 13272
rect 6856 13128 6920 13192
rect 6856 13048 6920 13112
rect 8268 13768 8332 13832
rect 8268 13688 8332 13752
rect 8268 13608 8332 13672
rect 8268 13528 8332 13592
rect 8268 13448 8332 13512
rect 8268 13368 8332 13432
rect 8268 13288 8332 13352
rect 8268 13208 8332 13272
rect 8268 13128 8332 13192
rect 8268 13048 8332 13112
rect 9680 13768 9744 13832
rect 9680 13688 9744 13752
rect 9680 13608 9744 13672
rect 9680 13528 9744 13592
rect 9680 13448 9744 13512
rect 9680 13368 9744 13432
rect 9680 13288 9744 13352
rect 9680 13208 9744 13272
rect 9680 13128 9744 13192
rect 9680 13048 9744 13112
rect 11092 13768 11156 13832
rect 11092 13688 11156 13752
rect 11092 13608 11156 13672
rect 11092 13528 11156 13592
rect 11092 13448 11156 13512
rect 11092 13368 11156 13432
rect 11092 13288 11156 13352
rect 11092 13208 11156 13272
rect 11092 13128 11156 13192
rect 11092 13048 11156 13112
rect 12504 13768 12568 13832
rect 12504 13688 12568 13752
rect 12504 13608 12568 13672
rect 12504 13528 12568 13592
rect 12504 13448 12568 13512
rect 12504 13368 12568 13432
rect 12504 13288 12568 13352
rect 12504 13208 12568 13272
rect 12504 13128 12568 13192
rect 12504 13048 12568 13112
rect 13916 13768 13980 13832
rect 13916 13688 13980 13752
rect 13916 13608 13980 13672
rect 13916 13528 13980 13592
rect 13916 13448 13980 13512
rect 13916 13368 13980 13432
rect 13916 13288 13980 13352
rect 13916 13208 13980 13272
rect 13916 13128 13980 13192
rect 13916 13048 13980 13112
rect 15328 13768 15392 13832
rect 15328 13688 15392 13752
rect 15328 13608 15392 13672
rect 15328 13528 15392 13592
rect 15328 13448 15392 13512
rect 15328 13368 15392 13432
rect 15328 13288 15392 13352
rect 15328 13208 15392 13272
rect 15328 13128 15392 13192
rect 15328 13048 15392 13112
rect 16740 13768 16804 13832
rect 16740 13688 16804 13752
rect 16740 13608 16804 13672
rect 16740 13528 16804 13592
rect 16740 13448 16804 13512
rect 16740 13368 16804 13432
rect 16740 13288 16804 13352
rect 16740 13208 16804 13272
rect 16740 13128 16804 13192
rect 16740 13048 16804 13112
rect 18152 13768 18216 13832
rect 18152 13688 18216 13752
rect 18152 13608 18216 13672
rect 18152 13528 18216 13592
rect 18152 13448 18216 13512
rect 18152 13368 18216 13432
rect 18152 13288 18216 13352
rect 18152 13208 18216 13272
rect 18152 13128 18216 13192
rect 18152 13048 18216 13112
rect 19564 13768 19628 13832
rect 19564 13688 19628 13752
rect 19564 13608 19628 13672
rect 19564 13528 19628 13592
rect 19564 13448 19628 13512
rect 19564 13368 19628 13432
rect 19564 13288 19628 13352
rect 19564 13208 19628 13272
rect 19564 13128 19628 13192
rect 19564 13048 19628 13112
rect 20976 13768 21040 13832
rect 20976 13688 21040 13752
rect 20976 13608 21040 13672
rect 20976 13528 21040 13592
rect 20976 13448 21040 13512
rect 20976 13368 21040 13432
rect 20976 13288 21040 13352
rect 20976 13208 21040 13272
rect 20976 13128 21040 13192
rect 20976 13048 21040 13112
rect 22388 13768 22452 13832
rect 22388 13688 22452 13752
rect 22388 13608 22452 13672
rect 22388 13528 22452 13592
rect 22388 13448 22452 13512
rect 22388 13368 22452 13432
rect 22388 13288 22452 13352
rect 22388 13208 22452 13272
rect 22388 13128 22452 13192
rect 22388 13048 22452 13112
rect 23800 13768 23864 13832
rect 23800 13688 23864 13752
rect 23800 13608 23864 13672
rect 23800 13528 23864 13592
rect 23800 13448 23864 13512
rect 23800 13368 23864 13432
rect 23800 13288 23864 13352
rect 23800 13208 23864 13272
rect 23800 13128 23864 13192
rect 23800 13048 23864 13112
rect -22796 12648 -22732 12712
rect -22796 12568 -22732 12632
rect -22796 12488 -22732 12552
rect -22796 12408 -22732 12472
rect -22796 12328 -22732 12392
rect -22796 12248 -22732 12312
rect -22796 12168 -22732 12232
rect -22796 12088 -22732 12152
rect -22796 12008 -22732 12072
rect -22796 11928 -22732 11992
rect -21384 12648 -21320 12712
rect -21384 12568 -21320 12632
rect -21384 12488 -21320 12552
rect -21384 12408 -21320 12472
rect -21384 12328 -21320 12392
rect -21384 12248 -21320 12312
rect -21384 12168 -21320 12232
rect -21384 12088 -21320 12152
rect -21384 12008 -21320 12072
rect -21384 11928 -21320 11992
rect -19972 12648 -19908 12712
rect -19972 12568 -19908 12632
rect -19972 12488 -19908 12552
rect -19972 12408 -19908 12472
rect -19972 12328 -19908 12392
rect -19972 12248 -19908 12312
rect -19972 12168 -19908 12232
rect -19972 12088 -19908 12152
rect -19972 12008 -19908 12072
rect -19972 11928 -19908 11992
rect -18560 12648 -18496 12712
rect -18560 12568 -18496 12632
rect -18560 12488 -18496 12552
rect -18560 12408 -18496 12472
rect -18560 12328 -18496 12392
rect -18560 12248 -18496 12312
rect -18560 12168 -18496 12232
rect -18560 12088 -18496 12152
rect -18560 12008 -18496 12072
rect -18560 11928 -18496 11992
rect -17148 12648 -17084 12712
rect -17148 12568 -17084 12632
rect -17148 12488 -17084 12552
rect -17148 12408 -17084 12472
rect -17148 12328 -17084 12392
rect -17148 12248 -17084 12312
rect -17148 12168 -17084 12232
rect -17148 12088 -17084 12152
rect -17148 12008 -17084 12072
rect -17148 11928 -17084 11992
rect -15736 12648 -15672 12712
rect -15736 12568 -15672 12632
rect -15736 12488 -15672 12552
rect -15736 12408 -15672 12472
rect -15736 12328 -15672 12392
rect -15736 12248 -15672 12312
rect -15736 12168 -15672 12232
rect -15736 12088 -15672 12152
rect -15736 12008 -15672 12072
rect -15736 11928 -15672 11992
rect -14324 12648 -14260 12712
rect -14324 12568 -14260 12632
rect -14324 12488 -14260 12552
rect -14324 12408 -14260 12472
rect -14324 12328 -14260 12392
rect -14324 12248 -14260 12312
rect -14324 12168 -14260 12232
rect -14324 12088 -14260 12152
rect -14324 12008 -14260 12072
rect -14324 11928 -14260 11992
rect -12912 12648 -12848 12712
rect -12912 12568 -12848 12632
rect -12912 12488 -12848 12552
rect -12912 12408 -12848 12472
rect -12912 12328 -12848 12392
rect -12912 12248 -12848 12312
rect -12912 12168 -12848 12232
rect -12912 12088 -12848 12152
rect -12912 12008 -12848 12072
rect -12912 11928 -12848 11992
rect -11500 12648 -11436 12712
rect -11500 12568 -11436 12632
rect -11500 12488 -11436 12552
rect -11500 12408 -11436 12472
rect -11500 12328 -11436 12392
rect -11500 12248 -11436 12312
rect -11500 12168 -11436 12232
rect -11500 12088 -11436 12152
rect -11500 12008 -11436 12072
rect -11500 11928 -11436 11992
rect -10088 12648 -10024 12712
rect -10088 12568 -10024 12632
rect -10088 12488 -10024 12552
rect -10088 12408 -10024 12472
rect -10088 12328 -10024 12392
rect -10088 12248 -10024 12312
rect -10088 12168 -10024 12232
rect -10088 12088 -10024 12152
rect -10088 12008 -10024 12072
rect -10088 11928 -10024 11992
rect -8676 12648 -8612 12712
rect -8676 12568 -8612 12632
rect -8676 12488 -8612 12552
rect -8676 12408 -8612 12472
rect -8676 12328 -8612 12392
rect -8676 12248 -8612 12312
rect -8676 12168 -8612 12232
rect -8676 12088 -8612 12152
rect -8676 12008 -8612 12072
rect -8676 11928 -8612 11992
rect -7264 12648 -7200 12712
rect -7264 12568 -7200 12632
rect -7264 12488 -7200 12552
rect -7264 12408 -7200 12472
rect -7264 12328 -7200 12392
rect -7264 12248 -7200 12312
rect -7264 12168 -7200 12232
rect -7264 12088 -7200 12152
rect -7264 12008 -7200 12072
rect -7264 11928 -7200 11992
rect -5852 12648 -5788 12712
rect -5852 12568 -5788 12632
rect -5852 12488 -5788 12552
rect -5852 12408 -5788 12472
rect -5852 12328 -5788 12392
rect -5852 12248 -5788 12312
rect -5852 12168 -5788 12232
rect -5852 12088 -5788 12152
rect -5852 12008 -5788 12072
rect -5852 11928 -5788 11992
rect -4440 12648 -4376 12712
rect -4440 12568 -4376 12632
rect -4440 12488 -4376 12552
rect -4440 12408 -4376 12472
rect -4440 12328 -4376 12392
rect -4440 12248 -4376 12312
rect -4440 12168 -4376 12232
rect -4440 12088 -4376 12152
rect -4440 12008 -4376 12072
rect -4440 11928 -4376 11992
rect -3028 12648 -2964 12712
rect -3028 12568 -2964 12632
rect -3028 12488 -2964 12552
rect -3028 12408 -2964 12472
rect -3028 12328 -2964 12392
rect -3028 12248 -2964 12312
rect -3028 12168 -2964 12232
rect -3028 12088 -2964 12152
rect -3028 12008 -2964 12072
rect -3028 11928 -2964 11992
rect -1616 12648 -1552 12712
rect -1616 12568 -1552 12632
rect -1616 12488 -1552 12552
rect -1616 12408 -1552 12472
rect -1616 12328 -1552 12392
rect -1616 12248 -1552 12312
rect -1616 12168 -1552 12232
rect -1616 12088 -1552 12152
rect -1616 12008 -1552 12072
rect -1616 11928 -1552 11992
rect -204 12648 -140 12712
rect -204 12568 -140 12632
rect -204 12488 -140 12552
rect -204 12408 -140 12472
rect -204 12328 -140 12392
rect -204 12248 -140 12312
rect -204 12168 -140 12232
rect -204 12088 -140 12152
rect -204 12008 -140 12072
rect -204 11928 -140 11992
rect 1208 12648 1272 12712
rect 1208 12568 1272 12632
rect 1208 12488 1272 12552
rect 1208 12408 1272 12472
rect 1208 12328 1272 12392
rect 1208 12248 1272 12312
rect 1208 12168 1272 12232
rect 1208 12088 1272 12152
rect 1208 12008 1272 12072
rect 1208 11928 1272 11992
rect 2620 12648 2684 12712
rect 2620 12568 2684 12632
rect 2620 12488 2684 12552
rect 2620 12408 2684 12472
rect 2620 12328 2684 12392
rect 2620 12248 2684 12312
rect 2620 12168 2684 12232
rect 2620 12088 2684 12152
rect 2620 12008 2684 12072
rect 2620 11928 2684 11992
rect 4032 12648 4096 12712
rect 4032 12568 4096 12632
rect 4032 12488 4096 12552
rect 4032 12408 4096 12472
rect 4032 12328 4096 12392
rect 4032 12248 4096 12312
rect 4032 12168 4096 12232
rect 4032 12088 4096 12152
rect 4032 12008 4096 12072
rect 4032 11928 4096 11992
rect 5444 12648 5508 12712
rect 5444 12568 5508 12632
rect 5444 12488 5508 12552
rect 5444 12408 5508 12472
rect 5444 12328 5508 12392
rect 5444 12248 5508 12312
rect 5444 12168 5508 12232
rect 5444 12088 5508 12152
rect 5444 12008 5508 12072
rect 5444 11928 5508 11992
rect 6856 12648 6920 12712
rect 6856 12568 6920 12632
rect 6856 12488 6920 12552
rect 6856 12408 6920 12472
rect 6856 12328 6920 12392
rect 6856 12248 6920 12312
rect 6856 12168 6920 12232
rect 6856 12088 6920 12152
rect 6856 12008 6920 12072
rect 6856 11928 6920 11992
rect 8268 12648 8332 12712
rect 8268 12568 8332 12632
rect 8268 12488 8332 12552
rect 8268 12408 8332 12472
rect 8268 12328 8332 12392
rect 8268 12248 8332 12312
rect 8268 12168 8332 12232
rect 8268 12088 8332 12152
rect 8268 12008 8332 12072
rect 8268 11928 8332 11992
rect 9680 12648 9744 12712
rect 9680 12568 9744 12632
rect 9680 12488 9744 12552
rect 9680 12408 9744 12472
rect 9680 12328 9744 12392
rect 9680 12248 9744 12312
rect 9680 12168 9744 12232
rect 9680 12088 9744 12152
rect 9680 12008 9744 12072
rect 9680 11928 9744 11992
rect 11092 12648 11156 12712
rect 11092 12568 11156 12632
rect 11092 12488 11156 12552
rect 11092 12408 11156 12472
rect 11092 12328 11156 12392
rect 11092 12248 11156 12312
rect 11092 12168 11156 12232
rect 11092 12088 11156 12152
rect 11092 12008 11156 12072
rect 11092 11928 11156 11992
rect 12504 12648 12568 12712
rect 12504 12568 12568 12632
rect 12504 12488 12568 12552
rect 12504 12408 12568 12472
rect 12504 12328 12568 12392
rect 12504 12248 12568 12312
rect 12504 12168 12568 12232
rect 12504 12088 12568 12152
rect 12504 12008 12568 12072
rect 12504 11928 12568 11992
rect 13916 12648 13980 12712
rect 13916 12568 13980 12632
rect 13916 12488 13980 12552
rect 13916 12408 13980 12472
rect 13916 12328 13980 12392
rect 13916 12248 13980 12312
rect 13916 12168 13980 12232
rect 13916 12088 13980 12152
rect 13916 12008 13980 12072
rect 13916 11928 13980 11992
rect 15328 12648 15392 12712
rect 15328 12568 15392 12632
rect 15328 12488 15392 12552
rect 15328 12408 15392 12472
rect 15328 12328 15392 12392
rect 15328 12248 15392 12312
rect 15328 12168 15392 12232
rect 15328 12088 15392 12152
rect 15328 12008 15392 12072
rect 15328 11928 15392 11992
rect 16740 12648 16804 12712
rect 16740 12568 16804 12632
rect 16740 12488 16804 12552
rect 16740 12408 16804 12472
rect 16740 12328 16804 12392
rect 16740 12248 16804 12312
rect 16740 12168 16804 12232
rect 16740 12088 16804 12152
rect 16740 12008 16804 12072
rect 16740 11928 16804 11992
rect 18152 12648 18216 12712
rect 18152 12568 18216 12632
rect 18152 12488 18216 12552
rect 18152 12408 18216 12472
rect 18152 12328 18216 12392
rect 18152 12248 18216 12312
rect 18152 12168 18216 12232
rect 18152 12088 18216 12152
rect 18152 12008 18216 12072
rect 18152 11928 18216 11992
rect 19564 12648 19628 12712
rect 19564 12568 19628 12632
rect 19564 12488 19628 12552
rect 19564 12408 19628 12472
rect 19564 12328 19628 12392
rect 19564 12248 19628 12312
rect 19564 12168 19628 12232
rect 19564 12088 19628 12152
rect 19564 12008 19628 12072
rect 19564 11928 19628 11992
rect 20976 12648 21040 12712
rect 20976 12568 21040 12632
rect 20976 12488 21040 12552
rect 20976 12408 21040 12472
rect 20976 12328 21040 12392
rect 20976 12248 21040 12312
rect 20976 12168 21040 12232
rect 20976 12088 21040 12152
rect 20976 12008 21040 12072
rect 20976 11928 21040 11992
rect 22388 12648 22452 12712
rect 22388 12568 22452 12632
rect 22388 12488 22452 12552
rect 22388 12408 22452 12472
rect 22388 12328 22452 12392
rect 22388 12248 22452 12312
rect 22388 12168 22452 12232
rect 22388 12088 22452 12152
rect 22388 12008 22452 12072
rect 22388 11928 22452 11992
rect 23800 12648 23864 12712
rect 23800 12568 23864 12632
rect 23800 12488 23864 12552
rect 23800 12408 23864 12472
rect 23800 12328 23864 12392
rect 23800 12248 23864 12312
rect 23800 12168 23864 12232
rect 23800 12088 23864 12152
rect 23800 12008 23864 12072
rect 23800 11928 23864 11992
rect -22796 11528 -22732 11592
rect -22796 11448 -22732 11512
rect -22796 11368 -22732 11432
rect -22796 11288 -22732 11352
rect -22796 11208 -22732 11272
rect -22796 11128 -22732 11192
rect -22796 11048 -22732 11112
rect -22796 10968 -22732 11032
rect -22796 10888 -22732 10952
rect -22796 10808 -22732 10872
rect -21384 11528 -21320 11592
rect -21384 11448 -21320 11512
rect -21384 11368 -21320 11432
rect -21384 11288 -21320 11352
rect -21384 11208 -21320 11272
rect -21384 11128 -21320 11192
rect -21384 11048 -21320 11112
rect -21384 10968 -21320 11032
rect -21384 10888 -21320 10952
rect -21384 10808 -21320 10872
rect -19972 11528 -19908 11592
rect -19972 11448 -19908 11512
rect -19972 11368 -19908 11432
rect -19972 11288 -19908 11352
rect -19972 11208 -19908 11272
rect -19972 11128 -19908 11192
rect -19972 11048 -19908 11112
rect -19972 10968 -19908 11032
rect -19972 10888 -19908 10952
rect -19972 10808 -19908 10872
rect -18560 11528 -18496 11592
rect -18560 11448 -18496 11512
rect -18560 11368 -18496 11432
rect -18560 11288 -18496 11352
rect -18560 11208 -18496 11272
rect -18560 11128 -18496 11192
rect -18560 11048 -18496 11112
rect -18560 10968 -18496 11032
rect -18560 10888 -18496 10952
rect -18560 10808 -18496 10872
rect -17148 11528 -17084 11592
rect -17148 11448 -17084 11512
rect -17148 11368 -17084 11432
rect -17148 11288 -17084 11352
rect -17148 11208 -17084 11272
rect -17148 11128 -17084 11192
rect -17148 11048 -17084 11112
rect -17148 10968 -17084 11032
rect -17148 10888 -17084 10952
rect -17148 10808 -17084 10872
rect -15736 11528 -15672 11592
rect -15736 11448 -15672 11512
rect -15736 11368 -15672 11432
rect -15736 11288 -15672 11352
rect -15736 11208 -15672 11272
rect -15736 11128 -15672 11192
rect -15736 11048 -15672 11112
rect -15736 10968 -15672 11032
rect -15736 10888 -15672 10952
rect -15736 10808 -15672 10872
rect -14324 11528 -14260 11592
rect -14324 11448 -14260 11512
rect -14324 11368 -14260 11432
rect -14324 11288 -14260 11352
rect -14324 11208 -14260 11272
rect -14324 11128 -14260 11192
rect -14324 11048 -14260 11112
rect -14324 10968 -14260 11032
rect -14324 10888 -14260 10952
rect -14324 10808 -14260 10872
rect -12912 11528 -12848 11592
rect -12912 11448 -12848 11512
rect -12912 11368 -12848 11432
rect -12912 11288 -12848 11352
rect -12912 11208 -12848 11272
rect -12912 11128 -12848 11192
rect -12912 11048 -12848 11112
rect -12912 10968 -12848 11032
rect -12912 10888 -12848 10952
rect -12912 10808 -12848 10872
rect -11500 11528 -11436 11592
rect -11500 11448 -11436 11512
rect -11500 11368 -11436 11432
rect -11500 11288 -11436 11352
rect -11500 11208 -11436 11272
rect -11500 11128 -11436 11192
rect -11500 11048 -11436 11112
rect -11500 10968 -11436 11032
rect -11500 10888 -11436 10952
rect -11500 10808 -11436 10872
rect -10088 11528 -10024 11592
rect -10088 11448 -10024 11512
rect -10088 11368 -10024 11432
rect -10088 11288 -10024 11352
rect -10088 11208 -10024 11272
rect -10088 11128 -10024 11192
rect -10088 11048 -10024 11112
rect -10088 10968 -10024 11032
rect -10088 10888 -10024 10952
rect -10088 10808 -10024 10872
rect -8676 11528 -8612 11592
rect -8676 11448 -8612 11512
rect -8676 11368 -8612 11432
rect -8676 11288 -8612 11352
rect -8676 11208 -8612 11272
rect -8676 11128 -8612 11192
rect -8676 11048 -8612 11112
rect -8676 10968 -8612 11032
rect -8676 10888 -8612 10952
rect -8676 10808 -8612 10872
rect -7264 11528 -7200 11592
rect -7264 11448 -7200 11512
rect -7264 11368 -7200 11432
rect -7264 11288 -7200 11352
rect -7264 11208 -7200 11272
rect -7264 11128 -7200 11192
rect -7264 11048 -7200 11112
rect -7264 10968 -7200 11032
rect -7264 10888 -7200 10952
rect -7264 10808 -7200 10872
rect -5852 11528 -5788 11592
rect -5852 11448 -5788 11512
rect -5852 11368 -5788 11432
rect -5852 11288 -5788 11352
rect -5852 11208 -5788 11272
rect -5852 11128 -5788 11192
rect -5852 11048 -5788 11112
rect -5852 10968 -5788 11032
rect -5852 10888 -5788 10952
rect -5852 10808 -5788 10872
rect -4440 11528 -4376 11592
rect -4440 11448 -4376 11512
rect -4440 11368 -4376 11432
rect -4440 11288 -4376 11352
rect -4440 11208 -4376 11272
rect -4440 11128 -4376 11192
rect -4440 11048 -4376 11112
rect -4440 10968 -4376 11032
rect -4440 10888 -4376 10952
rect -4440 10808 -4376 10872
rect -3028 11528 -2964 11592
rect -3028 11448 -2964 11512
rect -3028 11368 -2964 11432
rect -3028 11288 -2964 11352
rect -3028 11208 -2964 11272
rect -3028 11128 -2964 11192
rect -3028 11048 -2964 11112
rect -3028 10968 -2964 11032
rect -3028 10888 -2964 10952
rect -3028 10808 -2964 10872
rect -1616 11528 -1552 11592
rect -1616 11448 -1552 11512
rect -1616 11368 -1552 11432
rect -1616 11288 -1552 11352
rect -1616 11208 -1552 11272
rect -1616 11128 -1552 11192
rect -1616 11048 -1552 11112
rect -1616 10968 -1552 11032
rect -1616 10888 -1552 10952
rect -1616 10808 -1552 10872
rect -204 11528 -140 11592
rect -204 11448 -140 11512
rect -204 11368 -140 11432
rect -204 11288 -140 11352
rect -204 11208 -140 11272
rect -204 11128 -140 11192
rect -204 11048 -140 11112
rect -204 10968 -140 11032
rect -204 10888 -140 10952
rect -204 10808 -140 10872
rect 1208 11528 1272 11592
rect 1208 11448 1272 11512
rect 1208 11368 1272 11432
rect 1208 11288 1272 11352
rect 1208 11208 1272 11272
rect 1208 11128 1272 11192
rect 1208 11048 1272 11112
rect 1208 10968 1272 11032
rect 1208 10888 1272 10952
rect 1208 10808 1272 10872
rect 2620 11528 2684 11592
rect 2620 11448 2684 11512
rect 2620 11368 2684 11432
rect 2620 11288 2684 11352
rect 2620 11208 2684 11272
rect 2620 11128 2684 11192
rect 2620 11048 2684 11112
rect 2620 10968 2684 11032
rect 2620 10888 2684 10952
rect 2620 10808 2684 10872
rect 4032 11528 4096 11592
rect 4032 11448 4096 11512
rect 4032 11368 4096 11432
rect 4032 11288 4096 11352
rect 4032 11208 4096 11272
rect 4032 11128 4096 11192
rect 4032 11048 4096 11112
rect 4032 10968 4096 11032
rect 4032 10888 4096 10952
rect 4032 10808 4096 10872
rect 5444 11528 5508 11592
rect 5444 11448 5508 11512
rect 5444 11368 5508 11432
rect 5444 11288 5508 11352
rect 5444 11208 5508 11272
rect 5444 11128 5508 11192
rect 5444 11048 5508 11112
rect 5444 10968 5508 11032
rect 5444 10888 5508 10952
rect 5444 10808 5508 10872
rect 6856 11528 6920 11592
rect 6856 11448 6920 11512
rect 6856 11368 6920 11432
rect 6856 11288 6920 11352
rect 6856 11208 6920 11272
rect 6856 11128 6920 11192
rect 6856 11048 6920 11112
rect 6856 10968 6920 11032
rect 6856 10888 6920 10952
rect 6856 10808 6920 10872
rect 8268 11528 8332 11592
rect 8268 11448 8332 11512
rect 8268 11368 8332 11432
rect 8268 11288 8332 11352
rect 8268 11208 8332 11272
rect 8268 11128 8332 11192
rect 8268 11048 8332 11112
rect 8268 10968 8332 11032
rect 8268 10888 8332 10952
rect 8268 10808 8332 10872
rect 9680 11528 9744 11592
rect 9680 11448 9744 11512
rect 9680 11368 9744 11432
rect 9680 11288 9744 11352
rect 9680 11208 9744 11272
rect 9680 11128 9744 11192
rect 9680 11048 9744 11112
rect 9680 10968 9744 11032
rect 9680 10888 9744 10952
rect 9680 10808 9744 10872
rect 11092 11528 11156 11592
rect 11092 11448 11156 11512
rect 11092 11368 11156 11432
rect 11092 11288 11156 11352
rect 11092 11208 11156 11272
rect 11092 11128 11156 11192
rect 11092 11048 11156 11112
rect 11092 10968 11156 11032
rect 11092 10888 11156 10952
rect 11092 10808 11156 10872
rect 12504 11528 12568 11592
rect 12504 11448 12568 11512
rect 12504 11368 12568 11432
rect 12504 11288 12568 11352
rect 12504 11208 12568 11272
rect 12504 11128 12568 11192
rect 12504 11048 12568 11112
rect 12504 10968 12568 11032
rect 12504 10888 12568 10952
rect 12504 10808 12568 10872
rect 13916 11528 13980 11592
rect 13916 11448 13980 11512
rect 13916 11368 13980 11432
rect 13916 11288 13980 11352
rect 13916 11208 13980 11272
rect 13916 11128 13980 11192
rect 13916 11048 13980 11112
rect 13916 10968 13980 11032
rect 13916 10888 13980 10952
rect 13916 10808 13980 10872
rect 15328 11528 15392 11592
rect 15328 11448 15392 11512
rect 15328 11368 15392 11432
rect 15328 11288 15392 11352
rect 15328 11208 15392 11272
rect 15328 11128 15392 11192
rect 15328 11048 15392 11112
rect 15328 10968 15392 11032
rect 15328 10888 15392 10952
rect 15328 10808 15392 10872
rect 16740 11528 16804 11592
rect 16740 11448 16804 11512
rect 16740 11368 16804 11432
rect 16740 11288 16804 11352
rect 16740 11208 16804 11272
rect 16740 11128 16804 11192
rect 16740 11048 16804 11112
rect 16740 10968 16804 11032
rect 16740 10888 16804 10952
rect 16740 10808 16804 10872
rect 18152 11528 18216 11592
rect 18152 11448 18216 11512
rect 18152 11368 18216 11432
rect 18152 11288 18216 11352
rect 18152 11208 18216 11272
rect 18152 11128 18216 11192
rect 18152 11048 18216 11112
rect 18152 10968 18216 11032
rect 18152 10888 18216 10952
rect 18152 10808 18216 10872
rect 19564 11528 19628 11592
rect 19564 11448 19628 11512
rect 19564 11368 19628 11432
rect 19564 11288 19628 11352
rect 19564 11208 19628 11272
rect 19564 11128 19628 11192
rect 19564 11048 19628 11112
rect 19564 10968 19628 11032
rect 19564 10888 19628 10952
rect 19564 10808 19628 10872
rect 20976 11528 21040 11592
rect 20976 11448 21040 11512
rect 20976 11368 21040 11432
rect 20976 11288 21040 11352
rect 20976 11208 21040 11272
rect 20976 11128 21040 11192
rect 20976 11048 21040 11112
rect 20976 10968 21040 11032
rect 20976 10888 21040 10952
rect 20976 10808 21040 10872
rect 22388 11528 22452 11592
rect 22388 11448 22452 11512
rect 22388 11368 22452 11432
rect 22388 11288 22452 11352
rect 22388 11208 22452 11272
rect 22388 11128 22452 11192
rect 22388 11048 22452 11112
rect 22388 10968 22452 11032
rect 22388 10888 22452 10952
rect 22388 10808 22452 10872
rect 23800 11528 23864 11592
rect 23800 11448 23864 11512
rect 23800 11368 23864 11432
rect 23800 11288 23864 11352
rect 23800 11208 23864 11272
rect 23800 11128 23864 11192
rect 23800 11048 23864 11112
rect 23800 10968 23864 11032
rect 23800 10888 23864 10952
rect 23800 10808 23864 10872
rect -22796 10408 -22732 10472
rect -22796 10328 -22732 10392
rect -22796 10248 -22732 10312
rect -22796 10168 -22732 10232
rect -22796 10088 -22732 10152
rect -22796 10008 -22732 10072
rect -22796 9928 -22732 9992
rect -22796 9848 -22732 9912
rect -22796 9768 -22732 9832
rect -22796 9688 -22732 9752
rect -21384 10408 -21320 10472
rect -21384 10328 -21320 10392
rect -21384 10248 -21320 10312
rect -21384 10168 -21320 10232
rect -21384 10088 -21320 10152
rect -21384 10008 -21320 10072
rect -21384 9928 -21320 9992
rect -21384 9848 -21320 9912
rect -21384 9768 -21320 9832
rect -21384 9688 -21320 9752
rect -19972 10408 -19908 10472
rect -19972 10328 -19908 10392
rect -19972 10248 -19908 10312
rect -19972 10168 -19908 10232
rect -19972 10088 -19908 10152
rect -19972 10008 -19908 10072
rect -19972 9928 -19908 9992
rect -19972 9848 -19908 9912
rect -19972 9768 -19908 9832
rect -19972 9688 -19908 9752
rect -18560 10408 -18496 10472
rect -18560 10328 -18496 10392
rect -18560 10248 -18496 10312
rect -18560 10168 -18496 10232
rect -18560 10088 -18496 10152
rect -18560 10008 -18496 10072
rect -18560 9928 -18496 9992
rect -18560 9848 -18496 9912
rect -18560 9768 -18496 9832
rect -18560 9688 -18496 9752
rect -17148 10408 -17084 10472
rect -17148 10328 -17084 10392
rect -17148 10248 -17084 10312
rect -17148 10168 -17084 10232
rect -17148 10088 -17084 10152
rect -17148 10008 -17084 10072
rect -17148 9928 -17084 9992
rect -17148 9848 -17084 9912
rect -17148 9768 -17084 9832
rect -17148 9688 -17084 9752
rect -15736 10408 -15672 10472
rect -15736 10328 -15672 10392
rect -15736 10248 -15672 10312
rect -15736 10168 -15672 10232
rect -15736 10088 -15672 10152
rect -15736 10008 -15672 10072
rect -15736 9928 -15672 9992
rect -15736 9848 -15672 9912
rect -15736 9768 -15672 9832
rect -15736 9688 -15672 9752
rect -14324 10408 -14260 10472
rect -14324 10328 -14260 10392
rect -14324 10248 -14260 10312
rect -14324 10168 -14260 10232
rect -14324 10088 -14260 10152
rect -14324 10008 -14260 10072
rect -14324 9928 -14260 9992
rect -14324 9848 -14260 9912
rect -14324 9768 -14260 9832
rect -14324 9688 -14260 9752
rect -12912 10408 -12848 10472
rect -12912 10328 -12848 10392
rect -12912 10248 -12848 10312
rect -12912 10168 -12848 10232
rect -12912 10088 -12848 10152
rect -12912 10008 -12848 10072
rect -12912 9928 -12848 9992
rect -12912 9848 -12848 9912
rect -12912 9768 -12848 9832
rect -12912 9688 -12848 9752
rect -11500 10408 -11436 10472
rect -11500 10328 -11436 10392
rect -11500 10248 -11436 10312
rect -11500 10168 -11436 10232
rect -11500 10088 -11436 10152
rect -11500 10008 -11436 10072
rect -11500 9928 -11436 9992
rect -11500 9848 -11436 9912
rect -11500 9768 -11436 9832
rect -11500 9688 -11436 9752
rect -10088 10408 -10024 10472
rect -10088 10328 -10024 10392
rect -10088 10248 -10024 10312
rect -10088 10168 -10024 10232
rect -10088 10088 -10024 10152
rect -10088 10008 -10024 10072
rect -10088 9928 -10024 9992
rect -10088 9848 -10024 9912
rect -10088 9768 -10024 9832
rect -10088 9688 -10024 9752
rect -8676 10408 -8612 10472
rect -8676 10328 -8612 10392
rect -8676 10248 -8612 10312
rect -8676 10168 -8612 10232
rect -8676 10088 -8612 10152
rect -8676 10008 -8612 10072
rect -8676 9928 -8612 9992
rect -8676 9848 -8612 9912
rect -8676 9768 -8612 9832
rect -8676 9688 -8612 9752
rect -7264 10408 -7200 10472
rect -7264 10328 -7200 10392
rect -7264 10248 -7200 10312
rect -7264 10168 -7200 10232
rect -7264 10088 -7200 10152
rect -7264 10008 -7200 10072
rect -7264 9928 -7200 9992
rect -7264 9848 -7200 9912
rect -7264 9768 -7200 9832
rect -7264 9688 -7200 9752
rect -5852 10408 -5788 10472
rect -5852 10328 -5788 10392
rect -5852 10248 -5788 10312
rect -5852 10168 -5788 10232
rect -5852 10088 -5788 10152
rect -5852 10008 -5788 10072
rect -5852 9928 -5788 9992
rect -5852 9848 -5788 9912
rect -5852 9768 -5788 9832
rect -5852 9688 -5788 9752
rect -4440 10408 -4376 10472
rect -4440 10328 -4376 10392
rect -4440 10248 -4376 10312
rect -4440 10168 -4376 10232
rect -4440 10088 -4376 10152
rect -4440 10008 -4376 10072
rect -4440 9928 -4376 9992
rect -4440 9848 -4376 9912
rect -4440 9768 -4376 9832
rect -4440 9688 -4376 9752
rect -3028 10408 -2964 10472
rect -3028 10328 -2964 10392
rect -3028 10248 -2964 10312
rect -3028 10168 -2964 10232
rect -3028 10088 -2964 10152
rect -3028 10008 -2964 10072
rect -3028 9928 -2964 9992
rect -3028 9848 -2964 9912
rect -3028 9768 -2964 9832
rect -3028 9688 -2964 9752
rect -1616 10408 -1552 10472
rect -1616 10328 -1552 10392
rect -1616 10248 -1552 10312
rect -1616 10168 -1552 10232
rect -1616 10088 -1552 10152
rect -1616 10008 -1552 10072
rect -1616 9928 -1552 9992
rect -1616 9848 -1552 9912
rect -1616 9768 -1552 9832
rect -1616 9688 -1552 9752
rect -204 10408 -140 10472
rect -204 10328 -140 10392
rect -204 10248 -140 10312
rect -204 10168 -140 10232
rect -204 10088 -140 10152
rect -204 10008 -140 10072
rect -204 9928 -140 9992
rect -204 9848 -140 9912
rect -204 9768 -140 9832
rect -204 9688 -140 9752
rect 1208 10408 1272 10472
rect 1208 10328 1272 10392
rect 1208 10248 1272 10312
rect 1208 10168 1272 10232
rect 1208 10088 1272 10152
rect 1208 10008 1272 10072
rect 1208 9928 1272 9992
rect 1208 9848 1272 9912
rect 1208 9768 1272 9832
rect 1208 9688 1272 9752
rect 2620 10408 2684 10472
rect 2620 10328 2684 10392
rect 2620 10248 2684 10312
rect 2620 10168 2684 10232
rect 2620 10088 2684 10152
rect 2620 10008 2684 10072
rect 2620 9928 2684 9992
rect 2620 9848 2684 9912
rect 2620 9768 2684 9832
rect 2620 9688 2684 9752
rect 4032 10408 4096 10472
rect 4032 10328 4096 10392
rect 4032 10248 4096 10312
rect 4032 10168 4096 10232
rect 4032 10088 4096 10152
rect 4032 10008 4096 10072
rect 4032 9928 4096 9992
rect 4032 9848 4096 9912
rect 4032 9768 4096 9832
rect 4032 9688 4096 9752
rect 5444 10408 5508 10472
rect 5444 10328 5508 10392
rect 5444 10248 5508 10312
rect 5444 10168 5508 10232
rect 5444 10088 5508 10152
rect 5444 10008 5508 10072
rect 5444 9928 5508 9992
rect 5444 9848 5508 9912
rect 5444 9768 5508 9832
rect 5444 9688 5508 9752
rect 6856 10408 6920 10472
rect 6856 10328 6920 10392
rect 6856 10248 6920 10312
rect 6856 10168 6920 10232
rect 6856 10088 6920 10152
rect 6856 10008 6920 10072
rect 6856 9928 6920 9992
rect 6856 9848 6920 9912
rect 6856 9768 6920 9832
rect 6856 9688 6920 9752
rect 8268 10408 8332 10472
rect 8268 10328 8332 10392
rect 8268 10248 8332 10312
rect 8268 10168 8332 10232
rect 8268 10088 8332 10152
rect 8268 10008 8332 10072
rect 8268 9928 8332 9992
rect 8268 9848 8332 9912
rect 8268 9768 8332 9832
rect 8268 9688 8332 9752
rect 9680 10408 9744 10472
rect 9680 10328 9744 10392
rect 9680 10248 9744 10312
rect 9680 10168 9744 10232
rect 9680 10088 9744 10152
rect 9680 10008 9744 10072
rect 9680 9928 9744 9992
rect 9680 9848 9744 9912
rect 9680 9768 9744 9832
rect 9680 9688 9744 9752
rect 11092 10408 11156 10472
rect 11092 10328 11156 10392
rect 11092 10248 11156 10312
rect 11092 10168 11156 10232
rect 11092 10088 11156 10152
rect 11092 10008 11156 10072
rect 11092 9928 11156 9992
rect 11092 9848 11156 9912
rect 11092 9768 11156 9832
rect 11092 9688 11156 9752
rect 12504 10408 12568 10472
rect 12504 10328 12568 10392
rect 12504 10248 12568 10312
rect 12504 10168 12568 10232
rect 12504 10088 12568 10152
rect 12504 10008 12568 10072
rect 12504 9928 12568 9992
rect 12504 9848 12568 9912
rect 12504 9768 12568 9832
rect 12504 9688 12568 9752
rect 13916 10408 13980 10472
rect 13916 10328 13980 10392
rect 13916 10248 13980 10312
rect 13916 10168 13980 10232
rect 13916 10088 13980 10152
rect 13916 10008 13980 10072
rect 13916 9928 13980 9992
rect 13916 9848 13980 9912
rect 13916 9768 13980 9832
rect 13916 9688 13980 9752
rect 15328 10408 15392 10472
rect 15328 10328 15392 10392
rect 15328 10248 15392 10312
rect 15328 10168 15392 10232
rect 15328 10088 15392 10152
rect 15328 10008 15392 10072
rect 15328 9928 15392 9992
rect 15328 9848 15392 9912
rect 15328 9768 15392 9832
rect 15328 9688 15392 9752
rect 16740 10408 16804 10472
rect 16740 10328 16804 10392
rect 16740 10248 16804 10312
rect 16740 10168 16804 10232
rect 16740 10088 16804 10152
rect 16740 10008 16804 10072
rect 16740 9928 16804 9992
rect 16740 9848 16804 9912
rect 16740 9768 16804 9832
rect 16740 9688 16804 9752
rect 18152 10408 18216 10472
rect 18152 10328 18216 10392
rect 18152 10248 18216 10312
rect 18152 10168 18216 10232
rect 18152 10088 18216 10152
rect 18152 10008 18216 10072
rect 18152 9928 18216 9992
rect 18152 9848 18216 9912
rect 18152 9768 18216 9832
rect 18152 9688 18216 9752
rect 19564 10408 19628 10472
rect 19564 10328 19628 10392
rect 19564 10248 19628 10312
rect 19564 10168 19628 10232
rect 19564 10088 19628 10152
rect 19564 10008 19628 10072
rect 19564 9928 19628 9992
rect 19564 9848 19628 9912
rect 19564 9768 19628 9832
rect 19564 9688 19628 9752
rect 20976 10408 21040 10472
rect 20976 10328 21040 10392
rect 20976 10248 21040 10312
rect 20976 10168 21040 10232
rect 20976 10088 21040 10152
rect 20976 10008 21040 10072
rect 20976 9928 21040 9992
rect 20976 9848 21040 9912
rect 20976 9768 21040 9832
rect 20976 9688 21040 9752
rect 22388 10408 22452 10472
rect 22388 10328 22452 10392
rect 22388 10248 22452 10312
rect 22388 10168 22452 10232
rect 22388 10088 22452 10152
rect 22388 10008 22452 10072
rect 22388 9928 22452 9992
rect 22388 9848 22452 9912
rect 22388 9768 22452 9832
rect 22388 9688 22452 9752
rect 23800 10408 23864 10472
rect 23800 10328 23864 10392
rect 23800 10248 23864 10312
rect 23800 10168 23864 10232
rect 23800 10088 23864 10152
rect 23800 10008 23864 10072
rect 23800 9928 23864 9992
rect 23800 9848 23864 9912
rect 23800 9768 23864 9832
rect 23800 9688 23864 9752
rect -22796 9288 -22732 9352
rect -22796 9208 -22732 9272
rect -22796 9128 -22732 9192
rect -22796 9048 -22732 9112
rect -22796 8968 -22732 9032
rect -22796 8888 -22732 8952
rect -22796 8808 -22732 8872
rect -22796 8728 -22732 8792
rect -22796 8648 -22732 8712
rect -22796 8568 -22732 8632
rect -21384 9288 -21320 9352
rect -21384 9208 -21320 9272
rect -21384 9128 -21320 9192
rect -21384 9048 -21320 9112
rect -21384 8968 -21320 9032
rect -21384 8888 -21320 8952
rect -21384 8808 -21320 8872
rect -21384 8728 -21320 8792
rect -21384 8648 -21320 8712
rect -21384 8568 -21320 8632
rect -19972 9288 -19908 9352
rect -19972 9208 -19908 9272
rect -19972 9128 -19908 9192
rect -19972 9048 -19908 9112
rect -19972 8968 -19908 9032
rect -19972 8888 -19908 8952
rect -19972 8808 -19908 8872
rect -19972 8728 -19908 8792
rect -19972 8648 -19908 8712
rect -19972 8568 -19908 8632
rect -18560 9288 -18496 9352
rect -18560 9208 -18496 9272
rect -18560 9128 -18496 9192
rect -18560 9048 -18496 9112
rect -18560 8968 -18496 9032
rect -18560 8888 -18496 8952
rect -18560 8808 -18496 8872
rect -18560 8728 -18496 8792
rect -18560 8648 -18496 8712
rect -18560 8568 -18496 8632
rect -17148 9288 -17084 9352
rect -17148 9208 -17084 9272
rect -17148 9128 -17084 9192
rect -17148 9048 -17084 9112
rect -17148 8968 -17084 9032
rect -17148 8888 -17084 8952
rect -17148 8808 -17084 8872
rect -17148 8728 -17084 8792
rect -17148 8648 -17084 8712
rect -17148 8568 -17084 8632
rect -15736 9288 -15672 9352
rect -15736 9208 -15672 9272
rect -15736 9128 -15672 9192
rect -15736 9048 -15672 9112
rect -15736 8968 -15672 9032
rect -15736 8888 -15672 8952
rect -15736 8808 -15672 8872
rect -15736 8728 -15672 8792
rect -15736 8648 -15672 8712
rect -15736 8568 -15672 8632
rect -14324 9288 -14260 9352
rect -14324 9208 -14260 9272
rect -14324 9128 -14260 9192
rect -14324 9048 -14260 9112
rect -14324 8968 -14260 9032
rect -14324 8888 -14260 8952
rect -14324 8808 -14260 8872
rect -14324 8728 -14260 8792
rect -14324 8648 -14260 8712
rect -14324 8568 -14260 8632
rect -12912 9288 -12848 9352
rect -12912 9208 -12848 9272
rect -12912 9128 -12848 9192
rect -12912 9048 -12848 9112
rect -12912 8968 -12848 9032
rect -12912 8888 -12848 8952
rect -12912 8808 -12848 8872
rect -12912 8728 -12848 8792
rect -12912 8648 -12848 8712
rect -12912 8568 -12848 8632
rect -11500 9288 -11436 9352
rect -11500 9208 -11436 9272
rect -11500 9128 -11436 9192
rect -11500 9048 -11436 9112
rect -11500 8968 -11436 9032
rect -11500 8888 -11436 8952
rect -11500 8808 -11436 8872
rect -11500 8728 -11436 8792
rect -11500 8648 -11436 8712
rect -11500 8568 -11436 8632
rect -10088 9288 -10024 9352
rect -10088 9208 -10024 9272
rect -10088 9128 -10024 9192
rect -10088 9048 -10024 9112
rect -10088 8968 -10024 9032
rect -10088 8888 -10024 8952
rect -10088 8808 -10024 8872
rect -10088 8728 -10024 8792
rect -10088 8648 -10024 8712
rect -10088 8568 -10024 8632
rect -8676 9288 -8612 9352
rect -8676 9208 -8612 9272
rect -8676 9128 -8612 9192
rect -8676 9048 -8612 9112
rect -8676 8968 -8612 9032
rect -8676 8888 -8612 8952
rect -8676 8808 -8612 8872
rect -8676 8728 -8612 8792
rect -8676 8648 -8612 8712
rect -8676 8568 -8612 8632
rect -7264 9288 -7200 9352
rect -7264 9208 -7200 9272
rect -7264 9128 -7200 9192
rect -7264 9048 -7200 9112
rect -7264 8968 -7200 9032
rect -7264 8888 -7200 8952
rect -7264 8808 -7200 8872
rect -7264 8728 -7200 8792
rect -7264 8648 -7200 8712
rect -7264 8568 -7200 8632
rect -5852 9288 -5788 9352
rect -5852 9208 -5788 9272
rect -5852 9128 -5788 9192
rect -5852 9048 -5788 9112
rect -5852 8968 -5788 9032
rect -5852 8888 -5788 8952
rect -5852 8808 -5788 8872
rect -5852 8728 -5788 8792
rect -5852 8648 -5788 8712
rect -5852 8568 -5788 8632
rect -4440 9288 -4376 9352
rect -4440 9208 -4376 9272
rect -4440 9128 -4376 9192
rect -4440 9048 -4376 9112
rect -4440 8968 -4376 9032
rect -4440 8888 -4376 8952
rect -4440 8808 -4376 8872
rect -4440 8728 -4376 8792
rect -4440 8648 -4376 8712
rect -4440 8568 -4376 8632
rect -3028 9288 -2964 9352
rect -3028 9208 -2964 9272
rect -3028 9128 -2964 9192
rect -3028 9048 -2964 9112
rect -3028 8968 -2964 9032
rect -3028 8888 -2964 8952
rect -3028 8808 -2964 8872
rect -3028 8728 -2964 8792
rect -3028 8648 -2964 8712
rect -3028 8568 -2964 8632
rect -1616 9288 -1552 9352
rect -1616 9208 -1552 9272
rect -1616 9128 -1552 9192
rect -1616 9048 -1552 9112
rect -1616 8968 -1552 9032
rect -1616 8888 -1552 8952
rect -1616 8808 -1552 8872
rect -1616 8728 -1552 8792
rect -1616 8648 -1552 8712
rect -1616 8568 -1552 8632
rect -204 9288 -140 9352
rect -204 9208 -140 9272
rect -204 9128 -140 9192
rect -204 9048 -140 9112
rect -204 8968 -140 9032
rect -204 8888 -140 8952
rect -204 8808 -140 8872
rect -204 8728 -140 8792
rect -204 8648 -140 8712
rect -204 8568 -140 8632
rect 1208 9288 1272 9352
rect 1208 9208 1272 9272
rect 1208 9128 1272 9192
rect 1208 9048 1272 9112
rect 1208 8968 1272 9032
rect 1208 8888 1272 8952
rect 1208 8808 1272 8872
rect 1208 8728 1272 8792
rect 1208 8648 1272 8712
rect 1208 8568 1272 8632
rect 2620 9288 2684 9352
rect 2620 9208 2684 9272
rect 2620 9128 2684 9192
rect 2620 9048 2684 9112
rect 2620 8968 2684 9032
rect 2620 8888 2684 8952
rect 2620 8808 2684 8872
rect 2620 8728 2684 8792
rect 2620 8648 2684 8712
rect 2620 8568 2684 8632
rect 4032 9288 4096 9352
rect 4032 9208 4096 9272
rect 4032 9128 4096 9192
rect 4032 9048 4096 9112
rect 4032 8968 4096 9032
rect 4032 8888 4096 8952
rect 4032 8808 4096 8872
rect 4032 8728 4096 8792
rect 4032 8648 4096 8712
rect 4032 8568 4096 8632
rect 5444 9288 5508 9352
rect 5444 9208 5508 9272
rect 5444 9128 5508 9192
rect 5444 9048 5508 9112
rect 5444 8968 5508 9032
rect 5444 8888 5508 8952
rect 5444 8808 5508 8872
rect 5444 8728 5508 8792
rect 5444 8648 5508 8712
rect 5444 8568 5508 8632
rect 6856 9288 6920 9352
rect 6856 9208 6920 9272
rect 6856 9128 6920 9192
rect 6856 9048 6920 9112
rect 6856 8968 6920 9032
rect 6856 8888 6920 8952
rect 6856 8808 6920 8872
rect 6856 8728 6920 8792
rect 6856 8648 6920 8712
rect 6856 8568 6920 8632
rect 8268 9288 8332 9352
rect 8268 9208 8332 9272
rect 8268 9128 8332 9192
rect 8268 9048 8332 9112
rect 8268 8968 8332 9032
rect 8268 8888 8332 8952
rect 8268 8808 8332 8872
rect 8268 8728 8332 8792
rect 8268 8648 8332 8712
rect 8268 8568 8332 8632
rect 9680 9288 9744 9352
rect 9680 9208 9744 9272
rect 9680 9128 9744 9192
rect 9680 9048 9744 9112
rect 9680 8968 9744 9032
rect 9680 8888 9744 8952
rect 9680 8808 9744 8872
rect 9680 8728 9744 8792
rect 9680 8648 9744 8712
rect 9680 8568 9744 8632
rect 11092 9288 11156 9352
rect 11092 9208 11156 9272
rect 11092 9128 11156 9192
rect 11092 9048 11156 9112
rect 11092 8968 11156 9032
rect 11092 8888 11156 8952
rect 11092 8808 11156 8872
rect 11092 8728 11156 8792
rect 11092 8648 11156 8712
rect 11092 8568 11156 8632
rect 12504 9288 12568 9352
rect 12504 9208 12568 9272
rect 12504 9128 12568 9192
rect 12504 9048 12568 9112
rect 12504 8968 12568 9032
rect 12504 8888 12568 8952
rect 12504 8808 12568 8872
rect 12504 8728 12568 8792
rect 12504 8648 12568 8712
rect 12504 8568 12568 8632
rect 13916 9288 13980 9352
rect 13916 9208 13980 9272
rect 13916 9128 13980 9192
rect 13916 9048 13980 9112
rect 13916 8968 13980 9032
rect 13916 8888 13980 8952
rect 13916 8808 13980 8872
rect 13916 8728 13980 8792
rect 13916 8648 13980 8712
rect 13916 8568 13980 8632
rect 15328 9288 15392 9352
rect 15328 9208 15392 9272
rect 15328 9128 15392 9192
rect 15328 9048 15392 9112
rect 15328 8968 15392 9032
rect 15328 8888 15392 8952
rect 15328 8808 15392 8872
rect 15328 8728 15392 8792
rect 15328 8648 15392 8712
rect 15328 8568 15392 8632
rect 16740 9288 16804 9352
rect 16740 9208 16804 9272
rect 16740 9128 16804 9192
rect 16740 9048 16804 9112
rect 16740 8968 16804 9032
rect 16740 8888 16804 8952
rect 16740 8808 16804 8872
rect 16740 8728 16804 8792
rect 16740 8648 16804 8712
rect 16740 8568 16804 8632
rect 18152 9288 18216 9352
rect 18152 9208 18216 9272
rect 18152 9128 18216 9192
rect 18152 9048 18216 9112
rect 18152 8968 18216 9032
rect 18152 8888 18216 8952
rect 18152 8808 18216 8872
rect 18152 8728 18216 8792
rect 18152 8648 18216 8712
rect 18152 8568 18216 8632
rect 19564 9288 19628 9352
rect 19564 9208 19628 9272
rect 19564 9128 19628 9192
rect 19564 9048 19628 9112
rect 19564 8968 19628 9032
rect 19564 8888 19628 8952
rect 19564 8808 19628 8872
rect 19564 8728 19628 8792
rect 19564 8648 19628 8712
rect 19564 8568 19628 8632
rect 20976 9288 21040 9352
rect 20976 9208 21040 9272
rect 20976 9128 21040 9192
rect 20976 9048 21040 9112
rect 20976 8968 21040 9032
rect 20976 8888 21040 8952
rect 20976 8808 21040 8872
rect 20976 8728 21040 8792
rect 20976 8648 21040 8712
rect 20976 8568 21040 8632
rect 22388 9288 22452 9352
rect 22388 9208 22452 9272
rect 22388 9128 22452 9192
rect 22388 9048 22452 9112
rect 22388 8968 22452 9032
rect 22388 8888 22452 8952
rect 22388 8808 22452 8872
rect 22388 8728 22452 8792
rect 22388 8648 22452 8712
rect 22388 8568 22452 8632
rect 23800 9288 23864 9352
rect 23800 9208 23864 9272
rect 23800 9128 23864 9192
rect 23800 9048 23864 9112
rect 23800 8968 23864 9032
rect 23800 8888 23864 8952
rect 23800 8808 23864 8872
rect 23800 8728 23864 8792
rect 23800 8648 23864 8712
rect 23800 8568 23864 8632
rect -22796 8168 -22732 8232
rect -22796 8088 -22732 8152
rect -22796 8008 -22732 8072
rect -22796 7928 -22732 7992
rect -22796 7848 -22732 7912
rect -22796 7768 -22732 7832
rect -22796 7688 -22732 7752
rect -22796 7608 -22732 7672
rect -22796 7528 -22732 7592
rect -22796 7448 -22732 7512
rect -21384 8168 -21320 8232
rect -21384 8088 -21320 8152
rect -21384 8008 -21320 8072
rect -21384 7928 -21320 7992
rect -21384 7848 -21320 7912
rect -21384 7768 -21320 7832
rect -21384 7688 -21320 7752
rect -21384 7608 -21320 7672
rect -21384 7528 -21320 7592
rect -21384 7448 -21320 7512
rect -19972 8168 -19908 8232
rect -19972 8088 -19908 8152
rect -19972 8008 -19908 8072
rect -19972 7928 -19908 7992
rect -19972 7848 -19908 7912
rect -19972 7768 -19908 7832
rect -19972 7688 -19908 7752
rect -19972 7608 -19908 7672
rect -19972 7528 -19908 7592
rect -19972 7448 -19908 7512
rect -18560 8168 -18496 8232
rect -18560 8088 -18496 8152
rect -18560 8008 -18496 8072
rect -18560 7928 -18496 7992
rect -18560 7848 -18496 7912
rect -18560 7768 -18496 7832
rect -18560 7688 -18496 7752
rect -18560 7608 -18496 7672
rect -18560 7528 -18496 7592
rect -18560 7448 -18496 7512
rect -17148 8168 -17084 8232
rect -17148 8088 -17084 8152
rect -17148 8008 -17084 8072
rect -17148 7928 -17084 7992
rect -17148 7848 -17084 7912
rect -17148 7768 -17084 7832
rect -17148 7688 -17084 7752
rect -17148 7608 -17084 7672
rect -17148 7528 -17084 7592
rect -17148 7448 -17084 7512
rect -15736 8168 -15672 8232
rect -15736 8088 -15672 8152
rect -15736 8008 -15672 8072
rect -15736 7928 -15672 7992
rect -15736 7848 -15672 7912
rect -15736 7768 -15672 7832
rect -15736 7688 -15672 7752
rect -15736 7608 -15672 7672
rect -15736 7528 -15672 7592
rect -15736 7448 -15672 7512
rect -14324 8168 -14260 8232
rect -14324 8088 -14260 8152
rect -14324 8008 -14260 8072
rect -14324 7928 -14260 7992
rect -14324 7848 -14260 7912
rect -14324 7768 -14260 7832
rect -14324 7688 -14260 7752
rect -14324 7608 -14260 7672
rect -14324 7528 -14260 7592
rect -14324 7448 -14260 7512
rect -12912 8168 -12848 8232
rect -12912 8088 -12848 8152
rect -12912 8008 -12848 8072
rect -12912 7928 -12848 7992
rect -12912 7848 -12848 7912
rect -12912 7768 -12848 7832
rect -12912 7688 -12848 7752
rect -12912 7608 -12848 7672
rect -12912 7528 -12848 7592
rect -12912 7448 -12848 7512
rect -11500 8168 -11436 8232
rect -11500 8088 -11436 8152
rect -11500 8008 -11436 8072
rect -11500 7928 -11436 7992
rect -11500 7848 -11436 7912
rect -11500 7768 -11436 7832
rect -11500 7688 -11436 7752
rect -11500 7608 -11436 7672
rect -11500 7528 -11436 7592
rect -11500 7448 -11436 7512
rect -10088 8168 -10024 8232
rect -10088 8088 -10024 8152
rect -10088 8008 -10024 8072
rect -10088 7928 -10024 7992
rect -10088 7848 -10024 7912
rect -10088 7768 -10024 7832
rect -10088 7688 -10024 7752
rect -10088 7608 -10024 7672
rect -10088 7528 -10024 7592
rect -10088 7448 -10024 7512
rect -8676 8168 -8612 8232
rect -8676 8088 -8612 8152
rect -8676 8008 -8612 8072
rect -8676 7928 -8612 7992
rect -8676 7848 -8612 7912
rect -8676 7768 -8612 7832
rect -8676 7688 -8612 7752
rect -8676 7608 -8612 7672
rect -8676 7528 -8612 7592
rect -8676 7448 -8612 7512
rect -7264 8168 -7200 8232
rect -7264 8088 -7200 8152
rect -7264 8008 -7200 8072
rect -7264 7928 -7200 7992
rect -7264 7848 -7200 7912
rect -7264 7768 -7200 7832
rect -7264 7688 -7200 7752
rect -7264 7608 -7200 7672
rect -7264 7528 -7200 7592
rect -7264 7448 -7200 7512
rect -5852 8168 -5788 8232
rect -5852 8088 -5788 8152
rect -5852 8008 -5788 8072
rect -5852 7928 -5788 7992
rect -5852 7848 -5788 7912
rect -5852 7768 -5788 7832
rect -5852 7688 -5788 7752
rect -5852 7608 -5788 7672
rect -5852 7528 -5788 7592
rect -5852 7448 -5788 7512
rect -4440 8168 -4376 8232
rect -4440 8088 -4376 8152
rect -4440 8008 -4376 8072
rect -4440 7928 -4376 7992
rect -4440 7848 -4376 7912
rect -4440 7768 -4376 7832
rect -4440 7688 -4376 7752
rect -4440 7608 -4376 7672
rect -4440 7528 -4376 7592
rect -4440 7448 -4376 7512
rect -3028 8168 -2964 8232
rect -3028 8088 -2964 8152
rect -3028 8008 -2964 8072
rect -3028 7928 -2964 7992
rect -3028 7848 -2964 7912
rect -3028 7768 -2964 7832
rect -3028 7688 -2964 7752
rect -3028 7608 -2964 7672
rect -3028 7528 -2964 7592
rect -3028 7448 -2964 7512
rect -1616 8168 -1552 8232
rect -1616 8088 -1552 8152
rect -1616 8008 -1552 8072
rect -1616 7928 -1552 7992
rect -1616 7848 -1552 7912
rect -1616 7768 -1552 7832
rect -1616 7688 -1552 7752
rect -1616 7608 -1552 7672
rect -1616 7528 -1552 7592
rect -1616 7448 -1552 7512
rect -204 8168 -140 8232
rect -204 8088 -140 8152
rect -204 8008 -140 8072
rect -204 7928 -140 7992
rect -204 7848 -140 7912
rect -204 7768 -140 7832
rect -204 7688 -140 7752
rect -204 7608 -140 7672
rect -204 7528 -140 7592
rect -204 7448 -140 7512
rect 1208 8168 1272 8232
rect 1208 8088 1272 8152
rect 1208 8008 1272 8072
rect 1208 7928 1272 7992
rect 1208 7848 1272 7912
rect 1208 7768 1272 7832
rect 1208 7688 1272 7752
rect 1208 7608 1272 7672
rect 1208 7528 1272 7592
rect 1208 7448 1272 7512
rect 2620 8168 2684 8232
rect 2620 8088 2684 8152
rect 2620 8008 2684 8072
rect 2620 7928 2684 7992
rect 2620 7848 2684 7912
rect 2620 7768 2684 7832
rect 2620 7688 2684 7752
rect 2620 7608 2684 7672
rect 2620 7528 2684 7592
rect 2620 7448 2684 7512
rect 4032 8168 4096 8232
rect 4032 8088 4096 8152
rect 4032 8008 4096 8072
rect 4032 7928 4096 7992
rect 4032 7848 4096 7912
rect 4032 7768 4096 7832
rect 4032 7688 4096 7752
rect 4032 7608 4096 7672
rect 4032 7528 4096 7592
rect 4032 7448 4096 7512
rect 5444 8168 5508 8232
rect 5444 8088 5508 8152
rect 5444 8008 5508 8072
rect 5444 7928 5508 7992
rect 5444 7848 5508 7912
rect 5444 7768 5508 7832
rect 5444 7688 5508 7752
rect 5444 7608 5508 7672
rect 5444 7528 5508 7592
rect 5444 7448 5508 7512
rect 6856 8168 6920 8232
rect 6856 8088 6920 8152
rect 6856 8008 6920 8072
rect 6856 7928 6920 7992
rect 6856 7848 6920 7912
rect 6856 7768 6920 7832
rect 6856 7688 6920 7752
rect 6856 7608 6920 7672
rect 6856 7528 6920 7592
rect 6856 7448 6920 7512
rect 8268 8168 8332 8232
rect 8268 8088 8332 8152
rect 8268 8008 8332 8072
rect 8268 7928 8332 7992
rect 8268 7848 8332 7912
rect 8268 7768 8332 7832
rect 8268 7688 8332 7752
rect 8268 7608 8332 7672
rect 8268 7528 8332 7592
rect 8268 7448 8332 7512
rect 9680 8168 9744 8232
rect 9680 8088 9744 8152
rect 9680 8008 9744 8072
rect 9680 7928 9744 7992
rect 9680 7848 9744 7912
rect 9680 7768 9744 7832
rect 9680 7688 9744 7752
rect 9680 7608 9744 7672
rect 9680 7528 9744 7592
rect 9680 7448 9744 7512
rect 11092 8168 11156 8232
rect 11092 8088 11156 8152
rect 11092 8008 11156 8072
rect 11092 7928 11156 7992
rect 11092 7848 11156 7912
rect 11092 7768 11156 7832
rect 11092 7688 11156 7752
rect 11092 7608 11156 7672
rect 11092 7528 11156 7592
rect 11092 7448 11156 7512
rect 12504 8168 12568 8232
rect 12504 8088 12568 8152
rect 12504 8008 12568 8072
rect 12504 7928 12568 7992
rect 12504 7848 12568 7912
rect 12504 7768 12568 7832
rect 12504 7688 12568 7752
rect 12504 7608 12568 7672
rect 12504 7528 12568 7592
rect 12504 7448 12568 7512
rect 13916 8168 13980 8232
rect 13916 8088 13980 8152
rect 13916 8008 13980 8072
rect 13916 7928 13980 7992
rect 13916 7848 13980 7912
rect 13916 7768 13980 7832
rect 13916 7688 13980 7752
rect 13916 7608 13980 7672
rect 13916 7528 13980 7592
rect 13916 7448 13980 7512
rect 15328 8168 15392 8232
rect 15328 8088 15392 8152
rect 15328 8008 15392 8072
rect 15328 7928 15392 7992
rect 15328 7848 15392 7912
rect 15328 7768 15392 7832
rect 15328 7688 15392 7752
rect 15328 7608 15392 7672
rect 15328 7528 15392 7592
rect 15328 7448 15392 7512
rect 16740 8168 16804 8232
rect 16740 8088 16804 8152
rect 16740 8008 16804 8072
rect 16740 7928 16804 7992
rect 16740 7848 16804 7912
rect 16740 7768 16804 7832
rect 16740 7688 16804 7752
rect 16740 7608 16804 7672
rect 16740 7528 16804 7592
rect 16740 7448 16804 7512
rect 18152 8168 18216 8232
rect 18152 8088 18216 8152
rect 18152 8008 18216 8072
rect 18152 7928 18216 7992
rect 18152 7848 18216 7912
rect 18152 7768 18216 7832
rect 18152 7688 18216 7752
rect 18152 7608 18216 7672
rect 18152 7528 18216 7592
rect 18152 7448 18216 7512
rect 19564 8168 19628 8232
rect 19564 8088 19628 8152
rect 19564 8008 19628 8072
rect 19564 7928 19628 7992
rect 19564 7848 19628 7912
rect 19564 7768 19628 7832
rect 19564 7688 19628 7752
rect 19564 7608 19628 7672
rect 19564 7528 19628 7592
rect 19564 7448 19628 7512
rect 20976 8168 21040 8232
rect 20976 8088 21040 8152
rect 20976 8008 21040 8072
rect 20976 7928 21040 7992
rect 20976 7848 21040 7912
rect 20976 7768 21040 7832
rect 20976 7688 21040 7752
rect 20976 7608 21040 7672
rect 20976 7528 21040 7592
rect 20976 7448 21040 7512
rect 22388 8168 22452 8232
rect 22388 8088 22452 8152
rect 22388 8008 22452 8072
rect 22388 7928 22452 7992
rect 22388 7848 22452 7912
rect 22388 7768 22452 7832
rect 22388 7688 22452 7752
rect 22388 7608 22452 7672
rect 22388 7528 22452 7592
rect 22388 7448 22452 7512
rect 23800 8168 23864 8232
rect 23800 8088 23864 8152
rect 23800 8008 23864 8072
rect 23800 7928 23864 7992
rect 23800 7848 23864 7912
rect 23800 7768 23864 7832
rect 23800 7688 23864 7752
rect 23800 7608 23864 7672
rect 23800 7528 23864 7592
rect 23800 7448 23864 7512
rect -22796 7048 -22732 7112
rect -22796 6968 -22732 7032
rect -22796 6888 -22732 6952
rect -22796 6808 -22732 6872
rect -22796 6728 -22732 6792
rect -22796 6648 -22732 6712
rect -22796 6568 -22732 6632
rect -22796 6488 -22732 6552
rect -22796 6408 -22732 6472
rect -22796 6328 -22732 6392
rect -21384 7048 -21320 7112
rect -21384 6968 -21320 7032
rect -21384 6888 -21320 6952
rect -21384 6808 -21320 6872
rect -21384 6728 -21320 6792
rect -21384 6648 -21320 6712
rect -21384 6568 -21320 6632
rect -21384 6488 -21320 6552
rect -21384 6408 -21320 6472
rect -21384 6328 -21320 6392
rect -19972 7048 -19908 7112
rect -19972 6968 -19908 7032
rect -19972 6888 -19908 6952
rect -19972 6808 -19908 6872
rect -19972 6728 -19908 6792
rect -19972 6648 -19908 6712
rect -19972 6568 -19908 6632
rect -19972 6488 -19908 6552
rect -19972 6408 -19908 6472
rect -19972 6328 -19908 6392
rect -18560 7048 -18496 7112
rect -18560 6968 -18496 7032
rect -18560 6888 -18496 6952
rect -18560 6808 -18496 6872
rect -18560 6728 -18496 6792
rect -18560 6648 -18496 6712
rect -18560 6568 -18496 6632
rect -18560 6488 -18496 6552
rect -18560 6408 -18496 6472
rect -18560 6328 -18496 6392
rect -17148 7048 -17084 7112
rect -17148 6968 -17084 7032
rect -17148 6888 -17084 6952
rect -17148 6808 -17084 6872
rect -17148 6728 -17084 6792
rect -17148 6648 -17084 6712
rect -17148 6568 -17084 6632
rect -17148 6488 -17084 6552
rect -17148 6408 -17084 6472
rect -17148 6328 -17084 6392
rect -15736 7048 -15672 7112
rect -15736 6968 -15672 7032
rect -15736 6888 -15672 6952
rect -15736 6808 -15672 6872
rect -15736 6728 -15672 6792
rect -15736 6648 -15672 6712
rect -15736 6568 -15672 6632
rect -15736 6488 -15672 6552
rect -15736 6408 -15672 6472
rect -15736 6328 -15672 6392
rect -14324 7048 -14260 7112
rect -14324 6968 -14260 7032
rect -14324 6888 -14260 6952
rect -14324 6808 -14260 6872
rect -14324 6728 -14260 6792
rect -14324 6648 -14260 6712
rect -14324 6568 -14260 6632
rect -14324 6488 -14260 6552
rect -14324 6408 -14260 6472
rect -14324 6328 -14260 6392
rect -12912 7048 -12848 7112
rect -12912 6968 -12848 7032
rect -12912 6888 -12848 6952
rect -12912 6808 -12848 6872
rect -12912 6728 -12848 6792
rect -12912 6648 -12848 6712
rect -12912 6568 -12848 6632
rect -12912 6488 -12848 6552
rect -12912 6408 -12848 6472
rect -12912 6328 -12848 6392
rect -11500 7048 -11436 7112
rect -11500 6968 -11436 7032
rect -11500 6888 -11436 6952
rect -11500 6808 -11436 6872
rect -11500 6728 -11436 6792
rect -11500 6648 -11436 6712
rect -11500 6568 -11436 6632
rect -11500 6488 -11436 6552
rect -11500 6408 -11436 6472
rect -11500 6328 -11436 6392
rect -10088 7048 -10024 7112
rect -10088 6968 -10024 7032
rect -10088 6888 -10024 6952
rect -10088 6808 -10024 6872
rect -10088 6728 -10024 6792
rect -10088 6648 -10024 6712
rect -10088 6568 -10024 6632
rect -10088 6488 -10024 6552
rect -10088 6408 -10024 6472
rect -10088 6328 -10024 6392
rect -8676 7048 -8612 7112
rect -8676 6968 -8612 7032
rect -8676 6888 -8612 6952
rect -8676 6808 -8612 6872
rect -8676 6728 -8612 6792
rect -8676 6648 -8612 6712
rect -8676 6568 -8612 6632
rect -8676 6488 -8612 6552
rect -8676 6408 -8612 6472
rect -8676 6328 -8612 6392
rect -7264 7048 -7200 7112
rect -7264 6968 -7200 7032
rect -7264 6888 -7200 6952
rect -7264 6808 -7200 6872
rect -7264 6728 -7200 6792
rect -7264 6648 -7200 6712
rect -7264 6568 -7200 6632
rect -7264 6488 -7200 6552
rect -7264 6408 -7200 6472
rect -7264 6328 -7200 6392
rect -5852 7048 -5788 7112
rect -5852 6968 -5788 7032
rect -5852 6888 -5788 6952
rect -5852 6808 -5788 6872
rect -5852 6728 -5788 6792
rect -5852 6648 -5788 6712
rect -5852 6568 -5788 6632
rect -5852 6488 -5788 6552
rect -5852 6408 -5788 6472
rect -5852 6328 -5788 6392
rect -4440 7048 -4376 7112
rect -4440 6968 -4376 7032
rect -4440 6888 -4376 6952
rect -4440 6808 -4376 6872
rect -4440 6728 -4376 6792
rect -4440 6648 -4376 6712
rect -4440 6568 -4376 6632
rect -4440 6488 -4376 6552
rect -4440 6408 -4376 6472
rect -4440 6328 -4376 6392
rect -3028 7048 -2964 7112
rect -3028 6968 -2964 7032
rect -3028 6888 -2964 6952
rect -3028 6808 -2964 6872
rect -3028 6728 -2964 6792
rect -3028 6648 -2964 6712
rect -3028 6568 -2964 6632
rect -3028 6488 -2964 6552
rect -3028 6408 -2964 6472
rect -3028 6328 -2964 6392
rect -1616 7048 -1552 7112
rect -1616 6968 -1552 7032
rect -1616 6888 -1552 6952
rect -1616 6808 -1552 6872
rect -1616 6728 -1552 6792
rect -1616 6648 -1552 6712
rect -1616 6568 -1552 6632
rect -1616 6488 -1552 6552
rect -1616 6408 -1552 6472
rect -1616 6328 -1552 6392
rect -204 7048 -140 7112
rect -204 6968 -140 7032
rect -204 6888 -140 6952
rect -204 6808 -140 6872
rect -204 6728 -140 6792
rect -204 6648 -140 6712
rect -204 6568 -140 6632
rect -204 6488 -140 6552
rect -204 6408 -140 6472
rect -204 6328 -140 6392
rect 1208 7048 1272 7112
rect 1208 6968 1272 7032
rect 1208 6888 1272 6952
rect 1208 6808 1272 6872
rect 1208 6728 1272 6792
rect 1208 6648 1272 6712
rect 1208 6568 1272 6632
rect 1208 6488 1272 6552
rect 1208 6408 1272 6472
rect 1208 6328 1272 6392
rect 2620 7048 2684 7112
rect 2620 6968 2684 7032
rect 2620 6888 2684 6952
rect 2620 6808 2684 6872
rect 2620 6728 2684 6792
rect 2620 6648 2684 6712
rect 2620 6568 2684 6632
rect 2620 6488 2684 6552
rect 2620 6408 2684 6472
rect 2620 6328 2684 6392
rect 4032 7048 4096 7112
rect 4032 6968 4096 7032
rect 4032 6888 4096 6952
rect 4032 6808 4096 6872
rect 4032 6728 4096 6792
rect 4032 6648 4096 6712
rect 4032 6568 4096 6632
rect 4032 6488 4096 6552
rect 4032 6408 4096 6472
rect 4032 6328 4096 6392
rect 5444 7048 5508 7112
rect 5444 6968 5508 7032
rect 5444 6888 5508 6952
rect 5444 6808 5508 6872
rect 5444 6728 5508 6792
rect 5444 6648 5508 6712
rect 5444 6568 5508 6632
rect 5444 6488 5508 6552
rect 5444 6408 5508 6472
rect 5444 6328 5508 6392
rect 6856 7048 6920 7112
rect 6856 6968 6920 7032
rect 6856 6888 6920 6952
rect 6856 6808 6920 6872
rect 6856 6728 6920 6792
rect 6856 6648 6920 6712
rect 6856 6568 6920 6632
rect 6856 6488 6920 6552
rect 6856 6408 6920 6472
rect 6856 6328 6920 6392
rect 8268 7048 8332 7112
rect 8268 6968 8332 7032
rect 8268 6888 8332 6952
rect 8268 6808 8332 6872
rect 8268 6728 8332 6792
rect 8268 6648 8332 6712
rect 8268 6568 8332 6632
rect 8268 6488 8332 6552
rect 8268 6408 8332 6472
rect 8268 6328 8332 6392
rect 9680 7048 9744 7112
rect 9680 6968 9744 7032
rect 9680 6888 9744 6952
rect 9680 6808 9744 6872
rect 9680 6728 9744 6792
rect 9680 6648 9744 6712
rect 9680 6568 9744 6632
rect 9680 6488 9744 6552
rect 9680 6408 9744 6472
rect 9680 6328 9744 6392
rect 11092 7048 11156 7112
rect 11092 6968 11156 7032
rect 11092 6888 11156 6952
rect 11092 6808 11156 6872
rect 11092 6728 11156 6792
rect 11092 6648 11156 6712
rect 11092 6568 11156 6632
rect 11092 6488 11156 6552
rect 11092 6408 11156 6472
rect 11092 6328 11156 6392
rect 12504 7048 12568 7112
rect 12504 6968 12568 7032
rect 12504 6888 12568 6952
rect 12504 6808 12568 6872
rect 12504 6728 12568 6792
rect 12504 6648 12568 6712
rect 12504 6568 12568 6632
rect 12504 6488 12568 6552
rect 12504 6408 12568 6472
rect 12504 6328 12568 6392
rect 13916 7048 13980 7112
rect 13916 6968 13980 7032
rect 13916 6888 13980 6952
rect 13916 6808 13980 6872
rect 13916 6728 13980 6792
rect 13916 6648 13980 6712
rect 13916 6568 13980 6632
rect 13916 6488 13980 6552
rect 13916 6408 13980 6472
rect 13916 6328 13980 6392
rect 15328 7048 15392 7112
rect 15328 6968 15392 7032
rect 15328 6888 15392 6952
rect 15328 6808 15392 6872
rect 15328 6728 15392 6792
rect 15328 6648 15392 6712
rect 15328 6568 15392 6632
rect 15328 6488 15392 6552
rect 15328 6408 15392 6472
rect 15328 6328 15392 6392
rect 16740 7048 16804 7112
rect 16740 6968 16804 7032
rect 16740 6888 16804 6952
rect 16740 6808 16804 6872
rect 16740 6728 16804 6792
rect 16740 6648 16804 6712
rect 16740 6568 16804 6632
rect 16740 6488 16804 6552
rect 16740 6408 16804 6472
rect 16740 6328 16804 6392
rect 18152 7048 18216 7112
rect 18152 6968 18216 7032
rect 18152 6888 18216 6952
rect 18152 6808 18216 6872
rect 18152 6728 18216 6792
rect 18152 6648 18216 6712
rect 18152 6568 18216 6632
rect 18152 6488 18216 6552
rect 18152 6408 18216 6472
rect 18152 6328 18216 6392
rect 19564 7048 19628 7112
rect 19564 6968 19628 7032
rect 19564 6888 19628 6952
rect 19564 6808 19628 6872
rect 19564 6728 19628 6792
rect 19564 6648 19628 6712
rect 19564 6568 19628 6632
rect 19564 6488 19628 6552
rect 19564 6408 19628 6472
rect 19564 6328 19628 6392
rect 20976 7048 21040 7112
rect 20976 6968 21040 7032
rect 20976 6888 21040 6952
rect 20976 6808 21040 6872
rect 20976 6728 21040 6792
rect 20976 6648 21040 6712
rect 20976 6568 21040 6632
rect 20976 6488 21040 6552
rect 20976 6408 21040 6472
rect 20976 6328 21040 6392
rect 22388 7048 22452 7112
rect 22388 6968 22452 7032
rect 22388 6888 22452 6952
rect 22388 6808 22452 6872
rect 22388 6728 22452 6792
rect 22388 6648 22452 6712
rect 22388 6568 22452 6632
rect 22388 6488 22452 6552
rect 22388 6408 22452 6472
rect 22388 6328 22452 6392
rect 23800 7048 23864 7112
rect 23800 6968 23864 7032
rect 23800 6888 23864 6952
rect 23800 6808 23864 6872
rect 23800 6728 23864 6792
rect 23800 6648 23864 6712
rect 23800 6568 23864 6632
rect 23800 6488 23864 6552
rect 23800 6408 23864 6472
rect 23800 6328 23864 6392
rect -22796 5928 -22732 5992
rect -22796 5848 -22732 5912
rect -22796 5768 -22732 5832
rect -22796 5688 -22732 5752
rect -22796 5608 -22732 5672
rect -22796 5528 -22732 5592
rect -22796 5448 -22732 5512
rect -22796 5368 -22732 5432
rect -22796 5288 -22732 5352
rect -22796 5208 -22732 5272
rect -21384 5928 -21320 5992
rect -21384 5848 -21320 5912
rect -21384 5768 -21320 5832
rect -21384 5688 -21320 5752
rect -21384 5608 -21320 5672
rect -21384 5528 -21320 5592
rect -21384 5448 -21320 5512
rect -21384 5368 -21320 5432
rect -21384 5288 -21320 5352
rect -21384 5208 -21320 5272
rect -19972 5928 -19908 5992
rect -19972 5848 -19908 5912
rect -19972 5768 -19908 5832
rect -19972 5688 -19908 5752
rect -19972 5608 -19908 5672
rect -19972 5528 -19908 5592
rect -19972 5448 -19908 5512
rect -19972 5368 -19908 5432
rect -19972 5288 -19908 5352
rect -19972 5208 -19908 5272
rect -18560 5928 -18496 5992
rect -18560 5848 -18496 5912
rect -18560 5768 -18496 5832
rect -18560 5688 -18496 5752
rect -18560 5608 -18496 5672
rect -18560 5528 -18496 5592
rect -18560 5448 -18496 5512
rect -18560 5368 -18496 5432
rect -18560 5288 -18496 5352
rect -18560 5208 -18496 5272
rect -17148 5928 -17084 5992
rect -17148 5848 -17084 5912
rect -17148 5768 -17084 5832
rect -17148 5688 -17084 5752
rect -17148 5608 -17084 5672
rect -17148 5528 -17084 5592
rect -17148 5448 -17084 5512
rect -17148 5368 -17084 5432
rect -17148 5288 -17084 5352
rect -17148 5208 -17084 5272
rect -15736 5928 -15672 5992
rect -15736 5848 -15672 5912
rect -15736 5768 -15672 5832
rect -15736 5688 -15672 5752
rect -15736 5608 -15672 5672
rect -15736 5528 -15672 5592
rect -15736 5448 -15672 5512
rect -15736 5368 -15672 5432
rect -15736 5288 -15672 5352
rect -15736 5208 -15672 5272
rect -14324 5928 -14260 5992
rect -14324 5848 -14260 5912
rect -14324 5768 -14260 5832
rect -14324 5688 -14260 5752
rect -14324 5608 -14260 5672
rect -14324 5528 -14260 5592
rect -14324 5448 -14260 5512
rect -14324 5368 -14260 5432
rect -14324 5288 -14260 5352
rect -14324 5208 -14260 5272
rect -12912 5928 -12848 5992
rect -12912 5848 -12848 5912
rect -12912 5768 -12848 5832
rect -12912 5688 -12848 5752
rect -12912 5608 -12848 5672
rect -12912 5528 -12848 5592
rect -12912 5448 -12848 5512
rect -12912 5368 -12848 5432
rect -12912 5288 -12848 5352
rect -12912 5208 -12848 5272
rect -11500 5928 -11436 5992
rect -11500 5848 -11436 5912
rect -11500 5768 -11436 5832
rect -11500 5688 -11436 5752
rect -11500 5608 -11436 5672
rect -11500 5528 -11436 5592
rect -11500 5448 -11436 5512
rect -11500 5368 -11436 5432
rect -11500 5288 -11436 5352
rect -11500 5208 -11436 5272
rect -10088 5928 -10024 5992
rect -10088 5848 -10024 5912
rect -10088 5768 -10024 5832
rect -10088 5688 -10024 5752
rect -10088 5608 -10024 5672
rect -10088 5528 -10024 5592
rect -10088 5448 -10024 5512
rect -10088 5368 -10024 5432
rect -10088 5288 -10024 5352
rect -10088 5208 -10024 5272
rect -8676 5928 -8612 5992
rect -8676 5848 -8612 5912
rect -8676 5768 -8612 5832
rect -8676 5688 -8612 5752
rect -8676 5608 -8612 5672
rect -8676 5528 -8612 5592
rect -8676 5448 -8612 5512
rect -8676 5368 -8612 5432
rect -8676 5288 -8612 5352
rect -8676 5208 -8612 5272
rect -7264 5928 -7200 5992
rect -7264 5848 -7200 5912
rect -7264 5768 -7200 5832
rect -7264 5688 -7200 5752
rect -7264 5608 -7200 5672
rect -7264 5528 -7200 5592
rect -7264 5448 -7200 5512
rect -7264 5368 -7200 5432
rect -7264 5288 -7200 5352
rect -7264 5208 -7200 5272
rect -5852 5928 -5788 5992
rect -5852 5848 -5788 5912
rect -5852 5768 -5788 5832
rect -5852 5688 -5788 5752
rect -5852 5608 -5788 5672
rect -5852 5528 -5788 5592
rect -5852 5448 -5788 5512
rect -5852 5368 -5788 5432
rect -5852 5288 -5788 5352
rect -5852 5208 -5788 5272
rect -4440 5928 -4376 5992
rect -4440 5848 -4376 5912
rect -4440 5768 -4376 5832
rect -4440 5688 -4376 5752
rect -4440 5608 -4376 5672
rect -4440 5528 -4376 5592
rect -4440 5448 -4376 5512
rect -4440 5368 -4376 5432
rect -4440 5288 -4376 5352
rect -4440 5208 -4376 5272
rect -3028 5928 -2964 5992
rect -3028 5848 -2964 5912
rect -3028 5768 -2964 5832
rect -3028 5688 -2964 5752
rect -3028 5608 -2964 5672
rect -3028 5528 -2964 5592
rect -3028 5448 -2964 5512
rect -3028 5368 -2964 5432
rect -3028 5288 -2964 5352
rect -3028 5208 -2964 5272
rect -1616 5928 -1552 5992
rect -1616 5848 -1552 5912
rect -1616 5768 -1552 5832
rect -1616 5688 -1552 5752
rect -1616 5608 -1552 5672
rect -1616 5528 -1552 5592
rect -1616 5448 -1552 5512
rect -1616 5368 -1552 5432
rect -1616 5288 -1552 5352
rect -1616 5208 -1552 5272
rect -204 5928 -140 5992
rect -204 5848 -140 5912
rect -204 5768 -140 5832
rect -204 5688 -140 5752
rect -204 5608 -140 5672
rect -204 5528 -140 5592
rect -204 5448 -140 5512
rect -204 5368 -140 5432
rect -204 5288 -140 5352
rect -204 5208 -140 5272
rect 1208 5928 1272 5992
rect 1208 5848 1272 5912
rect 1208 5768 1272 5832
rect 1208 5688 1272 5752
rect 1208 5608 1272 5672
rect 1208 5528 1272 5592
rect 1208 5448 1272 5512
rect 1208 5368 1272 5432
rect 1208 5288 1272 5352
rect 1208 5208 1272 5272
rect 2620 5928 2684 5992
rect 2620 5848 2684 5912
rect 2620 5768 2684 5832
rect 2620 5688 2684 5752
rect 2620 5608 2684 5672
rect 2620 5528 2684 5592
rect 2620 5448 2684 5512
rect 2620 5368 2684 5432
rect 2620 5288 2684 5352
rect 2620 5208 2684 5272
rect 4032 5928 4096 5992
rect 4032 5848 4096 5912
rect 4032 5768 4096 5832
rect 4032 5688 4096 5752
rect 4032 5608 4096 5672
rect 4032 5528 4096 5592
rect 4032 5448 4096 5512
rect 4032 5368 4096 5432
rect 4032 5288 4096 5352
rect 4032 5208 4096 5272
rect 5444 5928 5508 5992
rect 5444 5848 5508 5912
rect 5444 5768 5508 5832
rect 5444 5688 5508 5752
rect 5444 5608 5508 5672
rect 5444 5528 5508 5592
rect 5444 5448 5508 5512
rect 5444 5368 5508 5432
rect 5444 5288 5508 5352
rect 5444 5208 5508 5272
rect 6856 5928 6920 5992
rect 6856 5848 6920 5912
rect 6856 5768 6920 5832
rect 6856 5688 6920 5752
rect 6856 5608 6920 5672
rect 6856 5528 6920 5592
rect 6856 5448 6920 5512
rect 6856 5368 6920 5432
rect 6856 5288 6920 5352
rect 6856 5208 6920 5272
rect 8268 5928 8332 5992
rect 8268 5848 8332 5912
rect 8268 5768 8332 5832
rect 8268 5688 8332 5752
rect 8268 5608 8332 5672
rect 8268 5528 8332 5592
rect 8268 5448 8332 5512
rect 8268 5368 8332 5432
rect 8268 5288 8332 5352
rect 8268 5208 8332 5272
rect 9680 5928 9744 5992
rect 9680 5848 9744 5912
rect 9680 5768 9744 5832
rect 9680 5688 9744 5752
rect 9680 5608 9744 5672
rect 9680 5528 9744 5592
rect 9680 5448 9744 5512
rect 9680 5368 9744 5432
rect 9680 5288 9744 5352
rect 9680 5208 9744 5272
rect 11092 5928 11156 5992
rect 11092 5848 11156 5912
rect 11092 5768 11156 5832
rect 11092 5688 11156 5752
rect 11092 5608 11156 5672
rect 11092 5528 11156 5592
rect 11092 5448 11156 5512
rect 11092 5368 11156 5432
rect 11092 5288 11156 5352
rect 11092 5208 11156 5272
rect 12504 5928 12568 5992
rect 12504 5848 12568 5912
rect 12504 5768 12568 5832
rect 12504 5688 12568 5752
rect 12504 5608 12568 5672
rect 12504 5528 12568 5592
rect 12504 5448 12568 5512
rect 12504 5368 12568 5432
rect 12504 5288 12568 5352
rect 12504 5208 12568 5272
rect 13916 5928 13980 5992
rect 13916 5848 13980 5912
rect 13916 5768 13980 5832
rect 13916 5688 13980 5752
rect 13916 5608 13980 5672
rect 13916 5528 13980 5592
rect 13916 5448 13980 5512
rect 13916 5368 13980 5432
rect 13916 5288 13980 5352
rect 13916 5208 13980 5272
rect 15328 5928 15392 5992
rect 15328 5848 15392 5912
rect 15328 5768 15392 5832
rect 15328 5688 15392 5752
rect 15328 5608 15392 5672
rect 15328 5528 15392 5592
rect 15328 5448 15392 5512
rect 15328 5368 15392 5432
rect 15328 5288 15392 5352
rect 15328 5208 15392 5272
rect 16740 5928 16804 5992
rect 16740 5848 16804 5912
rect 16740 5768 16804 5832
rect 16740 5688 16804 5752
rect 16740 5608 16804 5672
rect 16740 5528 16804 5592
rect 16740 5448 16804 5512
rect 16740 5368 16804 5432
rect 16740 5288 16804 5352
rect 16740 5208 16804 5272
rect 18152 5928 18216 5992
rect 18152 5848 18216 5912
rect 18152 5768 18216 5832
rect 18152 5688 18216 5752
rect 18152 5608 18216 5672
rect 18152 5528 18216 5592
rect 18152 5448 18216 5512
rect 18152 5368 18216 5432
rect 18152 5288 18216 5352
rect 18152 5208 18216 5272
rect 19564 5928 19628 5992
rect 19564 5848 19628 5912
rect 19564 5768 19628 5832
rect 19564 5688 19628 5752
rect 19564 5608 19628 5672
rect 19564 5528 19628 5592
rect 19564 5448 19628 5512
rect 19564 5368 19628 5432
rect 19564 5288 19628 5352
rect 19564 5208 19628 5272
rect 20976 5928 21040 5992
rect 20976 5848 21040 5912
rect 20976 5768 21040 5832
rect 20976 5688 21040 5752
rect 20976 5608 21040 5672
rect 20976 5528 21040 5592
rect 20976 5448 21040 5512
rect 20976 5368 21040 5432
rect 20976 5288 21040 5352
rect 20976 5208 21040 5272
rect 22388 5928 22452 5992
rect 22388 5848 22452 5912
rect 22388 5768 22452 5832
rect 22388 5688 22452 5752
rect 22388 5608 22452 5672
rect 22388 5528 22452 5592
rect 22388 5448 22452 5512
rect 22388 5368 22452 5432
rect 22388 5288 22452 5352
rect 22388 5208 22452 5272
rect 23800 5928 23864 5992
rect 23800 5848 23864 5912
rect 23800 5768 23864 5832
rect 23800 5688 23864 5752
rect 23800 5608 23864 5672
rect 23800 5528 23864 5592
rect 23800 5448 23864 5512
rect 23800 5368 23864 5432
rect 23800 5288 23864 5352
rect 23800 5208 23864 5272
rect -22796 4808 -22732 4872
rect -22796 4728 -22732 4792
rect -22796 4648 -22732 4712
rect -22796 4568 -22732 4632
rect -22796 4488 -22732 4552
rect -22796 4408 -22732 4472
rect -22796 4328 -22732 4392
rect -22796 4248 -22732 4312
rect -22796 4168 -22732 4232
rect -22796 4088 -22732 4152
rect -21384 4808 -21320 4872
rect -21384 4728 -21320 4792
rect -21384 4648 -21320 4712
rect -21384 4568 -21320 4632
rect -21384 4488 -21320 4552
rect -21384 4408 -21320 4472
rect -21384 4328 -21320 4392
rect -21384 4248 -21320 4312
rect -21384 4168 -21320 4232
rect -21384 4088 -21320 4152
rect -19972 4808 -19908 4872
rect -19972 4728 -19908 4792
rect -19972 4648 -19908 4712
rect -19972 4568 -19908 4632
rect -19972 4488 -19908 4552
rect -19972 4408 -19908 4472
rect -19972 4328 -19908 4392
rect -19972 4248 -19908 4312
rect -19972 4168 -19908 4232
rect -19972 4088 -19908 4152
rect -18560 4808 -18496 4872
rect -18560 4728 -18496 4792
rect -18560 4648 -18496 4712
rect -18560 4568 -18496 4632
rect -18560 4488 -18496 4552
rect -18560 4408 -18496 4472
rect -18560 4328 -18496 4392
rect -18560 4248 -18496 4312
rect -18560 4168 -18496 4232
rect -18560 4088 -18496 4152
rect -17148 4808 -17084 4872
rect -17148 4728 -17084 4792
rect -17148 4648 -17084 4712
rect -17148 4568 -17084 4632
rect -17148 4488 -17084 4552
rect -17148 4408 -17084 4472
rect -17148 4328 -17084 4392
rect -17148 4248 -17084 4312
rect -17148 4168 -17084 4232
rect -17148 4088 -17084 4152
rect -15736 4808 -15672 4872
rect -15736 4728 -15672 4792
rect -15736 4648 -15672 4712
rect -15736 4568 -15672 4632
rect -15736 4488 -15672 4552
rect -15736 4408 -15672 4472
rect -15736 4328 -15672 4392
rect -15736 4248 -15672 4312
rect -15736 4168 -15672 4232
rect -15736 4088 -15672 4152
rect -14324 4808 -14260 4872
rect -14324 4728 -14260 4792
rect -14324 4648 -14260 4712
rect -14324 4568 -14260 4632
rect -14324 4488 -14260 4552
rect -14324 4408 -14260 4472
rect -14324 4328 -14260 4392
rect -14324 4248 -14260 4312
rect -14324 4168 -14260 4232
rect -14324 4088 -14260 4152
rect -12912 4808 -12848 4872
rect -12912 4728 -12848 4792
rect -12912 4648 -12848 4712
rect -12912 4568 -12848 4632
rect -12912 4488 -12848 4552
rect -12912 4408 -12848 4472
rect -12912 4328 -12848 4392
rect -12912 4248 -12848 4312
rect -12912 4168 -12848 4232
rect -12912 4088 -12848 4152
rect -11500 4808 -11436 4872
rect -11500 4728 -11436 4792
rect -11500 4648 -11436 4712
rect -11500 4568 -11436 4632
rect -11500 4488 -11436 4552
rect -11500 4408 -11436 4472
rect -11500 4328 -11436 4392
rect -11500 4248 -11436 4312
rect -11500 4168 -11436 4232
rect -11500 4088 -11436 4152
rect -10088 4808 -10024 4872
rect -10088 4728 -10024 4792
rect -10088 4648 -10024 4712
rect -10088 4568 -10024 4632
rect -10088 4488 -10024 4552
rect -10088 4408 -10024 4472
rect -10088 4328 -10024 4392
rect -10088 4248 -10024 4312
rect -10088 4168 -10024 4232
rect -10088 4088 -10024 4152
rect -8676 4808 -8612 4872
rect -8676 4728 -8612 4792
rect -8676 4648 -8612 4712
rect -8676 4568 -8612 4632
rect -8676 4488 -8612 4552
rect -8676 4408 -8612 4472
rect -8676 4328 -8612 4392
rect -8676 4248 -8612 4312
rect -8676 4168 -8612 4232
rect -8676 4088 -8612 4152
rect -7264 4808 -7200 4872
rect -7264 4728 -7200 4792
rect -7264 4648 -7200 4712
rect -7264 4568 -7200 4632
rect -7264 4488 -7200 4552
rect -7264 4408 -7200 4472
rect -7264 4328 -7200 4392
rect -7264 4248 -7200 4312
rect -7264 4168 -7200 4232
rect -7264 4088 -7200 4152
rect -5852 4808 -5788 4872
rect -5852 4728 -5788 4792
rect -5852 4648 -5788 4712
rect -5852 4568 -5788 4632
rect -5852 4488 -5788 4552
rect -5852 4408 -5788 4472
rect -5852 4328 -5788 4392
rect -5852 4248 -5788 4312
rect -5852 4168 -5788 4232
rect -5852 4088 -5788 4152
rect -4440 4808 -4376 4872
rect -4440 4728 -4376 4792
rect -4440 4648 -4376 4712
rect -4440 4568 -4376 4632
rect -4440 4488 -4376 4552
rect -4440 4408 -4376 4472
rect -4440 4328 -4376 4392
rect -4440 4248 -4376 4312
rect -4440 4168 -4376 4232
rect -4440 4088 -4376 4152
rect -3028 4808 -2964 4872
rect -3028 4728 -2964 4792
rect -3028 4648 -2964 4712
rect -3028 4568 -2964 4632
rect -3028 4488 -2964 4552
rect -3028 4408 -2964 4472
rect -3028 4328 -2964 4392
rect -3028 4248 -2964 4312
rect -3028 4168 -2964 4232
rect -3028 4088 -2964 4152
rect -1616 4808 -1552 4872
rect -1616 4728 -1552 4792
rect -1616 4648 -1552 4712
rect -1616 4568 -1552 4632
rect -1616 4488 -1552 4552
rect -1616 4408 -1552 4472
rect -1616 4328 -1552 4392
rect -1616 4248 -1552 4312
rect -1616 4168 -1552 4232
rect -1616 4088 -1552 4152
rect -204 4808 -140 4872
rect -204 4728 -140 4792
rect -204 4648 -140 4712
rect -204 4568 -140 4632
rect -204 4488 -140 4552
rect -204 4408 -140 4472
rect -204 4328 -140 4392
rect -204 4248 -140 4312
rect -204 4168 -140 4232
rect -204 4088 -140 4152
rect 1208 4808 1272 4872
rect 1208 4728 1272 4792
rect 1208 4648 1272 4712
rect 1208 4568 1272 4632
rect 1208 4488 1272 4552
rect 1208 4408 1272 4472
rect 1208 4328 1272 4392
rect 1208 4248 1272 4312
rect 1208 4168 1272 4232
rect 1208 4088 1272 4152
rect 2620 4808 2684 4872
rect 2620 4728 2684 4792
rect 2620 4648 2684 4712
rect 2620 4568 2684 4632
rect 2620 4488 2684 4552
rect 2620 4408 2684 4472
rect 2620 4328 2684 4392
rect 2620 4248 2684 4312
rect 2620 4168 2684 4232
rect 2620 4088 2684 4152
rect 4032 4808 4096 4872
rect 4032 4728 4096 4792
rect 4032 4648 4096 4712
rect 4032 4568 4096 4632
rect 4032 4488 4096 4552
rect 4032 4408 4096 4472
rect 4032 4328 4096 4392
rect 4032 4248 4096 4312
rect 4032 4168 4096 4232
rect 4032 4088 4096 4152
rect 5444 4808 5508 4872
rect 5444 4728 5508 4792
rect 5444 4648 5508 4712
rect 5444 4568 5508 4632
rect 5444 4488 5508 4552
rect 5444 4408 5508 4472
rect 5444 4328 5508 4392
rect 5444 4248 5508 4312
rect 5444 4168 5508 4232
rect 5444 4088 5508 4152
rect 6856 4808 6920 4872
rect 6856 4728 6920 4792
rect 6856 4648 6920 4712
rect 6856 4568 6920 4632
rect 6856 4488 6920 4552
rect 6856 4408 6920 4472
rect 6856 4328 6920 4392
rect 6856 4248 6920 4312
rect 6856 4168 6920 4232
rect 6856 4088 6920 4152
rect 8268 4808 8332 4872
rect 8268 4728 8332 4792
rect 8268 4648 8332 4712
rect 8268 4568 8332 4632
rect 8268 4488 8332 4552
rect 8268 4408 8332 4472
rect 8268 4328 8332 4392
rect 8268 4248 8332 4312
rect 8268 4168 8332 4232
rect 8268 4088 8332 4152
rect 9680 4808 9744 4872
rect 9680 4728 9744 4792
rect 9680 4648 9744 4712
rect 9680 4568 9744 4632
rect 9680 4488 9744 4552
rect 9680 4408 9744 4472
rect 9680 4328 9744 4392
rect 9680 4248 9744 4312
rect 9680 4168 9744 4232
rect 9680 4088 9744 4152
rect 11092 4808 11156 4872
rect 11092 4728 11156 4792
rect 11092 4648 11156 4712
rect 11092 4568 11156 4632
rect 11092 4488 11156 4552
rect 11092 4408 11156 4472
rect 11092 4328 11156 4392
rect 11092 4248 11156 4312
rect 11092 4168 11156 4232
rect 11092 4088 11156 4152
rect 12504 4808 12568 4872
rect 12504 4728 12568 4792
rect 12504 4648 12568 4712
rect 12504 4568 12568 4632
rect 12504 4488 12568 4552
rect 12504 4408 12568 4472
rect 12504 4328 12568 4392
rect 12504 4248 12568 4312
rect 12504 4168 12568 4232
rect 12504 4088 12568 4152
rect 13916 4808 13980 4872
rect 13916 4728 13980 4792
rect 13916 4648 13980 4712
rect 13916 4568 13980 4632
rect 13916 4488 13980 4552
rect 13916 4408 13980 4472
rect 13916 4328 13980 4392
rect 13916 4248 13980 4312
rect 13916 4168 13980 4232
rect 13916 4088 13980 4152
rect 15328 4808 15392 4872
rect 15328 4728 15392 4792
rect 15328 4648 15392 4712
rect 15328 4568 15392 4632
rect 15328 4488 15392 4552
rect 15328 4408 15392 4472
rect 15328 4328 15392 4392
rect 15328 4248 15392 4312
rect 15328 4168 15392 4232
rect 15328 4088 15392 4152
rect 16740 4808 16804 4872
rect 16740 4728 16804 4792
rect 16740 4648 16804 4712
rect 16740 4568 16804 4632
rect 16740 4488 16804 4552
rect 16740 4408 16804 4472
rect 16740 4328 16804 4392
rect 16740 4248 16804 4312
rect 16740 4168 16804 4232
rect 16740 4088 16804 4152
rect 18152 4808 18216 4872
rect 18152 4728 18216 4792
rect 18152 4648 18216 4712
rect 18152 4568 18216 4632
rect 18152 4488 18216 4552
rect 18152 4408 18216 4472
rect 18152 4328 18216 4392
rect 18152 4248 18216 4312
rect 18152 4168 18216 4232
rect 18152 4088 18216 4152
rect 19564 4808 19628 4872
rect 19564 4728 19628 4792
rect 19564 4648 19628 4712
rect 19564 4568 19628 4632
rect 19564 4488 19628 4552
rect 19564 4408 19628 4472
rect 19564 4328 19628 4392
rect 19564 4248 19628 4312
rect 19564 4168 19628 4232
rect 19564 4088 19628 4152
rect 20976 4808 21040 4872
rect 20976 4728 21040 4792
rect 20976 4648 21040 4712
rect 20976 4568 21040 4632
rect 20976 4488 21040 4552
rect 20976 4408 21040 4472
rect 20976 4328 21040 4392
rect 20976 4248 21040 4312
rect 20976 4168 21040 4232
rect 20976 4088 21040 4152
rect 22388 4808 22452 4872
rect 22388 4728 22452 4792
rect 22388 4648 22452 4712
rect 22388 4568 22452 4632
rect 22388 4488 22452 4552
rect 22388 4408 22452 4472
rect 22388 4328 22452 4392
rect 22388 4248 22452 4312
rect 22388 4168 22452 4232
rect 22388 4088 22452 4152
rect 23800 4808 23864 4872
rect 23800 4728 23864 4792
rect 23800 4648 23864 4712
rect 23800 4568 23864 4632
rect 23800 4488 23864 4552
rect 23800 4408 23864 4472
rect 23800 4328 23864 4392
rect 23800 4248 23864 4312
rect 23800 4168 23864 4232
rect 23800 4088 23864 4152
rect -22796 3688 -22732 3752
rect -22796 3608 -22732 3672
rect -22796 3528 -22732 3592
rect -22796 3448 -22732 3512
rect -22796 3368 -22732 3432
rect -22796 3288 -22732 3352
rect -22796 3208 -22732 3272
rect -22796 3128 -22732 3192
rect -22796 3048 -22732 3112
rect -22796 2968 -22732 3032
rect -21384 3688 -21320 3752
rect -21384 3608 -21320 3672
rect -21384 3528 -21320 3592
rect -21384 3448 -21320 3512
rect -21384 3368 -21320 3432
rect -21384 3288 -21320 3352
rect -21384 3208 -21320 3272
rect -21384 3128 -21320 3192
rect -21384 3048 -21320 3112
rect -21384 2968 -21320 3032
rect -19972 3688 -19908 3752
rect -19972 3608 -19908 3672
rect -19972 3528 -19908 3592
rect -19972 3448 -19908 3512
rect -19972 3368 -19908 3432
rect -19972 3288 -19908 3352
rect -19972 3208 -19908 3272
rect -19972 3128 -19908 3192
rect -19972 3048 -19908 3112
rect -19972 2968 -19908 3032
rect -18560 3688 -18496 3752
rect -18560 3608 -18496 3672
rect -18560 3528 -18496 3592
rect -18560 3448 -18496 3512
rect -18560 3368 -18496 3432
rect -18560 3288 -18496 3352
rect -18560 3208 -18496 3272
rect -18560 3128 -18496 3192
rect -18560 3048 -18496 3112
rect -18560 2968 -18496 3032
rect -17148 3688 -17084 3752
rect -17148 3608 -17084 3672
rect -17148 3528 -17084 3592
rect -17148 3448 -17084 3512
rect -17148 3368 -17084 3432
rect -17148 3288 -17084 3352
rect -17148 3208 -17084 3272
rect -17148 3128 -17084 3192
rect -17148 3048 -17084 3112
rect -17148 2968 -17084 3032
rect -15736 3688 -15672 3752
rect -15736 3608 -15672 3672
rect -15736 3528 -15672 3592
rect -15736 3448 -15672 3512
rect -15736 3368 -15672 3432
rect -15736 3288 -15672 3352
rect -15736 3208 -15672 3272
rect -15736 3128 -15672 3192
rect -15736 3048 -15672 3112
rect -15736 2968 -15672 3032
rect -14324 3688 -14260 3752
rect -14324 3608 -14260 3672
rect -14324 3528 -14260 3592
rect -14324 3448 -14260 3512
rect -14324 3368 -14260 3432
rect -14324 3288 -14260 3352
rect -14324 3208 -14260 3272
rect -14324 3128 -14260 3192
rect -14324 3048 -14260 3112
rect -14324 2968 -14260 3032
rect -12912 3688 -12848 3752
rect -12912 3608 -12848 3672
rect -12912 3528 -12848 3592
rect -12912 3448 -12848 3512
rect -12912 3368 -12848 3432
rect -12912 3288 -12848 3352
rect -12912 3208 -12848 3272
rect -12912 3128 -12848 3192
rect -12912 3048 -12848 3112
rect -12912 2968 -12848 3032
rect -11500 3688 -11436 3752
rect -11500 3608 -11436 3672
rect -11500 3528 -11436 3592
rect -11500 3448 -11436 3512
rect -11500 3368 -11436 3432
rect -11500 3288 -11436 3352
rect -11500 3208 -11436 3272
rect -11500 3128 -11436 3192
rect -11500 3048 -11436 3112
rect -11500 2968 -11436 3032
rect -10088 3688 -10024 3752
rect -10088 3608 -10024 3672
rect -10088 3528 -10024 3592
rect -10088 3448 -10024 3512
rect -10088 3368 -10024 3432
rect -10088 3288 -10024 3352
rect -10088 3208 -10024 3272
rect -10088 3128 -10024 3192
rect -10088 3048 -10024 3112
rect -10088 2968 -10024 3032
rect -8676 3688 -8612 3752
rect -8676 3608 -8612 3672
rect -8676 3528 -8612 3592
rect -8676 3448 -8612 3512
rect -8676 3368 -8612 3432
rect -8676 3288 -8612 3352
rect -8676 3208 -8612 3272
rect -8676 3128 -8612 3192
rect -8676 3048 -8612 3112
rect -8676 2968 -8612 3032
rect -7264 3688 -7200 3752
rect -7264 3608 -7200 3672
rect -7264 3528 -7200 3592
rect -7264 3448 -7200 3512
rect -7264 3368 -7200 3432
rect -7264 3288 -7200 3352
rect -7264 3208 -7200 3272
rect -7264 3128 -7200 3192
rect -7264 3048 -7200 3112
rect -7264 2968 -7200 3032
rect -5852 3688 -5788 3752
rect -5852 3608 -5788 3672
rect -5852 3528 -5788 3592
rect -5852 3448 -5788 3512
rect -5852 3368 -5788 3432
rect -5852 3288 -5788 3352
rect -5852 3208 -5788 3272
rect -5852 3128 -5788 3192
rect -5852 3048 -5788 3112
rect -5852 2968 -5788 3032
rect -4440 3688 -4376 3752
rect -4440 3608 -4376 3672
rect -4440 3528 -4376 3592
rect -4440 3448 -4376 3512
rect -4440 3368 -4376 3432
rect -4440 3288 -4376 3352
rect -4440 3208 -4376 3272
rect -4440 3128 -4376 3192
rect -4440 3048 -4376 3112
rect -4440 2968 -4376 3032
rect -3028 3688 -2964 3752
rect -3028 3608 -2964 3672
rect -3028 3528 -2964 3592
rect -3028 3448 -2964 3512
rect -3028 3368 -2964 3432
rect -3028 3288 -2964 3352
rect -3028 3208 -2964 3272
rect -3028 3128 -2964 3192
rect -3028 3048 -2964 3112
rect -3028 2968 -2964 3032
rect -1616 3688 -1552 3752
rect -1616 3608 -1552 3672
rect -1616 3528 -1552 3592
rect -1616 3448 -1552 3512
rect -1616 3368 -1552 3432
rect -1616 3288 -1552 3352
rect -1616 3208 -1552 3272
rect -1616 3128 -1552 3192
rect -1616 3048 -1552 3112
rect -1616 2968 -1552 3032
rect -204 3688 -140 3752
rect -204 3608 -140 3672
rect -204 3528 -140 3592
rect -204 3448 -140 3512
rect -204 3368 -140 3432
rect -204 3288 -140 3352
rect -204 3208 -140 3272
rect -204 3128 -140 3192
rect -204 3048 -140 3112
rect -204 2968 -140 3032
rect 1208 3688 1272 3752
rect 1208 3608 1272 3672
rect 1208 3528 1272 3592
rect 1208 3448 1272 3512
rect 1208 3368 1272 3432
rect 1208 3288 1272 3352
rect 1208 3208 1272 3272
rect 1208 3128 1272 3192
rect 1208 3048 1272 3112
rect 1208 2968 1272 3032
rect 2620 3688 2684 3752
rect 2620 3608 2684 3672
rect 2620 3528 2684 3592
rect 2620 3448 2684 3512
rect 2620 3368 2684 3432
rect 2620 3288 2684 3352
rect 2620 3208 2684 3272
rect 2620 3128 2684 3192
rect 2620 3048 2684 3112
rect 2620 2968 2684 3032
rect 4032 3688 4096 3752
rect 4032 3608 4096 3672
rect 4032 3528 4096 3592
rect 4032 3448 4096 3512
rect 4032 3368 4096 3432
rect 4032 3288 4096 3352
rect 4032 3208 4096 3272
rect 4032 3128 4096 3192
rect 4032 3048 4096 3112
rect 4032 2968 4096 3032
rect 5444 3688 5508 3752
rect 5444 3608 5508 3672
rect 5444 3528 5508 3592
rect 5444 3448 5508 3512
rect 5444 3368 5508 3432
rect 5444 3288 5508 3352
rect 5444 3208 5508 3272
rect 5444 3128 5508 3192
rect 5444 3048 5508 3112
rect 5444 2968 5508 3032
rect 6856 3688 6920 3752
rect 6856 3608 6920 3672
rect 6856 3528 6920 3592
rect 6856 3448 6920 3512
rect 6856 3368 6920 3432
rect 6856 3288 6920 3352
rect 6856 3208 6920 3272
rect 6856 3128 6920 3192
rect 6856 3048 6920 3112
rect 6856 2968 6920 3032
rect 8268 3688 8332 3752
rect 8268 3608 8332 3672
rect 8268 3528 8332 3592
rect 8268 3448 8332 3512
rect 8268 3368 8332 3432
rect 8268 3288 8332 3352
rect 8268 3208 8332 3272
rect 8268 3128 8332 3192
rect 8268 3048 8332 3112
rect 8268 2968 8332 3032
rect 9680 3688 9744 3752
rect 9680 3608 9744 3672
rect 9680 3528 9744 3592
rect 9680 3448 9744 3512
rect 9680 3368 9744 3432
rect 9680 3288 9744 3352
rect 9680 3208 9744 3272
rect 9680 3128 9744 3192
rect 9680 3048 9744 3112
rect 9680 2968 9744 3032
rect 11092 3688 11156 3752
rect 11092 3608 11156 3672
rect 11092 3528 11156 3592
rect 11092 3448 11156 3512
rect 11092 3368 11156 3432
rect 11092 3288 11156 3352
rect 11092 3208 11156 3272
rect 11092 3128 11156 3192
rect 11092 3048 11156 3112
rect 11092 2968 11156 3032
rect 12504 3688 12568 3752
rect 12504 3608 12568 3672
rect 12504 3528 12568 3592
rect 12504 3448 12568 3512
rect 12504 3368 12568 3432
rect 12504 3288 12568 3352
rect 12504 3208 12568 3272
rect 12504 3128 12568 3192
rect 12504 3048 12568 3112
rect 12504 2968 12568 3032
rect 13916 3688 13980 3752
rect 13916 3608 13980 3672
rect 13916 3528 13980 3592
rect 13916 3448 13980 3512
rect 13916 3368 13980 3432
rect 13916 3288 13980 3352
rect 13916 3208 13980 3272
rect 13916 3128 13980 3192
rect 13916 3048 13980 3112
rect 13916 2968 13980 3032
rect 15328 3688 15392 3752
rect 15328 3608 15392 3672
rect 15328 3528 15392 3592
rect 15328 3448 15392 3512
rect 15328 3368 15392 3432
rect 15328 3288 15392 3352
rect 15328 3208 15392 3272
rect 15328 3128 15392 3192
rect 15328 3048 15392 3112
rect 15328 2968 15392 3032
rect 16740 3688 16804 3752
rect 16740 3608 16804 3672
rect 16740 3528 16804 3592
rect 16740 3448 16804 3512
rect 16740 3368 16804 3432
rect 16740 3288 16804 3352
rect 16740 3208 16804 3272
rect 16740 3128 16804 3192
rect 16740 3048 16804 3112
rect 16740 2968 16804 3032
rect 18152 3688 18216 3752
rect 18152 3608 18216 3672
rect 18152 3528 18216 3592
rect 18152 3448 18216 3512
rect 18152 3368 18216 3432
rect 18152 3288 18216 3352
rect 18152 3208 18216 3272
rect 18152 3128 18216 3192
rect 18152 3048 18216 3112
rect 18152 2968 18216 3032
rect 19564 3688 19628 3752
rect 19564 3608 19628 3672
rect 19564 3528 19628 3592
rect 19564 3448 19628 3512
rect 19564 3368 19628 3432
rect 19564 3288 19628 3352
rect 19564 3208 19628 3272
rect 19564 3128 19628 3192
rect 19564 3048 19628 3112
rect 19564 2968 19628 3032
rect 20976 3688 21040 3752
rect 20976 3608 21040 3672
rect 20976 3528 21040 3592
rect 20976 3448 21040 3512
rect 20976 3368 21040 3432
rect 20976 3288 21040 3352
rect 20976 3208 21040 3272
rect 20976 3128 21040 3192
rect 20976 3048 21040 3112
rect 20976 2968 21040 3032
rect 22388 3688 22452 3752
rect 22388 3608 22452 3672
rect 22388 3528 22452 3592
rect 22388 3448 22452 3512
rect 22388 3368 22452 3432
rect 22388 3288 22452 3352
rect 22388 3208 22452 3272
rect 22388 3128 22452 3192
rect 22388 3048 22452 3112
rect 22388 2968 22452 3032
rect 23800 3688 23864 3752
rect 23800 3608 23864 3672
rect 23800 3528 23864 3592
rect 23800 3448 23864 3512
rect 23800 3368 23864 3432
rect 23800 3288 23864 3352
rect 23800 3208 23864 3272
rect 23800 3128 23864 3192
rect 23800 3048 23864 3112
rect 23800 2968 23864 3032
rect -22796 2568 -22732 2632
rect -22796 2488 -22732 2552
rect -22796 2408 -22732 2472
rect -22796 2328 -22732 2392
rect -22796 2248 -22732 2312
rect -22796 2168 -22732 2232
rect -22796 2088 -22732 2152
rect -22796 2008 -22732 2072
rect -22796 1928 -22732 1992
rect -22796 1848 -22732 1912
rect -21384 2568 -21320 2632
rect -21384 2488 -21320 2552
rect -21384 2408 -21320 2472
rect -21384 2328 -21320 2392
rect -21384 2248 -21320 2312
rect -21384 2168 -21320 2232
rect -21384 2088 -21320 2152
rect -21384 2008 -21320 2072
rect -21384 1928 -21320 1992
rect -21384 1848 -21320 1912
rect -19972 2568 -19908 2632
rect -19972 2488 -19908 2552
rect -19972 2408 -19908 2472
rect -19972 2328 -19908 2392
rect -19972 2248 -19908 2312
rect -19972 2168 -19908 2232
rect -19972 2088 -19908 2152
rect -19972 2008 -19908 2072
rect -19972 1928 -19908 1992
rect -19972 1848 -19908 1912
rect -18560 2568 -18496 2632
rect -18560 2488 -18496 2552
rect -18560 2408 -18496 2472
rect -18560 2328 -18496 2392
rect -18560 2248 -18496 2312
rect -18560 2168 -18496 2232
rect -18560 2088 -18496 2152
rect -18560 2008 -18496 2072
rect -18560 1928 -18496 1992
rect -18560 1848 -18496 1912
rect -17148 2568 -17084 2632
rect -17148 2488 -17084 2552
rect -17148 2408 -17084 2472
rect -17148 2328 -17084 2392
rect -17148 2248 -17084 2312
rect -17148 2168 -17084 2232
rect -17148 2088 -17084 2152
rect -17148 2008 -17084 2072
rect -17148 1928 -17084 1992
rect -17148 1848 -17084 1912
rect -15736 2568 -15672 2632
rect -15736 2488 -15672 2552
rect -15736 2408 -15672 2472
rect -15736 2328 -15672 2392
rect -15736 2248 -15672 2312
rect -15736 2168 -15672 2232
rect -15736 2088 -15672 2152
rect -15736 2008 -15672 2072
rect -15736 1928 -15672 1992
rect -15736 1848 -15672 1912
rect -14324 2568 -14260 2632
rect -14324 2488 -14260 2552
rect -14324 2408 -14260 2472
rect -14324 2328 -14260 2392
rect -14324 2248 -14260 2312
rect -14324 2168 -14260 2232
rect -14324 2088 -14260 2152
rect -14324 2008 -14260 2072
rect -14324 1928 -14260 1992
rect -14324 1848 -14260 1912
rect -12912 2568 -12848 2632
rect -12912 2488 -12848 2552
rect -12912 2408 -12848 2472
rect -12912 2328 -12848 2392
rect -12912 2248 -12848 2312
rect -12912 2168 -12848 2232
rect -12912 2088 -12848 2152
rect -12912 2008 -12848 2072
rect -12912 1928 -12848 1992
rect -12912 1848 -12848 1912
rect -11500 2568 -11436 2632
rect -11500 2488 -11436 2552
rect -11500 2408 -11436 2472
rect -11500 2328 -11436 2392
rect -11500 2248 -11436 2312
rect -11500 2168 -11436 2232
rect -11500 2088 -11436 2152
rect -11500 2008 -11436 2072
rect -11500 1928 -11436 1992
rect -11500 1848 -11436 1912
rect -10088 2568 -10024 2632
rect -10088 2488 -10024 2552
rect -10088 2408 -10024 2472
rect -10088 2328 -10024 2392
rect -10088 2248 -10024 2312
rect -10088 2168 -10024 2232
rect -10088 2088 -10024 2152
rect -10088 2008 -10024 2072
rect -10088 1928 -10024 1992
rect -10088 1848 -10024 1912
rect -8676 2568 -8612 2632
rect -8676 2488 -8612 2552
rect -8676 2408 -8612 2472
rect -8676 2328 -8612 2392
rect -8676 2248 -8612 2312
rect -8676 2168 -8612 2232
rect -8676 2088 -8612 2152
rect -8676 2008 -8612 2072
rect -8676 1928 -8612 1992
rect -8676 1848 -8612 1912
rect -7264 2568 -7200 2632
rect -7264 2488 -7200 2552
rect -7264 2408 -7200 2472
rect -7264 2328 -7200 2392
rect -7264 2248 -7200 2312
rect -7264 2168 -7200 2232
rect -7264 2088 -7200 2152
rect -7264 2008 -7200 2072
rect -7264 1928 -7200 1992
rect -7264 1848 -7200 1912
rect -5852 2568 -5788 2632
rect -5852 2488 -5788 2552
rect -5852 2408 -5788 2472
rect -5852 2328 -5788 2392
rect -5852 2248 -5788 2312
rect -5852 2168 -5788 2232
rect -5852 2088 -5788 2152
rect -5852 2008 -5788 2072
rect -5852 1928 -5788 1992
rect -5852 1848 -5788 1912
rect -4440 2568 -4376 2632
rect -4440 2488 -4376 2552
rect -4440 2408 -4376 2472
rect -4440 2328 -4376 2392
rect -4440 2248 -4376 2312
rect -4440 2168 -4376 2232
rect -4440 2088 -4376 2152
rect -4440 2008 -4376 2072
rect -4440 1928 -4376 1992
rect -4440 1848 -4376 1912
rect -3028 2568 -2964 2632
rect -3028 2488 -2964 2552
rect -3028 2408 -2964 2472
rect -3028 2328 -2964 2392
rect -3028 2248 -2964 2312
rect -3028 2168 -2964 2232
rect -3028 2088 -2964 2152
rect -3028 2008 -2964 2072
rect -3028 1928 -2964 1992
rect -3028 1848 -2964 1912
rect -1616 2568 -1552 2632
rect -1616 2488 -1552 2552
rect -1616 2408 -1552 2472
rect -1616 2328 -1552 2392
rect -1616 2248 -1552 2312
rect -1616 2168 -1552 2232
rect -1616 2088 -1552 2152
rect -1616 2008 -1552 2072
rect -1616 1928 -1552 1992
rect -1616 1848 -1552 1912
rect -204 2568 -140 2632
rect -204 2488 -140 2552
rect -204 2408 -140 2472
rect -204 2328 -140 2392
rect -204 2248 -140 2312
rect -204 2168 -140 2232
rect -204 2088 -140 2152
rect -204 2008 -140 2072
rect -204 1928 -140 1992
rect -204 1848 -140 1912
rect 1208 2568 1272 2632
rect 1208 2488 1272 2552
rect 1208 2408 1272 2472
rect 1208 2328 1272 2392
rect 1208 2248 1272 2312
rect 1208 2168 1272 2232
rect 1208 2088 1272 2152
rect 1208 2008 1272 2072
rect 1208 1928 1272 1992
rect 1208 1848 1272 1912
rect 2620 2568 2684 2632
rect 2620 2488 2684 2552
rect 2620 2408 2684 2472
rect 2620 2328 2684 2392
rect 2620 2248 2684 2312
rect 2620 2168 2684 2232
rect 2620 2088 2684 2152
rect 2620 2008 2684 2072
rect 2620 1928 2684 1992
rect 2620 1848 2684 1912
rect 4032 2568 4096 2632
rect 4032 2488 4096 2552
rect 4032 2408 4096 2472
rect 4032 2328 4096 2392
rect 4032 2248 4096 2312
rect 4032 2168 4096 2232
rect 4032 2088 4096 2152
rect 4032 2008 4096 2072
rect 4032 1928 4096 1992
rect 4032 1848 4096 1912
rect 5444 2568 5508 2632
rect 5444 2488 5508 2552
rect 5444 2408 5508 2472
rect 5444 2328 5508 2392
rect 5444 2248 5508 2312
rect 5444 2168 5508 2232
rect 5444 2088 5508 2152
rect 5444 2008 5508 2072
rect 5444 1928 5508 1992
rect 5444 1848 5508 1912
rect 6856 2568 6920 2632
rect 6856 2488 6920 2552
rect 6856 2408 6920 2472
rect 6856 2328 6920 2392
rect 6856 2248 6920 2312
rect 6856 2168 6920 2232
rect 6856 2088 6920 2152
rect 6856 2008 6920 2072
rect 6856 1928 6920 1992
rect 6856 1848 6920 1912
rect 8268 2568 8332 2632
rect 8268 2488 8332 2552
rect 8268 2408 8332 2472
rect 8268 2328 8332 2392
rect 8268 2248 8332 2312
rect 8268 2168 8332 2232
rect 8268 2088 8332 2152
rect 8268 2008 8332 2072
rect 8268 1928 8332 1992
rect 8268 1848 8332 1912
rect 9680 2568 9744 2632
rect 9680 2488 9744 2552
rect 9680 2408 9744 2472
rect 9680 2328 9744 2392
rect 9680 2248 9744 2312
rect 9680 2168 9744 2232
rect 9680 2088 9744 2152
rect 9680 2008 9744 2072
rect 9680 1928 9744 1992
rect 9680 1848 9744 1912
rect 11092 2568 11156 2632
rect 11092 2488 11156 2552
rect 11092 2408 11156 2472
rect 11092 2328 11156 2392
rect 11092 2248 11156 2312
rect 11092 2168 11156 2232
rect 11092 2088 11156 2152
rect 11092 2008 11156 2072
rect 11092 1928 11156 1992
rect 11092 1848 11156 1912
rect 12504 2568 12568 2632
rect 12504 2488 12568 2552
rect 12504 2408 12568 2472
rect 12504 2328 12568 2392
rect 12504 2248 12568 2312
rect 12504 2168 12568 2232
rect 12504 2088 12568 2152
rect 12504 2008 12568 2072
rect 12504 1928 12568 1992
rect 12504 1848 12568 1912
rect 13916 2568 13980 2632
rect 13916 2488 13980 2552
rect 13916 2408 13980 2472
rect 13916 2328 13980 2392
rect 13916 2248 13980 2312
rect 13916 2168 13980 2232
rect 13916 2088 13980 2152
rect 13916 2008 13980 2072
rect 13916 1928 13980 1992
rect 13916 1848 13980 1912
rect 15328 2568 15392 2632
rect 15328 2488 15392 2552
rect 15328 2408 15392 2472
rect 15328 2328 15392 2392
rect 15328 2248 15392 2312
rect 15328 2168 15392 2232
rect 15328 2088 15392 2152
rect 15328 2008 15392 2072
rect 15328 1928 15392 1992
rect 15328 1848 15392 1912
rect 16740 2568 16804 2632
rect 16740 2488 16804 2552
rect 16740 2408 16804 2472
rect 16740 2328 16804 2392
rect 16740 2248 16804 2312
rect 16740 2168 16804 2232
rect 16740 2088 16804 2152
rect 16740 2008 16804 2072
rect 16740 1928 16804 1992
rect 16740 1848 16804 1912
rect 18152 2568 18216 2632
rect 18152 2488 18216 2552
rect 18152 2408 18216 2472
rect 18152 2328 18216 2392
rect 18152 2248 18216 2312
rect 18152 2168 18216 2232
rect 18152 2088 18216 2152
rect 18152 2008 18216 2072
rect 18152 1928 18216 1992
rect 18152 1848 18216 1912
rect 19564 2568 19628 2632
rect 19564 2488 19628 2552
rect 19564 2408 19628 2472
rect 19564 2328 19628 2392
rect 19564 2248 19628 2312
rect 19564 2168 19628 2232
rect 19564 2088 19628 2152
rect 19564 2008 19628 2072
rect 19564 1928 19628 1992
rect 19564 1848 19628 1912
rect 20976 2568 21040 2632
rect 20976 2488 21040 2552
rect 20976 2408 21040 2472
rect 20976 2328 21040 2392
rect 20976 2248 21040 2312
rect 20976 2168 21040 2232
rect 20976 2088 21040 2152
rect 20976 2008 21040 2072
rect 20976 1928 21040 1992
rect 20976 1848 21040 1912
rect 22388 2568 22452 2632
rect 22388 2488 22452 2552
rect 22388 2408 22452 2472
rect 22388 2328 22452 2392
rect 22388 2248 22452 2312
rect 22388 2168 22452 2232
rect 22388 2088 22452 2152
rect 22388 2008 22452 2072
rect 22388 1928 22452 1992
rect 22388 1848 22452 1912
rect 23800 2568 23864 2632
rect 23800 2488 23864 2552
rect 23800 2408 23864 2472
rect 23800 2328 23864 2392
rect 23800 2248 23864 2312
rect 23800 2168 23864 2232
rect 23800 2088 23864 2152
rect 23800 2008 23864 2072
rect 23800 1928 23864 1992
rect 23800 1848 23864 1912
rect -22796 1448 -22732 1512
rect -22796 1368 -22732 1432
rect -22796 1288 -22732 1352
rect -22796 1208 -22732 1272
rect -22796 1128 -22732 1192
rect -22796 1048 -22732 1112
rect -22796 968 -22732 1032
rect -22796 888 -22732 952
rect -22796 808 -22732 872
rect -22796 728 -22732 792
rect -21384 1448 -21320 1512
rect -21384 1368 -21320 1432
rect -21384 1288 -21320 1352
rect -21384 1208 -21320 1272
rect -21384 1128 -21320 1192
rect -21384 1048 -21320 1112
rect -21384 968 -21320 1032
rect -21384 888 -21320 952
rect -21384 808 -21320 872
rect -21384 728 -21320 792
rect -19972 1448 -19908 1512
rect -19972 1368 -19908 1432
rect -19972 1288 -19908 1352
rect -19972 1208 -19908 1272
rect -19972 1128 -19908 1192
rect -19972 1048 -19908 1112
rect -19972 968 -19908 1032
rect -19972 888 -19908 952
rect -19972 808 -19908 872
rect -19972 728 -19908 792
rect -18560 1448 -18496 1512
rect -18560 1368 -18496 1432
rect -18560 1288 -18496 1352
rect -18560 1208 -18496 1272
rect -18560 1128 -18496 1192
rect -18560 1048 -18496 1112
rect -18560 968 -18496 1032
rect -18560 888 -18496 952
rect -18560 808 -18496 872
rect -18560 728 -18496 792
rect -17148 1448 -17084 1512
rect -17148 1368 -17084 1432
rect -17148 1288 -17084 1352
rect -17148 1208 -17084 1272
rect -17148 1128 -17084 1192
rect -17148 1048 -17084 1112
rect -17148 968 -17084 1032
rect -17148 888 -17084 952
rect -17148 808 -17084 872
rect -17148 728 -17084 792
rect -15736 1448 -15672 1512
rect -15736 1368 -15672 1432
rect -15736 1288 -15672 1352
rect -15736 1208 -15672 1272
rect -15736 1128 -15672 1192
rect -15736 1048 -15672 1112
rect -15736 968 -15672 1032
rect -15736 888 -15672 952
rect -15736 808 -15672 872
rect -15736 728 -15672 792
rect -14324 1448 -14260 1512
rect -14324 1368 -14260 1432
rect -14324 1288 -14260 1352
rect -14324 1208 -14260 1272
rect -14324 1128 -14260 1192
rect -14324 1048 -14260 1112
rect -14324 968 -14260 1032
rect -14324 888 -14260 952
rect -14324 808 -14260 872
rect -14324 728 -14260 792
rect -12912 1448 -12848 1512
rect -12912 1368 -12848 1432
rect -12912 1288 -12848 1352
rect -12912 1208 -12848 1272
rect -12912 1128 -12848 1192
rect -12912 1048 -12848 1112
rect -12912 968 -12848 1032
rect -12912 888 -12848 952
rect -12912 808 -12848 872
rect -12912 728 -12848 792
rect -11500 1448 -11436 1512
rect -11500 1368 -11436 1432
rect -11500 1288 -11436 1352
rect -11500 1208 -11436 1272
rect -11500 1128 -11436 1192
rect -11500 1048 -11436 1112
rect -11500 968 -11436 1032
rect -11500 888 -11436 952
rect -11500 808 -11436 872
rect -11500 728 -11436 792
rect -10088 1448 -10024 1512
rect -10088 1368 -10024 1432
rect -10088 1288 -10024 1352
rect -10088 1208 -10024 1272
rect -10088 1128 -10024 1192
rect -10088 1048 -10024 1112
rect -10088 968 -10024 1032
rect -10088 888 -10024 952
rect -10088 808 -10024 872
rect -10088 728 -10024 792
rect -8676 1448 -8612 1512
rect -8676 1368 -8612 1432
rect -8676 1288 -8612 1352
rect -8676 1208 -8612 1272
rect -8676 1128 -8612 1192
rect -8676 1048 -8612 1112
rect -8676 968 -8612 1032
rect -8676 888 -8612 952
rect -8676 808 -8612 872
rect -8676 728 -8612 792
rect -7264 1448 -7200 1512
rect -7264 1368 -7200 1432
rect -7264 1288 -7200 1352
rect -7264 1208 -7200 1272
rect -7264 1128 -7200 1192
rect -7264 1048 -7200 1112
rect -7264 968 -7200 1032
rect -7264 888 -7200 952
rect -7264 808 -7200 872
rect -7264 728 -7200 792
rect -5852 1448 -5788 1512
rect -5852 1368 -5788 1432
rect -5852 1288 -5788 1352
rect -5852 1208 -5788 1272
rect -5852 1128 -5788 1192
rect -5852 1048 -5788 1112
rect -5852 968 -5788 1032
rect -5852 888 -5788 952
rect -5852 808 -5788 872
rect -5852 728 -5788 792
rect -4440 1448 -4376 1512
rect -4440 1368 -4376 1432
rect -4440 1288 -4376 1352
rect -4440 1208 -4376 1272
rect -4440 1128 -4376 1192
rect -4440 1048 -4376 1112
rect -4440 968 -4376 1032
rect -4440 888 -4376 952
rect -4440 808 -4376 872
rect -4440 728 -4376 792
rect -3028 1448 -2964 1512
rect -3028 1368 -2964 1432
rect -3028 1288 -2964 1352
rect -3028 1208 -2964 1272
rect -3028 1128 -2964 1192
rect -3028 1048 -2964 1112
rect -3028 968 -2964 1032
rect -3028 888 -2964 952
rect -3028 808 -2964 872
rect -3028 728 -2964 792
rect -1616 1448 -1552 1512
rect -1616 1368 -1552 1432
rect -1616 1288 -1552 1352
rect -1616 1208 -1552 1272
rect -1616 1128 -1552 1192
rect -1616 1048 -1552 1112
rect -1616 968 -1552 1032
rect -1616 888 -1552 952
rect -1616 808 -1552 872
rect -1616 728 -1552 792
rect -204 1448 -140 1512
rect -204 1368 -140 1432
rect -204 1288 -140 1352
rect -204 1208 -140 1272
rect -204 1128 -140 1192
rect -204 1048 -140 1112
rect -204 968 -140 1032
rect -204 888 -140 952
rect -204 808 -140 872
rect -204 728 -140 792
rect 1208 1448 1272 1512
rect 1208 1368 1272 1432
rect 1208 1288 1272 1352
rect 1208 1208 1272 1272
rect 1208 1128 1272 1192
rect 1208 1048 1272 1112
rect 1208 968 1272 1032
rect 1208 888 1272 952
rect 1208 808 1272 872
rect 1208 728 1272 792
rect 2620 1448 2684 1512
rect 2620 1368 2684 1432
rect 2620 1288 2684 1352
rect 2620 1208 2684 1272
rect 2620 1128 2684 1192
rect 2620 1048 2684 1112
rect 2620 968 2684 1032
rect 2620 888 2684 952
rect 2620 808 2684 872
rect 2620 728 2684 792
rect 4032 1448 4096 1512
rect 4032 1368 4096 1432
rect 4032 1288 4096 1352
rect 4032 1208 4096 1272
rect 4032 1128 4096 1192
rect 4032 1048 4096 1112
rect 4032 968 4096 1032
rect 4032 888 4096 952
rect 4032 808 4096 872
rect 4032 728 4096 792
rect 5444 1448 5508 1512
rect 5444 1368 5508 1432
rect 5444 1288 5508 1352
rect 5444 1208 5508 1272
rect 5444 1128 5508 1192
rect 5444 1048 5508 1112
rect 5444 968 5508 1032
rect 5444 888 5508 952
rect 5444 808 5508 872
rect 5444 728 5508 792
rect 6856 1448 6920 1512
rect 6856 1368 6920 1432
rect 6856 1288 6920 1352
rect 6856 1208 6920 1272
rect 6856 1128 6920 1192
rect 6856 1048 6920 1112
rect 6856 968 6920 1032
rect 6856 888 6920 952
rect 6856 808 6920 872
rect 6856 728 6920 792
rect 8268 1448 8332 1512
rect 8268 1368 8332 1432
rect 8268 1288 8332 1352
rect 8268 1208 8332 1272
rect 8268 1128 8332 1192
rect 8268 1048 8332 1112
rect 8268 968 8332 1032
rect 8268 888 8332 952
rect 8268 808 8332 872
rect 8268 728 8332 792
rect 9680 1448 9744 1512
rect 9680 1368 9744 1432
rect 9680 1288 9744 1352
rect 9680 1208 9744 1272
rect 9680 1128 9744 1192
rect 9680 1048 9744 1112
rect 9680 968 9744 1032
rect 9680 888 9744 952
rect 9680 808 9744 872
rect 9680 728 9744 792
rect 11092 1448 11156 1512
rect 11092 1368 11156 1432
rect 11092 1288 11156 1352
rect 11092 1208 11156 1272
rect 11092 1128 11156 1192
rect 11092 1048 11156 1112
rect 11092 968 11156 1032
rect 11092 888 11156 952
rect 11092 808 11156 872
rect 11092 728 11156 792
rect 12504 1448 12568 1512
rect 12504 1368 12568 1432
rect 12504 1288 12568 1352
rect 12504 1208 12568 1272
rect 12504 1128 12568 1192
rect 12504 1048 12568 1112
rect 12504 968 12568 1032
rect 12504 888 12568 952
rect 12504 808 12568 872
rect 12504 728 12568 792
rect 13916 1448 13980 1512
rect 13916 1368 13980 1432
rect 13916 1288 13980 1352
rect 13916 1208 13980 1272
rect 13916 1128 13980 1192
rect 13916 1048 13980 1112
rect 13916 968 13980 1032
rect 13916 888 13980 952
rect 13916 808 13980 872
rect 13916 728 13980 792
rect 15328 1448 15392 1512
rect 15328 1368 15392 1432
rect 15328 1288 15392 1352
rect 15328 1208 15392 1272
rect 15328 1128 15392 1192
rect 15328 1048 15392 1112
rect 15328 968 15392 1032
rect 15328 888 15392 952
rect 15328 808 15392 872
rect 15328 728 15392 792
rect 16740 1448 16804 1512
rect 16740 1368 16804 1432
rect 16740 1288 16804 1352
rect 16740 1208 16804 1272
rect 16740 1128 16804 1192
rect 16740 1048 16804 1112
rect 16740 968 16804 1032
rect 16740 888 16804 952
rect 16740 808 16804 872
rect 16740 728 16804 792
rect 18152 1448 18216 1512
rect 18152 1368 18216 1432
rect 18152 1288 18216 1352
rect 18152 1208 18216 1272
rect 18152 1128 18216 1192
rect 18152 1048 18216 1112
rect 18152 968 18216 1032
rect 18152 888 18216 952
rect 18152 808 18216 872
rect 18152 728 18216 792
rect 19564 1448 19628 1512
rect 19564 1368 19628 1432
rect 19564 1288 19628 1352
rect 19564 1208 19628 1272
rect 19564 1128 19628 1192
rect 19564 1048 19628 1112
rect 19564 968 19628 1032
rect 19564 888 19628 952
rect 19564 808 19628 872
rect 19564 728 19628 792
rect 20976 1448 21040 1512
rect 20976 1368 21040 1432
rect 20976 1288 21040 1352
rect 20976 1208 21040 1272
rect 20976 1128 21040 1192
rect 20976 1048 21040 1112
rect 20976 968 21040 1032
rect 20976 888 21040 952
rect 20976 808 21040 872
rect 20976 728 21040 792
rect 22388 1448 22452 1512
rect 22388 1368 22452 1432
rect 22388 1288 22452 1352
rect 22388 1208 22452 1272
rect 22388 1128 22452 1192
rect 22388 1048 22452 1112
rect 22388 968 22452 1032
rect 22388 888 22452 952
rect 22388 808 22452 872
rect 22388 728 22452 792
rect 23800 1448 23864 1512
rect 23800 1368 23864 1432
rect 23800 1288 23864 1352
rect 23800 1208 23864 1272
rect 23800 1128 23864 1192
rect 23800 1048 23864 1112
rect 23800 968 23864 1032
rect 23800 888 23864 952
rect 23800 808 23864 872
rect 23800 728 23864 792
rect -22796 328 -22732 392
rect -22796 248 -22732 312
rect -22796 168 -22732 232
rect -22796 88 -22732 152
rect -22796 8 -22732 72
rect -22796 -72 -22732 -8
rect -22796 -152 -22732 -88
rect -22796 -232 -22732 -168
rect -22796 -312 -22732 -248
rect -22796 -392 -22732 -328
rect -21384 328 -21320 392
rect -21384 248 -21320 312
rect -21384 168 -21320 232
rect -21384 88 -21320 152
rect -21384 8 -21320 72
rect -21384 -72 -21320 -8
rect -21384 -152 -21320 -88
rect -21384 -232 -21320 -168
rect -21384 -312 -21320 -248
rect -21384 -392 -21320 -328
rect -19972 328 -19908 392
rect -19972 248 -19908 312
rect -19972 168 -19908 232
rect -19972 88 -19908 152
rect -19972 8 -19908 72
rect -19972 -72 -19908 -8
rect -19972 -152 -19908 -88
rect -19972 -232 -19908 -168
rect -19972 -312 -19908 -248
rect -19972 -392 -19908 -328
rect -18560 328 -18496 392
rect -18560 248 -18496 312
rect -18560 168 -18496 232
rect -18560 88 -18496 152
rect -18560 8 -18496 72
rect -18560 -72 -18496 -8
rect -18560 -152 -18496 -88
rect -18560 -232 -18496 -168
rect -18560 -312 -18496 -248
rect -18560 -392 -18496 -328
rect -17148 328 -17084 392
rect -17148 248 -17084 312
rect -17148 168 -17084 232
rect -17148 88 -17084 152
rect -17148 8 -17084 72
rect -17148 -72 -17084 -8
rect -17148 -152 -17084 -88
rect -17148 -232 -17084 -168
rect -17148 -312 -17084 -248
rect -17148 -392 -17084 -328
rect -15736 328 -15672 392
rect -15736 248 -15672 312
rect -15736 168 -15672 232
rect -15736 88 -15672 152
rect -15736 8 -15672 72
rect -15736 -72 -15672 -8
rect -15736 -152 -15672 -88
rect -15736 -232 -15672 -168
rect -15736 -312 -15672 -248
rect -15736 -392 -15672 -328
rect -14324 328 -14260 392
rect -14324 248 -14260 312
rect -14324 168 -14260 232
rect -14324 88 -14260 152
rect -14324 8 -14260 72
rect -14324 -72 -14260 -8
rect -14324 -152 -14260 -88
rect -14324 -232 -14260 -168
rect -14324 -312 -14260 -248
rect -14324 -392 -14260 -328
rect -12912 328 -12848 392
rect -12912 248 -12848 312
rect -12912 168 -12848 232
rect -12912 88 -12848 152
rect -12912 8 -12848 72
rect -12912 -72 -12848 -8
rect -12912 -152 -12848 -88
rect -12912 -232 -12848 -168
rect -12912 -312 -12848 -248
rect -12912 -392 -12848 -328
rect -11500 328 -11436 392
rect -11500 248 -11436 312
rect -11500 168 -11436 232
rect -11500 88 -11436 152
rect -11500 8 -11436 72
rect -11500 -72 -11436 -8
rect -11500 -152 -11436 -88
rect -11500 -232 -11436 -168
rect -11500 -312 -11436 -248
rect -11500 -392 -11436 -328
rect -10088 328 -10024 392
rect -10088 248 -10024 312
rect -10088 168 -10024 232
rect -10088 88 -10024 152
rect -10088 8 -10024 72
rect -10088 -72 -10024 -8
rect -10088 -152 -10024 -88
rect -10088 -232 -10024 -168
rect -10088 -312 -10024 -248
rect -10088 -392 -10024 -328
rect -8676 328 -8612 392
rect -8676 248 -8612 312
rect -8676 168 -8612 232
rect -8676 88 -8612 152
rect -8676 8 -8612 72
rect -8676 -72 -8612 -8
rect -8676 -152 -8612 -88
rect -8676 -232 -8612 -168
rect -8676 -312 -8612 -248
rect -8676 -392 -8612 -328
rect -7264 328 -7200 392
rect -7264 248 -7200 312
rect -7264 168 -7200 232
rect -7264 88 -7200 152
rect -7264 8 -7200 72
rect -7264 -72 -7200 -8
rect -7264 -152 -7200 -88
rect -7264 -232 -7200 -168
rect -7264 -312 -7200 -248
rect -7264 -392 -7200 -328
rect -5852 328 -5788 392
rect -5852 248 -5788 312
rect -5852 168 -5788 232
rect -5852 88 -5788 152
rect -5852 8 -5788 72
rect -5852 -72 -5788 -8
rect -5852 -152 -5788 -88
rect -5852 -232 -5788 -168
rect -5852 -312 -5788 -248
rect -5852 -392 -5788 -328
rect -4440 328 -4376 392
rect -4440 248 -4376 312
rect -4440 168 -4376 232
rect -4440 88 -4376 152
rect -4440 8 -4376 72
rect -4440 -72 -4376 -8
rect -4440 -152 -4376 -88
rect -4440 -232 -4376 -168
rect -4440 -312 -4376 -248
rect -4440 -392 -4376 -328
rect -3028 328 -2964 392
rect -3028 248 -2964 312
rect -3028 168 -2964 232
rect -3028 88 -2964 152
rect -3028 8 -2964 72
rect -3028 -72 -2964 -8
rect -3028 -152 -2964 -88
rect -3028 -232 -2964 -168
rect -3028 -312 -2964 -248
rect -3028 -392 -2964 -328
rect -1616 328 -1552 392
rect -1616 248 -1552 312
rect -1616 168 -1552 232
rect -1616 88 -1552 152
rect -1616 8 -1552 72
rect -1616 -72 -1552 -8
rect -1616 -152 -1552 -88
rect -1616 -232 -1552 -168
rect -1616 -312 -1552 -248
rect -1616 -392 -1552 -328
rect -204 328 -140 392
rect -204 248 -140 312
rect -204 168 -140 232
rect -204 88 -140 152
rect -204 8 -140 72
rect -204 -72 -140 -8
rect -204 -152 -140 -88
rect -204 -232 -140 -168
rect -204 -312 -140 -248
rect -204 -392 -140 -328
rect 1208 328 1272 392
rect 1208 248 1272 312
rect 1208 168 1272 232
rect 1208 88 1272 152
rect 1208 8 1272 72
rect 1208 -72 1272 -8
rect 1208 -152 1272 -88
rect 1208 -232 1272 -168
rect 1208 -312 1272 -248
rect 1208 -392 1272 -328
rect 2620 328 2684 392
rect 2620 248 2684 312
rect 2620 168 2684 232
rect 2620 88 2684 152
rect 2620 8 2684 72
rect 2620 -72 2684 -8
rect 2620 -152 2684 -88
rect 2620 -232 2684 -168
rect 2620 -312 2684 -248
rect 2620 -392 2684 -328
rect 4032 328 4096 392
rect 4032 248 4096 312
rect 4032 168 4096 232
rect 4032 88 4096 152
rect 4032 8 4096 72
rect 4032 -72 4096 -8
rect 4032 -152 4096 -88
rect 4032 -232 4096 -168
rect 4032 -312 4096 -248
rect 4032 -392 4096 -328
rect 5444 328 5508 392
rect 5444 248 5508 312
rect 5444 168 5508 232
rect 5444 88 5508 152
rect 5444 8 5508 72
rect 5444 -72 5508 -8
rect 5444 -152 5508 -88
rect 5444 -232 5508 -168
rect 5444 -312 5508 -248
rect 5444 -392 5508 -328
rect 6856 328 6920 392
rect 6856 248 6920 312
rect 6856 168 6920 232
rect 6856 88 6920 152
rect 6856 8 6920 72
rect 6856 -72 6920 -8
rect 6856 -152 6920 -88
rect 6856 -232 6920 -168
rect 6856 -312 6920 -248
rect 6856 -392 6920 -328
rect 8268 328 8332 392
rect 8268 248 8332 312
rect 8268 168 8332 232
rect 8268 88 8332 152
rect 8268 8 8332 72
rect 8268 -72 8332 -8
rect 8268 -152 8332 -88
rect 8268 -232 8332 -168
rect 8268 -312 8332 -248
rect 8268 -392 8332 -328
rect 9680 328 9744 392
rect 9680 248 9744 312
rect 9680 168 9744 232
rect 9680 88 9744 152
rect 9680 8 9744 72
rect 9680 -72 9744 -8
rect 9680 -152 9744 -88
rect 9680 -232 9744 -168
rect 9680 -312 9744 -248
rect 9680 -392 9744 -328
rect 11092 328 11156 392
rect 11092 248 11156 312
rect 11092 168 11156 232
rect 11092 88 11156 152
rect 11092 8 11156 72
rect 11092 -72 11156 -8
rect 11092 -152 11156 -88
rect 11092 -232 11156 -168
rect 11092 -312 11156 -248
rect 11092 -392 11156 -328
rect 12504 328 12568 392
rect 12504 248 12568 312
rect 12504 168 12568 232
rect 12504 88 12568 152
rect 12504 8 12568 72
rect 12504 -72 12568 -8
rect 12504 -152 12568 -88
rect 12504 -232 12568 -168
rect 12504 -312 12568 -248
rect 12504 -392 12568 -328
rect 13916 328 13980 392
rect 13916 248 13980 312
rect 13916 168 13980 232
rect 13916 88 13980 152
rect 13916 8 13980 72
rect 13916 -72 13980 -8
rect 13916 -152 13980 -88
rect 13916 -232 13980 -168
rect 13916 -312 13980 -248
rect 13916 -392 13980 -328
rect 15328 328 15392 392
rect 15328 248 15392 312
rect 15328 168 15392 232
rect 15328 88 15392 152
rect 15328 8 15392 72
rect 15328 -72 15392 -8
rect 15328 -152 15392 -88
rect 15328 -232 15392 -168
rect 15328 -312 15392 -248
rect 15328 -392 15392 -328
rect 16740 328 16804 392
rect 16740 248 16804 312
rect 16740 168 16804 232
rect 16740 88 16804 152
rect 16740 8 16804 72
rect 16740 -72 16804 -8
rect 16740 -152 16804 -88
rect 16740 -232 16804 -168
rect 16740 -312 16804 -248
rect 16740 -392 16804 -328
rect 18152 328 18216 392
rect 18152 248 18216 312
rect 18152 168 18216 232
rect 18152 88 18216 152
rect 18152 8 18216 72
rect 18152 -72 18216 -8
rect 18152 -152 18216 -88
rect 18152 -232 18216 -168
rect 18152 -312 18216 -248
rect 18152 -392 18216 -328
rect 19564 328 19628 392
rect 19564 248 19628 312
rect 19564 168 19628 232
rect 19564 88 19628 152
rect 19564 8 19628 72
rect 19564 -72 19628 -8
rect 19564 -152 19628 -88
rect 19564 -232 19628 -168
rect 19564 -312 19628 -248
rect 19564 -392 19628 -328
rect 20976 328 21040 392
rect 20976 248 21040 312
rect 20976 168 21040 232
rect 20976 88 21040 152
rect 20976 8 21040 72
rect 20976 -72 21040 -8
rect 20976 -152 21040 -88
rect 20976 -232 21040 -168
rect 20976 -312 21040 -248
rect 20976 -392 21040 -328
rect 22388 328 22452 392
rect 22388 248 22452 312
rect 22388 168 22452 232
rect 22388 88 22452 152
rect 22388 8 22452 72
rect 22388 -72 22452 -8
rect 22388 -152 22452 -88
rect 22388 -232 22452 -168
rect 22388 -312 22452 -248
rect 22388 -392 22452 -328
rect 23800 328 23864 392
rect 23800 248 23864 312
rect 23800 168 23864 232
rect 23800 88 23864 152
rect 23800 8 23864 72
rect 23800 -72 23864 -8
rect 23800 -152 23864 -88
rect 23800 -232 23864 -168
rect 23800 -312 23864 -248
rect 23800 -392 23864 -328
rect -22796 -792 -22732 -728
rect -22796 -872 -22732 -808
rect -22796 -952 -22732 -888
rect -22796 -1032 -22732 -968
rect -22796 -1112 -22732 -1048
rect -22796 -1192 -22732 -1128
rect -22796 -1272 -22732 -1208
rect -22796 -1352 -22732 -1288
rect -22796 -1432 -22732 -1368
rect -22796 -1512 -22732 -1448
rect -21384 -792 -21320 -728
rect -21384 -872 -21320 -808
rect -21384 -952 -21320 -888
rect -21384 -1032 -21320 -968
rect -21384 -1112 -21320 -1048
rect -21384 -1192 -21320 -1128
rect -21384 -1272 -21320 -1208
rect -21384 -1352 -21320 -1288
rect -21384 -1432 -21320 -1368
rect -21384 -1512 -21320 -1448
rect -19972 -792 -19908 -728
rect -19972 -872 -19908 -808
rect -19972 -952 -19908 -888
rect -19972 -1032 -19908 -968
rect -19972 -1112 -19908 -1048
rect -19972 -1192 -19908 -1128
rect -19972 -1272 -19908 -1208
rect -19972 -1352 -19908 -1288
rect -19972 -1432 -19908 -1368
rect -19972 -1512 -19908 -1448
rect -18560 -792 -18496 -728
rect -18560 -872 -18496 -808
rect -18560 -952 -18496 -888
rect -18560 -1032 -18496 -968
rect -18560 -1112 -18496 -1048
rect -18560 -1192 -18496 -1128
rect -18560 -1272 -18496 -1208
rect -18560 -1352 -18496 -1288
rect -18560 -1432 -18496 -1368
rect -18560 -1512 -18496 -1448
rect -17148 -792 -17084 -728
rect -17148 -872 -17084 -808
rect -17148 -952 -17084 -888
rect -17148 -1032 -17084 -968
rect -17148 -1112 -17084 -1048
rect -17148 -1192 -17084 -1128
rect -17148 -1272 -17084 -1208
rect -17148 -1352 -17084 -1288
rect -17148 -1432 -17084 -1368
rect -17148 -1512 -17084 -1448
rect -15736 -792 -15672 -728
rect -15736 -872 -15672 -808
rect -15736 -952 -15672 -888
rect -15736 -1032 -15672 -968
rect -15736 -1112 -15672 -1048
rect -15736 -1192 -15672 -1128
rect -15736 -1272 -15672 -1208
rect -15736 -1352 -15672 -1288
rect -15736 -1432 -15672 -1368
rect -15736 -1512 -15672 -1448
rect -14324 -792 -14260 -728
rect -14324 -872 -14260 -808
rect -14324 -952 -14260 -888
rect -14324 -1032 -14260 -968
rect -14324 -1112 -14260 -1048
rect -14324 -1192 -14260 -1128
rect -14324 -1272 -14260 -1208
rect -14324 -1352 -14260 -1288
rect -14324 -1432 -14260 -1368
rect -14324 -1512 -14260 -1448
rect -12912 -792 -12848 -728
rect -12912 -872 -12848 -808
rect -12912 -952 -12848 -888
rect -12912 -1032 -12848 -968
rect -12912 -1112 -12848 -1048
rect -12912 -1192 -12848 -1128
rect -12912 -1272 -12848 -1208
rect -12912 -1352 -12848 -1288
rect -12912 -1432 -12848 -1368
rect -12912 -1512 -12848 -1448
rect -11500 -792 -11436 -728
rect -11500 -872 -11436 -808
rect -11500 -952 -11436 -888
rect -11500 -1032 -11436 -968
rect -11500 -1112 -11436 -1048
rect -11500 -1192 -11436 -1128
rect -11500 -1272 -11436 -1208
rect -11500 -1352 -11436 -1288
rect -11500 -1432 -11436 -1368
rect -11500 -1512 -11436 -1448
rect -10088 -792 -10024 -728
rect -10088 -872 -10024 -808
rect -10088 -952 -10024 -888
rect -10088 -1032 -10024 -968
rect -10088 -1112 -10024 -1048
rect -10088 -1192 -10024 -1128
rect -10088 -1272 -10024 -1208
rect -10088 -1352 -10024 -1288
rect -10088 -1432 -10024 -1368
rect -10088 -1512 -10024 -1448
rect -8676 -792 -8612 -728
rect -8676 -872 -8612 -808
rect -8676 -952 -8612 -888
rect -8676 -1032 -8612 -968
rect -8676 -1112 -8612 -1048
rect -8676 -1192 -8612 -1128
rect -8676 -1272 -8612 -1208
rect -8676 -1352 -8612 -1288
rect -8676 -1432 -8612 -1368
rect -8676 -1512 -8612 -1448
rect -7264 -792 -7200 -728
rect -7264 -872 -7200 -808
rect -7264 -952 -7200 -888
rect -7264 -1032 -7200 -968
rect -7264 -1112 -7200 -1048
rect -7264 -1192 -7200 -1128
rect -7264 -1272 -7200 -1208
rect -7264 -1352 -7200 -1288
rect -7264 -1432 -7200 -1368
rect -7264 -1512 -7200 -1448
rect -5852 -792 -5788 -728
rect -5852 -872 -5788 -808
rect -5852 -952 -5788 -888
rect -5852 -1032 -5788 -968
rect -5852 -1112 -5788 -1048
rect -5852 -1192 -5788 -1128
rect -5852 -1272 -5788 -1208
rect -5852 -1352 -5788 -1288
rect -5852 -1432 -5788 -1368
rect -5852 -1512 -5788 -1448
rect -4440 -792 -4376 -728
rect -4440 -872 -4376 -808
rect -4440 -952 -4376 -888
rect -4440 -1032 -4376 -968
rect -4440 -1112 -4376 -1048
rect -4440 -1192 -4376 -1128
rect -4440 -1272 -4376 -1208
rect -4440 -1352 -4376 -1288
rect -4440 -1432 -4376 -1368
rect -4440 -1512 -4376 -1448
rect -3028 -792 -2964 -728
rect -3028 -872 -2964 -808
rect -3028 -952 -2964 -888
rect -3028 -1032 -2964 -968
rect -3028 -1112 -2964 -1048
rect -3028 -1192 -2964 -1128
rect -3028 -1272 -2964 -1208
rect -3028 -1352 -2964 -1288
rect -3028 -1432 -2964 -1368
rect -3028 -1512 -2964 -1448
rect -1616 -792 -1552 -728
rect -1616 -872 -1552 -808
rect -1616 -952 -1552 -888
rect -1616 -1032 -1552 -968
rect -1616 -1112 -1552 -1048
rect -1616 -1192 -1552 -1128
rect -1616 -1272 -1552 -1208
rect -1616 -1352 -1552 -1288
rect -1616 -1432 -1552 -1368
rect -1616 -1512 -1552 -1448
rect -204 -792 -140 -728
rect -204 -872 -140 -808
rect -204 -952 -140 -888
rect -204 -1032 -140 -968
rect -204 -1112 -140 -1048
rect -204 -1192 -140 -1128
rect -204 -1272 -140 -1208
rect -204 -1352 -140 -1288
rect -204 -1432 -140 -1368
rect -204 -1512 -140 -1448
rect 1208 -792 1272 -728
rect 1208 -872 1272 -808
rect 1208 -952 1272 -888
rect 1208 -1032 1272 -968
rect 1208 -1112 1272 -1048
rect 1208 -1192 1272 -1128
rect 1208 -1272 1272 -1208
rect 1208 -1352 1272 -1288
rect 1208 -1432 1272 -1368
rect 1208 -1512 1272 -1448
rect 2620 -792 2684 -728
rect 2620 -872 2684 -808
rect 2620 -952 2684 -888
rect 2620 -1032 2684 -968
rect 2620 -1112 2684 -1048
rect 2620 -1192 2684 -1128
rect 2620 -1272 2684 -1208
rect 2620 -1352 2684 -1288
rect 2620 -1432 2684 -1368
rect 2620 -1512 2684 -1448
rect 4032 -792 4096 -728
rect 4032 -872 4096 -808
rect 4032 -952 4096 -888
rect 4032 -1032 4096 -968
rect 4032 -1112 4096 -1048
rect 4032 -1192 4096 -1128
rect 4032 -1272 4096 -1208
rect 4032 -1352 4096 -1288
rect 4032 -1432 4096 -1368
rect 4032 -1512 4096 -1448
rect 5444 -792 5508 -728
rect 5444 -872 5508 -808
rect 5444 -952 5508 -888
rect 5444 -1032 5508 -968
rect 5444 -1112 5508 -1048
rect 5444 -1192 5508 -1128
rect 5444 -1272 5508 -1208
rect 5444 -1352 5508 -1288
rect 5444 -1432 5508 -1368
rect 5444 -1512 5508 -1448
rect 6856 -792 6920 -728
rect 6856 -872 6920 -808
rect 6856 -952 6920 -888
rect 6856 -1032 6920 -968
rect 6856 -1112 6920 -1048
rect 6856 -1192 6920 -1128
rect 6856 -1272 6920 -1208
rect 6856 -1352 6920 -1288
rect 6856 -1432 6920 -1368
rect 6856 -1512 6920 -1448
rect 8268 -792 8332 -728
rect 8268 -872 8332 -808
rect 8268 -952 8332 -888
rect 8268 -1032 8332 -968
rect 8268 -1112 8332 -1048
rect 8268 -1192 8332 -1128
rect 8268 -1272 8332 -1208
rect 8268 -1352 8332 -1288
rect 8268 -1432 8332 -1368
rect 8268 -1512 8332 -1448
rect 9680 -792 9744 -728
rect 9680 -872 9744 -808
rect 9680 -952 9744 -888
rect 9680 -1032 9744 -968
rect 9680 -1112 9744 -1048
rect 9680 -1192 9744 -1128
rect 9680 -1272 9744 -1208
rect 9680 -1352 9744 -1288
rect 9680 -1432 9744 -1368
rect 9680 -1512 9744 -1448
rect 11092 -792 11156 -728
rect 11092 -872 11156 -808
rect 11092 -952 11156 -888
rect 11092 -1032 11156 -968
rect 11092 -1112 11156 -1048
rect 11092 -1192 11156 -1128
rect 11092 -1272 11156 -1208
rect 11092 -1352 11156 -1288
rect 11092 -1432 11156 -1368
rect 11092 -1512 11156 -1448
rect 12504 -792 12568 -728
rect 12504 -872 12568 -808
rect 12504 -952 12568 -888
rect 12504 -1032 12568 -968
rect 12504 -1112 12568 -1048
rect 12504 -1192 12568 -1128
rect 12504 -1272 12568 -1208
rect 12504 -1352 12568 -1288
rect 12504 -1432 12568 -1368
rect 12504 -1512 12568 -1448
rect 13916 -792 13980 -728
rect 13916 -872 13980 -808
rect 13916 -952 13980 -888
rect 13916 -1032 13980 -968
rect 13916 -1112 13980 -1048
rect 13916 -1192 13980 -1128
rect 13916 -1272 13980 -1208
rect 13916 -1352 13980 -1288
rect 13916 -1432 13980 -1368
rect 13916 -1512 13980 -1448
rect 15328 -792 15392 -728
rect 15328 -872 15392 -808
rect 15328 -952 15392 -888
rect 15328 -1032 15392 -968
rect 15328 -1112 15392 -1048
rect 15328 -1192 15392 -1128
rect 15328 -1272 15392 -1208
rect 15328 -1352 15392 -1288
rect 15328 -1432 15392 -1368
rect 15328 -1512 15392 -1448
rect 16740 -792 16804 -728
rect 16740 -872 16804 -808
rect 16740 -952 16804 -888
rect 16740 -1032 16804 -968
rect 16740 -1112 16804 -1048
rect 16740 -1192 16804 -1128
rect 16740 -1272 16804 -1208
rect 16740 -1352 16804 -1288
rect 16740 -1432 16804 -1368
rect 16740 -1512 16804 -1448
rect 18152 -792 18216 -728
rect 18152 -872 18216 -808
rect 18152 -952 18216 -888
rect 18152 -1032 18216 -968
rect 18152 -1112 18216 -1048
rect 18152 -1192 18216 -1128
rect 18152 -1272 18216 -1208
rect 18152 -1352 18216 -1288
rect 18152 -1432 18216 -1368
rect 18152 -1512 18216 -1448
rect 19564 -792 19628 -728
rect 19564 -872 19628 -808
rect 19564 -952 19628 -888
rect 19564 -1032 19628 -968
rect 19564 -1112 19628 -1048
rect 19564 -1192 19628 -1128
rect 19564 -1272 19628 -1208
rect 19564 -1352 19628 -1288
rect 19564 -1432 19628 -1368
rect 19564 -1512 19628 -1448
rect 20976 -792 21040 -728
rect 20976 -872 21040 -808
rect 20976 -952 21040 -888
rect 20976 -1032 21040 -968
rect 20976 -1112 21040 -1048
rect 20976 -1192 21040 -1128
rect 20976 -1272 21040 -1208
rect 20976 -1352 21040 -1288
rect 20976 -1432 21040 -1368
rect 20976 -1512 21040 -1448
rect 22388 -792 22452 -728
rect 22388 -872 22452 -808
rect 22388 -952 22452 -888
rect 22388 -1032 22452 -968
rect 22388 -1112 22452 -1048
rect 22388 -1192 22452 -1128
rect 22388 -1272 22452 -1208
rect 22388 -1352 22452 -1288
rect 22388 -1432 22452 -1368
rect 22388 -1512 22452 -1448
rect 23800 -792 23864 -728
rect 23800 -872 23864 -808
rect 23800 -952 23864 -888
rect 23800 -1032 23864 -968
rect 23800 -1112 23864 -1048
rect 23800 -1192 23864 -1128
rect 23800 -1272 23864 -1208
rect 23800 -1352 23864 -1288
rect 23800 -1432 23864 -1368
rect 23800 -1512 23864 -1448
rect -22796 -1912 -22732 -1848
rect -22796 -1992 -22732 -1928
rect -22796 -2072 -22732 -2008
rect -22796 -2152 -22732 -2088
rect -22796 -2232 -22732 -2168
rect -22796 -2312 -22732 -2248
rect -22796 -2392 -22732 -2328
rect -22796 -2472 -22732 -2408
rect -22796 -2552 -22732 -2488
rect -22796 -2632 -22732 -2568
rect -21384 -1912 -21320 -1848
rect -21384 -1992 -21320 -1928
rect -21384 -2072 -21320 -2008
rect -21384 -2152 -21320 -2088
rect -21384 -2232 -21320 -2168
rect -21384 -2312 -21320 -2248
rect -21384 -2392 -21320 -2328
rect -21384 -2472 -21320 -2408
rect -21384 -2552 -21320 -2488
rect -21384 -2632 -21320 -2568
rect -19972 -1912 -19908 -1848
rect -19972 -1992 -19908 -1928
rect -19972 -2072 -19908 -2008
rect -19972 -2152 -19908 -2088
rect -19972 -2232 -19908 -2168
rect -19972 -2312 -19908 -2248
rect -19972 -2392 -19908 -2328
rect -19972 -2472 -19908 -2408
rect -19972 -2552 -19908 -2488
rect -19972 -2632 -19908 -2568
rect -18560 -1912 -18496 -1848
rect -18560 -1992 -18496 -1928
rect -18560 -2072 -18496 -2008
rect -18560 -2152 -18496 -2088
rect -18560 -2232 -18496 -2168
rect -18560 -2312 -18496 -2248
rect -18560 -2392 -18496 -2328
rect -18560 -2472 -18496 -2408
rect -18560 -2552 -18496 -2488
rect -18560 -2632 -18496 -2568
rect -17148 -1912 -17084 -1848
rect -17148 -1992 -17084 -1928
rect -17148 -2072 -17084 -2008
rect -17148 -2152 -17084 -2088
rect -17148 -2232 -17084 -2168
rect -17148 -2312 -17084 -2248
rect -17148 -2392 -17084 -2328
rect -17148 -2472 -17084 -2408
rect -17148 -2552 -17084 -2488
rect -17148 -2632 -17084 -2568
rect -15736 -1912 -15672 -1848
rect -15736 -1992 -15672 -1928
rect -15736 -2072 -15672 -2008
rect -15736 -2152 -15672 -2088
rect -15736 -2232 -15672 -2168
rect -15736 -2312 -15672 -2248
rect -15736 -2392 -15672 -2328
rect -15736 -2472 -15672 -2408
rect -15736 -2552 -15672 -2488
rect -15736 -2632 -15672 -2568
rect -14324 -1912 -14260 -1848
rect -14324 -1992 -14260 -1928
rect -14324 -2072 -14260 -2008
rect -14324 -2152 -14260 -2088
rect -14324 -2232 -14260 -2168
rect -14324 -2312 -14260 -2248
rect -14324 -2392 -14260 -2328
rect -14324 -2472 -14260 -2408
rect -14324 -2552 -14260 -2488
rect -14324 -2632 -14260 -2568
rect -12912 -1912 -12848 -1848
rect -12912 -1992 -12848 -1928
rect -12912 -2072 -12848 -2008
rect -12912 -2152 -12848 -2088
rect -12912 -2232 -12848 -2168
rect -12912 -2312 -12848 -2248
rect -12912 -2392 -12848 -2328
rect -12912 -2472 -12848 -2408
rect -12912 -2552 -12848 -2488
rect -12912 -2632 -12848 -2568
rect -11500 -1912 -11436 -1848
rect -11500 -1992 -11436 -1928
rect -11500 -2072 -11436 -2008
rect -11500 -2152 -11436 -2088
rect -11500 -2232 -11436 -2168
rect -11500 -2312 -11436 -2248
rect -11500 -2392 -11436 -2328
rect -11500 -2472 -11436 -2408
rect -11500 -2552 -11436 -2488
rect -11500 -2632 -11436 -2568
rect -10088 -1912 -10024 -1848
rect -10088 -1992 -10024 -1928
rect -10088 -2072 -10024 -2008
rect -10088 -2152 -10024 -2088
rect -10088 -2232 -10024 -2168
rect -10088 -2312 -10024 -2248
rect -10088 -2392 -10024 -2328
rect -10088 -2472 -10024 -2408
rect -10088 -2552 -10024 -2488
rect -10088 -2632 -10024 -2568
rect -8676 -1912 -8612 -1848
rect -8676 -1992 -8612 -1928
rect -8676 -2072 -8612 -2008
rect -8676 -2152 -8612 -2088
rect -8676 -2232 -8612 -2168
rect -8676 -2312 -8612 -2248
rect -8676 -2392 -8612 -2328
rect -8676 -2472 -8612 -2408
rect -8676 -2552 -8612 -2488
rect -8676 -2632 -8612 -2568
rect -7264 -1912 -7200 -1848
rect -7264 -1992 -7200 -1928
rect -7264 -2072 -7200 -2008
rect -7264 -2152 -7200 -2088
rect -7264 -2232 -7200 -2168
rect -7264 -2312 -7200 -2248
rect -7264 -2392 -7200 -2328
rect -7264 -2472 -7200 -2408
rect -7264 -2552 -7200 -2488
rect -7264 -2632 -7200 -2568
rect -5852 -1912 -5788 -1848
rect -5852 -1992 -5788 -1928
rect -5852 -2072 -5788 -2008
rect -5852 -2152 -5788 -2088
rect -5852 -2232 -5788 -2168
rect -5852 -2312 -5788 -2248
rect -5852 -2392 -5788 -2328
rect -5852 -2472 -5788 -2408
rect -5852 -2552 -5788 -2488
rect -5852 -2632 -5788 -2568
rect -4440 -1912 -4376 -1848
rect -4440 -1992 -4376 -1928
rect -4440 -2072 -4376 -2008
rect -4440 -2152 -4376 -2088
rect -4440 -2232 -4376 -2168
rect -4440 -2312 -4376 -2248
rect -4440 -2392 -4376 -2328
rect -4440 -2472 -4376 -2408
rect -4440 -2552 -4376 -2488
rect -4440 -2632 -4376 -2568
rect -3028 -1912 -2964 -1848
rect -3028 -1992 -2964 -1928
rect -3028 -2072 -2964 -2008
rect -3028 -2152 -2964 -2088
rect -3028 -2232 -2964 -2168
rect -3028 -2312 -2964 -2248
rect -3028 -2392 -2964 -2328
rect -3028 -2472 -2964 -2408
rect -3028 -2552 -2964 -2488
rect -3028 -2632 -2964 -2568
rect -1616 -1912 -1552 -1848
rect -1616 -1992 -1552 -1928
rect -1616 -2072 -1552 -2008
rect -1616 -2152 -1552 -2088
rect -1616 -2232 -1552 -2168
rect -1616 -2312 -1552 -2248
rect -1616 -2392 -1552 -2328
rect -1616 -2472 -1552 -2408
rect -1616 -2552 -1552 -2488
rect -1616 -2632 -1552 -2568
rect -204 -1912 -140 -1848
rect -204 -1992 -140 -1928
rect -204 -2072 -140 -2008
rect -204 -2152 -140 -2088
rect -204 -2232 -140 -2168
rect -204 -2312 -140 -2248
rect -204 -2392 -140 -2328
rect -204 -2472 -140 -2408
rect -204 -2552 -140 -2488
rect -204 -2632 -140 -2568
rect 1208 -1912 1272 -1848
rect 1208 -1992 1272 -1928
rect 1208 -2072 1272 -2008
rect 1208 -2152 1272 -2088
rect 1208 -2232 1272 -2168
rect 1208 -2312 1272 -2248
rect 1208 -2392 1272 -2328
rect 1208 -2472 1272 -2408
rect 1208 -2552 1272 -2488
rect 1208 -2632 1272 -2568
rect 2620 -1912 2684 -1848
rect 2620 -1992 2684 -1928
rect 2620 -2072 2684 -2008
rect 2620 -2152 2684 -2088
rect 2620 -2232 2684 -2168
rect 2620 -2312 2684 -2248
rect 2620 -2392 2684 -2328
rect 2620 -2472 2684 -2408
rect 2620 -2552 2684 -2488
rect 2620 -2632 2684 -2568
rect 4032 -1912 4096 -1848
rect 4032 -1992 4096 -1928
rect 4032 -2072 4096 -2008
rect 4032 -2152 4096 -2088
rect 4032 -2232 4096 -2168
rect 4032 -2312 4096 -2248
rect 4032 -2392 4096 -2328
rect 4032 -2472 4096 -2408
rect 4032 -2552 4096 -2488
rect 4032 -2632 4096 -2568
rect 5444 -1912 5508 -1848
rect 5444 -1992 5508 -1928
rect 5444 -2072 5508 -2008
rect 5444 -2152 5508 -2088
rect 5444 -2232 5508 -2168
rect 5444 -2312 5508 -2248
rect 5444 -2392 5508 -2328
rect 5444 -2472 5508 -2408
rect 5444 -2552 5508 -2488
rect 5444 -2632 5508 -2568
rect 6856 -1912 6920 -1848
rect 6856 -1992 6920 -1928
rect 6856 -2072 6920 -2008
rect 6856 -2152 6920 -2088
rect 6856 -2232 6920 -2168
rect 6856 -2312 6920 -2248
rect 6856 -2392 6920 -2328
rect 6856 -2472 6920 -2408
rect 6856 -2552 6920 -2488
rect 6856 -2632 6920 -2568
rect 8268 -1912 8332 -1848
rect 8268 -1992 8332 -1928
rect 8268 -2072 8332 -2008
rect 8268 -2152 8332 -2088
rect 8268 -2232 8332 -2168
rect 8268 -2312 8332 -2248
rect 8268 -2392 8332 -2328
rect 8268 -2472 8332 -2408
rect 8268 -2552 8332 -2488
rect 8268 -2632 8332 -2568
rect 9680 -1912 9744 -1848
rect 9680 -1992 9744 -1928
rect 9680 -2072 9744 -2008
rect 9680 -2152 9744 -2088
rect 9680 -2232 9744 -2168
rect 9680 -2312 9744 -2248
rect 9680 -2392 9744 -2328
rect 9680 -2472 9744 -2408
rect 9680 -2552 9744 -2488
rect 9680 -2632 9744 -2568
rect 11092 -1912 11156 -1848
rect 11092 -1992 11156 -1928
rect 11092 -2072 11156 -2008
rect 11092 -2152 11156 -2088
rect 11092 -2232 11156 -2168
rect 11092 -2312 11156 -2248
rect 11092 -2392 11156 -2328
rect 11092 -2472 11156 -2408
rect 11092 -2552 11156 -2488
rect 11092 -2632 11156 -2568
rect 12504 -1912 12568 -1848
rect 12504 -1992 12568 -1928
rect 12504 -2072 12568 -2008
rect 12504 -2152 12568 -2088
rect 12504 -2232 12568 -2168
rect 12504 -2312 12568 -2248
rect 12504 -2392 12568 -2328
rect 12504 -2472 12568 -2408
rect 12504 -2552 12568 -2488
rect 12504 -2632 12568 -2568
rect 13916 -1912 13980 -1848
rect 13916 -1992 13980 -1928
rect 13916 -2072 13980 -2008
rect 13916 -2152 13980 -2088
rect 13916 -2232 13980 -2168
rect 13916 -2312 13980 -2248
rect 13916 -2392 13980 -2328
rect 13916 -2472 13980 -2408
rect 13916 -2552 13980 -2488
rect 13916 -2632 13980 -2568
rect 15328 -1912 15392 -1848
rect 15328 -1992 15392 -1928
rect 15328 -2072 15392 -2008
rect 15328 -2152 15392 -2088
rect 15328 -2232 15392 -2168
rect 15328 -2312 15392 -2248
rect 15328 -2392 15392 -2328
rect 15328 -2472 15392 -2408
rect 15328 -2552 15392 -2488
rect 15328 -2632 15392 -2568
rect 16740 -1912 16804 -1848
rect 16740 -1992 16804 -1928
rect 16740 -2072 16804 -2008
rect 16740 -2152 16804 -2088
rect 16740 -2232 16804 -2168
rect 16740 -2312 16804 -2248
rect 16740 -2392 16804 -2328
rect 16740 -2472 16804 -2408
rect 16740 -2552 16804 -2488
rect 16740 -2632 16804 -2568
rect 18152 -1912 18216 -1848
rect 18152 -1992 18216 -1928
rect 18152 -2072 18216 -2008
rect 18152 -2152 18216 -2088
rect 18152 -2232 18216 -2168
rect 18152 -2312 18216 -2248
rect 18152 -2392 18216 -2328
rect 18152 -2472 18216 -2408
rect 18152 -2552 18216 -2488
rect 18152 -2632 18216 -2568
rect 19564 -1912 19628 -1848
rect 19564 -1992 19628 -1928
rect 19564 -2072 19628 -2008
rect 19564 -2152 19628 -2088
rect 19564 -2232 19628 -2168
rect 19564 -2312 19628 -2248
rect 19564 -2392 19628 -2328
rect 19564 -2472 19628 -2408
rect 19564 -2552 19628 -2488
rect 19564 -2632 19628 -2568
rect 20976 -1912 21040 -1848
rect 20976 -1992 21040 -1928
rect 20976 -2072 21040 -2008
rect 20976 -2152 21040 -2088
rect 20976 -2232 21040 -2168
rect 20976 -2312 21040 -2248
rect 20976 -2392 21040 -2328
rect 20976 -2472 21040 -2408
rect 20976 -2552 21040 -2488
rect 20976 -2632 21040 -2568
rect 22388 -1912 22452 -1848
rect 22388 -1992 22452 -1928
rect 22388 -2072 22452 -2008
rect 22388 -2152 22452 -2088
rect 22388 -2232 22452 -2168
rect 22388 -2312 22452 -2248
rect 22388 -2392 22452 -2328
rect 22388 -2472 22452 -2408
rect 22388 -2552 22452 -2488
rect 22388 -2632 22452 -2568
rect 23800 -1912 23864 -1848
rect 23800 -1992 23864 -1928
rect 23800 -2072 23864 -2008
rect 23800 -2152 23864 -2088
rect 23800 -2232 23864 -2168
rect 23800 -2312 23864 -2248
rect 23800 -2392 23864 -2328
rect 23800 -2472 23864 -2408
rect 23800 -2552 23864 -2488
rect 23800 -2632 23864 -2568
rect -22796 -3032 -22732 -2968
rect -22796 -3112 -22732 -3048
rect -22796 -3192 -22732 -3128
rect -22796 -3272 -22732 -3208
rect -22796 -3352 -22732 -3288
rect -22796 -3432 -22732 -3368
rect -22796 -3512 -22732 -3448
rect -22796 -3592 -22732 -3528
rect -22796 -3672 -22732 -3608
rect -22796 -3752 -22732 -3688
rect -21384 -3032 -21320 -2968
rect -21384 -3112 -21320 -3048
rect -21384 -3192 -21320 -3128
rect -21384 -3272 -21320 -3208
rect -21384 -3352 -21320 -3288
rect -21384 -3432 -21320 -3368
rect -21384 -3512 -21320 -3448
rect -21384 -3592 -21320 -3528
rect -21384 -3672 -21320 -3608
rect -21384 -3752 -21320 -3688
rect -19972 -3032 -19908 -2968
rect -19972 -3112 -19908 -3048
rect -19972 -3192 -19908 -3128
rect -19972 -3272 -19908 -3208
rect -19972 -3352 -19908 -3288
rect -19972 -3432 -19908 -3368
rect -19972 -3512 -19908 -3448
rect -19972 -3592 -19908 -3528
rect -19972 -3672 -19908 -3608
rect -19972 -3752 -19908 -3688
rect -18560 -3032 -18496 -2968
rect -18560 -3112 -18496 -3048
rect -18560 -3192 -18496 -3128
rect -18560 -3272 -18496 -3208
rect -18560 -3352 -18496 -3288
rect -18560 -3432 -18496 -3368
rect -18560 -3512 -18496 -3448
rect -18560 -3592 -18496 -3528
rect -18560 -3672 -18496 -3608
rect -18560 -3752 -18496 -3688
rect -17148 -3032 -17084 -2968
rect -17148 -3112 -17084 -3048
rect -17148 -3192 -17084 -3128
rect -17148 -3272 -17084 -3208
rect -17148 -3352 -17084 -3288
rect -17148 -3432 -17084 -3368
rect -17148 -3512 -17084 -3448
rect -17148 -3592 -17084 -3528
rect -17148 -3672 -17084 -3608
rect -17148 -3752 -17084 -3688
rect -15736 -3032 -15672 -2968
rect -15736 -3112 -15672 -3048
rect -15736 -3192 -15672 -3128
rect -15736 -3272 -15672 -3208
rect -15736 -3352 -15672 -3288
rect -15736 -3432 -15672 -3368
rect -15736 -3512 -15672 -3448
rect -15736 -3592 -15672 -3528
rect -15736 -3672 -15672 -3608
rect -15736 -3752 -15672 -3688
rect -14324 -3032 -14260 -2968
rect -14324 -3112 -14260 -3048
rect -14324 -3192 -14260 -3128
rect -14324 -3272 -14260 -3208
rect -14324 -3352 -14260 -3288
rect -14324 -3432 -14260 -3368
rect -14324 -3512 -14260 -3448
rect -14324 -3592 -14260 -3528
rect -14324 -3672 -14260 -3608
rect -14324 -3752 -14260 -3688
rect -12912 -3032 -12848 -2968
rect -12912 -3112 -12848 -3048
rect -12912 -3192 -12848 -3128
rect -12912 -3272 -12848 -3208
rect -12912 -3352 -12848 -3288
rect -12912 -3432 -12848 -3368
rect -12912 -3512 -12848 -3448
rect -12912 -3592 -12848 -3528
rect -12912 -3672 -12848 -3608
rect -12912 -3752 -12848 -3688
rect -11500 -3032 -11436 -2968
rect -11500 -3112 -11436 -3048
rect -11500 -3192 -11436 -3128
rect -11500 -3272 -11436 -3208
rect -11500 -3352 -11436 -3288
rect -11500 -3432 -11436 -3368
rect -11500 -3512 -11436 -3448
rect -11500 -3592 -11436 -3528
rect -11500 -3672 -11436 -3608
rect -11500 -3752 -11436 -3688
rect -10088 -3032 -10024 -2968
rect -10088 -3112 -10024 -3048
rect -10088 -3192 -10024 -3128
rect -10088 -3272 -10024 -3208
rect -10088 -3352 -10024 -3288
rect -10088 -3432 -10024 -3368
rect -10088 -3512 -10024 -3448
rect -10088 -3592 -10024 -3528
rect -10088 -3672 -10024 -3608
rect -10088 -3752 -10024 -3688
rect -8676 -3032 -8612 -2968
rect -8676 -3112 -8612 -3048
rect -8676 -3192 -8612 -3128
rect -8676 -3272 -8612 -3208
rect -8676 -3352 -8612 -3288
rect -8676 -3432 -8612 -3368
rect -8676 -3512 -8612 -3448
rect -8676 -3592 -8612 -3528
rect -8676 -3672 -8612 -3608
rect -8676 -3752 -8612 -3688
rect -7264 -3032 -7200 -2968
rect -7264 -3112 -7200 -3048
rect -7264 -3192 -7200 -3128
rect -7264 -3272 -7200 -3208
rect -7264 -3352 -7200 -3288
rect -7264 -3432 -7200 -3368
rect -7264 -3512 -7200 -3448
rect -7264 -3592 -7200 -3528
rect -7264 -3672 -7200 -3608
rect -7264 -3752 -7200 -3688
rect -5852 -3032 -5788 -2968
rect -5852 -3112 -5788 -3048
rect -5852 -3192 -5788 -3128
rect -5852 -3272 -5788 -3208
rect -5852 -3352 -5788 -3288
rect -5852 -3432 -5788 -3368
rect -5852 -3512 -5788 -3448
rect -5852 -3592 -5788 -3528
rect -5852 -3672 -5788 -3608
rect -5852 -3752 -5788 -3688
rect -4440 -3032 -4376 -2968
rect -4440 -3112 -4376 -3048
rect -4440 -3192 -4376 -3128
rect -4440 -3272 -4376 -3208
rect -4440 -3352 -4376 -3288
rect -4440 -3432 -4376 -3368
rect -4440 -3512 -4376 -3448
rect -4440 -3592 -4376 -3528
rect -4440 -3672 -4376 -3608
rect -4440 -3752 -4376 -3688
rect -3028 -3032 -2964 -2968
rect -3028 -3112 -2964 -3048
rect -3028 -3192 -2964 -3128
rect -3028 -3272 -2964 -3208
rect -3028 -3352 -2964 -3288
rect -3028 -3432 -2964 -3368
rect -3028 -3512 -2964 -3448
rect -3028 -3592 -2964 -3528
rect -3028 -3672 -2964 -3608
rect -3028 -3752 -2964 -3688
rect -1616 -3032 -1552 -2968
rect -1616 -3112 -1552 -3048
rect -1616 -3192 -1552 -3128
rect -1616 -3272 -1552 -3208
rect -1616 -3352 -1552 -3288
rect -1616 -3432 -1552 -3368
rect -1616 -3512 -1552 -3448
rect -1616 -3592 -1552 -3528
rect -1616 -3672 -1552 -3608
rect -1616 -3752 -1552 -3688
rect -204 -3032 -140 -2968
rect -204 -3112 -140 -3048
rect -204 -3192 -140 -3128
rect -204 -3272 -140 -3208
rect -204 -3352 -140 -3288
rect -204 -3432 -140 -3368
rect -204 -3512 -140 -3448
rect -204 -3592 -140 -3528
rect -204 -3672 -140 -3608
rect -204 -3752 -140 -3688
rect 1208 -3032 1272 -2968
rect 1208 -3112 1272 -3048
rect 1208 -3192 1272 -3128
rect 1208 -3272 1272 -3208
rect 1208 -3352 1272 -3288
rect 1208 -3432 1272 -3368
rect 1208 -3512 1272 -3448
rect 1208 -3592 1272 -3528
rect 1208 -3672 1272 -3608
rect 1208 -3752 1272 -3688
rect 2620 -3032 2684 -2968
rect 2620 -3112 2684 -3048
rect 2620 -3192 2684 -3128
rect 2620 -3272 2684 -3208
rect 2620 -3352 2684 -3288
rect 2620 -3432 2684 -3368
rect 2620 -3512 2684 -3448
rect 2620 -3592 2684 -3528
rect 2620 -3672 2684 -3608
rect 2620 -3752 2684 -3688
rect 4032 -3032 4096 -2968
rect 4032 -3112 4096 -3048
rect 4032 -3192 4096 -3128
rect 4032 -3272 4096 -3208
rect 4032 -3352 4096 -3288
rect 4032 -3432 4096 -3368
rect 4032 -3512 4096 -3448
rect 4032 -3592 4096 -3528
rect 4032 -3672 4096 -3608
rect 4032 -3752 4096 -3688
rect 5444 -3032 5508 -2968
rect 5444 -3112 5508 -3048
rect 5444 -3192 5508 -3128
rect 5444 -3272 5508 -3208
rect 5444 -3352 5508 -3288
rect 5444 -3432 5508 -3368
rect 5444 -3512 5508 -3448
rect 5444 -3592 5508 -3528
rect 5444 -3672 5508 -3608
rect 5444 -3752 5508 -3688
rect 6856 -3032 6920 -2968
rect 6856 -3112 6920 -3048
rect 6856 -3192 6920 -3128
rect 6856 -3272 6920 -3208
rect 6856 -3352 6920 -3288
rect 6856 -3432 6920 -3368
rect 6856 -3512 6920 -3448
rect 6856 -3592 6920 -3528
rect 6856 -3672 6920 -3608
rect 6856 -3752 6920 -3688
rect 8268 -3032 8332 -2968
rect 8268 -3112 8332 -3048
rect 8268 -3192 8332 -3128
rect 8268 -3272 8332 -3208
rect 8268 -3352 8332 -3288
rect 8268 -3432 8332 -3368
rect 8268 -3512 8332 -3448
rect 8268 -3592 8332 -3528
rect 8268 -3672 8332 -3608
rect 8268 -3752 8332 -3688
rect 9680 -3032 9744 -2968
rect 9680 -3112 9744 -3048
rect 9680 -3192 9744 -3128
rect 9680 -3272 9744 -3208
rect 9680 -3352 9744 -3288
rect 9680 -3432 9744 -3368
rect 9680 -3512 9744 -3448
rect 9680 -3592 9744 -3528
rect 9680 -3672 9744 -3608
rect 9680 -3752 9744 -3688
rect 11092 -3032 11156 -2968
rect 11092 -3112 11156 -3048
rect 11092 -3192 11156 -3128
rect 11092 -3272 11156 -3208
rect 11092 -3352 11156 -3288
rect 11092 -3432 11156 -3368
rect 11092 -3512 11156 -3448
rect 11092 -3592 11156 -3528
rect 11092 -3672 11156 -3608
rect 11092 -3752 11156 -3688
rect 12504 -3032 12568 -2968
rect 12504 -3112 12568 -3048
rect 12504 -3192 12568 -3128
rect 12504 -3272 12568 -3208
rect 12504 -3352 12568 -3288
rect 12504 -3432 12568 -3368
rect 12504 -3512 12568 -3448
rect 12504 -3592 12568 -3528
rect 12504 -3672 12568 -3608
rect 12504 -3752 12568 -3688
rect 13916 -3032 13980 -2968
rect 13916 -3112 13980 -3048
rect 13916 -3192 13980 -3128
rect 13916 -3272 13980 -3208
rect 13916 -3352 13980 -3288
rect 13916 -3432 13980 -3368
rect 13916 -3512 13980 -3448
rect 13916 -3592 13980 -3528
rect 13916 -3672 13980 -3608
rect 13916 -3752 13980 -3688
rect 15328 -3032 15392 -2968
rect 15328 -3112 15392 -3048
rect 15328 -3192 15392 -3128
rect 15328 -3272 15392 -3208
rect 15328 -3352 15392 -3288
rect 15328 -3432 15392 -3368
rect 15328 -3512 15392 -3448
rect 15328 -3592 15392 -3528
rect 15328 -3672 15392 -3608
rect 15328 -3752 15392 -3688
rect 16740 -3032 16804 -2968
rect 16740 -3112 16804 -3048
rect 16740 -3192 16804 -3128
rect 16740 -3272 16804 -3208
rect 16740 -3352 16804 -3288
rect 16740 -3432 16804 -3368
rect 16740 -3512 16804 -3448
rect 16740 -3592 16804 -3528
rect 16740 -3672 16804 -3608
rect 16740 -3752 16804 -3688
rect 18152 -3032 18216 -2968
rect 18152 -3112 18216 -3048
rect 18152 -3192 18216 -3128
rect 18152 -3272 18216 -3208
rect 18152 -3352 18216 -3288
rect 18152 -3432 18216 -3368
rect 18152 -3512 18216 -3448
rect 18152 -3592 18216 -3528
rect 18152 -3672 18216 -3608
rect 18152 -3752 18216 -3688
rect 19564 -3032 19628 -2968
rect 19564 -3112 19628 -3048
rect 19564 -3192 19628 -3128
rect 19564 -3272 19628 -3208
rect 19564 -3352 19628 -3288
rect 19564 -3432 19628 -3368
rect 19564 -3512 19628 -3448
rect 19564 -3592 19628 -3528
rect 19564 -3672 19628 -3608
rect 19564 -3752 19628 -3688
rect 20976 -3032 21040 -2968
rect 20976 -3112 21040 -3048
rect 20976 -3192 21040 -3128
rect 20976 -3272 21040 -3208
rect 20976 -3352 21040 -3288
rect 20976 -3432 21040 -3368
rect 20976 -3512 21040 -3448
rect 20976 -3592 21040 -3528
rect 20976 -3672 21040 -3608
rect 20976 -3752 21040 -3688
rect 22388 -3032 22452 -2968
rect 22388 -3112 22452 -3048
rect 22388 -3192 22452 -3128
rect 22388 -3272 22452 -3208
rect 22388 -3352 22452 -3288
rect 22388 -3432 22452 -3368
rect 22388 -3512 22452 -3448
rect 22388 -3592 22452 -3528
rect 22388 -3672 22452 -3608
rect 22388 -3752 22452 -3688
rect 23800 -3032 23864 -2968
rect 23800 -3112 23864 -3048
rect 23800 -3192 23864 -3128
rect 23800 -3272 23864 -3208
rect 23800 -3352 23864 -3288
rect 23800 -3432 23864 -3368
rect 23800 -3512 23864 -3448
rect 23800 -3592 23864 -3528
rect 23800 -3672 23864 -3608
rect 23800 -3752 23864 -3688
rect -22796 -4152 -22732 -4088
rect -22796 -4232 -22732 -4168
rect -22796 -4312 -22732 -4248
rect -22796 -4392 -22732 -4328
rect -22796 -4472 -22732 -4408
rect -22796 -4552 -22732 -4488
rect -22796 -4632 -22732 -4568
rect -22796 -4712 -22732 -4648
rect -22796 -4792 -22732 -4728
rect -22796 -4872 -22732 -4808
rect -21384 -4152 -21320 -4088
rect -21384 -4232 -21320 -4168
rect -21384 -4312 -21320 -4248
rect -21384 -4392 -21320 -4328
rect -21384 -4472 -21320 -4408
rect -21384 -4552 -21320 -4488
rect -21384 -4632 -21320 -4568
rect -21384 -4712 -21320 -4648
rect -21384 -4792 -21320 -4728
rect -21384 -4872 -21320 -4808
rect -19972 -4152 -19908 -4088
rect -19972 -4232 -19908 -4168
rect -19972 -4312 -19908 -4248
rect -19972 -4392 -19908 -4328
rect -19972 -4472 -19908 -4408
rect -19972 -4552 -19908 -4488
rect -19972 -4632 -19908 -4568
rect -19972 -4712 -19908 -4648
rect -19972 -4792 -19908 -4728
rect -19972 -4872 -19908 -4808
rect -18560 -4152 -18496 -4088
rect -18560 -4232 -18496 -4168
rect -18560 -4312 -18496 -4248
rect -18560 -4392 -18496 -4328
rect -18560 -4472 -18496 -4408
rect -18560 -4552 -18496 -4488
rect -18560 -4632 -18496 -4568
rect -18560 -4712 -18496 -4648
rect -18560 -4792 -18496 -4728
rect -18560 -4872 -18496 -4808
rect -17148 -4152 -17084 -4088
rect -17148 -4232 -17084 -4168
rect -17148 -4312 -17084 -4248
rect -17148 -4392 -17084 -4328
rect -17148 -4472 -17084 -4408
rect -17148 -4552 -17084 -4488
rect -17148 -4632 -17084 -4568
rect -17148 -4712 -17084 -4648
rect -17148 -4792 -17084 -4728
rect -17148 -4872 -17084 -4808
rect -15736 -4152 -15672 -4088
rect -15736 -4232 -15672 -4168
rect -15736 -4312 -15672 -4248
rect -15736 -4392 -15672 -4328
rect -15736 -4472 -15672 -4408
rect -15736 -4552 -15672 -4488
rect -15736 -4632 -15672 -4568
rect -15736 -4712 -15672 -4648
rect -15736 -4792 -15672 -4728
rect -15736 -4872 -15672 -4808
rect -14324 -4152 -14260 -4088
rect -14324 -4232 -14260 -4168
rect -14324 -4312 -14260 -4248
rect -14324 -4392 -14260 -4328
rect -14324 -4472 -14260 -4408
rect -14324 -4552 -14260 -4488
rect -14324 -4632 -14260 -4568
rect -14324 -4712 -14260 -4648
rect -14324 -4792 -14260 -4728
rect -14324 -4872 -14260 -4808
rect -12912 -4152 -12848 -4088
rect -12912 -4232 -12848 -4168
rect -12912 -4312 -12848 -4248
rect -12912 -4392 -12848 -4328
rect -12912 -4472 -12848 -4408
rect -12912 -4552 -12848 -4488
rect -12912 -4632 -12848 -4568
rect -12912 -4712 -12848 -4648
rect -12912 -4792 -12848 -4728
rect -12912 -4872 -12848 -4808
rect -11500 -4152 -11436 -4088
rect -11500 -4232 -11436 -4168
rect -11500 -4312 -11436 -4248
rect -11500 -4392 -11436 -4328
rect -11500 -4472 -11436 -4408
rect -11500 -4552 -11436 -4488
rect -11500 -4632 -11436 -4568
rect -11500 -4712 -11436 -4648
rect -11500 -4792 -11436 -4728
rect -11500 -4872 -11436 -4808
rect -10088 -4152 -10024 -4088
rect -10088 -4232 -10024 -4168
rect -10088 -4312 -10024 -4248
rect -10088 -4392 -10024 -4328
rect -10088 -4472 -10024 -4408
rect -10088 -4552 -10024 -4488
rect -10088 -4632 -10024 -4568
rect -10088 -4712 -10024 -4648
rect -10088 -4792 -10024 -4728
rect -10088 -4872 -10024 -4808
rect -8676 -4152 -8612 -4088
rect -8676 -4232 -8612 -4168
rect -8676 -4312 -8612 -4248
rect -8676 -4392 -8612 -4328
rect -8676 -4472 -8612 -4408
rect -8676 -4552 -8612 -4488
rect -8676 -4632 -8612 -4568
rect -8676 -4712 -8612 -4648
rect -8676 -4792 -8612 -4728
rect -8676 -4872 -8612 -4808
rect -7264 -4152 -7200 -4088
rect -7264 -4232 -7200 -4168
rect -7264 -4312 -7200 -4248
rect -7264 -4392 -7200 -4328
rect -7264 -4472 -7200 -4408
rect -7264 -4552 -7200 -4488
rect -7264 -4632 -7200 -4568
rect -7264 -4712 -7200 -4648
rect -7264 -4792 -7200 -4728
rect -7264 -4872 -7200 -4808
rect -5852 -4152 -5788 -4088
rect -5852 -4232 -5788 -4168
rect -5852 -4312 -5788 -4248
rect -5852 -4392 -5788 -4328
rect -5852 -4472 -5788 -4408
rect -5852 -4552 -5788 -4488
rect -5852 -4632 -5788 -4568
rect -5852 -4712 -5788 -4648
rect -5852 -4792 -5788 -4728
rect -5852 -4872 -5788 -4808
rect -4440 -4152 -4376 -4088
rect -4440 -4232 -4376 -4168
rect -4440 -4312 -4376 -4248
rect -4440 -4392 -4376 -4328
rect -4440 -4472 -4376 -4408
rect -4440 -4552 -4376 -4488
rect -4440 -4632 -4376 -4568
rect -4440 -4712 -4376 -4648
rect -4440 -4792 -4376 -4728
rect -4440 -4872 -4376 -4808
rect -3028 -4152 -2964 -4088
rect -3028 -4232 -2964 -4168
rect -3028 -4312 -2964 -4248
rect -3028 -4392 -2964 -4328
rect -3028 -4472 -2964 -4408
rect -3028 -4552 -2964 -4488
rect -3028 -4632 -2964 -4568
rect -3028 -4712 -2964 -4648
rect -3028 -4792 -2964 -4728
rect -3028 -4872 -2964 -4808
rect -1616 -4152 -1552 -4088
rect -1616 -4232 -1552 -4168
rect -1616 -4312 -1552 -4248
rect -1616 -4392 -1552 -4328
rect -1616 -4472 -1552 -4408
rect -1616 -4552 -1552 -4488
rect -1616 -4632 -1552 -4568
rect -1616 -4712 -1552 -4648
rect -1616 -4792 -1552 -4728
rect -1616 -4872 -1552 -4808
rect -204 -4152 -140 -4088
rect -204 -4232 -140 -4168
rect -204 -4312 -140 -4248
rect -204 -4392 -140 -4328
rect -204 -4472 -140 -4408
rect -204 -4552 -140 -4488
rect -204 -4632 -140 -4568
rect -204 -4712 -140 -4648
rect -204 -4792 -140 -4728
rect -204 -4872 -140 -4808
rect 1208 -4152 1272 -4088
rect 1208 -4232 1272 -4168
rect 1208 -4312 1272 -4248
rect 1208 -4392 1272 -4328
rect 1208 -4472 1272 -4408
rect 1208 -4552 1272 -4488
rect 1208 -4632 1272 -4568
rect 1208 -4712 1272 -4648
rect 1208 -4792 1272 -4728
rect 1208 -4872 1272 -4808
rect 2620 -4152 2684 -4088
rect 2620 -4232 2684 -4168
rect 2620 -4312 2684 -4248
rect 2620 -4392 2684 -4328
rect 2620 -4472 2684 -4408
rect 2620 -4552 2684 -4488
rect 2620 -4632 2684 -4568
rect 2620 -4712 2684 -4648
rect 2620 -4792 2684 -4728
rect 2620 -4872 2684 -4808
rect 4032 -4152 4096 -4088
rect 4032 -4232 4096 -4168
rect 4032 -4312 4096 -4248
rect 4032 -4392 4096 -4328
rect 4032 -4472 4096 -4408
rect 4032 -4552 4096 -4488
rect 4032 -4632 4096 -4568
rect 4032 -4712 4096 -4648
rect 4032 -4792 4096 -4728
rect 4032 -4872 4096 -4808
rect 5444 -4152 5508 -4088
rect 5444 -4232 5508 -4168
rect 5444 -4312 5508 -4248
rect 5444 -4392 5508 -4328
rect 5444 -4472 5508 -4408
rect 5444 -4552 5508 -4488
rect 5444 -4632 5508 -4568
rect 5444 -4712 5508 -4648
rect 5444 -4792 5508 -4728
rect 5444 -4872 5508 -4808
rect 6856 -4152 6920 -4088
rect 6856 -4232 6920 -4168
rect 6856 -4312 6920 -4248
rect 6856 -4392 6920 -4328
rect 6856 -4472 6920 -4408
rect 6856 -4552 6920 -4488
rect 6856 -4632 6920 -4568
rect 6856 -4712 6920 -4648
rect 6856 -4792 6920 -4728
rect 6856 -4872 6920 -4808
rect 8268 -4152 8332 -4088
rect 8268 -4232 8332 -4168
rect 8268 -4312 8332 -4248
rect 8268 -4392 8332 -4328
rect 8268 -4472 8332 -4408
rect 8268 -4552 8332 -4488
rect 8268 -4632 8332 -4568
rect 8268 -4712 8332 -4648
rect 8268 -4792 8332 -4728
rect 8268 -4872 8332 -4808
rect 9680 -4152 9744 -4088
rect 9680 -4232 9744 -4168
rect 9680 -4312 9744 -4248
rect 9680 -4392 9744 -4328
rect 9680 -4472 9744 -4408
rect 9680 -4552 9744 -4488
rect 9680 -4632 9744 -4568
rect 9680 -4712 9744 -4648
rect 9680 -4792 9744 -4728
rect 9680 -4872 9744 -4808
rect 11092 -4152 11156 -4088
rect 11092 -4232 11156 -4168
rect 11092 -4312 11156 -4248
rect 11092 -4392 11156 -4328
rect 11092 -4472 11156 -4408
rect 11092 -4552 11156 -4488
rect 11092 -4632 11156 -4568
rect 11092 -4712 11156 -4648
rect 11092 -4792 11156 -4728
rect 11092 -4872 11156 -4808
rect 12504 -4152 12568 -4088
rect 12504 -4232 12568 -4168
rect 12504 -4312 12568 -4248
rect 12504 -4392 12568 -4328
rect 12504 -4472 12568 -4408
rect 12504 -4552 12568 -4488
rect 12504 -4632 12568 -4568
rect 12504 -4712 12568 -4648
rect 12504 -4792 12568 -4728
rect 12504 -4872 12568 -4808
rect 13916 -4152 13980 -4088
rect 13916 -4232 13980 -4168
rect 13916 -4312 13980 -4248
rect 13916 -4392 13980 -4328
rect 13916 -4472 13980 -4408
rect 13916 -4552 13980 -4488
rect 13916 -4632 13980 -4568
rect 13916 -4712 13980 -4648
rect 13916 -4792 13980 -4728
rect 13916 -4872 13980 -4808
rect 15328 -4152 15392 -4088
rect 15328 -4232 15392 -4168
rect 15328 -4312 15392 -4248
rect 15328 -4392 15392 -4328
rect 15328 -4472 15392 -4408
rect 15328 -4552 15392 -4488
rect 15328 -4632 15392 -4568
rect 15328 -4712 15392 -4648
rect 15328 -4792 15392 -4728
rect 15328 -4872 15392 -4808
rect 16740 -4152 16804 -4088
rect 16740 -4232 16804 -4168
rect 16740 -4312 16804 -4248
rect 16740 -4392 16804 -4328
rect 16740 -4472 16804 -4408
rect 16740 -4552 16804 -4488
rect 16740 -4632 16804 -4568
rect 16740 -4712 16804 -4648
rect 16740 -4792 16804 -4728
rect 16740 -4872 16804 -4808
rect 18152 -4152 18216 -4088
rect 18152 -4232 18216 -4168
rect 18152 -4312 18216 -4248
rect 18152 -4392 18216 -4328
rect 18152 -4472 18216 -4408
rect 18152 -4552 18216 -4488
rect 18152 -4632 18216 -4568
rect 18152 -4712 18216 -4648
rect 18152 -4792 18216 -4728
rect 18152 -4872 18216 -4808
rect 19564 -4152 19628 -4088
rect 19564 -4232 19628 -4168
rect 19564 -4312 19628 -4248
rect 19564 -4392 19628 -4328
rect 19564 -4472 19628 -4408
rect 19564 -4552 19628 -4488
rect 19564 -4632 19628 -4568
rect 19564 -4712 19628 -4648
rect 19564 -4792 19628 -4728
rect 19564 -4872 19628 -4808
rect 20976 -4152 21040 -4088
rect 20976 -4232 21040 -4168
rect 20976 -4312 21040 -4248
rect 20976 -4392 21040 -4328
rect 20976 -4472 21040 -4408
rect 20976 -4552 21040 -4488
rect 20976 -4632 21040 -4568
rect 20976 -4712 21040 -4648
rect 20976 -4792 21040 -4728
rect 20976 -4872 21040 -4808
rect 22388 -4152 22452 -4088
rect 22388 -4232 22452 -4168
rect 22388 -4312 22452 -4248
rect 22388 -4392 22452 -4328
rect 22388 -4472 22452 -4408
rect 22388 -4552 22452 -4488
rect 22388 -4632 22452 -4568
rect 22388 -4712 22452 -4648
rect 22388 -4792 22452 -4728
rect 22388 -4872 22452 -4808
rect 23800 -4152 23864 -4088
rect 23800 -4232 23864 -4168
rect 23800 -4312 23864 -4248
rect 23800 -4392 23864 -4328
rect 23800 -4472 23864 -4408
rect 23800 -4552 23864 -4488
rect 23800 -4632 23864 -4568
rect 23800 -4712 23864 -4648
rect 23800 -4792 23864 -4728
rect 23800 -4872 23864 -4808
rect -22796 -5272 -22732 -5208
rect -22796 -5352 -22732 -5288
rect -22796 -5432 -22732 -5368
rect -22796 -5512 -22732 -5448
rect -22796 -5592 -22732 -5528
rect -22796 -5672 -22732 -5608
rect -22796 -5752 -22732 -5688
rect -22796 -5832 -22732 -5768
rect -22796 -5912 -22732 -5848
rect -22796 -5992 -22732 -5928
rect -21384 -5272 -21320 -5208
rect -21384 -5352 -21320 -5288
rect -21384 -5432 -21320 -5368
rect -21384 -5512 -21320 -5448
rect -21384 -5592 -21320 -5528
rect -21384 -5672 -21320 -5608
rect -21384 -5752 -21320 -5688
rect -21384 -5832 -21320 -5768
rect -21384 -5912 -21320 -5848
rect -21384 -5992 -21320 -5928
rect -19972 -5272 -19908 -5208
rect -19972 -5352 -19908 -5288
rect -19972 -5432 -19908 -5368
rect -19972 -5512 -19908 -5448
rect -19972 -5592 -19908 -5528
rect -19972 -5672 -19908 -5608
rect -19972 -5752 -19908 -5688
rect -19972 -5832 -19908 -5768
rect -19972 -5912 -19908 -5848
rect -19972 -5992 -19908 -5928
rect -18560 -5272 -18496 -5208
rect -18560 -5352 -18496 -5288
rect -18560 -5432 -18496 -5368
rect -18560 -5512 -18496 -5448
rect -18560 -5592 -18496 -5528
rect -18560 -5672 -18496 -5608
rect -18560 -5752 -18496 -5688
rect -18560 -5832 -18496 -5768
rect -18560 -5912 -18496 -5848
rect -18560 -5992 -18496 -5928
rect -17148 -5272 -17084 -5208
rect -17148 -5352 -17084 -5288
rect -17148 -5432 -17084 -5368
rect -17148 -5512 -17084 -5448
rect -17148 -5592 -17084 -5528
rect -17148 -5672 -17084 -5608
rect -17148 -5752 -17084 -5688
rect -17148 -5832 -17084 -5768
rect -17148 -5912 -17084 -5848
rect -17148 -5992 -17084 -5928
rect -15736 -5272 -15672 -5208
rect -15736 -5352 -15672 -5288
rect -15736 -5432 -15672 -5368
rect -15736 -5512 -15672 -5448
rect -15736 -5592 -15672 -5528
rect -15736 -5672 -15672 -5608
rect -15736 -5752 -15672 -5688
rect -15736 -5832 -15672 -5768
rect -15736 -5912 -15672 -5848
rect -15736 -5992 -15672 -5928
rect -14324 -5272 -14260 -5208
rect -14324 -5352 -14260 -5288
rect -14324 -5432 -14260 -5368
rect -14324 -5512 -14260 -5448
rect -14324 -5592 -14260 -5528
rect -14324 -5672 -14260 -5608
rect -14324 -5752 -14260 -5688
rect -14324 -5832 -14260 -5768
rect -14324 -5912 -14260 -5848
rect -14324 -5992 -14260 -5928
rect -12912 -5272 -12848 -5208
rect -12912 -5352 -12848 -5288
rect -12912 -5432 -12848 -5368
rect -12912 -5512 -12848 -5448
rect -12912 -5592 -12848 -5528
rect -12912 -5672 -12848 -5608
rect -12912 -5752 -12848 -5688
rect -12912 -5832 -12848 -5768
rect -12912 -5912 -12848 -5848
rect -12912 -5992 -12848 -5928
rect -11500 -5272 -11436 -5208
rect -11500 -5352 -11436 -5288
rect -11500 -5432 -11436 -5368
rect -11500 -5512 -11436 -5448
rect -11500 -5592 -11436 -5528
rect -11500 -5672 -11436 -5608
rect -11500 -5752 -11436 -5688
rect -11500 -5832 -11436 -5768
rect -11500 -5912 -11436 -5848
rect -11500 -5992 -11436 -5928
rect -10088 -5272 -10024 -5208
rect -10088 -5352 -10024 -5288
rect -10088 -5432 -10024 -5368
rect -10088 -5512 -10024 -5448
rect -10088 -5592 -10024 -5528
rect -10088 -5672 -10024 -5608
rect -10088 -5752 -10024 -5688
rect -10088 -5832 -10024 -5768
rect -10088 -5912 -10024 -5848
rect -10088 -5992 -10024 -5928
rect -8676 -5272 -8612 -5208
rect -8676 -5352 -8612 -5288
rect -8676 -5432 -8612 -5368
rect -8676 -5512 -8612 -5448
rect -8676 -5592 -8612 -5528
rect -8676 -5672 -8612 -5608
rect -8676 -5752 -8612 -5688
rect -8676 -5832 -8612 -5768
rect -8676 -5912 -8612 -5848
rect -8676 -5992 -8612 -5928
rect -7264 -5272 -7200 -5208
rect -7264 -5352 -7200 -5288
rect -7264 -5432 -7200 -5368
rect -7264 -5512 -7200 -5448
rect -7264 -5592 -7200 -5528
rect -7264 -5672 -7200 -5608
rect -7264 -5752 -7200 -5688
rect -7264 -5832 -7200 -5768
rect -7264 -5912 -7200 -5848
rect -7264 -5992 -7200 -5928
rect -5852 -5272 -5788 -5208
rect -5852 -5352 -5788 -5288
rect -5852 -5432 -5788 -5368
rect -5852 -5512 -5788 -5448
rect -5852 -5592 -5788 -5528
rect -5852 -5672 -5788 -5608
rect -5852 -5752 -5788 -5688
rect -5852 -5832 -5788 -5768
rect -5852 -5912 -5788 -5848
rect -5852 -5992 -5788 -5928
rect -4440 -5272 -4376 -5208
rect -4440 -5352 -4376 -5288
rect -4440 -5432 -4376 -5368
rect -4440 -5512 -4376 -5448
rect -4440 -5592 -4376 -5528
rect -4440 -5672 -4376 -5608
rect -4440 -5752 -4376 -5688
rect -4440 -5832 -4376 -5768
rect -4440 -5912 -4376 -5848
rect -4440 -5992 -4376 -5928
rect -3028 -5272 -2964 -5208
rect -3028 -5352 -2964 -5288
rect -3028 -5432 -2964 -5368
rect -3028 -5512 -2964 -5448
rect -3028 -5592 -2964 -5528
rect -3028 -5672 -2964 -5608
rect -3028 -5752 -2964 -5688
rect -3028 -5832 -2964 -5768
rect -3028 -5912 -2964 -5848
rect -3028 -5992 -2964 -5928
rect -1616 -5272 -1552 -5208
rect -1616 -5352 -1552 -5288
rect -1616 -5432 -1552 -5368
rect -1616 -5512 -1552 -5448
rect -1616 -5592 -1552 -5528
rect -1616 -5672 -1552 -5608
rect -1616 -5752 -1552 -5688
rect -1616 -5832 -1552 -5768
rect -1616 -5912 -1552 -5848
rect -1616 -5992 -1552 -5928
rect -204 -5272 -140 -5208
rect -204 -5352 -140 -5288
rect -204 -5432 -140 -5368
rect -204 -5512 -140 -5448
rect -204 -5592 -140 -5528
rect -204 -5672 -140 -5608
rect -204 -5752 -140 -5688
rect -204 -5832 -140 -5768
rect -204 -5912 -140 -5848
rect -204 -5992 -140 -5928
rect 1208 -5272 1272 -5208
rect 1208 -5352 1272 -5288
rect 1208 -5432 1272 -5368
rect 1208 -5512 1272 -5448
rect 1208 -5592 1272 -5528
rect 1208 -5672 1272 -5608
rect 1208 -5752 1272 -5688
rect 1208 -5832 1272 -5768
rect 1208 -5912 1272 -5848
rect 1208 -5992 1272 -5928
rect 2620 -5272 2684 -5208
rect 2620 -5352 2684 -5288
rect 2620 -5432 2684 -5368
rect 2620 -5512 2684 -5448
rect 2620 -5592 2684 -5528
rect 2620 -5672 2684 -5608
rect 2620 -5752 2684 -5688
rect 2620 -5832 2684 -5768
rect 2620 -5912 2684 -5848
rect 2620 -5992 2684 -5928
rect 4032 -5272 4096 -5208
rect 4032 -5352 4096 -5288
rect 4032 -5432 4096 -5368
rect 4032 -5512 4096 -5448
rect 4032 -5592 4096 -5528
rect 4032 -5672 4096 -5608
rect 4032 -5752 4096 -5688
rect 4032 -5832 4096 -5768
rect 4032 -5912 4096 -5848
rect 4032 -5992 4096 -5928
rect 5444 -5272 5508 -5208
rect 5444 -5352 5508 -5288
rect 5444 -5432 5508 -5368
rect 5444 -5512 5508 -5448
rect 5444 -5592 5508 -5528
rect 5444 -5672 5508 -5608
rect 5444 -5752 5508 -5688
rect 5444 -5832 5508 -5768
rect 5444 -5912 5508 -5848
rect 5444 -5992 5508 -5928
rect 6856 -5272 6920 -5208
rect 6856 -5352 6920 -5288
rect 6856 -5432 6920 -5368
rect 6856 -5512 6920 -5448
rect 6856 -5592 6920 -5528
rect 6856 -5672 6920 -5608
rect 6856 -5752 6920 -5688
rect 6856 -5832 6920 -5768
rect 6856 -5912 6920 -5848
rect 6856 -5992 6920 -5928
rect 8268 -5272 8332 -5208
rect 8268 -5352 8332 -5288
rect 8268 -5432 8332 -5368
rect 8268 -5512 8332 -5448
rect 8268 -5592 8332 -5528
rect 8268 -5672 8332 -5608
rect 8268 -5752 8332 -5688
rect 8268 -5832 8332 -5768
rect 8268 -5912 8332 -5848
rect 8268 -5992 8332 -5928
rect 9680 -5272 9744 -5208
rect 9680 -5352 9744 -5288
rect 9680 -5432 9744 -5368
rect 9680 -5512 9744 -5448
rect 9680 -5592 9744 -5528
rect 9680 -5672 9744 -5608
rect 9680 -5752 9744 -5688
rect 9680 -5832 9744 -5768
rect 9680 -5912 9744 -5848
rect 9680 -5992 9744 -5928
rect 11092 -5272 11156 -5208
rect 11092 -5352 11156 -5288
rect 11092 -5432 11156 -5368
rect 11092 -5512 11156 -5448
rect 11092 -5592 11156 -5528
rect 11092 -5672 11156 -5608
rect 11092 -5752 11156 -5688
rect 11092 -5832 11156 -5768
rect 11092 -5912 11156 -5848
rect 11092 -5992 11156 -5928
rect 12504 -5272 12568 -5208
rect 12504 -5352 12568 -5288
rect 12504 -5432 12568 -5368
rect 12504 -5512 12568 -5448
rect 12504 -5592 12568 -5528
rect 12504 -5672 12568 -5608
rect 12504 -5752 12568 -5688
rect 12504 -5832 12568 -5768
rect 12504 -5912 12568 -5848
rect 12504 -5992 12568 -5928
rect 13916 -5272 13980 -5208
rect 13916 -5352 13980 -5288
rect 13916 -5432 13980 -5368
rect 13916 -5512 13980 -5448
rect 13916 -5592 13980 -5528
rect 13916 -5672 13980 -5608
rect 13916 -5752 13980 -5688
rect 13916 -5832 13980 -5768
rect 13916 -5912 13980 -5848
rect 13916 -5992 13980 -5928
rect 15328 -5272 15392 -5208
rect 15328 -5352 15392 -5288
rect 15328 -5432 15392 -5368
rect 15328 -5512 15392 -5448
rect 15328 -5592 15392 -5528
rect 15328 -5672 15392 -5608
rect 15328 -5752 15392 -5688
rect 15328 -5832 15392 -5768
rect 15328 -5912 15392 -5848
rect 15328 -5992 15392 -5928
rect 16740 -5272 16804 -5208
rect 16740 -5352 16804 -5288
rect 16740 -5432 16804 -5368
rect 16740 -5512 16804 -5448
rect 16740 -5592 16804 -5528
rect 16740 -5672 16804 -5608
rect 16740 -5752 16804 -5688
rect 16740 -5832 16804 -5768
rect 16740 -5912 16804 -5848
rect 16740 -5992 16804 -5928
rect 18152 -5272 18216 -5208
rect 18152 -5352 18216 -5288
rect 18152 -5432 18216 -5368
rect 18152 -5512 18216 -5448
rect 18152 -5592 18216 -5528
rect 18152 -5672 18216 -5608
rect 18152 -5752 18216 -5688
rect 18152 -5832 18216 -5768
rect 18152 -5912 18216 -5848
rect 18152 -5992 18216 -5928
rect 19564 -5272 19628 -5208
rect 19564 -5352 19628 -5288
rect 19564 -5432 19628 -5368
rect 19564 -5512 19628 -5448
rect 19564 -5592 19628 -5528
rect 19564 -5672 19628 -5608
rect 19564 -5752 19628 -5688
rect 19564 -5832 19628 -5768
rect 19564 -5912 19628 -5848
rect 19564 -5992 19628 -5928
rect 20976 -5272 21040 -5208
rect 20976 -5352 21040 -5288
rect 20976 -5432 21040 -5368
rect 20976 -5512 21040 -5448
rect 20976 -5592 21040 -5528
rect 20976 -5672 21040 -5608
rect 20976 -5752 21040 -5688
rect 20976 -5832 21040 -5768
rect 20976 -5912 21040 -5848
rect 20976 -5992 21040 -5928
rect 22388 -5272 22452 -5208
rect 22388 -5352 22452 -5288
rect 22388 -5432 22452 -5368
rect 22388 -5512 22452 -5448
rect 22388 -5592 22452 -5528
rect 22388 -5672 22452 -5608
rect 22388 -5752 22452 -5688
rect 22388 -5832 22452 -5768
rect 22388 -5912 22452 -5848
rect 22388 -5992 22452 -5928
rect 23800 -5272 23864 -5208
rect 23800 -5352 23864 -5288
rect 23800 -5432 23864 -5368
rect 23800 -5512 23864 -5448
rect 23800 -5592 23864 -5528
rect 23800 -5672 23864 -5608
rect 23800 -5752 23864 -5688
rect 23800 -5832 23864 -5768
rect 23800 -5912 23864 -5848
rect 23800 -5992 23864 -5928
rect -22796 -6392 -22732 -6328
rect -22796 -6472 -22732 -6408
rect -22796 -6552 -22732 -6488
rect -22796 -6632 -22732 -6568
rect -22796 -6712 -22732 -6648
rect -22796 -6792 -22732 -6728
rect -22796 -6872 -22732 -6808
rect -22796 -6952 -22732 -6888
rect -22796 -7032 -22732 -6968
rect -22796 -7112 -22732 -7048
rect -21384 -6392 -21320 -6328
rect -21384 -6472 -21320 -6408
rect -21384 -6552 -21320 -6488
rect -21384 -6632 -21320 -6568
rect -21384 -6712 -21320 -6648
rect -21384 -6792 -21320 -6728
rect -21384 -6872 -21320 -6808
rect -21384 -6952 -21320 -6888
rect -21384 -7032 -21320 -6968
rect -21384 -7112 -21320 -7048
rect -19972 -6392 -19908 -6328
rect -19972 -6472 -19908 -6408
rect -19972 -6552 -19908 -6488
rect -19972 -6632 -19908 -6568
rect -19972 -6712 -19908 -6648
rect -19972 -6792 -19908 -6728
rect -19972 -6872 -19908 -6808
rect -19972 -6952 -19908 -6888
rect -19972 -7032 -19908 -6968
rect -19972 -7112 -19908 -7048
rect -18560 -6392 -18496 -6328
rect -18560 -6472 -18496 -6408
rect -18560 -6552 -18496 -6488
rect -18560 -6632 -18496 -6568
rect -18560 -6712 -18496 -6648
rect -18560 -6792 -18496 -6728
rect -18560 -6872 -18496 -6808
rect -18560 -6952 -18496 -6888
rect -18560 -7032 -18496 -6968
rect -18560 -7112 -18496 -7048
rect -17148 -6392 -17084 -6328
rect -17148 -6472 -17084 -6408
rect -17148 -6552 -17084 -6488
rect -17148 -6632 -17084 -6568
rect -17148 -6712 -17084 -6648
rect -17148 -6792 -17084 -6728
rect -17148 -6872 -17084 -6808
rect -17148 -6952 -17084 -6888
rect -17148 -7032 -17084 -6968
rect -17148 -7112 -17084 -7048
rect -15736 -6392 -15672 -6328
rect -15736 -6472 -15672 -6408
rect -15736 -6552 -15672 -6488
rect -15736 -6632 -15672 -6568
rect -15736 -6712 -15672 -6648
rect -15736 -6792 -15672 -6728
rect -15736 -6872 -15672 -6808
rect -15736 -6952 -15672 -6888
rect -15736 -7032 -15672 -6968
rect -15736 -7112 -15672 -7048
rect -14324 -6392 -14260 -6328
rect -14324 -6472 -14260 -6408
rect -14324 -6552 -14260 -6488
rect -14324 -6632 -14260 -6568
rect -14324 -6712 -14260 -6648
rect -14324 -6792 -14260 -6728
rect -14324 -6872 -14260 -6808
rect -14324 -6952 -14260 -6888
rect -14324 -7032 -14260 -6968
rect -14324 -7112 -14260 -7048
rect -12912 -6392 -12848 -6328
rect -12912 -6472 -12848 -6408
rect -12912 -6552 -12848 -6488
rect -12912 -6632 -12848 -6568
rect -12912 -6712 -12848 -6648
rect -12912 -6792 -12848 -6728
rect -12912 -6872 -12848 -6808
rect -12912 -6952 -12848 -6888
rect -12912 -7032 -12848 -6968
rect -12912 -7112 -12848 -7048
rect -11500 -6392 -11436 -6328
rect -11500 -6472 -11436 -6408
rect -11500 -6552 -11436 -6488
rect -11500 -6632 -11436 -6568
rect -11500 -6712 -11436 -6648
rect -11500 -6792 -11436 -6728
rect -11500 -6872 -11436 -6808
rect -11500 -6952 -11436 -6888
rect -11500 -7032 -11436 -6968
rect -11500 -7112 -11436 -7048
rect -10088 -6392 -10024 -6328
rect -10088 -6472 -10024 -6408
rect -10088 -6552 -10024 -6488
rect -10088 -6632 -10024 -6568
rect -10088 -6712 -10024 -6648
rect -10088 -6792 -10024 -6728
rect -10088 -6872 -10024 -6808
rect -10088 -6952 -10024 -6888
rect -10088 -7032 -10024 -6968
rect -10088 -7112 -10024 -7048
rect -8676 -6392 -8612 -6328
rect -8676 -6472 -8612 -6408
rect -8676 -6552 -8612 -6488
rect -8676 -6632 -8612 -6568
rect -8676 -6712 -8612 -6648
rect -8676 -6792 -8612 -6728
rect -8676 -6872 -8612 -6808
rect -8676 -6952 -8612 -6888
rect -8676 -7032 -8612 -6968
rect -8676 -7112 -8612 -7048
rect -7264 -6392 -7200 -6328
rect -7264 -6472 -7200 -6408
rect -7264 -6552 -7200 -6488
rect -7264 -6632 -7200 -6568
rect -7264 -6712 -7200 -6648
rect -7264 -6792 -7200 -6728
rect -7264 -6872 -7200 -6808
rect -7264 -6952 -7200 -6888
rect -7264 -7032 -7200 -6968
rect -7264 -7112 -7200 -7048
rect -5852 -6392 -5788 -6328
rect -5852 -6472 -5788 -6408
rect -5852 -6552 -5788 -6488
rect -5852 -6632 -5788 -6568
rect -5852 -6712 -5788 -6648
rect -5852 -6792 -5788 -6728
rect -5852 -6872 -5788 -6808
rect -5852 -6952 -5788 -6888
rect -5852 -7032 -5788 -6968
rect -5852 -7112 -5788 -7048
rect -4440 -6392 -4376 -6328
rect -4440 -6472 -4376 -6408
rect -4440 -6552 -4376 -6488
rect -4440 -6632 -4376 -6568
rect -4440 -6712 -4376 -6648
rect -4440 -6792 -4376 -6728
rect -4440 -6872 -4376 -6808
rect -4440 -6952 -4376 -6888
rect -4440 -7032 -4376 -6968
rect -4440 -7112 -4376 -7048
rect -3028 -6392 -2964 -6328
rect -3028 -6472 -2964 -6408
rect -3028 -6552 -2964 -6488
rect -3028 -6632 -2964 -6568
rect -3028 -6712 -2964 -6648
rect -3028 -6792 -2964 -6728
rect -3028 -6872 -2964 -6808
rect -3028 -6952 -2964 -6888
rect -3028 -7032 -2964 -6968
rect -3028 -7112 -2964 -7048
rect -1616 -6392 -1552 -6328
rect -1616 -6472 -1552 -6408
rect -1616 -6552 -1552 -6488
rect -1616 -6632 -1552 -6568
rect -1616 -6712 -1552 -6648
rect -1616 -6792 -1552 -6728
rect -1616 -6872 -1552 -6808
rect -1616 -6952 -1552 -6888
rect -1616 -7032 -1552 -6968
rect -1616 -7112 -1552 -7048
rect -204 -6392 -140 -6328
rect -204 -6472 -140 -6408
rect -204 -6552 -140 -6488
rect -204 -6632 -140 -6568
rect -204 -6712 -140 -6648
rect -204 -6792 -140 -6728
rect -204 -6872 -140 -6808
rect -204 -6952 -140 -6888
rect -204 -7032 -140 -6968
rect -204 -7112 -140 -7048
rect 1208 -6392 1272 -6328
rect 1208 -6472 1272 -6408
rect 1208 -6552 1272 -6488
rect 1208 -6632 1272 -6568
rect 1208 -6712 1272 -6648
rect 1208 -6792 1272 -6728
rect 1208 -6872 1272 -6808
rect 1208 -6952 1272 -6888
rect 1208 -7032 1272 -6968
rect 1208 -7112 1272 -7048
rect 2620 -6392 2684 -6328
rect 2620 -6472 2684 -6408
rect 2620 -6552 2684 -6488
rect 2620 -6632 2684 -6568
rect 2620 -6712 2684 -6648
rect 2620 -6792 2684 -6728
rect 2620 -6872 2684 -6808
rect 2620 -6952 2684 -6888
rect 2620 -7032 2684 -6968
rect 2620 -7112 2684 -7048
rect 4032 -6392 4096 -6328
rect 4032 -6472 4096 -6408
rect 4032 -6552 4096 -6488
rect 4032 -6632 4096 -6568
rect 4032 -6712 4096 -6648
rect 4032 -6792 4096 -6728
rect 4032 -6872 4096 -6808
rect 4032 -6952 4096 -6888
rect 4032 -7032 4096 -6968
rect 4032 -7112 4096 -7048
rect 5444 -6392 5508 -6328
rect 5444 -6472 5508 -6408
rect 5444 -6552 5508 -6488
rect 5444 -6632 5508 -6568
rect 5444 -6712 5508 -6648
rect 5444 -6792 5508 -6728
rect 5444 -6872 5508 -6808
rect 5444 -6952 5508 -6888
rect 5444 -7032 5508 -6968
rect 5444 -7112 5508 -7048
rect 6856 -6392 6920 -6328
rect 6856 -6472 6920 -6408
rect 6856 -6552 6920 -6488
rect 6856 -6632 6920 -6568
rect 6856 -6712 6920 -6648
rect 6856 -6792 6920 -6728
rect 6856 -6872 6920 -6808
rect 6856 -6952 6920 -6888
rect 6856 -7032 6920 -6968
rect 6856 -7112 6920 -7048
rect 8268 -6392 8332 -6328
rect 8268 -6472 8332 -6408
rect 8268 -6552 8332 -6488
rect 8268 -6632 8332 -6568
rect 8268 -6712 8332 -6648
rect 8268 -6792 8332 -6728
rect 8268 -6872 8332 -6808
rect 8268 -6952 8332 -6888
rect 8268 -7032 8332 -6968
rect 8268 -7112 8332 -7048
rect 9680 -6392 9744 -6328
rect 9680 -6472 9744 -6408
rect 9680 -6552 9744 -6488
rect 9680 -6632 9744 -6568
rect 9680 -6712 9744 -6648
rect 9680 -6792 9744 -6728
rect 9680 -6872 9744 -6808
rect 9680 -6952 9744 -6888
rect 9680 -7032 9744 -6968
rect 9680 -7112 9744 -7048
rect 11092 -6392 11156 -6328
rect 11092 -6472 11156 -6408
rect 11092 -6552 11156 -6488
rect 11092 -6632 11156 -6568
rect 11092 -6712 11156 -6648
rect 11092 -6792 11156 -6728
rect 11092 -6872 11156 -6808
rect 11092 -6952 11156 -6888
rect 11092 -7032 11156 -6968
rect 11092 -7112 11156 -7048
rect 12504 -6392 12568 -6328
rect 12504 -6472 12568 -6408
rect 12504 -6552 12568 -6488
rect 12504 -6632 12568 -6568
rect 12504 -6712 12568 -6648
rect 12504 -6792 12568 -6728
rect 12504 -6872 12568 -6808
rect 12504 -6952 12568 -6888
rect 12504 -7032 12568 -6968
rect 12504 -7112 12568 -7048
rect 13916 -6392 13980 -6328
rect 13916 -6472 13980 -6408
rect 13916 -6552 13980 -6488
rect 13916 -6632 13980 -6568
rect 13916 -6712 13980 -6648
rect 13916 -6792 13980 -6728
rect 13916 -6872 13980 -6808
rect 13916 -6952 13980 -6888
rect 13916 -7032 13980 -6968
rect 13916 -7112 13980 -7048
rect 15328 -6392 15392 -6328
rect 15328 -6472 15392 -6408
rect 15328 -6552 15392 -6488
rect 15328 -6632 15392 -6568
rect 15328 -6712 15392 -6648
rect 15328 -6792 15392 -6728
rect 15328 -6872 15392 -6808
rect 15328 -6952 15392 -6888
rect 15328 -7032 15392 -6968
rect 15328 -7112 15392 -7048
rect 16740 -6392 16804 -6328
rect 16740 -6472 16804 -6408
rect 16740 -6552 16804 -6488
rect 16740 -6632 16804 -6568
rect 16740 -6712 16804 -6648
rect 16740 -6792 16804 -6728
rect 16740 -6872 16804 -6808
rect 16740 -6952 16804 -6888
rect 16740 -7032 16804 -6968
rect 16740 -7112 16804 -7048
rect 18152 -6392 18216 -6328
rect 18152 -6472 18216 -6408
rect 18152 -6552 18216 -6488
rect 18152 -6632 18216 -6568
rect 18152 -6712 18216 -6648
rect 18152 -6792 18216 -6728
rect 18152 -6872 18216 -6808
rect 18152 -6952 18216 -6888
rect 18152 -7032 18216 -6968
rect 18152 -7112 18216 -7048
rect 19564 -6392 19628 -6328
rect 19564 -6472 19628 -6408
rect 19564 -6552 19628 -6488
rect 19564 -6632 19628 -6568
rect 19564 -6712 19628 -6648
rect 19564 -6792 19628 -6728
rect 19564 -6872 19628 -6808
rect 19564 -6952 19628 -6888
rect 19564 -7032 19628 -6968
rect 19564 -7112 19628 -7048
rect 20976 -6392 21040 -6328
rect 20976 -6472 21040 -6408
rect 20976 -6552 21040 -6488
rect 20976 -6632 21040 -6568
rect 20976 -6712 21040 -6648
rect 20976 -6792 21040 -6728
rect 20976 -6872 21040 -6808
rect 20976 -6952 21040 -6888
rect 20976 -7032 21040 -6968
rect 20976 -7112 21040 -7048
rect 22388 -6392 22452 -6328
rect 22388 -6472 22452 -6408
rect 22388 -6552 22452 -6488
rect 22388 -6632 22452 -6568
rect 22388 -6712 22452 -6648
rect 22388 -6792 22452 -6728
rect 22388 -6872 22452 -6808
rect 22388 -6952 22452 -6888
rect 22388 -7032 22452 -6968
rect 22388 -7112 22452 -7048
rect 23800 -6392 23864 -6328
rect 23800 -6472 23864 -6408
rect 23800 -6552 23864 -6488
rect 23800 -6632 23864 -6568
rect 23800 -6712 23864 -6648
rect 23800 -6792 23864 -6728
rect 23800 -6872 23864 -6808
rect 23800 -6952 23864 -6888
rect 23800 -7032 23864 -6968
rect 23800 -7112 23864 -7048
rect -22796 -7512 -22732 -7448
rect -22796 -7592 -22732 -7528
rect -22796 -7672 -22732 -7608
rect -22796 -7752 -22732 -7688
rect -22796 -7832 -22732 -7768
rect -22796 -7912 -22732 -7848
rect -22796 -7992 -22732 -7928
rect -22796 -8072 -22732 -8008
rect -22796 -8152 -22732 -8088
rect -22796 -8232 -22732 -8168
rect -21384 -7512 -21320 -7448
rect -21384 -7592 -21320 -7528
rect -21384 -7672 -21320 -7608
rect -21384 -7752 -21320 -7688
rect -21384 -7832 -21320 -7768
rect -21384 -7912 -21320 -7848
rect -21384 -7992 -21320 -7928
rect -21384 -8072 -21320 -8008
rect -21384 -8152 -21320 -8088
rect -21384 -8232 -21320 -8168
rect -19972 -7512 -19908 -7448
rect -19972 -7592 -19908 -7528
rect -19972 -7672 -19908 -7608
rect -19972 -7752 -19908 -7688
rect -19972 -7832 -19908 -7768
rect -19972 -7912 -19908 -7848
rect -19972 -7992 -19908 -7928
rect -19972 -8072 -19908 -8008
rect -19972 -8152 -19908 -8088
rect -19972 -8232 -19908 -8168
rect -18560 -7512 -18496 -7448
rect -18560 -7592 -18496 -7528
rect -18560 -7672 -18496 -7608
rect -18560 -7752 -18496 -7688
rect -18560 -7832 -18496 -7768
rect -18560 -7912 -18496 -7848
rect -18560 -7992 -18496 -7928
rect -18560 -8072 -18496 -8008
rect -18560 -8152 -18496 -8088
rect -18560 -8232 -18496 -8168
rect -17148 -7512 -17084 -7448
rect -17148 -7592 -17084 -7528
rect -17148 -7672 -17084 -7608
rect -17148 -7752 -17084 -7688
rect -17148 -7832 -17084 -7768
rect -17148 -7912 -17084 -7848
rect -17148 -7992 -17084 -7928
rect -17148 -8072 -17084 -8008
rect -17148 -8152 -17084 -8088
rect -17148 -8232 -17084 -8168
rect -15736 -7512 -15672 -7448
rect -15736 -7592 -15672 -7528
rect -15736 -7672 -15672 -7608
rect -15736 -7752 -15672 -7688
rect -15736 -7832 -15672 -7768
rect -15736 -7912 -15672 -7848
rect -15736 -7992 -15672 -7928
rect -15736 -8072 -15672 -8008
rect -15736 -8152 -15672 -8088
rect -15736 -8232 -15672 -8168
rect -14324 -7512 -14260 -7448
rect -14324 -7592 -14260 -7528
rect -14324 -7672 -14260 -7608
rect -14324 -7752 -14260 -7688
rect -14324 -7832 -14260 -7768
rect -14324 -7912 -14260 -7848
rect -14324 -7992 -14260 -7928
rect -14324 -8072 -14260 -8008
rect -14324 -8152 -14260 -8088
rect -14324 -8232 -14260 -8168
rect -12912 -7512 -12848 -7448
rect -12912 -7592 -12848 -7528
rect -12912 -7672 -12848 -7608
rect -12912 -7752 -12848 -7688
rect -12912 -7832 -12848 -7768
rect -12912 -7912 -12848 -7848
rect -12912 -7992 -12848 -7928
rect -12912 -8072 -12848 -8008
rect -12912 -8152 -12848 -8088
rect -12912 -8232 -12848 -8168
rect -11500 -7512 -11436 -7448
rect -11500 -7592 -11436 -7528
rect -11500 -7672 -11436 -7608
rect -11500 -7752 -11436 -7688
rect -11500 -7832 -11436 -7768
rect -11500 -7912 -11436 -7848
rect -11500 -7992 -11436 -7928
rect -11500 -8072 -11436 -8008
rect -11500 -8152 -11436 -8088
rect -11500 -8232 -11436 -8168
rect -10088 -7512 -10024 -7448
rect -10088 -7592 -10024 -7528
rect -10088 -7672 -10024 -7608
rect -10088 -7752 -10024 -7688
rect -10088 -7832 -10024 -7768
rect -10088 -7912 -10024 -7848
rect -10088 -7992 -10024 -7928
rect -10088 -8072 -10024 -8008
rect -10088 -8152 -10024 -8088
rect -10088 -8232 -10024 -8168
rect -8676 -7512 -8612 -7448
rect -8676 -7592 -8612 -7528
rect -8676 -7672 -8612 -7608
rect -8676 -7752 -8612 -7688
rect -8676 -7832 -8612 -7768
rect -8676 -7912 -8612 -7848
rect -8676 -7992 -8612 -7928
rect -8676 -8072 -8612 -8008
rect -8676 -8152 -8612 -8088
rect -8676 -8232 -8612 -8168
rect -7264 -7512 -7200 -7448
rect -7264 -7592 -7200 -7528
rect -7264 -7672 -7200 -7608
rect -7264 -7752 -7200 -7688
rect -7264 -7832 -7200 -7768
rect -7264 -7912 -7200 -7848
rect -7264 -7992 -7200 -7928
rect -7264 -8072 -7200 -8008
rect -7264 -8152 -7200 -8088
rect -7264 -8232 -7200 -8168
rect -5852 -7512 -5788 -7448
rect -5852 -7592 -5788 -7528
rect -5852 -7672 -5788 -7608
rect -5852 -7752 -5788 -7688
rect -5852 -7832 -5788 -7768
rect -5852 -7912 -5788 -7848
rect -5852 -7992 -5788 -7928
rect -5852 -8072 -5788 -8008
rect -5852 -8152 -5788 -8088
rect -5852 -8232 -5788 -8168
rect -4440 -7512 -4376 -7448
rect -4440 -7592 -4376 -7528
rect -4440 -7672 -4376 -7608
rect -4440 -7752 -4376 -7688
rect -4440 -7832 -4376 -7768
rect -4440 -7912 -4376 -7848
rect -4440 -7992 -4376 -7928
rect -4440 -8072 -4376 -8008
rect -4440 -8152 -4376 -8088
rect -4440 -8232 -4376 -8168
rect -3028 -7512 -2964 -7448
rect -3028 -7592 -2964 -7528
rect -3028 -7672 -2964 -7608
rect -3028 -7752 -2964 -7688
rect -3028 -7832 -2964 -7768
rect -3028 -7912 -2964 -7848
rect -3028 -7992 -2964 -7928
rect -3028 -8072 -2964 -8008
rect -3028 -8152 -2964 -8088
rect -3028 -8232 -2964 -8168
rect -1616 -7512 -1552 -7448
rect -1616 -7592 -1552 -7528
rect -1616 -7672 -1552 -7608
rect -1616 -7752 -1552 -7688
rect -1616 -7832 -1552 -7768
rect -1616 -7912 -1552 -7848
rect -1616 -7992 -1552 -7928
rect -1616 -8072 -1552 -8008
rect -1616 -8152 -1552 -8088
rect -1616 -8232 -1552 -8168
rect -204 -7512 -140 -7448
rect -204 -7592 -140 -7528
rect -204 -7672 -140 -7608
rect -204 -7752 -140 -7688
rect -204 -7832 -140 -7768
rect -204 -7912 -140 -7848
rect -204 -7992 -140 -7928
rect -204 -8072 -140 -8008
rect -204 -8152 -140 -8088
rect -204 -8232 -140 -8168
rect 1208 -7512 1272 -7448
rect 1208 -7592 1272 -7528
rect 1208 -7672 1272 -7608
rect 1208 -7752 1272 -7688
rect 1208 -7832 1272 -7768
rect 1208 -7912 1272 -7848
rect 1208 -7992 1272 -7928
rect 1208 -8072 1272 -8008
rect 1208 -8152 1272 -8088
rect 1208 -8232 1272 -8168
rect 2620 -7512 2684 -7448
rect 2620 -7592 2684 -7528
rect 2620 -7672 2684 -7608
rect 2620 -7752 2684 -7688
rect 2620 -7832 2684 -7768
rect 2620 -7912 2684 -7848
rect 2620 -7992 2684 -7928
rect 2620 -8072 2684 -8008
rect 2620 -8152 2684 -8088
rect 2620 -8232 2684 -8168
rect 4032 -7512 4096 -7448
rect 4032 -7592 4096 -7528
rect 4032 -7672 4096 -7608
rect 4032 -7752 4096 -7688
rect 4032 -7832 4096 -7768
rect 4032 -7912 4096 -7848
rect 4032 -7992 4096 -7928
rect 4032 -8072 4096 -8008
rect 4032 -8152 4096 -8088
rect 4032 -8232 4096 -8168
rect 5444 -7512 5508 -7448
rect 5444 -7592 5508 -7528
rect 5444 -7672 5508 -7608
rect 5444 -7752 5508 -7688
rect 5444 -7832 5508 -7768
rect 5444 -7912 5508 -7848
rect 5444 -7992 5508 -7928
rect 5444 -8072 5508 -8008
rect 5444 -8152 5508 -8088
rect 5444 -8232 5508 -8168
rect 6856 -7512 6920 -7448
rect 6856 -7592 6920 -7528
rect 6856 -7672 6920 -7608
rect 6856 -7752 6920 -7688
rect 6856 -7832 6920 -7768
rect 6856 -7912 6920 -7848
rect 6856 -7992 6920 -7928
rect 6856 -8072 6920 -8008
rect 6856 -8152 6920 -8088
rect 6856 -8232 6920 -8168
rect 8268 -7512 8332 -7448
rect 8268 -7592 8332 -7528
rect 8268 -7672 8332 -7608
rect 8268 -7752 8332 -7688
rect 8268 -7832 8332 -7768
rect 8268 -7912 8332 -7848
rect 8268 -7992 8332 -7928
rect 8268 -8072 8332 -8008
rect 8268 -8152 8332 -8088
rect 8268 -8232 8332 -8168
rect 9680 -7512 9744 -7448
rect 9680 -7592 9744 -7528
rect 9680 -7672 9744 -7608
rect 9680 -7752 9744 -7688
rect 9680 -7832 9744 -7768
rect 9680 -7912 9744 -7848
rect 9680 -7992 9744 -7928
rect 9680 -8072 9744 -8008
rect 9680 -8152 9744 -8088
rect 9680 -8232 9744 -8168
rect 11092 -7512 11156 -7448
rect 11092 -7592 11156 -7528
rect 11092 -7672 11156 -7608
rect 11092 -7752 11156 -7688
rect 11092 -7832 11156 -7768
rect 11092 -7912 11156 -7848
rect 11092 -7992 11156 -7928
rect 11092 -8072 11156 -8008
rect 11092 -8152 11156 -8088
rect 11092 -8232 11156 -8168
rect 12504 -7512 12568 -7448
rect 12504 -7592 12568 -7528
rect 12504 -7672 12568 -7608
rect 12504 -7752 12568 -7688
rect 12504 -7832 12568 -7768
rect 12504 -7912 12568 -7848
rect 12504 -7992 12568 -7928
rect 12504 -8072 12568 -8008
rect 12504 -8152 12568 -8088
rect 12504 -8232 12568 -8168
rect 13916 -7512 13980 -7448
rect 13916 -7592 13980 -7528
rect 13916 -7672 13980 -7608
rect 13916 -7752 13980 -7688
rect 13916 -7832 13980 -7768
rect 13916 -7912 13980 -7848
rect 13916 -7992 13980 -7928
rect 13916 -8072 13980 -8008
rect 13916 -8152 13980 -8088
rect 13916 -8232 13980 -8168
rect 15328 -7512 15392 -7448
rect 15328 -7592 15392 -7528
rect 15328 -7672 15392 -7608
rect 15328 -7752 15392 -7688
rect 15328 -7832 15392 -7768
rect 15328 -7912 15392 -7848
rect 15328 -7992 15392 -7928
rect 15328 -8072 15392 -8008
rect 15328 -8152 15392 -8088
rect 15328 -8232 15392 -8168
rect 16740 -7512 16804 -7448
rect 16740 -7592 16804 -7528
rect 16740 -7672 16804 -7608
rect 16740 -7752 16804 -7688
rect 16740 -7832 16804 -7768
rect 16740 -7912 16804 -7848
rect 16740 -7992 16804 -7928
rect 16740 -8072 16804 -8008
rect 16740 -8152 16804 -8088
rect 16740 -8232 16804 -8168
rect 18152 -7512 18216 -7448
rect 18152 -7592 18216 -7528
rect 18152 -7672 18216 -7608
rect 18152 -7752 18216 -7688
rect 18152 -7832 18216 -7768
rect 18152 -7912 18216 -7848
rect 18152 -7992 18216 -7928
rect 18152 -8072 18216 -8008
rect 18152 -8152 18216 -8088
rect 18152 -8232 18216 -8168
rect 19564 -7512 19628 -7448
rect 19564 -7592 19628 -7528
rect 19564 -7672 19628 -7608
rect 19564 -7752 19628 -7688
rect 19564 -7832 19628 -7768
rect 19564 -7912 19628 -7848
rect 19564 -7992 19628 -7928
rect 19564 -8072 19628 -8008
rect 19564 -8152 19628 -8088
rect 19564 -8232 19628 -8168
rect 20976 -7512 21040 -7448
rect 20976 -7592 21040 -7528
rect 20976 -7672 21040 -7608
rect 20976 -7752 21040 -7688
rect 20976 -7832 21040 -7768
rect 20976 -7912 21040 -7848
rect 20976 -7992 21040 -7928
rect 20976 -8072 21040 -8008
rect 20976 -8152 21040 -8088
rect 20976 -8232 21040 -8168
rect 22388 -7512 22452 -7448
rect 22388 -7592 22452 -7528
rect 22388 -7672 22452 -7608
rect 22388 -7752 22452 -7688
rect 22388 -7832 22452 -7768
rect 22388 -7912 22452 -7848
rect 22388 -7992 22452 -7928
rect 22388 -8072 22452 -8008
rect 22388 -8152 22452 -8088
rect 22388 -8232 22452 -8168
rect 23800 -7512 23864 -7448
rect 23800 -7592 23864 -7528
rect 23800 -7672 23864 -7608
rect 23800 -7752 23864 -7688
rect 23800 -7832 23864 -7768
rect 23800 -7912 23864 -7848
rect 23800 -7992 23864 -7928
rect 23800 -8072 23864 -8008
rect 23800 -8152 23864 -8088
rect 23800 -8232 23864 -8168
rect -22796 -8632 -22732 -8568
rect -22796 -8712 -22732 -8648
rect -22796 -8792 -22732 -8728
rect -22796 -8872 -22732 -8808
rect -22796 -8952 -22732 -8888
rect -22796 -9032 -22732 -8968
rect -22796 -9112 -22732 -9048
rect -22796 -9192 -22732 -9128
rect -22796 -9272 -22732 -9208
rect -22796 -9352 -22732 -9288
rect -21384 -8632 -21320 -8568
rect -21384 -8712 -21320 -8648
rect -21384 -8792 -21320 -8728
rect -21384 -8872 -21320 -8808
rect -21384 -8952 -21320 -8888
rect -21384 -9032 -21320 -8968
rect -21384 -9112 -21320 -9048
rect -21384 -9192 -21320 -9128
rect -21384 -9272 -21320 -9208
rect -21384 -9352 -21320 -9288
rect -19972 -8632 -19908 -8568
rect -19972 -8712 -19908 -8648
rect -19972 -8792 -19908 -8728
rect -19972 -8872 -19908 -8808
rect -19972 -8952 -19908 -8888
rect -19972 -9032 -19908 -8968
rect -19972 -9112 -19908 -9048
rect -19972 -9192 -19908 -9128
rect -19972 -9272 -19908 -9208
rect -19972 -9352 -19908 -9288
rect -18560 -8632 -18496 -8568
rect -18560 -8712 -18496 -8648
rect -18560 -8792 -18496 -8728
rect -18560 -8872 -18496 -8808
rect -18560 -8952 -18496 -8888
rect -18560 -9032 -18496 -8968
rect -18560 -9112 -18496 -9048
rect -18560 -9192 -18496 -9128
rect -18560 -9272 -18496 -9208
rect -18560 -9352 -18496 -9288
rect -17148 -8632 -17084 -8568
rect -17148 -8712 -17084 -8648
rect -17148 -8792 -17084 -8728
rect -17148 -8872 -17084 -8808
rect -17148 -8952 -17084 -8888
rect -17148 -9032 -17084 -8968
rect -17148 -9112 -17084 -9048
rect -17148 -9192 -17084 -9128
rect -17148 -9272 -17084 -9208
rect -17148 -9352 -17084 -9288
rect -15736 -8632 -15672 -8568
rect -15736 -8712 -15672 -8648
rect -15736 -8792 -15672 -8728
rect -15736 -8872 -15672 -8808
rect -15736 -8952 -15672 -8888
rect -15736 -9032 -15672 -8968
rect -15736 -9112 -15672 -9048
rect -15736 -9192 -15672 -9128
rect -15736 -9272 -15672 -9208
rect -15736 -9352 -15672 -9288
rect -14324 -8632 -14260 -8568
rect -14324 -8712 -14260 -8648
rect -14324 -8792 -14260 -8728
rect -14324 -8872 -14260 -8808
rect -14324 -8952 -14260 -8888
rect -14324 -9032 -14260 -8968
rect -14324 -9112 -14260 -9048
rect -14324 -9192 -14260 -9128
rect -14324 -9272 -14260 -9208
rect -14324 -9352 -14260 -9288
rect -12912 -8632 -12848 -8568
rect -12912 -8712 -12848 -8648
rect -12912 -8792 -12848 -8728
rect -12912 -8872 -12848 -8808
rect -12912 -8952 -12848 -8888
rect -12912 -9032 -12848 -8968
rect -12912 -9112 -12848 -9048
rect -12912 -9192 -12848 -9128
rect -12912 -9272 -12848 -9208
rect -12912 -9352 -12848 -9288
rect -11500 -8632 -11436 -8568
rect -11500 -8712 -11436 -8648
rect -11500 -8792 -11436 -8728
rect -11500 -8872 -11436 -8808
rect -11500 -8952 -11436 -8888
rect -11500 -9032 -11436 -8968
rect -11500 -9112 -11436 -9048
rect -11500 -9192 -11436 -9128
rect -11500 -9272 -11436 -9208
rect -11500 -9352 -11436 -9288
rect -10088 -8632 -10024 -8568
rect -10088 -8712 -10024 -8648
rect -10088 -8792 -10024 -8728
rect -10088 -8872 -10024 -8808
rect -10088 -8952 -10024 -8888
rect -10088 -9032 -10024 -8968
rect -10088 -9112 -10024 -9048
rect -10088 -9192 -10024 -9128
rect -10088 -9272 -10024 -9208
rect -10088 -9352 -10024 -9288
rect -8676 -8632 -8612 -8568
rect -8676 -8712 -8612 -8648
rect -8676 -8792 -8612 -8728
rect -8676 -8872 -8612 -8808
rect -8676 -8952 -8612 -8888
rect -8676 -9032 -8612 -8968
rect -8676 -9112 -8612 -9048
rect -8676 -9192 -8612 -9128
rect -8676 -9272 -8612 -9208
rect -8676 -9352 -8612 -9288
rect -7264 -8632 -7200 -8568
rect -7264 -8712 -7200 -8648
rect -7264 -8792 -7200 -8728
rect -7264 -8872 -7200 -8808
rect -7264 -8952 -7200 -8888
rect -7264 -9032 -7200 -8968
rect -7264 -9112 -7200 -9048
rect -7264 -9192 -7200 -9128
rect -7264 -9272 -7200 -9208
rect -7264 -9352 -7200 -9288
rect -5852 -8632 -5788 -8568
rect -5852 -8712 -5788 -8648
rect -5852 -8792 -5788 -8728
rect -5852 -8872 -5788 -8808
rect -5852 -8952 -5788 -8888
rect -5852 -9032 -5788 -8968
rect -5852 -9112 -5788 -9048
rect -5852 -9192 -5788 -9128
rect -5852 -9272 -5788 -9208
rect -5852 -9352 -5788 -9288
rect -4440 -8632 -4376 -8568
rect -4440 -8712 -4376 -8648
rect -4440 -8792 -4376 -8728
rect -4440 -8872 -4376 -8808
rect -4440 -8952 -4376 -8888
rect -4440 -9032 -4376 -8968
rect -4440 -9112 -4376 -9048
rect -4440 -9192 -4376 -9128
rect -4440 -9272 -4376 -9208
rect -4440 -9352 -4376 -9288
rect -3028 -8632 -2964 -8568
rect -3028 -8712 -2964 -8648
rect -3028 -8792 -2964 -8728
rect -3028 -8872 -2964 -8808
rect -3028 -8952 -2964 -8888
rect -3028 -9032 -2964 -8968
rect -3028 -9112 -2964 -9048
rect -3028 -9192 -2964 -9128
rect -3028 -9272 -2964 -9208
rect -3028 -9352 -2964 -9288
rect -1616 -8632 -1552 -8568
rect -1616 -8712 -1552 -8648
rect -1616 -8792 -1552 -8728
rect -1616 -8872 -1552 -8808
rect -1616 -8952 -1552 -8888
rect -1616 -9032 -1552 -8968
rect -1616 -9112 -1552 -9048
rect -1616 -9192 -1552 -9128
rect -1616 -9272 -1552 -9208
rect -1616 -9352 -1552 -9288
rect -204 -8632 -140 -8568
rect -204 -8712 -140 -8648
rect -204 -8792 -140 -8728
rect -204 -8872 -140 -8808
rect -204 -8952 -140 -8888
rect -204 -9032 -140 -8968
rect -204 -9112 -140 -9048
rect -204 -9192 -140 -9128
rect -204 -9272 -140 -9208
rect -204 -9352 -140 -9288
rect 1208 -8632 1272 -8568
rect 1208 -8712 1272 -8648
rect 1208 -8792 1272 -8728
rect 1208 -8872 1272 -8808
rect 1208 -8952 1272 -8888
rect 1208 -9032 1272 -8968
rect 1208 -9112 1272 -9048
rect 1208 -9192 1272 -9128
rect 1208 -9272 1272 -9208
rect 1208 -9352 1272 -9288
rect 2620 -8632 2684 -8568
rect 2620 -8712 2684 -8648
rect 2620 -8792 2684 -8728
rect 2620 -8872 2684 -8808
rect 2620 -8952 2684 -8888
rect 2620 -9032 2684 -8968
rect 2620 -9112 2684 -9048
rect 2620 -9192 2684 -9128
rect 2620 -9272 2684 -9208
rect 2620 -9352 2684 -9288
rect 4032 -8632 4096 -8568
rect 4032 -8712 4096 -8648
rect 4032 -8792 4096 -8728
rect 4032 -8872 4096 -8808
rect 4032 -8952 4096 -8888
rect 4032 -9032 4096 -8968
rect 4032 -9112 4096 -9048
rect 4032 -9192 4096 -9128
rect 4032 -9272 4096 -9208
rect 4032 -9352 4096 -9288
rect 5444 -8632 5508 -8568
rect 5444 -8712 5508 -8648
rect 5444 -8792 5508 -8728
rect 5444 -8872 5508 -8808
rect 5444 -8952 5508 -8888
rect 5444 -9032 5508 -8968
rect 5444 -9112 5508 -9048
rect 5444 -9192 5508 -9128
rect 5444 -9272 5508 -9208
rect 5444 -9352 5508 -9288
rect 6856 -8632 6920 -8568
rect 6856 -8712 6920 -8648
rect 6856 -8792 6920 -8728
rect 6856 -8872 6920 -8808
rect 6856 -8952 6920 -8888
rect 6856 -9032 6920 -8968
rect 6856 -9112 6920 -9048
rect 6856 -9192 6920 -9128
rect 6856 -9272 6920 -9208
rect 6856 -9352 6920 -9288
rect 8268 -8632 8332 -8568
rect 8268 -8712 8332 -8648
rect 8268 -8792 8332 -8728
rect 8268 -8872 8332 -8808
rect 8268 -8952 8332 -8888
rect 8268 -9032 8332 -8968
rect 8268 -9112 8332 -9048
rect 8268 -9192 8332 -9128
rect 8268 -9272 8332 -9208
rect 8268 -9352 8332 -9288
rect 9680 -8632 9744 -8568
rect 9680 -8712 9744 -8648
rect 9680 -8792 9744 -8728
rect 9680 -8872 9744 -8808
rect 9680 -8952 9744 -8888
rect 9680 -9032 9744 -8968
rect 9680 -9112 9744 -9048
rect 9680 -9192 9744 -9128
rect 9680 -9272 9744 -9208
rect 9680 -9352 9744 -9288
rect 11092 -8632 11156 -8568
rect 11092 -8712 11156 -8648
rect 11092 -8792 11156 -8728
rect 11092 -8872 11156 -8808
rect 11092 -8952 11156 -8888
rect 11092 -9032 11156 -8968
rect 11092 -9112 11156 -9048
rect 11092 -9192 11156 -9128
rect 11092 -9272 11156 -9208
rect 11092 -9352 11156 -9288
rect 12504 -8632 12568 -8568
rect 12504 -8712 12568 -8648
rect 12504 -8792 12568 -8728
rect 12504 -8872 12568 -8808
rect 12504 -8952 12568 -8888
rect 12504 -9032 12568 -8968
rect 12504 -9112 12568 -9048
rect 12504 -9192 12568 -9128
rect 12504 -9272 12568 -9208
rect 12504 -9352 12568 -9288
rect 13916 -8632 13980 -8568
rect 13916 -8712 13980 -8648
rect 13916 -8792 13980 -8728
rect 13916 -8872 13980 -8808
rect 13916 -8952 13980 -8888
rect 13916 -9032 13980 -8968
rect 13916 -9112 13980 -9048
rect 13916 -9192 13980 -9128
rect 13916 -9272 13980 -9208
rect 13916 -9352 13980 -9288
rect 15328 -8632 15392 -8568
rect 15328 -8712 15392 -8648
rect 15328 -8792 15392 -8728
rect 15328 -8872 15392 -8808
rect 15328 -8952 15392 -8888
rect 15328 -9032 15392 -8968
rect 15328 -9112 15392 -9048
rect 15328 -9192 15392 -9128
rect 15328 -9272 15392 -9208
rect 15328 -9352 15392 -9288
rect 16740 -8632 16804 -8568
rect 16740 -8712 16804 -8648
rect 16740 -8792 16804 -8728
rect 16740 -8872 16804 -8808
rect 16740 -8952 16804 -8888
rect 16740 -9032 16804 -8968
rect 16740 -9112 16804 -9048
rect 16740 -9192 16804 -9128
rect 16740 -9272 16804 -9208
rect 16740 -9352 16804 -9288
rect 18152 -8632 18216 -8568
rect 18152 -8712 18216 -8648
rect 18152 -8792 18216 -8728
rect 18152 -8872 18216 -8808
rect 18152 -8952 18216 -8888
rect 18152 -9032 18216 -8968
rect 18152 -9112 18216 -9048
rect 18152 -9192 18216 -9128
rect 18152 -9272 18216 -9208
rect 18152 -9352 18216 -9288
rect 19564 -8632 19628 -8568
rect 19564 -8712 19628 -8648
rect 19564 -8792 19628 -8728
rect 19564 -8872 19628 -8808
rect 19564 -8952 19628 -8888
rect 19564 -9032 19628 -8968
rect 19564 -9112 19628 -9048
rect 19564 -9192 19628 -9128
rect 19564 -9272 19628 -9208
rect 19564 -9352 19628 -9288
rect 20976 -8632 21040 -8568
rect 20976 -8712 21040 -8648
rect 20976 -8792 21040 -8728
rect 20976 -8872 21040 -8808
rect 20976 -8952 21040 -8888
rect 20976 -9032 21040 -8968
rect 20976 -9112 21040 -9048
rect 20976 -9192 21040 -9128
rect 20976 -9272 21040 -9208
rect 20976 -9352 21040 -9288
rect 22388 -8632 22452 -8568
rect 22388 -8712 22452 -8648
rect 22388 -8792 22452 -8728
rect 22388 -8872 22452 -8808
rect 22388 -8952 22452 -8888
rect 22388 -9032 22452 -8968
rect 22388 -9112 22452 -9048
rect 22388 -9192 22452 -9128
rect 22388 -9272 22452 -9208
rect 22388 -9352 22452 -9288
rect 23800 -8632 23864 -8568
rect 23800 -8712 23864 -8648
rect 23800 -8792 23864 -8728
rect 23800 -8872 23864 -8808
rect 23800 -8952 23864 -8888
rect 23800 -9032 23864 -8968
rect 23800 -9112 23864 -9048
rect 23800 -9192 23864 -9128
rect 23800 -9272 23864 -9208
rect 23800 -9352 23864 -9288
rect -22796 -9752 -22732 -9688
rect -22796 -9832 -22732 -9768
rect -22796 -9912 -22732 -9848
rect -22796 -9992 -22732 -9928
rect -22796 -10072 -22732 -10008
rect -22796 -10152 -22732 -10088
rect -22796 -10232 -22732 -10168
rect -22796 -10312 -22732 -10248
rect -22796 -10392 -22732 -10328
rect -22796 -10472 -22732 -10408
rect -21384 -9752 -21320 -9688
rect -21384 -9832 -21320 -9768
rect -21384 -9912 -21320 -9848
rect -21384 -9992 -21320 -9928
rect -21384 -10072 -21320 -10008
rect -21384 -10152 -21320 -10088
rect -21384 -10232 -21320 -10168
rect -21384 -10312 -21320 -10248
rect -21384 -10392 -21320 -10328
rect -21384 -10472 -21320 -10408
rect -19972 -9752 -19908 -9688
rect -19972 -9832 -19908 -9768
rect -19972 -9912 -19908 -9848
rect -19972 -9992 -19908 -9928
rect -19972 -10072 -19908 -10008
rect -19972 -10152 -19908 -10088
rect -19972 -10232 -19908 -10168
rect -19972 -10312 -19908 -10248
rect -19972 -10392 -19908 -10328
rect -19972 -10472 -19908 -10408
rect -18560 -9752 -18496 -9688
rect -18560 -9832 -18496 -9768
rect -18560 -9912 -18496 -9848
rect -18560 -9992 -18496 -9928
rect -18560 -10072 -18496 -10008
rect -18560 -10152 -18496 -10088
rect -18560 -10232 -18496 -10168
rect -18560 -10312 -18496 -10248
rect -18560 -10392 -18496 -10328
rect -18560 -10472 -18496 -10408
rect -17148 -9752 -17084 -9688
rect -17148 -9832 -17084 -9768
rect -17148 -9912 -17084 -9848
rect -17148 -9992 -17084 -9928
rect -17148 -10072 -17084 -10008
rect -17148 -10152 -17084 -10088
rect -17148 -10232 -17084 -10168
rect -17148 -10312 -17084 -10248
rect -17148 -10392 -17084 -10328
rect -17148 -10472 -17084 -10408
rect -15736 -9752 -15672 -9688
rect -15736 -9832 -15672 -9768
rect -15736 -9912 -15672 -9848
rect -15736 -9992 -15672 -9928
rect -15736 -10072 -15672 -10008
rect -15736 -10152 -15672 -10088
rect -15736 -10232 -15672 -10168
rect -15736 -10312 -15672 -10248
rect -15736 -10392 -15672 -10328
rect -15736 -10472 -15672 -10408
rect -14324 -9752 -14260 -9688
rect -14324 -9832 -14260 -9768
rect -14324 -9912 -14260 -9848
rect -14324 -9992 -14260 -9928
rect -14324 -10072 -14260 -10008
rect -14324 -10152 -14260 -10088
rect -14324 -10232 -14260 -10168
rect -14324 -10312 -14260 -10248
rect -14324 -10392 -14260 -10328
rect -14324 -10472 -14260 -10408
rect -12912 -9752 -12848 -9688
rect -12912 -9832 -12848 -9768
rect -12912 -9912 -12848 -9848
rect -12912 -9992 -12848 -9928
rect -12912 -10072 -12848 -10008
rect -12912 -10152 -12848 -10088
rect -12912 -10232 -12848 -10168
rect -12912 -10312 -12848 -10248
rect -12912 -10392 -12848 -10328
rect -12912 -10472 -12848 -10408
rect -11500 -9752 -11436 -9688
rect -11500 -9832 -11436 -9768
rect -11500 -9912 -11436 -9848
rect -11500 -9992 -11436 -9928
rect -11500 -10072 -11436 -10008
rect -11500 -10152 -11436 -10088
rect -11500 -10232 -11436 -10168
rect -11500 -10312 -11436 -10248
rect -11500 -10392 -11436 -10328
rect -11500 -10472 -11436 -10408
rect -10088 -9752 -10024 -9688
rect -10088 -9832 -10024 -9768
rect -10088 -9912 -10024 -9848
rect -10088 -9992 -10024 -9928
rect -10088 -10072 -10024 -10008
rect -10088 -10152 -10024 -10088
rect -10088 -10232 -10024 -10168
rect -10088 -10312 -10024 -10248
rect -10088 -10392 -10024 -10328
rect -10088 -10472 -10024 -10408
rect -8676 -9752 -8612 -9688
rect -8676 -9832 -8612 -9768
rect -8676 -9912 -8612 -9848
rect -8676 -9992 -8612 -9928
rect -8676 -10072 -8612 -10008
rect -8676 -10152 -8612 -10088
rect -8676 -10232 -8612 -10168
rect -8676 -10312 -8612 -10248
rect -8676 -10392 -8612 -10328
rect -8676 -10472 -8612 -10408
rect -7264 -9752 -7200 -9688
rect -7264 -9832 -7200 -9768
rect -7264 -9912 -7200 -9848
rect -7264 -9992 -7200 -9928
rect -7264 -10072 -7200 -10008
rect -7264 -10152 -7200 -10088
rect -7264 -10232 -7200 -10168
rect -7264 -10312 -7200 -10248
rect -7264 -10392 -7200 -10328
rect -7264 -10472 -7200 -10408
rect -5852 -9752 -5788 -9688
rect -5852 -9832 -5788 -9768
rect -5852 -9912 -5788 -9848
rect -5852 -9992 -5788 -9928
rect -5852 -10072 -5788 -10008
rect -5852 -10152 -5788 -10088
rect -5852 -10232 -5788 -10168
rect -5852 -10312 -5788 -10248
rect -5852 -10392 -5788 -10328
rect -5852 -10472 -5788 -10408
rect -4440 -9752 -4376 -9688
rect -4440 -9832 -4376 -9768
rect -4440 -9912 -4376 -9848
rect -4440 -9992 -4376 -9928
rect -4440 -10072 -4376 -10008
rect -4440 -10152 -4376 -10088
rect -4440 -10232 -4376 -10168
rect -4440 -10312 -4376 -10248
rect -4440 -10392 -4376 -10328
rect -4440 -10472 -4376 -10408
rect -3028 -9752 -2964 -9688
rect -3028 -9832 -2964 -9768
rect -3028 -9912 -2964 -9848
rect -3028 -9992 -2964 -9928
rect -3028 -10072 -2964 -10008
rect -3028 -10152 -2964 -10088
rect -3028 -10232 -2964 -10168
rect -3028 -10312 -2964 -10248
rect -3028 -10392 -2964 -10328
rect -3028 -10472 -2964 -10408
rect -1616 -9752 -1552 -9688
rect -1616 -9832 -1552 -9768
rect -1616 -9912 -1552 -9848
rect -1616 -9992 -1552 -9928
rect -1616 -10072 -1552 -10008
rect -1616 -10152 -1552 -10088
rect -1616 -10232 -1552 -10168
rect -1616 -10312 -1552 -10248
rect -1616 -10392 -1552 -10328
rect -1616 -10472 -1552 -10408
rect -204 -9752 -140 -9688
rect -204 -9832 -140 -9768
rect -204 -9912 -140 -9848
rect -204 -9992 -140 -9928
rect -204 -10072 -140 -10008
rect -204 -10152 -140 -10088
rect -204 -10232 -140 -10168
rect -204 -10312 -140 -10248
rect -204 -10392 -140 -10328
rect -204 -10472 -140 -10408
rect 1208 -9752 1272 -9688
rect 1208 -9832 1272 -9768
rect 1208 -9912 1272 -9848
rect 1208 -9992 1272 -9928
rect 1208 -10072 1272 -10008
rect 1208 -10152 1272 -10088
rect 1208 -10232 1272 -10168
rect 1208 -10312 1272 -10248
rect 1208 -10392 1272 -10328
rect 1208 -10472 1272 -10408
rect 2620 -9752 2684 -9688
rect 2620 -9832 2684 -9768
rect 2620 -9912 2684 -9848
rect 2620 -9992 2684 -9928
rect 2620 -10072 2684 -10008
rect 2620 -10152 2684 -10088
rect 2620 -10232 2684 -10168
rect 2620 -10312 2684 -10248
rect 2620 -10392 2684 -10328
rect 2620 -10472 2684 -10408
rect 4032 -9752 4096 -9688
rect 4032 -9832 4096 -9768
rect 4032 -9912 4096 -9848
rect 4032 -9992 4096 -9928
rect 4032 -10072 4096 -10008
rect 4032 -10152 4096 -10088
rect 4032 -10232 4096 -10168
rect 4032 -10312 4096 -10248
rect 4032 -10392 4096 -10328
rect 4032 -10472 4096 -10408
rect 5444 -9752 5508 -9688
rect 5444 -9832 5508 -9768
rect 5444 -9912 5508 -9848
rect 5444 -9992 5508 -9928
rect 5444 -10072 5508 -10008
rect 5444 -10152 5508 -10088
rect 5444 -10232 5508 -10168
rect 5444 -10312 5508 -10248
rect 5444 -10392 5508 -10328
rect 5444 -10472 5508 -10408
rect 6856 -9752 6920 -9688
rect 6856 -9832 6920 -9768
rect 6856 -9912 6920 -9848
rect 6856 -9992 6920 -9928
rect 6856 -10072 6920 -10008
rect 6856 -10152 6920 -10088
rect 6856 -10232 6920 -10168
rect 6856 -10312 6920 -10248
rect 6856 -10392 6920 -10328
rect 6856 -10472 6920 -10408
rect 8268 -9752 8332 -9688
rect 8268 -9832 8332 -9768
rect 8268 -9912 8332 -9848
rect 8268 -9992 8332 -9928
rect 8268 -10072 8332 -10008
rect 8268 -10152 8332 -10088
rect 8268 -10232 8332 -10168
rect 8268 -10312 8332 -10248
rect 8268 -10392 8332 -10328
rect 8268 -10472 8332 -10408
rect 9680 -9752 9744 -9688
rect 9680 -9832 9744 -9768
rect 9680 -9912 9744 -9848
rect 9680 -9992 9744 -9928
rect 9680 -10072 9744 -10008
rect 9680 -10152 9744 -10088
rect 9680 -10232 9744 -10168
rect 9680 -10312 9744 -10248
rect 9680 -10392 9744 -10328
rect 9680 -10472 9744 -10408
rect 11092 -9752 11156 -9688
rect 11092 -9832 11156 -9768
rect 11092 -9912 11156 -9848
rect 11092 -9992 11156 -9928
rect 11092 -10072 11156 -10008
rect 11092 -10152 11156 -10088
rect 11092 -10232 11156 -10168
rect 11092 -10312 11156 -10248
rect 11092 -10392 11156 -10328
rect 11092 -10472 11156 -10408
rect 12504 -9752 12568 -9688
rect 12504 -9832 12568 -9768
rect 12504 -9912 12568 -9848
rect 12504 -9992 12568 -9928
rect 12504 -10072 12568 -10008
rect 12504 -10152 12568 -10088
rect 12504 -10232 12568 -10168
rect 12504 -10312 12568 -10248
rect 12504 -10392 12568 -10328
rect 12504 -10472 12568 -10408
rect 13916 -9752 13980 -9688
rect 13916 -9832 13980 -9768
rect 13916 -9912 13980 -9848
rect 13916 -9992 13980 -9928
rect 13916 -10072 13980 -10008
rect 13916 -10152 13980 -10088
rect 13916 -10232 13980 -10168
rect 13916 -10312 13980 -10248
rect 13916 -10392 13980 -10328
rect 13916 -10472 13980 -10408
rect 15328 -9752 15392 -9688
rect 15328 -9832 15392 -9768
rect 15328 -9912 15392 -9848
rect 15328 -9992 15392 -9928
rect 15328 -10072 15392 -10008
rect 15328 -10152 15392 -10088
rect 15328 -10232 15392 -10168
rect 15328 -10312 15392 -10248
rect 15328 -10392 15392 -10328
rect 15328 -10472 15392 -10408
rect 16740 -9752 16804 -9688
rect 16740 -9832 16804 -9768
rect 16740 -9912 16804 -9848
rect 16740 -9992 16804 -9928
rect 16740 -10072 16804 -10008
rect 16740 -10152 16804 -10088
rect 16740 -10232 16804 -10168
rect 16740 -10312 16804 -10248
rect 16740 -10392 16804 -10328
rect 16740 -10472 16804 -10408
rect 18152 -9752 18216 -9688
rect 18152 -9832 18216 -9768
rect 18152 -9912 18216 -9848
rect 18152 -9992 18216 -9928
rect 18152 -10072 18216 -10008
rect 18152 -10152 18216 -10088
rect 18152 -10232 18216 -10168
rect 18152 -10312 18216 -10248
rect 18152 -10392 18216 -10328
rect 18152 -10472 18216 -10408
rect 19564 -9752 19628 -9688
rect 19564 -9832 19628 -9768
rect 19564 -9912 19628 -9848
rect 19564 -9992 19628 -9928
rect 19564 -10072 19628 -10008
rect 19564 -10152 19628 -10088
rect 19564 -10232 19628 -10168
rect 19564 -10312 19628 -10248
rect 19564 -10392 19628 -10328
rect 19564 -10472 19628 -10408
rect 20976 -9752 21040 -9688
rect 20976 -9832 21040 -9768
rect 20976 -9912 21040 -9848
rect 20976 -9992 21040 -9928
rect 20976 -10072 21040 -10008
rect 20976 -10152 21040 -10088
rect 20976 -10232 21040 -10168
rect 20976 -10312 21040 -10248
rect 20976 -10392 21040 -10328
rect 20976 -10472 21040 -10408
rect 22388 -9752 22452 -9688
rect 22388 -9832 22452 -9768
rect 22388 -9912 22452 -9848
rect 22388 -9992 22452 -9928
rect 22388 -10072 22452 -10008
rect 22388 -10152 22452 -10088
rect 22388 -10232 22452 -10168
rect 22388 -10312 22452 -10248
rect 22388 -10392 22452 -10328
rect 22388 -10472 22452 -10408
rect 23800 -9752 23864 -9688
rect 23800 -9832 23864 -9768
rect 23800 -9912 23864 -9848
rect 23800 -9992 23864 -9928
rect 23800 -10072 23864 -10008
rect 23800 -10152 23864 -10088
rect 23800 -10232 23864 -10168
rect 23800 -10312 23864 -10248
rect 23800 -10392 23864 -10328
rect 23800 -10472 23864 -10408
rect -22796 -10872 -22732 -10808
rect -22796 -10952 -22732 -10888
rect -22796 -11032 -22732 -10968
rect -22796 -11112 -22732 -11048
rect -22796 -11192 -22732 -11128
rect -22796 -11272 -22732 -11208
rect -22796 -11352 -22732 -11288
rect -22796 -11432 -22732 -11368
rect -22796 -11512 -22732 -11448
rect -22796 -11592 -22732 -11528
rect -21384 -10872 -21320 -10808
rect -21384 -10952 -21320 -10888
rect -21384 -11032 -21320 -10968
rect -21384 -11112 -21320 -11048
rect -21384 -11192 -21320 -11128
rect -21384 -11272 -21320 -11208
rect -21384 -11352 -21320 -11288
rect -21384 -11432 -21320 -11368
rect -21384 -11512 -21320 -11448
rect -21384 -11592 -21320 -11528
rect -19972 -10872 -19908 -10808
rect -19972 -10952 -19908 -10888
rect -19972 -11032 -19908 -10968
rect -19972 -11112 -19908 -11048
rect -19972 -11192 -19908 -11128
rect -19972 -11272 -19908 -11208
rect -19972 -11352 -19908 -11288
rect -19972 -11432 -19908 -11368
rect -19972 -11512 -19908 -11448
rect -19972 -11592 -19908 -11528
rect -18560 -10872 -18496 -10808
rect -18560 -10952 -18496 -10888
rect -18560 -11032 -18496 -10968
rect -18560 -11112 -18496 -11048
rect -18560 -11192 -18496 -11128
rect -18560 -11272 -18496 -11208
rect -18560 -11352 -18496 -11288
rect -18560 -11432 -18496 -11368
rect -18560 -11512 -18496 -11448
rect -18560 -11592 -18496 -11528
rect -17148 -10872 -17084 -10808
rect -17148 -10952 -17084 -10888
rect -17148 -11032 -17084 -10968
rect -17148 -11112 -17084 -11048
rect -17148 -11192 -17084 -11128
rect -17148 -11272 -17084 -11208
rect -17148 -11352 -17084 -11288
rect -17148 -11432 -17084 -11368
rect -17148 -11512 -17084 -11448
rect -17148 -11592 -17084 -11528
rect -15736 -10872 -15672 -10808
rect -15736 -10952 -15672 -10888
rect -15736 -11032 -15672 -10968
rect -15736 -11112 -15672 -11048
rect -15736 -11192 -15672 -11128
rect -15736 -11272 -15672 -11208
rect -15736 -11352 -15672 -11288
rect -15736 -11432 -15672 -11368
rect -15736 -11512 -15672 -11448
rect -15736 -11592 -15672 -11528
rect -14324 -10872 -14260 -10808
rect -14324 -10952 -14260 -10888
rect -14324 -11032 -14260 -10968
rect -14324 -11112 -14260 -11048
rect -14324 -11192 -14260 -11128
rect -14324 -11272 -14260 -11208
rect -14324 -11352 -14260 -11288
rect -14324 -11432 -14260 -11368
rect -14324 -11512 -14260 -11448
rect -14324 -11592 -14260 -11528
rect -12912 -10872 -12848 -10808
rect -12912 -10952 -12848 -10888
rect -12912 -11032 -12848 -10968
rect -12912 -11112 -12848 -11048
rect -12912 -11192 -12848 -11128
rect -12912 -11272 -12848 -11208
rect -12912 -11352 -12848 -11288
rect -12912 -11432 -12848 -11368
rect -12912 -11512 -12848 -11448
rect -12912 -11592 -12848 -11528
rect -11500 -10872 -11436 -10808
rect -11500 -10952 -11436 -10888
rect -11500 -11032 -11436 -10968
rect -11500 -11112 -11436 -11048
rect -11500 -11192 -11436 -11128
rect -11500 -11272 -11436 -11208
rect -11500 -11352 -11436 -11288
rect -11500 -11432 -11436 -11368
rect -11500 -11512 -11436 -11448
rect -11500 -11592 -11436 -11528
rect -10088 -10872 -10024 -10808
rect -10088 -10952 -10024 -10888
rect -10088 -11032 -10024 -10968
rect -10088 -11112 -10024 -11048
rect -10088 -11192 -10024 -11128
rect -10088 -11272 -10024 -11208
rect -10088 -11352 -10024 -11288
rect -10088 -11432 -10024 -11368
rect -10088 -11512 -10024 -11448
rect -10088 -11592 -10024 -11528
rect -8676 -10872 -8612 -10808
rect -8676 -10952 -8612 -10888
rect -8676 -11032 -8612 -10968
rect -8676 -11112 -8612 -11048
rect -8676 -11192 -8612 -11128
rect -8676 -11272 -8612 -11208
rect -8676 -11352 -8612 -11288
rect -8676 -11432 -8612 -11368
rect -8676 -11512 -8612 -11448
rect -8676 -11592 -8612 -11528
rect -7264 -10872 -7200 -10808
rect -7264 -10952 -7200 -10888
rect -7264 -11032 -7200 -10968
rect -7264 -11112 -7200 -11048
rect -7264 -11192 -7200 -11128
rect -7264 -11272 -7200 -11208
rect -7264 -11352 -7200 -11288
rect -7264 -11432 -7200 -11368
rect -7264 -11512 -7200 -11448
rect -7264 -11592 -7200 -11528
rect -5852 -10872 -5788 -10808
rect -5852 -10952 -5788 -10888
rect -5852 -11032 -5788 -10968
rect -5852 -11112 -5788 -11048
rect -5852 -11192 -5788 -11128
rect -5852 -11272 -5788 -11208
rect -5852 -11352 -5788 -11288
rect -5852 -11432 -5788 -11368
rect -5852 -11512 -5788 -11448
rect -5852 -11592 -5788 -11528
rect -4440 -10872 -4376 -10808
rect -4440 -10952 -4376 -10888
rect -4440 -11032 -4376 -10968
rect -4440 -11112 -4376 -11048
rect -4440 -11192 -4376 -11128
rect -4440 -11272 -4376 -11208
rect -4440 -11352 -4376 -11288
rect -4440 -11432 -4376 -11368
rect -4440 -11512 -4376 -11448
rect -4440 -11592 -4376 -11528
rect -3028 -10872 -2964 -10808
rect -3028 -10952 -2964 -10888
rect -3028 -11032 -2964 -10968
rect -3028 -11112 -2964 -11048
rect -3028 -11192 -2964 -11128
rect -3028 -11272 -2964 -11208
rect -3028 -11352 -2964 -11288
rect -3028 -11432 -2964 -11368
rect -3028 -11512 -2964 -11448
rect -3028 -11592 -2964 -11528
rect -1616 -10872 -1552 -10808
rect -1616 -10952 -1552 -10888
rect -1616 -11032 -1552 -10968
rect -1616 -11112 -1552 -11048
rect -1616 -11192 -1552 -11128
rect -1616 -11272 -1552 -11208
rect -1616 -11352 -1552 -11288
rect -1616 -11432 -1552 -11368
rect -1616 -11512 -1552 -11448
rect -1616 -11592 -1552 -11528
rect -204 -10872 -140 -10808
rect -204 -10952 -140 -10888
rect -204 -11032 -140 -10968
rect -204 -11112 -140 -11048
rect -204 -11192 -140 -11128
rect -204 -11272 -140 -11208
rect -204 -11352 -140 -11288
rect -204 -11432 -140 -11368
rect -204 -11512 -140 -11448
rect -204 -11592 -140 -11528
rect 1208 -10872 1272 -10808
rect 1208 -10952 1272 -10888
rect 1208 -11032 1272 -10968
rect 1208 -11112 1272 -11048
rect 1208 -11192 1272 -11128
rect 1208 -11272 1272 -11208
rect 1208 -11352 1272 -11288
rect 1208 -11432 1272 -11368
rect 1208 -11512 1272 -11448
rect 1208 -11592 1272 -11528
rect 2620 -10872 2684 -10808
rect 2620 -10952 2684 -10888
rect 2620 -11032 2684 -10968
rect 2620 -11112 2684 -11048
rect 2620 -11192 2684 -11128
rect 2620 -11272 2684 -11208
rect 2620 -11352 2684 -11288
rect 2620 -11432 2684 -11368
rect 2620 -11512 2684 -11448
rect 2620 -11592 2684 -11528
rect 4032 -10872 4096 -10808
rect 4032 -10952 4096 -10888
rect 4032 -11032 4096 -10968
rect 4032 -11112 4096 -11048
rect 4032 -11192 4096 -11128
rect 4032 -11272 4096 -11208
rect 4032 -11352 4096 -11288
rect 4032 -11432 4096 -11368
rect 4032 -11512 4096 -11448
rect 4032 -11592 4096 -11528
rect 5444 -10872 5508 -10808
rect 5444 -10952 5508 -10888
rect 5444 -11032 5508 -10968
rect 5444 -11112 5508 -11048
rect 5444 -11192 5508 -11128
rect 5444 -11272 5508 -11208
rect 5444 -11352 5508 -11288
rect 5444 -11432 5508 -11368
rect 5444 -11512 5508 -11448
rect 5444 -11592 5508 -11528
rect 6856 -10872 6920 -10808
rect 6856 -10952 6920 -10888
rect 6856 -11032 6920 -10968
rect 6856 -11112 6920 -11048
rect 6856 -11192 6920 -11128
rect 6856 -11272 6920 -11208
rect 6856 -11352 6920 -11288
rect 6856 -11432 6920 -11368
rect 6856 -11512 6920 -11448
rect 6856 -11592 6920 -11528
rect 8268 -10872 8332 -10808
rect 8268 -10952 8332 -10888
rect 8268 -11032 8332 -10968
rect 8268 -11112 8332 -11048
rect 8268 -11192 8332 -11128
rect 8268 -11272 8332 -11208
rect 8268 -11352 8332 -11288
rect 8268 -11432 8332 -11368
rect 8268 -11512 8332 -11448
rect 8268 -11592 8332 -11528
rect 9680 -10872 9744 -10808
rect 9680 -10952 9744 -10888
rect 9680 -11032 9744 -10968
rect 9680 -11112 9744 -11048
rect 9680 -11192 9744 -11128
rect 9680 -11272 9744 -11208
rect 9680 -11352 9744 -11288
rect 9680 -11432 9744 -11368
rect 9680 -11512 9744 -11448
rect 9680 -11592 9744 -11528
rect 11092 -10872 11156 -10808
rect 11092 -10952 11156 -10888
rect 11092 -11032 11156 -10968
rect 11092 -11112 11156 -11048
rect 11092 -11192 11156 -11128
rect 11092 -11272 11156 -11208
rect 11092 -11352 11156 -11288
rect 11092 -11432 11156 -11368
rect 11092 -11512 11156 -11448
rect 11092 -11592 11156 -11528
rect 12504 -10872 12568 -10808
rect 12504 -10952 12568 -10888
rect 12504 -11032 12568 -10968
rect 12504 -11112 12568 -11048
rect 12504 -11192 12568 -11128
rect 12504 -11272 12568 -11208
rect 12504 -11352 12568 -11288
rect 12504 -11432 12568 -11368
rect 12504 -11512 12568 -11448
rect 12504 -11592 12568 -11528
rect 13916 -10872 13980 -10808
rect 13916 -10952 13980 -10888
rect 13916 -11032 13980 -10968
rect 13916 -11112 13980 -11048
rect 13916 -11192 13980 -11128
rect 13916 -11272 13980 -11208
rect 13916 -11352 13980 -11288
rect 13916 -11432 13980 -11368
rect 13916 -11512 13980 -11448
rect 13916 -11592 13980 -11528
rect 15328 -10872 15392 -10808
rect 15328 -10952 15392 -10888
rect 15328 -11032 15392 -10968
rect 15328 -11112 15392 -11048
rect 15328 -11192 15392 -11128
rect 15328 -11272 15392 -11208
rect 15328 -11352 15392 -11288
rect 15328 -11432 15392 -11368
rect 15328 -11512 15392 -11448
rect 15328 -11592 15392 -11528
rect 16740 -10872 16804 -10808
rect 16740 -10952 16804 -10888
rect 16740 -11032 16804 -10968
rect 16740 -11112 16804 -11048
rect 16740 -11192 16804 -11128
rect 16740 -11272 16804 -11208
rect 16740 -11352 16804 -11288
rect 16740 -11432 16804 -11368
rect 16740 -11512 16804 -11448
rect 16740 -11592 16804 -11528
rect 18152 -10872 18216 -10808
rect 18152 -10952 18216 -10888
rect 18152 -11032 18216 -10968
rect 18152 -11112 18216 -11048
rect 18152 -11192 18216 -11128
rect 18152 -11272 18216 -11208
rect 18152 -11352 18216 -11288
rect 18152 -11432 18216 -11368
rect 18152 -11512 18216 -11448
rect 18152 -11592 18216 -11528
rect 19564 -10872 19628 -10808
rect 19564 -10952 19628 -10888
rect 19564 -11032 19628 -10968
rect 19564 -11112 19628 -11048
rect 19564 -11192 19628 -11128
rect 19564 -11272 19628 -11208
rect 19564 -11352 19628 -11288
rect 19564 -11432 19628 -11368
rect 19564 -11512 19628 -11448
rect 19564 -11592 19628 -11528
rect 20976 -10872 21040 -10808
rect 20976 -10952 21040 -10888
rect 20976 -11032 21040 -10968
rect 20976 -11112 21040 -11048
rect 20976 -11192 21040 -11128
rect 20976 -11272 21040 -11208
rect 20976 -11352 21040 -11288
rect 20976 -11432 21040 -11368
rect 20976 -11512 21040 -11448
rect 20976 -11592 21040 -11528
rect 22388 -10872 22452 -10808
rect 22388 -10952 22452 -10888
rect 22388 -11032 22452 -10968
rect 22388 -11112 22452 -11048
rect 22388 -11192 22452 -11128
rect 22388 -11272 22452 -11208
rect 22388 -11352 22452 -11288
rect 22388 -11432 22452 -11368
rect 22388 -11512 22452 -11448
rect 22388 -11592 22452 -11528
rect 23800 -10872 23864 -10808
rect 23800 -10952 23864 -10888
rect 23800 -11032 23864 -10968
rect 23800 -11112 23864 -11048
rect 23800 -11192 23864 -11128
rect 23800 -11272 23864 -11208
rect 23800 -11352 23864 -11288
rect 23800 -11432 23864 -11368
rect 23800 -11512 23864 -11448
rect 23800 -11592 23864 -11528
rect -22796 -11992 -22732 -11928
rect -22796 -12072 -22732 -12008
rect -22796 -12152 -22732 -12088
rect -22796 -12232 -22732 -12168
rect -22796 -12312 -22732 -12248
rect -22796 -12392 -22732 -12328
rect -22796 -12472 -22732 -12408
rect -22796 -12552 -22732 -12488
rect -22796 -12632 -22732 -12568
rect -22796 -12712 -22732 -12648
rect -21384 -11992 -21320 -11928
rect -21384 -12072 -21320 -12008
rect -21384 -12152 -21320 -12088
rect -21384 -12232 -21320 -12168
rect -21384 -12312 -21320 -12248
rect -21384 -12392 -21320 -12328
rect -21384 -12472 -21320 -12408
rect -21384 -12552 -21320 -12488
rect -21384 -12632 -21320 -12568
rect -21384 -12712 -21320 -12648
rect -19972 -11992 -19908 -11928
rect -19972 -12072 -19908 -12008
rect -19972 -12152 -19908 -12088
rect -19972 -12232 -19908 -12168
rect -19972 -12312 -19908 -12248
rect -19972 -12392 -19908 -12328
rect -19972 -12472 -19908 -12408
rect -19972 -12552 -19908 -12488
rect -19972 -12632 -19908 -12568
rect -19972 -12712 -19908 -12648
rect -18560 -11992 -18496 -11928
rect -18560 -12072 -18496 -12008
rect -18560 -12152 -18496 -12088
rect -18560 -12232 -18496 -12168
rect -18560 -12312 -18496 -12248
rect -18560 -12392 -18496 -12328
rect -18560 -12472 -18496 -12408
rect -18560 -12552 -18496 -12488
rect -18560 -12632 -18496 -12568
rect -18560 -12712 -18496 -12648
rect -17148 -11992 -17084 -11928
rect -17148 -12072 -17084 -12008
rect -17148 -12152 -17084 -12088
rect -17148 -12232 -17084 -12168
rect -17148 -12312 -17084 -12248
rect -17148 -12392 -17084 -12328
rect -17148 -12472 -17084 -12408
rect -17148 -12552 -17084 -12488
rect -17148 -12632 -17084 -12568
rect -17148 -12712 -17084 -12648
rect -15736 -11992 -15672 -11928
rect -15736 -12072 -15672 -12008
rect -15736 -12152 -15672 -12088
rect -15736 -12232 -15672 -12168
rect -15736 -12312 -15672 -12248
rect -15736 -12392 -15672 -12328
rect -15736 -12472 -15672 -12408
rect -15736 -12552 -15672 -12488
rect -15736 -12632 -15672 -12568
rect -15736 -12712 -15672 -12648
rect -14324 -11992 -14260 -11928
rect -14324 -12072 -14260 -12008
rect -14324 -12152 -14260 -12088
rect -14324 -12232 -14260 -12168
rect -14324 -12312 -14260 -12248
rect -14324 -12392 -14260 -12328
rect -14324 -12472 -14260 -12408
rect -14324 -12552 -14260 -12488
rect -14324 -12632 -14260 -12568
rect -14324 -12712 -14260 -12648
rect -12912 -11992 -12848 -11928
rect -12912 -12072 -12848 -12008
rect -12912 -12152 -12848 -12088
rect -12912 -12232 -12848 -12168
rect -12912 -12312 -12848 -12248
rect -12912 -12392 -12848 -12328
rect -12912 -12472 -12848 -12408
rect -12912 -12552 -12848 -12488
rect -12912 -12632 -12848 -12568
rect -12912 -12712 -12848 -12648
rect -11500 -11992 -11436 -11928
rect -11500 -12072 -11436 -12008
rect -11500 -12152 -11436 -12088
rect -11500 -12232 -11436 -12168
rect -11500 -12312 -11436 -12248
rect -11500 -12392 -11436 -12328
rect -11500 -12472 -11436 -12408
rect -11500 -12552 -11436 -12488
rect -11500 -12632 -11436 -12568
rect -11500 -12712 -11436 -12648
rect -10088 -11992 -10024 -11928
rect -10088 -12072 -10024 -12008
rect -10088 -12152 -10024 -12088
rect -10088 -12232 -10024 -12168
rect -10088 -12312 -10024 -12248
rect -10088 -12392 -10024 -12328
rect -10088 -12472 -10024 -12408
rect -10088 -12552 -10024 -12488
rect -10088 -12632 -10024 -12568
rect -10088 -12712 -10024 -12648
rect -8676 -11992 -8612 -11928
rect -8676 -12072 -8612 -12008
rect -8676 -12152 -8612 -12088
rect -8676 -12232 -8612 -12168
rect -8676 -12312 -8612 -12248
rect -8676 -12392 -8612 -12328
rect -8676 -12472 -8612 -12408
rect -8676 -12552 -8612 -12488
rect -8676 -12632 -8612 -12568
rect -8676 -12712 -8612 -12648
rect -7264 -11992 -7200 -11928
rect -7264 -12072 -7200 -12008
rect -7264 -12152 -7200 -12088
rect -7264 -12232 -7200 -12168
rect -7264 -12312 -7200 -12248
rect -7264 -12392 -7200 -12328
rect -7264 -12472 -7200 -12408
rect -7264 -12552 -7200 -12488
rect -7264 -12632 -7200 -12568
rect -7264 -12712 -7200 -12648
rect -5852 -11992 -5788 -11928
rect -5852 -12072 -5788 -12008
rect -5852 -12152 -5788 -12088
rect -5852 -12232 -5788 -12168
rect -5852 -12312 -5788 -12248
rect -5852 -12392 -5788 -12328
rect -5852 -12472 -5788 -12408
rect -5852 -12552 -5788 -12488
rect -5852 -12632 -5788 -12568
rect -5852 -12712 -5788 -12648
rect -4440 -11992 -4376 -11928
rect -4440 -12072 -4376 -12008
rect -4440 -12152 -4376 -12088
rect -4440 -12232 -4376 -12168
rect -4440 -12312 -4376 -12248
rect -4440 -12392 -4376 -12328
rect -4440 -12472 -4376 -12408
rect -4440 -12552 -4376 -12488
rect -4440 -12632 -4376 -12568
rect -4440 -12712 -4376 -12648
rect -3028 -11992 -2964 -11928
rect -3028 -12072 -2964 -12008
rect -3028 -12152 -2964 -12088
rect -3028 -12232 -2964 -12168
rect -3028 -12312 -2964 -12248
rect -3028 -12392 -2964 -12328
rect -3028 -12472 -2964 -12408
rect -3028 -12552 -2964 -12488
rect -3028 -12632 -2964 -12568
rect -3028 -12712 -2964 -12648
rect -1616 -11992 -1552 -11928
rect -1616 -12072 -1552 -12008
rect -1616 -12152 -1552 -12088
rect -1616 -12232 -1552 -12168
rect -1616 -12312 -1552 -12248
rect -1616 -12392 -1552 -12328
rect -1616 -12472 -1552 -12408
rect -1616 -12552 -1552 -12488
rect -1616 -12632 -1552 -12568
rect -1616 -12712 -1552 -12648
rect -204 -11992 -140 -11928
rect -204 -12072 -140 -12008
rect -204 -12152 -140 -12088
rect -204 -12232 -140 -12168
rect -204 -12312 -140 -12248
rect -204 -12392 -140 -12328
rect -204 -12472 -140 -12408
rect -204 -12552 -140 -12488
rect -204 -12632 -140 -12568
rect -204 -12712 -140 -12648
rect 1208 -11992 1272 -11928
rect 1208 -12072 1272 -12008
rect 1208 -12152 1272 -12088
rect 1208 -12232 1272 -12168
rect 1208 -12312 1272 -12248
rect 1208 -12392 1272 -12328
rect 1208 -12472 1272 -12408
rect 1208 -12552 1272 -12488
rect 1208 -12632 1272 -12568
rect 1208 -12712 1272 -12648
rect 2620 -11992 2684 -11928
rect 2620 -12072 2684 -12008
rect 2620 -12152 2684 -12088
rect 2620 -12232 2684 -12168
rect 2620 -12312 2684 -12248
rect 2620 -12392 2684 -12328
rect 2620 -12472 2684 -12408
rect 2620 -12552 2684 -12488
rect 2620 -12632 2684 -12568
rect 2620 -12712 2684 -12648
rect 4032 -11992 4096 -11928
rect 4032 -12072 4096 -12008
rect 4032 -12152 4096 -12088
rect 4032 -12232 4096 -12168
rect 4032 -12312 4096 -12248
rect 4032 -12392 4096 -12328
rect 4032 -12472 4096 -12408
rect 4032 -12552 4096 -12488
rect 4032 -12632 4096 -12568
rect 4032 -12712 4096 -12648
rect 5444 -11992 5508 -11928
rect 5444 -12072 5508 -12008
rect 5444 -12152 5508 -12088
rect 5444 -12232 5508 -12168
rect 5444 -12312 5508 -12248
rect 5444 -12392 5508 -12328
rect 5444 -12472 5508 -12408
rect 5444 -12552 5508 -12488
rect 5444 -12632 5508 -12568
rect 5444 -12712 5508 -12648
rect 6856 -11992 6920 -11928
rect 6856 -12072 6920 -12008
rect 6856 -12152 6920 -12088
rect 6856 -12232 6920 -12168
rect 6856 -12312 6920 -12248
rect 6856 -12392 6920 -12328
rect 6856 -12472 6920 -12408
rect 6856 -12552 6920 -12488
rect 6856 -12632 6920 -12568
rect 6856 -12712 6920 -12648
rect 8268 -11992 8332 -11928
rect 8268 -12072 8332 -12008
rect 8268 -12152 8332 -12088
rect 8268 -12232 8332 -12168
rect 8268 -12312 8332 -12248
rect 8268 -12392 8332 -12328
rect 8268 -12472 8332 -12408
rect 8268 -12552 8332 -12488
rect 8268 -12632 8332 -12568
rect 8268 -12712 8332 -12648
rect 9680 -11992 9744 -11928
rect 9680 -12072 9744 -12008
rect 9680 -12152 9744 -12088
rect 9680 -12232 9744 -12168
rect 9680 -12312 9744 -12248
rect 9680 -12392 9744 -12328
rect 9680 -12472 9744 -12408
rect 9680 -12552 9744 -12488
rect 9680 -12632 9744 -12568
rect 9680 -12712 9744 -12648
rect 11092 -11992 11156 -11928
rect 11092 -12072 11156 -12008
rect 11092 -12152 11156 -12088
rect 11092 -12232 11156 -12168
rect 11092 -12312 11156 -12248
rect 11092 -12392 11156 -12328
rect 11092 -12472 11156 -12408
rect 11092 -12552 11156 -12488
rect 11092 -12632 11156 -12568
rect 11092 -12712 11156 -12648
rect 12504 -11992 12568 -11928
rect 12504 -12072 12568 -12008
rect 12504 -12152 12568 -12088
rect 12504 -12232 12568 -12168
rect 12504 -12312 12568 -12248
rect 12504 -12392 12568 -12328
rect 12504 -12472 12568 -12408
rect 12504 -12552 12568 -12488
rect 12504 -12632 12568 -12568
rect 12504 -12712 12568 -12648
rect 13916 -11992 13980 -11928
rect 13916 -12072 13980 -12008
rect 13916 -12152 13980 -12088
rect 13916 -12232 13980 -12168
rect 13916 -12312 13980 -12248
rect 13916 -12392 13980 -12328
rect 13916 -12472 13980 -12408
rect 13916 -12552 13980 -12488
rect 13916 -12632 13980 -12568
rect 13916 -12712 13980 -12648
rect 15328 -11992 15392 -11928
rect 15328 -12072 15392 -12008
rect 15328 -12152 15392 -12088
rect 15328 -12232 15392 -12168
rect 15328 -12312 15392 -12248
rect 15328 -12392 15392 -12328
rect 15328 -12472 15392 -12408
rect 15328 -12552 15392 -12488
rect 15328 -12632 15392 -12568
rect 15328 -12712 15392 -12648
rect 16740 -11992 16804 -11928
rect 16740 -12072 16804 -12008
rect 16740 -12152 16804 -12088
rect 16740 -12232 16804 -12168
rect 16740 -12312 16804 -12248
rect 16740 -12392 16804 -12328
rect 16740 -12472 16804 -12408
rect 16740 -12552 16804 -12488
rect 16740 -12632 16804 -12568
rect 16740 -12712 16804 -12648
rect 18152 -11992 18216 -11928
rect 18152 -12072 18216 -12008
rect 18152 -12152 18216 -12088
rect 18152 -12232 18216 -12168
rect 18152 -12312 18216 -12248
rect 18152 -12392 18216 -12328
rect 18152 -12472 18216 -12408
rect 18152 -12552 18216 -12488
rect 18152 -12632 18216 -12568
rect 18152 -12712 18216 -12648
rect 19564 -11992 19628 -11928
rect 19564 -12072 19628 -12008
rect 19564 -12152 19628 -12088
rect 19564 -12232 19628 -12168
rect 19564 -12312 19628 -12248
rect 19564 -12392 19628 -12328
rect 19564 -12472 19628 -12408
rect 19564 -12552 19628 -12488
rect 19564 -12632 19628 -12568
rect 19564 -12712 19628 -12648
rect 20976 -11992 21040 -11928
rect 20976 -12072 21040 -12008
rect 20976 -12152 21040 -12088
rect 20976 -12232 21040 -12168
rect 20976 -12312 21040 -12248
rect 20976 -12392 21040 -12328
rect 20976 -12472 21040 -12408
rect 20976 -12552 21040 -12488
rect 20976 -12632 21040 -12568
rect 20976 -12712 21040 -12648
rect 22388 -11992 22452 -11928
rect 22388 -12072 22452 -12008
rect 22388 -12152 22452 -12088
rect 22388 -12232 22452 -12168
rect 22388 -12312 22452 -12248
rect 22388 -12392 22452 -12328
rect 22388 -12472 22452 -12408
rect 22388 -12552 22452 -12488
rect 22388 -12632 22452 -12568
rect 22388 -12712 22452 -12648
rect 23800 -11992 23864 -11928
rect 23800 -12072 23864 -12008
rect 23800 -12152 23864 -12088
rect 23800 -12232 23864 -12168
rect 23800 -12312 23864 -12248
rect 23800 -12392 23864 -12328
rect 23800 -12472 23864 -12408
rect 23800 -12552 23864 -12488
rect 23800 -12632 23864 -12568
rect 23800 -12712 23864 -12648
rect -22796 -13112 -22732 -13048
rect -22796 -13192 -22732 -13128
rect -22796 -13272 -22732 -13208
rect -22796 -13352 -22732 -13288
rect -22796 -13432 -22732 -13368
rect -22796 -13512 -22732 -13448
rect -22796 -13592 -22732 -13528
rect -22796 -13672 -22732 -13608
rect -22796 -13752 -22732 -13688
rect -22796 -13832 -22732 -13768
rect -21384 -13112 -21320 -13048
rect -21384 -13192 -21320 -13128
rect -21384 -13272 -21320 -13208
rect -21384 -13352 -21320 -13288
rect -21384 -13432 -21320 -13368
rect -21384 -13512 -21320 -13448
rect -21384 -13592 -21320 -13528
rect -21384 -13672 -21320 -13608
rect -21384 -13752 -21320 -13688
rect -21384 -13832 -21320 -13768
rect -19972 -13112 -19908 -13048
rect -19972 -13192 -19908 -13128
rect -19972 -13272 -19908 -13208
rect -19972 -13352 -19908 -13288
rect -19972 -13432 -19908 -13368
rect -19972 -13512 -19908 -13448
rect -19972 -13592 -19908 -13528
rect -19972 -13672 -19908 -13608
rect -19972 -13752 -19908 -13688
rect -19972 -13832 -19908 -13768
rect -18560 -13112 -18496 -13048
rect -18560 -13192 -18496 -13128
rect -18560 -13272 -18496 -13208
rect -18560 -13352 -18496 -13288
rect -18560 -13432 -18496 -13368
rect -18560 -13512 -18496 -13448
rect -18560 -13592 -18496 -13528
rect -18560 -13672 -18496 -13608
rect -18560 -13752 -18496 -13688
rect -18560 -13832 -18496 -13768
rect -17148 -13112 -17084 -13048
rect -17148 -13192 -17084 -13128
rect -17148 -13272 -17084 -13208
rect -17148 -13352 -17084 -13288
rect -17148 -13432 -17084 -13368
rect -17148 -13512 -17084 -13448
rect -17148 -13592 -17084 -13528
rect -17148 -13672 -17084 -13608
rect -17148 -13752 -17084 -13688
rect -17148 -13832 -17084 -13768
rect -15736 -13112 -15672 -13048
rect -15736 -13192 -15672 -13128
rect -15736 -13272 -15672 -13208
rect -15736 -13352 -15672 -13288
rect -15736 -13432 -15672 -13368
rect -15736 -13512 -15672 -13448
rect -15736 -13592 -15672 -13528
rect -15736 -13672 -15672 -13608
rect -15736 -13752 -15672 -13688
rect -15736 -13832 -15672 -13768
rect -14324 -13112 -14260 -13048
rect -14324 -13192 -14260 -13128
rect -14324 -13272 -14260 -13208
rect -14324 -13352 -14260 -13288
rect -14324 -13432 -14260 -13368
rect -14324 -13512 -14260 -13448
rect -14324 -13592 -14260 -13528
rect -14324 -13672 -14260 -13608
rect -14324 -13752 -14260 -13688
rect -14324 -13832 -14260 -13768
rect -12912 -13112 -12848 -13048
rect -12912 -13192 -12848 -13128
rect -12912 -13272 -12848 -13208
rect -12912 -13352 -12848 -13288
rect -12912 -13432 -12848 -13368
rect -12912 -13512 -12848 -13448
rect -12912 -13592 -12848 -13528
rect -12912 -13672 -12848 -13608
rect -12912 -13752 -12848 -13688
rect -12912 -13832 -12848 -13768
rect -11500 -13112 -11436 -13048
rect -11500 -13192 -11436 -13128
rect -11500 -13272 -11436 -13208
rect -11500 -13352 -11436 -13288
rect -11500 -13432 -11436 -13368
rect -11500 -13512 -11436 -13448
rect -11500 -13592 -11436 -13528
rect -11500 -13672 -11436 -13608
rect -11500 -13752 -11436 -13688
rect -11500 -13832 -11436 -13768
rect -10088 -13112 -10024 -13048
rect -10088 -13192 -10024 -13128
rect -10088 -13272 -10024 -13208
rect -10088 -13352 -10024 -13288
rect -10088 -13432 -10024 -13368
rect -10088 -13512 -10024 -13448
rect -10088 -13592 -10024 -13528
rect -10088 -13672 -10024 -13608
rect -10088 -13752 -10024 -13688
rect -10088 -13832 -10024 -13768
rect -8676 -13112 -8612 -13048
rect -8676 -13192 -8612 -13128
rect -8676 -13272 -8612 -13208
rect -8676 -13352 -8612 -13288
rect -8676 -13432 -8612 -13368
rect -8676 -13512 -8612 -13448
rect -8676 -13592 -8612 -13528
rect -8676 -13672 -8612 -13608
rect -8676 -13752 -8612 -13688
rect -8676 -13832 -8612 -13768
rect -7264 -13112 -7200 -13048
rect -7264 -13192 -7200 -13128
rect -7264 -13272 -7200 -13208
rect -7264 -13352 -7200 -13288
rect -7264 -13432 -7200 -13368
rect -7264 -13512 -7200 -13448
rect -7264 -13592 -7200 -13528
rect -7264 -13672 -7200 -13608
rect -7264 -13752 -7200 -13688
rect -7264 -13832 -7200 -13768
rect -5852 -13112 -5788 -13048
rect -5852 -13192 -5788 -13128
rect -5852 -13272 -5788 -13208
rect -5852 -13352 -5788 -13288
rect -5852 -13432 -5788 -13368
rect -5852 -13512 -5788 -13448
rect -5852 -13592 -5788 -13528
rect -5852 -13672 -5788 -13608
rect -5852 -13752 -5788 -13688
rect -5852 -13832 -5788 -13768
rect -4440 -13112 -4376 -13048
rect -4440 -13192 -4376 -13128
rect -4440 -13272 -4376 -13208
rect -4440 -13352 -4376 -13288
rect -4440 -13432 -4376 -13368
rect -4440 -13512 -4376 -13448
rect -4440 -13592 -4376 -13528
rect -4440 -13672 -4376 -13608
rect -4440 -13752 -4376 -13688
rect -4440 -13832 -4376 -13768
rect -3028 -13112 -2964 -13048
rect -3028 -13192 -2964 -13128
rect -3028 -13272 -2964 -13208
rect -3028 -13352 -2964 -13288
rect -3028 -13432 -2964 -13368
rect -3028 -13512 -2964 -13448
rect -3028 -13592 -2964 -13528
rect -3028 -13672 -2964 -13608
rect -3028 -13752 -2964 -13688
rect -3028 -13832 -2964 -13768
rect -1616 -13112 -1552 -13048
rect -1616 -13192 -1552 -13128
rect -1616 -13272 -1552 -13208
rect -1616 -13352 -1552 -13288
rect -1616 -13432 -1552 -13368
rect -1616 -13512 -1552 -13448
rect -1616 -13592 -1552 -13528
rect -1616 -13672 -1552 -13608
rect -1616 -13752 -1552 -13688
rect -1616 -13832 -1552 -13768
rect -204 -13112 -140 -13048
rect -204 -13192 -140 -13128
rect -204 -13272 -140 -13208
rect -204 -13352 -140 -13288
rect -204 -13432 -140 -13368
rect -204 -13512 -140 -13448
rect -204 -13592 -140 -13528
rect -204 -13672 -140 -13608
rect -204 -13752 -140 -13688
rect -204 -13832 -140 -13768
rect 1208 -13112 1272 -13048
rect 1208 -13192 1272 -13128
rect 1208 -13272 1272 -13208
rect 1208 -13352 1272 -13288
rect 1208 -13432 1272 -13368
rect 1208 -13512 1272 -13448
rect 1208 -13592 1272 -13528
rect 1208 -13672 1272 -13608
rect 1208 -13752 1272 -13688
rect 1208 -13832 1272 -13768
rect 2620 -13112 2684 -13048
rect 2620 -13192 2684 -13128
rect 2620 -13272 2684 -13208
rect 2620 -13352 2684 -13288
rect 2620 -13432 2684 -13368
rect 2620 -13512 2684 -13448
rect 2620 -13592 2684 -13528
rect 2620 -13672 2684 -13608
rect 2620 -13752 2684 -13688
rect 2620 -13832 2684 -13768
rect 4032 -13112 4096 -13048
rect 4032 -13192 4096 -13128
rect 4032 -13272 4096 -13208
rect 4032 -13352 4096 -13288
rect 4032 -13432 4096 -13368
rect 4032 -13512 4096 -13448
rect 4032 -13592 4096 -13528
rect 4032 -13672 4096 -13608
rect 4032 -13752 4096 -13688
rect 4032 -13832 4096 -13768
rect 5444 -13112 5508 -13048
rect 5444 -13192 5508 -13128
rect 5444 -13272 5508 -13208
rect 5444 -13352 5508 -13288
rect 5444 -13432 5508 -13368
rect 5444 -13512 5508 -13448
rect 5444 -13592 5508 -13528
rect 5444 -13672 5508 -13608
rect 5444 -13752 5508 -13688
rect 5444 -13832 5508 -13768
rect 6856 -13112 6920 -13048
rect 6856 -13192 6920 -13128
rect 6856 -13272 6920 -13208
rect 6856 -13352 6920 -13288
rect 6856 -13432 6920 -13368
rect 6856 -13512 6920 -13448
rect 6856 -13592 6920 -13528
rect 6856 -13672 6920 -13608
rect 6856 -13752 6920 -13688
rect 6856 -13832 6920 -13768
rect 8268 -13112 8332 -13048
rect 8268 -13192 8332 -13128
rect 8268 -13272 8332 -13208
rect 8268 -13352 8332 -13288
rect 8268 -13432 8332 -13368
rect 8268 -13512 8332 -13448
rect 8268 -13592 8332 -13528
rect 8268 -13672 8332 -13608
rect 8268 -13752 8332 -13688
rect 8268 -13832 8332 -13768
rect 9680 -13112 9744 -13048
rect 9680 -13192 9744 -13128
rect 9680 -13272 9744 -13208
rect 9680 -13352 9744 -13288
rect 9680 -13432 9744 -13368
rect 9680 -13512 9744 -13448
rect 9680 -13592 9744 -13528
rect 9680 -13672 9744 -13608
rect 9680 -13752 9744 -13688
rect 9680 -13832 9744 -13768
rect 11092 -13112 11156 -13048
rect 11092 -13192 11156 -13128
rect 11092 -13272 11156 -13208
rect 11092 -13352 11156 -13288
rect 11092 -13432 11156 -13368
rect 11092 -13512 11156 -13448
rect 11092 -13592 11156 -13528
rect 11092 -13672 11156 -13608
rect 11092 -13752 11156 -13688
rect 11092 -13832 11156 -13768
rect 12504 -13112 12568 -13048
rect 12504 -13192 12568 -13128
rect 12504 -13272 12568 -13208
rect 12504 -13352 12568 -13288
rect 12504 -13432 12568 -13368
rect 12504 -13512 12568 -13448
rect 12504 -13592 12568 -13528
rect 12504 -13672 12568 -13608
rect 12504 -13752 12568 -13688
rect 12504 -13832 12568 -13768
rect 13916 -13112 13980 -13048
rect 13916 -13192 13980 -13128
rect 13916 -13272 13980 -13208
rect 13916 -13352 13980 -13288
rect 13916 -13432 13980 -13368
rect 13916 -13512 13980 -13448
rect 13916 -13592 13980 -13528
rect 13916 -13672 13980 -13608
rect 13916 -13752 13980 -13688
rect 13916 -13832 13980 -13768
rect 15328 -13112 15392 -13048
rect 15328 -13192 15392 -13128
rect 15328 -13272 15392 -13208
rect 15328 -13352 15392 -13288
rect 15328 -13432 15392 -13368
rect 15328 -13512 15392 -13448
rect 15328 -13592 15392 -13528
rect 15328 -13672 15392 -13608
rect 15328 -13752 15392 -13688
rect 15328 -13832 15392 -13768
rect 16740 -13112 16804 -13048
rect 16740 -13192 16804 -13128
rect 16740 -13272 16804 -13208
rect 16740 -13352 16804 -13288
rect 16740 -13432 16804 -13368
rect 16740 -13512 16804 -13448
rect 16740 -13592 16804 -13528
rect 16740 -13672 16804 -13608
rect 16740 -13752 16804 -13688
rect 16740 -13832 16804 -13768
rect 18152 -13112 18216 -13048
rect 18152 -13192 18216 -13128
rect 18152 -13272 18216 -13208
rect 18152 -13352 18216 -13288
rect 18152 -13432 18216 -13368
rect 18152 -13512 18216 -13448
rect 18152 -13592 18216 -13528
rect 18152 -13672 18216 -13608
rect 18152 -13752 18216 -13688
rect 18152 -13832 18216 -13768
rect 19564 -13112 19628 -13048
rect 19564 -13192 19628 -13128
rect 19564 -13272 19628 -13208
rect 19564 -13352 19628 -13288
rect 19564 -13432 19628 -13368
rect 19564 -13512 19628 -13448
rect 19564 -13592 19628 -13528
rect 19564 -13672 19628 -13608
rect 19564 -13752 19628 -13688
rect 19564 -13832 19628 -13768
rect 20976 -13112 21040 -13048
rect 20976 -13192 21040 -13128
rect 20976 -13272 21040 -13208
rect 20976 -13352 21040 -13288
rect 20976 -13432 21040 -13368
rect 20976 -13512 21040 -13448
rect 20976 -13592 21040 -13528
rect 20976 -13672 21040 -13608
rect 20976 -13752 21040 -13688
rect 20976 -13832 21040 -13768
rect 22388 -13112 22452 -13048
rect 22388 -13192 22452 -13128
rect 22388 -13272 22452 -13208
rect 22388 -13352 22452 -13288
rect 22388 -13432 22452 -13368
rect 22388 -13512 22452 -13448
rect 22388 -13592 22452 -13528
rect 22388 -13672 22452 -13608
rect 22388 -13752 22452 -13688
rect 22388 -13832 22452 -13768
rect 23800 -13112 23864 -13048
rect 23800 -13192 23864 -13128
rect 23800 -13272 23864 -13208
rect 23800 -13352 23864 -13288
rect 23800 -13432 23864 -13368
rect 23800 -13512 23864 -13448
rect 23800 -13592 23864 -13528
rect 23800 -13672 23864 -13608
rect 23800 -13752 23864 -13688
rect 23800 -13832 23864 -13768
rect -22796 -14232 -22732 -14168
rect -22796 -14312 -22732 -14248
rect -22796 -14392 -22732 -14328
rect -22796 -14472 -22732 -14408
rect -22796 -14552 -22732 -14488
rect -22796 -14632 -22732 -14568
rect -22796 -14712 -22732 -14648
rect -22796 -14792 -22732 -14728
rect -22796 -14872 -22732 -14808
rect -22796 -14952 -22732 -14888
rect -21384 -14232 -21320 -14168
rect -21384 -14312 -21320 -14248
rect -21384 -14392 -21320 -14328
rect -21384 -14472 -21320 -14408
rect -21384 -14552 -21320 -14488
rect -21384 -14632 -21320 -14568
rect -21384 -14712 -21320 -14648
rect -21384 -14792 -21320 -14728
rect -21384 -14872 -21320 -14808
rect -21384 -14952 -21320 -14888
rect -19972 -14232 -19908 -14168
rect -19972 -14312 -19908 -14248
rect -19972 -14392 -19908 -14328
rect -19972 -14472 -19908 -14408
rect -19972 -14552 -19908 -14488
rect -19972 -14632 -19908 -14568
rect -19972 -14712 -19908 -14648
rect -19972 -14792 -19908 -14728
rect -19972 -14872 -19908 -14808
rect -19972 -14952 -19908 -14888
rect -18560 -14232 -18496 -14168
rect -18560 -14312 -18496 -14248
rect -18560 -14392 -18496 -14328
rect -18560 -14472 -18496 -14408
rect -18560 -14552 -18496 -14488
rect -18560 -14632 -18496 -14568
rect -18560 -14712 -18496 -14648
rect -18560 -14792 -18496 -14728
rect -18560 -14872 -18496 -14808
rect -18560 -14952 -18496 -14888
rect -17148 -14232 -17084 -14168
rect -17148 -14312 -17084 -14248
rect -17148 -14392 -17084 -14328
rect -17148 -14472 -17084 -14408
rect -17148 -14552 -17084 -14488
rect -17148 -14632 -17084 -14568
rect -17148 -14712 -17084 -14648
rect -17148 -14792 -17084 -14728
rect -17148 -14872 -17084 -14808
rect -17148 -14952 -17084 -14888
rect -15736 -14232 -15672 -14168
rect -15736 -14312 -15672 -14248
rect -15736 -14392 -15672 -14328
rect -15736 -14472 -15672 -14408
rect -15736 -14552 -15672 -14488
rect -15736 -14632 -15672 -14568
rect -15736 -14712 -15672 -14648
rect -15736 -14792 -15672 -14728
rect -15736 -14872 -15672 -14808
rect -15736 -14952 -15672 -14888
rect -14324 -14232 -14260 -14168
rect -14324 -14312 -14260 -14248
rect -14324 -14392 -14260 -14328
rect -14324 -14472 -14260 -14408
rect -14324 -14552 -14260 -14488
rect -14324 -14632 -14260 -14568
rect -14324 -14712 -14260 -14648
rect -14324 -14792 -14260 -14728
rect -14324 -14872 -14260 -14808
rect -14324 -14952 -14260 -14888
rect -12912 -14232 -12848 -14168
rect -12912 -14312 -12848 -14248
rect -12912 -14392 -12848 -14328
rect -12912 -14472 -12848 -14408
rect -12912 -14552 -12848 -14488
rect -12912 -14632 -12848 -14568
rect -12912 -14712 -12848 -14648
rect -12912 -14792 -12848 -14728
rect -12912 -14872 -12848 -14808
rect -12912 -14952 -12848 -14888
rect -11500 -14232 -11436 -14168
rect -11500 -14312 -11436 -14248
rect -11500 -14392 -11436 -14328
rect -11500 -14472 -11436 -14408
rect -11500 -14552 -11436 -14488
rect -11500 -14632 -11436 -14568
rect -11500 -14712 -11436 -14648
rect -11500 -14792 -11436 -14728
rect -11500 -14872 -11436 -14808
rect -11500 -14952 -11436 -14888
rect -10088 -14232 -10024 -14168
rect -10088 -14312 -10024 -14248
rect -10088 -14392 -10024 -14328
rect -10088 -14472 -10024 -14408
rect -10088 -14552 -10024 -14488
rect -10088 -14632 -10024 -14568
rect -10088 -14712 -10024 -14648
rect -10088 -14792 -10024 -14728
rect -10088 -14872 -10024 -14808
rect -10088 -14952 -10024 -14888
rect -8676 -14232 -8612 -14168
rect -8676 -14312 -8612 -14248
rect -8676 -14392 -8612 -14328
rect -8676 -14472 -8612 -14408
rect -8676 -14552 -8612 -14488
rect -8676 -14632 -8612 -14568
rect -8676 -14712 -8612 -14648
rect -8676 -14792 -8612 -14728
rect -8676 -14872 -8612 -14808
rect -8676 -14952 -8612 -14888
rect -7264 -14232 -7200 -14168
rect -7264 -14312 -7200 -14248
rect -7264 -14392 -7200 -14328
rect -7264 -14472 -7200 -14408
rect -7264 -14552 -7200 -14488
rect -7264 -14632 -7200 -14568
rect -7264 -14712 -7200 -14648
rect -7264 -14792 -7200 -14728
rect -7264 -14872 -7200 -14808
rect -7264 -14952 -7200 -14888
rect -5852 -14232 -5788 -14168
rect -5852 -14312 -5788 -14248
rect -5852 -14392 -5788 -14328
rect -5852 -14472 -5788 -14408
rect -5852 -14552 -5788 -14488
rect -5852 -14632 -5788 -14568
rect -5852 -14712 -5788 -14648
rect -5852 -14792 -5788 -14728
rect -5852 -14872 -5788 -14808
rect -5852 -14952 -5788 -14888
rect -4440 -14232 -4376 -14168
rect -4440 -14312 -4376 -14248
rect -4440 -14392 -4376 -14328
rect -4440 -14472 -4376 -14408
rect -4440 -14552 -4376 -14488
rect -4440 -14632 -4376 -14568
rect -4440 -14712 -4376 -14648
rect -4440 -14792 -4376 -14728
rect -4440 -14872 -4376 -14808
rect -4440 -14952 -4376 -14888
rect -3028 -14232 -2964 -14168
rect -3028 -14312 -2964 -14248
rect -3028 -14392 -2964 -14328
rect -3028 -14472 -2964 -14408
rect -3028 -14552 -2964 -14488
rect -3028 -14632 -2964 -14568
rect -3028 -14712 -2964 -14648
rect -3028 -14792 -2964 -14728
rect -3028 -14872 -2964 -14808
rect -3028 -14952 -2964 -14888
rect -1616 -14232 -1552 -14168
rect -1616 -14312 -1552 -14248
rect -1616 -14392 -1552 -14328
rect -1616 -14472 -1552 -14408
rect -1616 -14552 -1552 -14488
rect -1616 -14632 -1552 -14568
rect -1616 -14712 -1552 -14648
rect -1616 -14792 -1552 -14728
rect -1616 -14872 -1552 -14808
rect -1616 -14952 -1552 -14888
rect -204 -14232 -140 -14168
rect -204 -14312 -140 -14248
rect -204 -14392 -140 -14328
rect -204 -14472 -140 -14408
rect -204 -14552 -140 -14488
rect -204 -14632 -140 -14568
rect -204 -14712 -140 -14648
rect -204 -14792 -140 -14728
rect -204 -14872 -140 -14808
rect -204 -14952 -140 -14888
rect 1208 -14232 1272 -14168
rect 1208 -14312 1272 -14248
rect 1208 -14392 1272 -14328
rect 1208 -14472 1272 -14408
rect 1208 -14552 1272 -14488
rect 1208 -14632 1272 -14568
rect 1208 -14712 1272 -14648
rect 1208 -14792 1272 -14728
rect 1208 -14872 1272 -14808
rect 1208 -14952 1272 -14888
rect 2620 -14232 2684 -14168
rect 2620 -14312 2684 -14248
rect 2620 -14392 2684 -14328
rect 2620 -14472 2684 -14408
rect 2620 -14552 2684 -14488
rect 2620 -14632 2684 -14568
rect 2620 -14712 2684 -14648
rect 2620 -14792 2684 -14728
rect 2620 -14872 2684 -14808
rect 2620 -14952 2684 -14888
rect 4032 -14232 4096 -14168
rect 4032 -14312 4096 -14248
rect 4032 -14392 4096 -14328
rect 4032 -14472 4096 -14408
rect 4032 -14552 4096 -14488
rect 4032 -14632 4096 -14568
rect 4032 -14712 4096 -14648
rect 4032 -14792 4096 -14728
rect 4032 -14872 4096 -14808
rect 4032 -14952 4096 -14888
rect 5444 -14232 5508 -14168
rect 5444 -14312 5508 -14248
rect 5444 -14392 5508 -14328
rect 5444 -14472 5508 -14408
rect 5444 -14552 5508 -14488
rect 5444 -14632 5508 -14568
rect 5444 -14712 5508 -14648
rect 5444 -14792 5508 -14728
rect 5444 -14872 5508 -14808
rect 5444 -14952 5508 -14888
rect 6856 -14232 6920 -14168
rect 6856 -14312 6920 -14248
rect 6856 -14392 6920 -14328
rect 6856 -14472 6920 -14408
rect 6856 -14552 6920 -14488
rect 6856 -14632 6920 -14568
rect 6856 -14712 6920 -14648
rect 6856 -14792 6920 -14728
rect 6856 -14872 6920 -14808
rect 6856 -14952 6920 -14888
rect 8268 -14232 8332 -14168
rect 8268 -14312 8332 -14248
rect 8268 -14392 8332 -14328
rect 8268 -14472 8332 -14408
rect 8268 -14552 8332 -14488
rect 8268 -14632 8332 -14568
rect 8268 -14712 8332 -14648
rect 8268 -14792 8332 -14728
rect 8268 -14872 8332 -14808
rect 8268 -14952 8332 -14888
rect 9680 -14232 9744 -14168
rect 9680 -14312 9744 -14248
rect 9680 -14392 9744 -14328
rect 9680 -14472 9744 -14408
rect 9680 -14552 9744 -14488
rect 9680 -14632 9744 -14568
rect 9680 -14712 9744 -14648
rect 9680 -14792 9744 -14728
rect 9680 -14872 9744 -14808
rect 9680 -14952 9744 -14888
rect 11092 -14232 11156 -14168
rect 11092 -14312 11156 -14248
rect 11092 -14392 11156 -14328
rect 11092 -14472 11156 -14408
rect 11092 -14552 11156 -14488
rect 11092 -14632 11156 -14568
rect 11092 -14712 11156 -14648
rect 11092 -14792 11156 -14728
rect 11092 -14872 11156 -14808
rect 11092 -14952 11156 -14888
rect 12504 -14232 12568 -14168
rect 12504 -14312 12568 -14248
rect 12504 -14392 12568 -14328
rect 12504 -14472 12568 -14408
rect 12504 -14552 12568 -14488
rect 12504 -14632 12568 -14568
rect 12504 -14712 12568 -14648
rect 12504 -14792 12568 -14728
rect 12504 -14872 12568 -14808
rect 12504 -14952 12568 -14888
rect 13916 -14232 13980 -14168
rect 13916 -14312 13980 -14248
rect 13916 -14392 13980 -14328
rect 13916 -14472 13980 -14408
rect 13916 -14552 13980 -14488
rect 13916 -14632 13980 -14568
rect 13916 -14712 13980 -14648
rect 13916 -14792 13980 -14728
rect 13916 -14872 13980 -14808
rect 13916 -14952 13980 -14888
rect 15328 -14232 15392 -14168
rect 15328 -14312 15392 -14248
rect 15328 -14392 15392 -14328
rect 15328 -14472 15392 -14408
rect 15328 -14552 15392 -14488
rect 15328 -14632 15392 -14568
rect 15328 -14712 15392 -14648
rect 15328 -14792 15392 -14728
rect 15328 -14872 15392 -14808
rect 15328 -14952 15392 -14888
rect 16740 -14232 16804 -14168
rect 16740 -14312 16804 -14248
rect 16740 -14392 16804 -14328
rect 16740 -14472 16804 -14408
rect 16740 -14552 16804 -14488
rect 16740 -14632 16804 -14568
rect 16740 -14712 16804 -14648
rect 16740 -14792 16804 -14728
rect 16740 -14872 16804 -14808
rect 16740 -14952 16804 -14888
rect 18152 -14232 18216 -14168
rect 18152 -14312 18216 -14248
rect 18152 -14392 18216 -14328
rect 18152 -14472 18216 -14408
rect 18152 -14552 18216 -14488
rect 18152 -14632 18216 -14568
rect 18152 -14712 18216 -14648
rect 18152 -14792 18216 -14728
rect 18152 -14872 18216 -14808
rect 18152 -14952 18216 -14888
rect 19564 -14232 19628 -14168
rect 19564 -14312 19628 -14248
rect 19564 -14392 19628 -14328
rect 19564 -14472 19628 -14408
rect 19564 -14552 19628 -14488
rect 19564 -14632 19628 -14568
rect 19564 -14712 19628 -14648
rect 19564 -14792 19628 -14728
rect 19564 -14872 19628 -14808
rect 19564 -14952 19628 -14888
rect 20976 -14232 21040 -14168
rect 20976 -14312 21040 -14248
rect 20976 -14392 21040 -14328
rect 20976 -14472 21040 -14408
rect 20976 -14552 21040 -14488
rect 20976 -14632 21040 -14568
rect 20976 -14712 21040 -14648
rect 20976 -14792 21040 -14728
rect 20976 -14872 21040 -14808
rect 20976 -14952 21040 -14888
rect 22388 -14232 22452 -14168
rect 22388 -14312 22452 -14248
rect 22388 -14392 22452 -14328
rect 22388 -14472 22452 -14408
rect 22388 -14552 22452 -14488
rect 22388 -14632 22452 -14568
rect 22388 -14712 22452 -14648
rect 22388 -14792 22452 -14728
rect 22388 -14872 22452 -14808
rect 22388 -14952 22452 -14888
rect 23800 -14232 23864 -14168
rect 23800 -14312 23864 -14248
rect 23800 -14392 23864 -14328
rect 23800 -14472 23864 -14408
rect 23800 -14552 23864 -14488
rect 23800 -14632 23864 -14568
rect 23800 -14712 23864 -14648
rect 23800 -14792 23864 -14728
rect 23800 -14872 23864 -14808
rect 23800 -14952 23864 -14888
rect -22796 -15352 -22732 -15288
rect -22796 -15432 -22732 -15368
rect -22796 -15512 -22732 -15448
rect -22796 -15592 -22732 -15528
rect -22796 -15672 -22732 -15608
rect -22796 -15752 -22732 -15688
rect -22796 -15832 -22732 -15768
rect -22796 -15912 -22732 -15848
rect -22796 -15992 -22732 -15928
rect -22796 -16072 -22732 -16008
rect -21384 -15352 -21320 -15288
rect -21384 -15432 -21320 -15368
rect -21384 -15512 -21320 -15448
rect -21384 -15592 -21320 -15528
rect -21384 -15672 -21320 -15608
rect -21384 -15752 -21320 -15688
rect -21384 -15832 -21320 -15768
rect -21384 -15912 -21320 -15848
rect -21384 -15992 -21320 -15928
rect -21384 -16072 -21320 -16008
rect -19972 -15352 -19908 -15288
rect -19972 -15432 -19908 -15368
rect -19972 -15512 -19908 -15448
rect -19972 -15592 -19908 -15528
rect -19972 -15672 -19908 -15608
rect -19972 -15752 -19908 -15688
rect -19972 -15832 -19908 -15768
rect -19972 -15912 -19908 -15848
rect -19972 -15992 -19908 -15928
rect -19972 -16072 -19908 -16008
rect -18560 -15352 -18496 -15288
rect -18560 -15432 -18496 -15368
rect -18560 -15512 -18496 -15448
rect -18560 -15592 -18496 -15528
rect -18560 -15672 -18496 -15608
rect -18560 -15752 -18496 -15688
rect -18560 -15832 -18496 -15768
rect -18560 -15912 -18496 -15848
rect -18560 -15992 -18496 -15928
rect -18560 -16072 -18496 -16008
rect -17148 -15352 -17084 -15288
rect -17148 -15432 -17084 -15368
rect -17148 -15512 -17084 -15448
rect -17148 -15592 -17084 -15528
rect -17148 -15672 -17084 -15608
rect -17148 -15752 -17084 -15688
rect -17148 -15832 -17084 -15768
rect -17148 -15912 -17084 -15848
rect -17148 -15992 -17084 -15928
rect -17148 -16072 -17084 -16008
rect -15736 -15352 -15672 -15288
rect -15736 -15432 -15672 -15368
rect -15736 -15512 -15672 -15448
rect -15736 -15592 -15672 -15528
rect -15736 -15672 -15672 -15608
rect -15736 -15752 -15672 -15688
rect -15736 -15832 -15672 -15768
rect -15736 -15912 -15672 -15848
rect -15736 -15992 -15672 -15928
rect -15736 -16072 -15672 -16008
rect -14324 -15352 -14260 -15288
rect -14324 -15432 -14260 -15368
rect -14324 -15512 -14260 -15448
rect -14324 -15592 -14260 -15528
rect -14324 -15672 -14260 -15608
rect -14324 -15752 -14260 -15688
rect -14324 -15832 -14260 -15768
rect -14324 -15912 -14260 -15848
rect -14324 -15992 -14260 -15928
rect -14324 -16072 -14260 -16008
rect -12912 -15352 -12848 -15288
rect -12912 -15432 -12848 -15368
rect -12912 -15512 -12848 -15448
rect -12912 -15592 -12848 -15528
rect -12912 -15672 -12848 -15608
rect -12912 -15752 -12848 -15688
rect -12912 -15832 -12848 -15768
rect -12912 -15912 -12848 -15848
rect -12912 -15992 -12848 -15928
rect -12912 -16072 -12848 -16008
rect -11500 -15352 -11436 -15288
rect -11500 -15432 -11436 -15368
rect -11500 -15512 -11436 -15448
rect -11500 -15592 -11436 -15528
rect -11500 -15672 -11436 -15608
rect -11500 -15752 -11436 -15688
rect -11500 -15832 -11436 -15768
rect -11500 -15912 -11436 -15848
rect -11500 -15992 -11436 -15928
rect -11500 -16072 -11436 -16008
rect -10088 -15352 -10024 -15288
rect -10088 -15432 -10024 -15368
rect -10088 -15512 -10024 -15448
rect -10088 -15592 -10024 -15528
rect -10088 -15672 -10024 -15608
rect -10088 -15752 -10024 -15688
rect -10088 -15832 -10024 -15768
rect -10088 -15912 -10024 -15848
rect -10088 -15992 -10024 -15928
rect -10088 -16072 -10024 -16008
rect -8676 -15352 -8612 -15288
rect -8676 -15432 -8612 -15368
rect -8676 -15512 -8612 -15448
rect -8676 -15592 -8612 -15528
rect -8676 -15672 -8612 -15608
rect -8676 -15752 -8612 -15688
rect -8676 -15832 -8612 -15768
rect -8676 -15912 -8612 -15848
rect -8676 -15992 -8612 -15928
rect -8676 -16072 -8612 -16008
rect -7264 -15352 -7200 -15288
rect -7264 -15432 -7200 -15368
rect -7264 -15512 -7200 -15448
rect -7264 -15592 -7200 -15528
rect -7264 -15672 -7200 -15608
rect -7264 -15752 -7200 -15688
rect -7264 -15832 -7200 -15768
rect -7264 -15912 -7200 -15848
rect -7264 -15992 -7200 -15928
rect -7264 -16072 -7200 -16008
rect -5852 -15352 -5788 -15288
rect -5852 -15432 -5788 -15368
rect -5852 -15512 -5788 -15448
rect -5852 -15592 -5788 -15528
rect -5852 -15672 -5788 -15608
rect -5852 -15752 -5788 -15688
rect -5852 -15832 -5788 -15768
rect -5852 -15912 -5788 -15848
rect -5852 -15992 -5788 -15928
rect -5852 -16072 -5788 -16008
rect -4440 -15352 -4376 -15288
rect -4440 -15432 -4376 -15368
rect -4440 -15512 -4376 -15448
rect -4440 -15592 -4376 -15528
rect -4440 -15672 -4376 -15608
rect -4440 -15752 -4376 -15688
rect -4440 -15832 -4376 -15768
rect -4440 -15912 -4376 -15848
rect -4440 -15992 -4376 -15928
rect -4440 -16072 -4376 -16008
rect -3028 -15352 -2964 -15288
rect -3028 -15432 -2964 -15368
rect -3028 -15512 -2964 -15448
rect -3028 -15592 -2964 -15528
rect -3028 -15672 -2964 -15608
rect -3028 -15752 -2964 -15688
rect -3028 -15832 -2964 -15768
rect -3028 -15912 -2964 -15848
rect -3028 -15992 -2964 -15928
rect -3028 -16072 -2964 -16008
rect -1616 -15352 -1552 -15288
rect -1616 -15432 -1552 -15368
rect -1616 -15512 -1552 -15448
rect -1616 -15592 -1552 -15528
rect -1616 -15672 -1552 -15608
rect -1616 -15752 -1552 -15688
rect -1616 -15832 -1552 -15768
rect -1616 -15912 -1552 -15848
rect -1616 -15992 -1552 -15928
rect -1616 -16072 -1552 -16008
rect -204 -15352 -140 -15288
rect -204 -15432 -140 -15368
rect -204 -15512 -140 -15448
rect -204 -15592 -140 -15528
rect -204 -15672 -140 -15608
rect -204 -15752 -140 -15688
rect -204 -15832 -140 -15768
rect -204 -15912 -140 -15848
rect -204 -15992 -140 -15928
rect -204 -16072 -140 -16008
rect 1208 -15352 1272 -15288
rect 1208 -15432 1272 -15368
rect 1208 -15512 1272 -15448
rect 1208 -15592 1272 -15528
rect 1208 -15672 1272 -15608
rect 1208 -15752 1272 -15688
rect 1208 -15832 1272 -15768
rect 1208 -15912 1272 -15848
rect 1208 -15992 1272 -15928
rect 1208 -16072 1272 -16008
rect 2620 -15352 2684 -15288
rect 2620 -15432 2684 -15368
rect 2620 -15512 2684 -15448
rect 2620 -15592 2684 -15528
rect 2620 -15672 2684 -15608
rect 2620 -15752 2684 -15688
rect 2620 -15832 2684 -15768
rect 2620 -15912 2684 -15848
rect 2620 -15992 2684 -15928
rect 2620 -16072 2684 -16008
rect 4032 -15352 4096 -15288
rect 4032 -15432 4096 -15368
rect 4032 -15512 4096 -15448
rect 4032 -15592 4096 -15528
rect 4032 -15672 4096 -15608
rect 4032 -15752 4096 -15688
rect 4032 -15832 4096 -15768
rect 4032 -15912 4096 -15848
rect 4032 -15992 4096 -15928
rect 4032 -16072 4096 -16008
rect 5444 -15352 5508 -15288
rect 5444 -15432 5508 -15368
rect 5444 -15512 5508 -15448
rect 5444 -15592 5508 -15528
rect 5444 -15672 5508 -15608
rect 5444 -15752 5508 -15688
rect 5444 -15832 5508 -15768
rect 5444 -15912 5508 -15848
rect 5444 -15992 5508 -15928
rect 5444 -16072 5508 -16008
rect 6856 -15352 6920 -15288
rect 6856 -15432 6920 -15368
rect 6856 -15512 6920 -15448
rect 6856 -15592 6920 -15528
rect 6856 -15672 6920 -15608
rect 6856 -15752 6920 -15688
rect 6856 -15832 6920 -15768
rect 6856 -15912 6920 -15848
rect 6856 -15992 6920 -15928
rect 6856 -16072 6920 -16008
rect 8268 -15352 8332 -15288
rect 8268 -15432 8332 -15368
rect 8268 -15512 8332 -15448
rect 8268 -15592 8332 -15528
rect 8268 -15672 8332 -15608
rect 8268 -15752 8332 -15688
rect 8268 -15832 8332 -15768
rect 8268 -15912 8332 -15848
rect 8268 -15992 8332 -15928
rect 8268 -16072 8332 -16008
rect 9680 -15352 9744 -15288
rect 9680 -15432 9744 -15368
rect 9680 -15512 9744 -15448
rect 9680 -15592 9744 -15528
rect 9680 -15672 9744 -15608
rect 9680 -15752 9744 -15688
rect 9680 -15832 9744 -15768
rect 9680 -15912 9744 -15848
rect 9680 -15992 9744 -15928
rect 9680 -16072 9744 -16008
rect 11092 -15352 11156 -15288
rect 11092 -15432 11156 -15368
rect 11092 -15512 11156 -15448
rect 11092 -15592 11156 -15528
rect 11092 -15672 11156 -15608
rect 11092 -15752 11156 -15688
rect 11092 -15832 11156 -15768
rect 11092 -15912 11156 -15848
rect 11092 -15992 11156 -15928
rect 11092 -16072 11156 -16008
rect 12504 -15352 12568 -15288
rect 12504 -15432 12568 -15368
rect 12504 -15512 12568 -15448
rect 12504 -15592 12568 -15528
rect 12504 -15672 12568 -15608
rect 12504 -15752 12568 -15688
rect 12504 -15832 12568 -15768
rect 12504 -15912 12568 -15848
rect 12504 -15992 12568 -15928
rect 12504 -16072 12568 -16008
rect 13916 -15352 13980 -15288
rect 13916 -15432 13980 -15368
rect 13916 -15512 13980 -15448
rect 13916 -15592 13980 -15528
rect 13916 -15672 13980 -15608
rect 13916 -15752 13980 -15688
rect 13916 -15832 13980 -15768
rect 13916 -15912 13980 -15848
rect 13916 -15992 13980 -15928
rect 13916 -16072 13980 -16008
rect 15328 -15352 15392 -15288
rect 15328 -15432 15392 -15368
rect 15328 -15512 15392 -15448
rect 15328 -15592 15392 -15528
rect 15328 -15672 15392 -15608
rect 15328 -15752 15392 -15688
rect 15328 -15832 15392 -15768
rect 15328 -15912 15392 -15848
rect 15328 -15992 15392 -15928
rect 15328 -16072 15392 -16008
rect 16740 -15352 16804 -15288
rect 16740 -15432 16804 -15368
rect 16740 -15512 16804 -15448
rect 16740 -15592 16804 -15528
rect 16740 -15672 16804 -15608
rect 16740 -15752 16804 -15688
rect 16740 -15832 16804 -15768
rect 16740 -15912 16804 -15848
rect 16740 -15992 16804 -15928
rect 16740 -16072 16804 -16008
rect 18152 -15352 18216 -15288
rect 18152 -15432 18216 -15368
rect 18152 -15512 18216 -15448
rect 18152 -15592 18216 -15528
rect 18152 -15672 18216 -15608
rect 18152 -15752 18216 -15688
rect 18152 -15832 18216 -15768
rect 18152 -15912 18216 -15848
rect 18152 -15992 18216 -15928
rect 18152 -16072 18216 -16008
rect 19564 -15352 19628 -15288
rect 19564 -15432 19628 -15368
rect 19564 -15512 19628 -15448
rect 19564 -15592 19628 -15528
rect 19564 -15672 19628 -15608
rect 19564 -15752 19628 -15688
rect 19564 -15832 19628 -15768
rect 19564 -15912 19628 -15848
rect 19564 -15992 19628 -15928
rect 19564 -16072 19628 -16008
rect 20976 -15352 21040 -15288
rect 20976 -15432 21040 -15368
rect 20976 -15512 21040 -15448
rect 20976 -15592 21040 -15528
rect 20976 -15672 21040 -15608
rect 20976 -15752 21040 -15688
rect 20976 -15832 21040 -15768
rect 20976 -15912 21040 -15848
rect 20976 -15992 21040 -15928
rect 20976 -16072 21040 -16008
rect 22388 -15352 22452 -15288
rect 22388 -15432 22452 -15368
rect 22388 -15512 22452 -15448
rect 22388 -15592 22452 -15528
rect 22388 -15672 22452 -15608
rect 22388 -15752 22452 -15688
rect 22388 -15832 22452 -15768
rect 22388 -15912 22452 -15848
rect 22388 -15992 22452 -15928
rect 22388 -16072 22452 -16008
rect 23800 -15352 23864 -15288
rect 23800 -15432 23864 -15368
rect 23800 -15512 23864 -15448
rect 23800 -15592 23864 -15528
rect 23800 -15672 23864 -15608
rect 23800 -15752 23864 -15688
rect 23800 -15832 23864 -15768
rect 23800 -15912 23864 -15848
rect 23800 -15992 23864 -15928
rect 23800 -16072 23864 -16008
rect -22796 -16472 -22732 -16408
rect -22796 -16552 -22732 -16488
rect -22796 -16632 -22732 -16568
rect -22796 -16712 -22732 -16648
rect -22796 -16792 -22732 -16728
rect -22796 -16872 -22732 -16808
rect -22796 -16952 -22732 -16888
rect -22796 -17032 -22732 -16968
rect -22796 -17112 -22732 -17048
rect -22796 -17192 -22732 -17128
rect -21384 -16472 -21320 -16408
rect -21384 -16552 -21320 -16488
rect -21384 -16632 -21320 -16568
rect -21384 -16712 -21320 -16648
rect -21384 -16792 -21320 -16728
rect -21384 -16872 -21320 -16808
rect -21384 -16952 -21320 -16888
rect -21384 -17032 -21320 -16968
rect -21384 -17112 -21320 -17048
rect -21384 -17192 -21320 -17128
rect -19972 -16472 -19908 -16408
rect -19972 -16552 -19908 -16488
rect -19972 -16632 -19908 -16568
rect -19972 -16712 -19908 -16648
rect -19972 -16792 -19908 -16728
rect -19972 -16872 -19908 -16808
rect -19972 -16952 -19908 -16888
rect -19972 -17032 -19908 -16968
rect -19972 -17112 -19908 -17048
rect -19972 -17192 -19908 -17128
rect -18560 -16472 -18496 -16408
rect -18560 -16552 -18496 -16488
rect -18560 -16632 -18496 -16568
rect -18560 -16712 -18496 -16648
rect -18560 -16792 -18496 -16728
rect -18560 -16872 -18496 -16808
rect -18560 -16952 -18496 -16888
rect -18560 -17032 -18496 -16968
rect -18560 -17112 -18496 -17048
rect -18560 -17192 -18496 -17128
rect -17148 -16472 -17084 -16408
rect -17148 -16552 -17084 -16488
rect -17148 -16632 -17084 -16568
rect -17148 -16712 -17084 -16648
rect -17148 -16792 -17084 -16728
rect -17148 -16872 -17084 -16808
rect -17148 -16952 -17084 -16888
rect -17148 -17032 -17084 -16968
rect -17148 -17112 -17084 -17048
rect -17148 -17192 -17084 -17128
rect -15736 -16472 -15672 -16408
rect -15736 -16552 -15672 -16488
rect -15736 -16632 -15672 -16568
rect -15736 -16712 -15672 -16648
rect -15736 -16792 -15672 -16728
rect -15736 -16872 -15672 -16808
rect -15736 -16952 -15672 -16888
rect -15736 -17032 -15672 -16968
rect -15736 -17112 -15672 -17048
rect -15736 -17192 -15672 -17128
rect -14324 -16472 -14260 -16408
rect -14324 -16552 -14260 -16488
rect -14324 -16632 -14260 -16568
rect -14324 -16712 -14260 -16648
rect -14324 -16792 -14260 -16728
rect -14324 -16872 -14260 -16808
rect -14324 -16952 -14260 -16888
rect -14324 -17032 -14260 -16968
rect -14324 -17112 -14260 -17048
rect -14324 -17192 -14260 -17128
rect -12912 -16472 -12848 -16408
rect -12912 -16552 -12848 -16488
rect -12912 -16632 -12848 -16568
rect -12912 -16712 -12848 -16648
rect -12912 -16792 -12848 -16728
rect -12912 -16872 -12848 -16808
rect -12912 -16952 -12848 -16888
rect -12912 -17032 -12848 -16968
rect -12912 -17112 -12848 -17048
rect -12912 -17192 -12848 -17128
rect -11500 -16472 -11436 -16408
rect -11500 -16552 -11436 -16488
rect -11500 -16632 -11436 -16568
rect -11500 -16712 -11436 -16648
rect -11500 -16792 -11436 -16728
rect -11500 -16872 -11436 -16808
rect -11500 -16952 -11436 -16888
rect -11500 -17032 -11436 -16968
rect -11500 -17112 -11436 -17048
rect -11500 -17192 -11436 -17128
rect -10088 -16472 -10024 -16408
rect -10088 -16552 -10024 -16488
rect -10088 -16632 -10024 -16568
rect -10088 -16712 -10024 -16648
rect -10088 -16792 -10024 -16728
rect -10088 -16872 -10024 -16808
rect -10088 -16952 -10024 -16888
rect -10088 -17032 -10024 -16968
rect -10088 -17112 -10024 -17048
rect -10088 -17192 -10024 -17128
rect -8676 -16472 -8612 -16408
rect -8676 -16552 -8612 -16488
rect -8676 -16632 -8612 -16568
rect -8676 -16712 -8612 -16648
rect -8676 -16792 -8612 -16728
rect -8676 -16872 -8612 -16808
rect -8676 -16952 -8612 -16888
rect -8676 -17032 -8612 -16968
rect -8676 -17112 -8612 -17048
rect -8676 -17192 -8612 -17128
rect -7264 -16472 -7200 -16408
rect -7264 -16552 -7200 -16488
rect -7264 -16632 -7200 -16568
rect -7264 -16712 -7200 -16648
rect -7264 -16792 -7200 -16728
rect -7264 -16872 -7200 -16808
rect -7264 -16952 -7200 -16888
rect -7264 -17032 -7200 -16968
rect -7264 -17112 -7200 -17048
rect -7264 -17192 -7200 -17128
rect -5852 -16472 -5788 -16408
rect -5852 -16552 -5788 -16488
rect -5852 -16632 -5788 -16568
rect -5852 -16712 -5788 -16648
rect -5852 -16792 -5788 -16728
rect -5852 -16872 -5788 -16808
rect -5852 -16952 -5788 -16888
rect -5852 -17032 -5788 -16968
rect -5852 -17112 -5788 -17048
rect -5852 -17192 -5788 -17128
rect -4440 -16472 -4376 -16408
rect -4440 -16552 -4376 -16488
rect -4440 -16632 -4376 -16568
rect -4440 -16712 -4376 -16648
rect -4440 -16792 -4376 -16728
rect -4440 -16872 -4376 -16808
rect -4440 -16952 -4376 -16888
rect -4440 -17032 -4376 -16968
rect -4440 -17112 -4376 -17048
rect -4440 -17192 -4376 -17128
rect -3028 -16472 -2964 -16408
rect -3028 -16552 -2964 -16488
rect -3028 -16632 -2964 -16568
rect -3028 -16712 -2964 -16648
rect -3028 -16792 -2964 -16728
rect -3028 -16872 -2964 -16808
rect -3028 -16952 -2964 -16888
rect -3028 -17032 -2964 -16968
rect -3028 -17112 -2964 -17048
rect -3028 -17192 -2964 -17128
rect -1616 -16472 -1552 -16408
rect -1616 -16552 -1552 -16488
rect -1616 -16632 -1552 -16568
rect -1616 -16712 -1552 -16648
rect -1616 -16792 -1552 -16728
rect -1616 -16872 -1552 -16808
rect -1616 -16952 -1552 -16888
rect -1616 -17032 -1552 -16968
rect -1616 -17112 -1552 -17048
rect -1616 -17192 -1552 -17128
rect -204 -16472 -140 -16408
rect -204 -16552 -140 -16488
rect -204 -16632 -140 -16568
rect -204 -16712 -140 -16648
rect -204 -16792 -140 -16728
rect -204 -16872 -140 -16808
rect -204 -16952 -140 -16888
rect -204 -17032 -140 -16968
rect -204 -17112 -140 -17048
rect -204 -17192 -140 -17128
rect 1208 -16472 1272 -16408
rect 1208 -16552 1272 -16488
rect 1208 -16632 1272 -16568
rect 1208 -16712 1272 -16648
rect 1208 -16792 1272 -16728
rect 1208 -16872 1272 -16808
rect 1208 -16952 1272 -16888
rect 1208 -17032 1272 -16968
rect 1208 -17112 1272 -17048
rect 1208 -17192 1272 -17128
rect 2620 -16472 2684 -16408
rect 2620 -16552 2684 -16488
rect 2620 -16632 2684 -16568
rect 2620 -16712 2684 -16648
rect 2620 -16792 2684 -16728
rect 2620 -16872 2684 -16808
rect 2620 -16952 2684 -16888
rect 2620 -17032 2684 -16968
rect 2620 -17112 2684 -17048
rect 2620 -17192 2684 -17128
rect 4032 -16472 4096 -16408
rect 4032 -16552 4096 -16488
rect 4032 -16632 4096 -16568
rect 4032 -16712 4096 -16648
rect 4032 -16792 4096 -16728
rect 4032 -16872 4096 -16808
rect 4032 -16952 4096 -16888
rect 4032 -17032 4096 -16968
rect 4032 -17112 4096 -17048
rect 4032 -17192 4096 -17128
rect 5444 -16472 5508 -16408
rect 5444 -16552 5508 -16488
rect 5444 -16632 5508 -16568
rect 5444 -16712 5508 -16648
rect 5444 -16792 5508 -16728
rect 5444 -16872 5508 -16808
rect 5444 -16952 5508 -16888
rect 5444 -17032 5508 -16968
rect 5444 -17112 5508 -17048
rect 5444 -17192 5508 -17128
rect 6856 -16472 6920 -16408
rect 6856 -16552 6920 -16488
rect 6856 -16632 6920 -16568
rect 6856 -16712 6920 -16648
rect 6856 -16792 6920 -16728
rect 6856 -16872 6920 -16808
rect 6856 -16952 6920 -16888
rect 6856 -17032 6920 -16968
rect 6856 -17112 6920 -17048
rect 6856 -17192 6920 -17128
rect 8268 -16472 8332 -16408
rect 8268 -16552 8332 -16488
rect 8268 -16632 8332 -16568
rect 8268 -16712 8332 -16648
rect 8268 -16792 8332 -16728
rect 8268 -16872 8332 -16808
rect 8268 -16952 8332 -16888
rect 8268 -17032 8332 -16968
rect 8268 -17112 8332 -17048
rect 8268 -17192 8332 -17128
rect 9680 -16472 9744 -16408
rect 9680 -16552 9744 -16488
rect 9680 -16632 9744 -16568
rect 9680 -16712 9744 -16648
rect 9680 -16792 9744 -16728
rect 9680 -16872 9744 -16808
rect 9680 -16952 9744 -16888
rect 9680 -17032 9744 -16968
rect 9680 -17112 9744 -17048
rect 9680 -17192 9744 -17128
rect 11092 -16472 11156 -16408
rect 11092 -16552 11156 -16488
rect 11092 -16632 11156 -16568
rect 11092 -16712 11156 -16648
rect 11092 -16792 11156 -16728
rect 11092 -16872 11156 -16808
rect 11092 -16952 11156 -16888
rect 11092 -17032 11156 -16968
rect 11092 -17112 11156 -17048
rect 11092 -17192 11156 -17128
rect 12504 -16472 12568 -16408
rect 12504 -16552 12568 -16488
rect 12504 -16632 12568 -16568
rect 12504 -16712 12568 -16648
rect 12504 -16792 12568 -16728
rect 12504 -16872 12568 -16808
rect 12504 -16952 12568 -16888
rect 12504 -17032 12568 -16968
rect 12504 -17112 12568 -17048
rect 12504 -17192 12568 -17128
rect 13916 -16472 13980 -16408
rect 13916 -16552 13980 -16488
rect 13916 -16632 13980 -16568
rect 13916 -16712 13980 -16648
rect 13916 -16792 13980 -16728
rect 13916 -16872 13980 -16808
rect 13916 -16952 13980 -16888
rect 13916 -17032 13980 -16968
rect 13916 -17112 13980 -17048
rect 13916 -17192 13980 -17128
rect 15328 -16472 15392 -16408
rect 15328 -16552 15392 -16488
rect 15328 -16632 15392 -16568
rect 15328 -16712 15392 -16648
rect 15328 -16792 15392 -16728
rect 15328 -16872 15392 -16808
rect 15328 -16952 15392 -16888
rect 15328 -17032 15392 -16968
rect 15328 -17112 15392 -17048
rect 15328 -17192 15392 -17128
rect 16740 -16472 16804 -16408
rect 16740 -16552 16804 -16488
rect 16740 -16632 16804 -16568
rect 16740 -16712 16804 -16648
rect 16740 -16792 16804 -16728
rect 16740 -16872 16804 -16808
rect 16740 -16952 16804 -16888
rect 16740 -17032 16804 -16968
rect 16740 -17112 16804 -17048
rect 16740 -17192 16804 -17128
rect 18152 -16472 18216 -16408
rect 18152 -16552 18216 -16488
rect 18152 -16632 18216 -16568
rect 18152 -16712 18216 -16648
rect 18152 -16792 18216 -16728
rect 18152 -16872 18216 -16808
rect 18152 -16952 18216 -16888
rect 18152 -17032 18216 -16968
rect 18152 -17112 18216 -17048
rect 18152 -17192 18216 -17128
rect 19564 -16472 19628 -16408
rect 19564 -16552 19628 -16488
rect 19564 -16632 19628 -16568
rect 19564 -16712 19628 -16648
rect 19564 -16792 19628 -16728
rect 19564 -16872 19628 -16808
rect 19564 -16952 19628 -16888
rect 19564 -17032 19628 -16968
rect 19564 -17112 19628 -17048
rect 19564 -17192 19628 -17128
rect 20976 -16472 21040 -16408
rect 20976 -16552 21040 -16488
rect 20976 -16632 21040 -16568
rect 20976 -16712 21040 -16648
rect 20976 -16792 21040 -16728
rect 20976 -16872 21040 -16808
rect 20976 -16952 21040 -16888
rect 20976 -17032 21040 -16968
rect 20976 -17112 21040 -17048
rect 20976 -17192 21040 -17128
rect 22388 -16472 22452 -16408
rect 22388 -16552 22452 -16488
rect 22388 -16632 22452 -16568
rect 22388 -16712 22452 -16648
rect 22388 -16792 22452 -16728
rect 22388 -16872 22452 -16808
rect 22388 -16952 22452 -16888
rect 22388 -17032 22452 -16968
rect 22388 -17112 22452 -17048
rect 22388 -17192 22452 -17128
rect 23800 -16472 23864 -16408
rect 23800 -16552 23864 -16488
rect 23800 -16632 23864 -16568
rect 23800 -16712 23864 -16648
rect 23800 -16792 23864 -16728
rect 23800 -16872 23864 -16808
rect 23800 -16952 23864 -16888
rect 23800 -17032 23864 -16968
rect 23800 -17112 23864 -17048
rect 23800 -17192 23864 -17128
rect -22796 -17592 -22732 -17528
rect -22796 -17672 -22732 -17608
rect -22796 -17752 -22732 -17688
rect -22796 -17832 -22732 -17768
rect -22796 -17912 -22732 -17848
rect -22796 -17992 -22732 -17928
rect -22796 -18072 -22732 -18008
rect -22796 -18152 -22732 -18088
rect -22796 -18232 -22732 -18168
rect -22796 -18312 -22732 -18248
rect -21384 -17592 -21320 -17528
rect -21384 -17672 -21320 -17608
rect -21384 -17752 -21320 -17688
rect -21384 -17832 -21320 -17768
rect -21384 -17912 -21320 -17848
rect -21384 -17992 -21320 -17928
rect -21384 -18072 -21320 -18008
rect -21384 -18152 -21320 -18088
rect -21384 -18232 -21320 -18168
rect -21384 -18312 -21320 -18248
rect -19972 -17592 -19908 -17528
rect -19972 -17672 -19908 -17608
rect -19972 -17752 -19908 -17688
rect -19972 -17832 -19908 -17768
rect -19972 -17912 -19908 -17848
rect -19972 -17992 -19908 -17928
rect -19972 -18072 -19908 -18008
rect -19972 -18152 -19908 -18088
rect -19972 -18232 -19908 -18168
rect -19972 -18312 -19908 -18248
rect -18560 -17592 -18496 -17528
rect -18560 -17672 -18496 -17608
rect -18560 -17752 -18496 -17688
rect -18560 -17832 -18496 -17768
rect -18560 -17912 -18496 -17848
rect -18560 -17992 -18496 -17928
rect -18560 -18072 -18496 -18008
rect -18560 -18152 -18496 -18088
rect -18560 -18232 -18496 -18168
rect -18560 -18312 -18496 -18248
rect -17148 -17592 -17084 -17528
rect -17148 -17672 -17084 -17608
rect -17148 -17752 -17084 -17688
rect -17148 -17832 -17084 -17768
rect -17148 -17912 -17084 -17848
rect -17148 -17992 -17084 -17928
rect -17148 -18072 -17084 -18008
rect -17148 -18152 -17084 -18088
rect -17148 -18232 -17084 -18168
rect -17148 -18312 -17084 -18248
rect -15736 -17592 -15672 -17528
rect -15736 -17672 -15672 -17608
rect -15736 -17752 -15672 -17688
rect -15736 -17832 -15672 -17768
rect -15736 -17912 -15672 -17848
rect -15736 -17992 -15672 -17928
rect -15736 -18072 -15672 -18008
rect -15736 -18152 -15672 -18088
rect -15736 -18232 -15672 -18168
rect -15736 -18312 -15672 -18248
rect -14324 -17592 -14260 -17528
rect -14324 -17672 -14260 -17608
rect -14324 -17752 -14260 -17688
rect -14324 -17832 -14260 -17768
rect -14324 -17912 -14260 -17848
rect -14324 -17992 -14260 -17928
rect -14324 -18072 -14260 -18008
rect -14324 -18152 -14260 -18088
rect -14324 -18232 -14260 -18168
rect -14324 -18312 -14260 -18248
rect -12912 -17592 -12848 -17528
rect -12912 -17672 -12848 -17608
rect -12912 -17752 -12848 -17688
rect -12912 -17832 -12848 -17768
rect -12912 -17912 -12848 -17848
rect -12912 -17992 -12848 -17928
rect -12912 -18072 -12848 -18008
rect -12912 -18152 -12848 -18088
rect -12912 -18232 -12848 -18168
rect -12912 -18312 -12848 -18248
rect -11500 -17592 -11436 -17528
rect -11500 -17672 -11436 -17608
rect -11500 -17752 -11436 -17688
rect -11500 -17832 -11436 -17768
rect -11500 -17912 -11436 -17848
rect -11500 -17992 -11436 -17928
rect -11500 -18072 -11436 -18008
rect -11500 -18152 -11436 -18088
rect -11500 -18232 -11436 -18168
rect -11500 -18312 -11436 -18248
rect -10088 -17592 -10024 -17528
rect -10088 -17672 -10024 -17608
rect -10088 -17752 -10024 -17688
rect -10088 -17832 -10024 -17768
rect -10088 -17912 -10024 -17848
rect -10088 -17992 -10024 -17928
rect -10088 -18072 -10024 -18008
rect -10088 -18152 -10024 -18088
rect -10088 -18232 -10024 -18168
rect -10088 -18312 -10024 -18248
rect -8676 -17592 -8612 -17528
rect -8676 -17672 -8612 -17608
rect -8676 -17752 -8612 -17688
rect -8676 -17832 -8612 -17768
rect -8676 -17912 -8612 -17848
rect -8676 -17992 -8612 -17928
rect -8676 -18072 -8612 -18008
rect -8676 -18152 -8612 -18088
rect -8676 -18232 -8612 -18168
rect -8676 -18312 -8612 -18248
rect -7264 -17592 -7200 -17528
rect -7264 -17672 -7200 -17608
rect -7264 -17752 -7200 -17688
rect -7264 -17832 -7200 -17768
rect -7264 -17912 -7200 -17848
rect -7264 -17992 -7200 -17928
rect -7264 -18072 -7200 -18008
rect -7264 -18152 -7200 -18088
rect -7264 -18232 -7200 -18168
rect -7264 -18312 -7200 -18248
rect -5852 -17592 -5788 -17528
rect -5852 -17672 -5788 -17608
rect -5852 -17752 -5788 -17688
rect -5852 -17832 -5788 -17768
rect -5852 -17912 -5788 -17848
rect -5852 -17992 -5788 -17928
rect -5852 -18072 -5788 -18008
rect -5852 -18152 -5788 -18088
rect -5852 -18232 -5788 -18168
rect -5852 -18312 -5788 -18248
rect -4440 -17592 -4376 -17528
rect -4440 -17672 -4376 -17608
rect -4440 -17752 -4376 -17688
rect -4440 -17832 -4376 -17768
rect -4440 -17912 -4376 -17848
rect -4440 -17992 -4376 -17928
rect -4440 -18072 -4376 -18008
rect -4440 -18152 -4376 -18088
rect -4440 -18232 -4376 -18168
rect -4440 -18312 -4376 -18248
rect -3028 -17592 -2964 -17528
rect -3028 -17672 -2964 -17608
rect -3028 -17752 -2964 -17688
rect -3028 -17832 -2964 -17768
rect -3028 -17912 -2964 -17848
rect -3028 -17992 -2964 -17928
rect -3028 -18072 -2964 -18008
rect -3028 -18152 -2964 -18088
rect -3028 -18232 -2964 -18168
rect -3028 -18312 -2964 -18248
rect -1616 -17592 -1552 -17528
rect -1616 -17672 -1552 -17608
rect -1616 -17752 -1552 -17688
rect -1616 -17832 -1552 -17768
rect -1616 -17912 -1552 -17848
rect -1616 -17992 -1552 -17928
rect -1616 -18072 -1552 -18008
rect -1616 -18152 -1552 -18088
rect -1616 -18232 -1552 -18168
rect -1616 -18312 -1552 -18248
rect -204 -17592 -140 -17528
rect -204 -17672 -140 -17608
rect -204 -17752 -140 -17688
rect -204 -17832 -140 -17768
rect -204 -17912 -140 -17848
rect -204 -17992 -140 -17928
rect -204 -18072 -140 -18008
rect -204 -18152 -140 -18088
rect -204 -18232 -140 -18168
rect -204 -18312 -140 -18248
rect 1208 -17592 1272 -17528
rect 1208 -17672 1272 -17608
rect 1208 -17752 1272 -17688
rect 1208 -17832 1272 -17768
rect 1208 -17912 1272 -17848
rect 1208 -17992 1272 -17928
rect 1208 -18072 1272 -18008
rect 1208 -18152 1272 -18088
rect 1208 -18232 1272 -18168
rect 1208 -18312 1272 -18248
rect 2620 -17592 2684 -17528
rect 2620 -17672 2684 -17608
rect 2620 -17752 2684 -17688
rect 2620 -17832 2684 -17768
rect 2620 -17912 2684 -17848
rect 2620 -17992 2684 -17928
rect 2620 -18072 2684 -18008
rect 2620 -18152 2684 -18088
rect 2620 -18232 2684 -18168
rect 2620 -18312 2684 -18248
rect 4032 -17592 4096 -17528
rect 4032 -17672 4096 -17608
rect 4032 -17752 4096 -17688
rect 4032 -17832 4096 -17768
rect 4032 -17912 4096 -17848
rect 4032 -17992 4096 -17928
rect 4032 -18072 4096 -18008
rect 4032 -18152 4096 -18088
rect 4032 -18232 4096 -18168
rect 4032 -18312 4096 -18248
rect 5444 -17592 5508 -17528
rect 5444 -17672 5508 -17608
rect 5444 -17752 5508 -17688
rect 5444 -17832 5508 -17768
rect 5444 -17912 5508 -17848
rect 5444 -17992 5508 -17928
rect 5444 -18072 5508 -18008
rect 5444 -18152 5508 -18088
rect 5444 -18232 5508 -18168
rect 5444 -18312 5508 -18248
rect 6856 -17592 6920 -17528
rect 6856 -17672 6920 -17608
rect 6856 -17752 6920 -17688
rect 6856 -17832 6920 -17768
rect 6856 -17912 6920 -17848
rect 6856 -17992 6920 -17928
rect 6856 -18072 6920 -18008
rect 6856 -18152 6920 -18088
rect 6856 -18232 6920 -18168
rect 6856 -18312 6920 -18248
rect 8268 -17592 8332 -17528
rect 8268 -17672 8332 -17608
rect 8268 -17752 8332 -17688
rect 8268 -17832 8332 -17768
rect 8268 -17912 8332 -17848
rect 8268 -17992 8332 -17928
rect 8268 -18072 8332 -18008
rect 8268 -18152 8332 -18088
rect 8268 -18232 8332 -18168
rect 8268 -18312 8332 -18248
rect 9680 -17592 9744 -17528
rect 9680 -17672 9744 -17608
rect 9680 -17752 9744 -17688
rect 9680 -17832 9744 -17768
rect 9680 -17912 9744 -17848
rect 9680 -17992 9744 -17928
rect 9680 -18072 9744 -18008
rect 9680 -18152 9744 -18088
rect 9680 -18232 9744 -18168
rect 9680 -18312 9744 -18248
rect 11092 -17592 11156 -17528
rect 11092 -17672 11156 -17608
rect 11092 -17752 11156 -17688
rect 11092 -17832 11156 -17768
rect 11092 -17912 11156 -17848
rect 11092 -17992 11156 -17928
rect 11092 -18072 11156 -18008
rect 11092 -18152 11156 -18088
rect 11092 -18232 11156 -18168
rect 11092 -18312 11156 -18248
rect 12504 -17592 12568 -17528
rect 12504 -17672 12568 -17608
rect 12504 -17752 12568 -17688
rect 12504 -17832 12568 -17768
rect 12504 -17912 12568 -17848
rect 12504 -17992 12568 -17928
rect 12504 -18072 12568 -18008
rect 12504 -18152 12568 -18088
rect 12504 -18232 12568 -18168
rect 12504 -18312 12568 -18248
rect 13916 -17592 13980 -17528
rect 13916 -17672 13980 -17608
rect 13916 -17752 13980 -17688
rect 13916 -17832 13980 -17768
rect 13916 -17912 13980 -17848
rect 13916 -17992 13980 -17928
rect 13916 -18072 13980 -18008
rect 13916 -18152 13980 -18088
rect 13916 -18232 13980 -18168
rect 13916 -18312 13980 -18248
rect 15328 -17592 15392 -17528
rect 15328 -17672 15392 -17608
rect 15328 -17752 15392 -17688
rect 15328 -17832 15392 -17768
rect 15328 -17912 15392 -17848
rect 15328 -17992 15392 -17928
rect 15328 -18072 15392 -18008
rect 15328 -18152 15392 -18088
rect 15328 -18232 15392 -18168
rect 15328 -18312 15392 -18248
rect 16740 -17592 16804 -17528
rect 16740 -17672 16804 -17608
rect 16740 -17752 16804 -17688
rect 16740 -17832 16804 -17768
rect 16740 -17912 16804 -17848
rect 16740 -17992 16804 -17928
rect 16740 -18072 16804 -18008
rect 16740 -18152 16804 -18088
rect 16740 -18232 16804 -18168
rect 16740 -18312 16804 -18248
rect 18152 -17592 18216 -17528
rect 18152 -17672 18216 -17608
rect 18152 -17752 18216 -17688
rect 18152 -17832 18216 -17768
rect 18152 -17912 18216 -17848
rect 18152 -17992 18216 -17928
rect 18152 -18072 18216 -18008
rect 18152 -18152 18216 -18088
rect 18152 -18232 18216 -18168
rect 18152 -18312 18216 -18248
rect 19564 -17592 19628 -17528
rect 19564 -17672 19628 -17608
rect 19564 -17752 19628 -17688
rect 19564 -17832 19628 -17768
rect 19564 -17912 19628 -17848
rect 19564 -17992 19628 -17928
rect 19564 -18072 19628 -18008
rect 19564 -18152 19628 -18088
rect 19564 -18232 19628 -18168
rect 19564 -18312 19628 -18248
rect 20976 -17592 21040 -17528
rect 20976 -17672 21040 -17608
rect 20976 -17752 21040 -17688
rect 20976 -17832 21040 -17768
rect 20976 -17912 21040 -17848
rect 20976 -17992 21040 -17928
rect 20976 -18072 21040 -18008
rect 20976 -18152 21040 -18088
rect 20976 -18232 21040 -18168
rect 20976 -18312 21040 -18248
rect 22388 -17592 22452 -17528
rect 22388 -17672 22452 -17608
rect 22388 -17752 22452 -17688
rect 22388 -17832 22452 -17768
rect 22388 -17912 22452 -17848
rect 22388 -17992 22452 -17928
rect 22388 -18072 22452 -18008
rect 22388 -18152 22452 -18088
rect 22388 -18232 22452 -18168
rect 22388 -18312 22452 -18248
rect 23800 -17592 23864 -17528
rect 23800 -17672 23864 -17608
rect 23800 -17752 23864 -17688
rect 23800 -17832 23864 -17768
rect 23800 -17912 23864 -17848
rect 23800 -17992 23864 -17928
rect 23800 -18072 23864 -18008
rect 23800 -18152 23864 -18088
rect 23800 -18232 23864 -18168
rect 23800 -18312 23864 -18248
<< mimcap >>
rect -23844 18272 -23044 18320
rect -23844 17568 -23796 18272
rect -23092 17568 -23044 18272
rect -23844 17520 -23044 17568
rect -22432 18272 -21632 18320
rect -22432 17568 -22384 18272
rect -21680 17568 -21632 18272
rect -22432 17520 -21632 17568
rect -21020 18272 -20220 18320
rect -21020 17568 -20972 18272
rect -20268 17568 -20220 18272
rect -21020 17520 -20220 17568
rect -19608 18272 -18808 18320
rect -19608 17568 -19560 18272
rect -18856 17568 -18808 18272
rect -19608 17520 -18808 17568
rect -18196 18272 -17396 18320
rect -18196 17568 -18148 18272
rect -17444 17568 -17396 18272
rect -18196 17520 -17396 17568
rect -16784 18272 -15984 18320
rect -16784 17568 -16736 18272
rect -16032 17568 -15984 18272
rect -16784 17520 -15984 17568
rect -15372 18272 -14572 18320
rect -15372 17568 -15324 18272
rect -14620 17568 -14572 18272
rect -15372 17520 -14572 17568
rect -13960 18272 -13160 18320
rect -13960 17568 -13912 18272
rect -13208 17568 -13160 18272
rect -13960 17520 -13160 17568
rect -12548 18272 -11748 18320
rect -12548 17568 -12500 18272
rect -11796 17568 -11748 18272
rect -12548 17520 -11748 17568
rect -11136 18272 -10336 18320
rect -11136 17568 -11088 18272
rect -10384 17568 -10336 18272
rect -11136 17520 -10336 17568
rect -9724 18272 -8924 18320
rect -9724 17568 -9676 18272
rect -8972 17568 -8924 18272
rect -9724 17520 -8924 17568
rect -8312 18272 -7512 18320
rect -8312 17568 -8264 18272
rect -7560 17568 -7512 18272
rect -8312 17520 -7512 17568
rect -6900 18272 -6100 18320
rect -6900 17568 -6852 18272
rect -6148 17568 -6100 18272
rect -6900 17520 -6100 17568
rect -5488 18272 -4688 18320
rect -5488 17568 -5440 18272
rect -4736 17568 -4688 18272
rect -5488 17520 -4688 17568
rect -4076 18272 -3276 18320
rect -4076 17568 -4028 18272
rect -3324 17568 -3276 18272
rect -4076 17520 -3276 17568
rect -2664 18272 -1864 18320
rect -2664 17568 -2616 18272
rect -1912 17568 -1864 18272
rect -2664 17520 -1864 17568
rect -1252 18272 -452 18320
rect -1252 17568 -1204 18272
rect -500 17568 -452 18272
rect -1252 17520 -452 17568
rect 160 18272 960 18320
rect 160 17568 208 18272
rect 912 17568 960 18272
rect 160 17520 960 17568
rect 1572 18272 2372 18320
rect 1572 17568 1620 18272
rect 2324 17568 2372 18272
rect 1572 17520 2372 17568
rect 2984 18272 3784 18320
rect 2984 17568 3032 18272
rect 3736 17568 3784 18272
rect 2984 17520 3784 17568
rect 4396 18272 5196 18320
rect 4396 17568 4444 18272
rect 5148 17568 5196 18272
rect 4396 17520 5196 17568
rect 5808 18272 6608 18320
rect 5808 17568 5856 18272
rect 6560 17568 6608 18272
rect 5808 17520 6608 17568
rect 7220 18272 8020 18320
rect 7220 17568 7268 18272
rect 7972 17568 8020 18272
rect 7220 17520 8020 17568
rect 8632 18272 9432 18320
rect 8632 17568 8680 18272
rect 9384 17568 9432 18272
rect 8632 17520 9432 17568
rect 10044 18272 10844 18320
rect 10044 17568 10092 18272
rect 10796 17568 10844 18272
rect 10044 17520 10844 17568
rect 11456 18272 12256 18320
rect 11456 17568 11504 18272
rect 12208 17568 12256 18272
rect 11456 17520 12256 17568
rect 12868 18272 13668 18320
rect 12868 17568 12916 18272
rect 13620 17568 13668 18272
rect 12868 17520 13668 17568
rect 14280 18272 15080 18320
rect 14280 17568 14328 18272
rect 15032 17568 15080 18272
rect 14280 17520 15080 17568
rect 15692 18272 16492 18320
rect 15692 17568 15740 18272
rect 16444 17568 16492 18272
rect 15692 17520 16492 17568
rect 17104 18272 17904 18320
rect 17104 17568 17152 18272
rect 17856 17568 17904 18272
rect 17104 17520 17904 17568
rect 18516 18272 19316 18320
rect 18516 17568 18564 18272
rect 19268 17568 19316 18272
rect 18516 17520 19316 17568
rect 19928 18272 20728 18320
rect 19928 17568 19976 18272
rect 20680 17568 20728 18272
rect 19928 17520 20728 17568
rect 21340 18272 22140 18320
rect 21340 17568 21388 18272
rect 22092 17568 22140 18272
rect 21340 17520 22140 17568
rect 22752 18272 23552 18320
rect 22752 17568 22800 18272
rect 23504 17568 23552 18272
rect 22752 17520 23552 17568
rect -23844 17152 -23044 17200
rect -23844 16448 -23796 17152
rect -23092 16448 -23044 17152
rect -23844 16400 -23044 16448
rect -22432 17152 -21632 17200
rect -22432 16448 -22384 17152
rect -21680 16448 -21632 17152
rect -22432 16400 -21632 16448
rect -21020 17152 -20220 17200
rect -21020 16448 -20972 17152
rect -20268 16448 -20220 17152
rect -21020 16400 -20220 16448
rect -19608 17152 -18808 17200
rect -19608 16448 -19560 17152
rect -18856 16448 -18808 17152
rect -19608 16400 -18808 16448
rect -18196 17152 -17396 17200
rect -18196 16448 -18148 17152
rect -17444 16448 -17396 17152
rect -18196 16400 -17396 16448
rect -16784 17152 -15984 17200
rect -16784 16448 -16736 17152
rect -16032 16448 -15984 17152
rect -16784 16400 -15984 16448
rect -15372 17152 -14572 17200
rect -15372 16448 -15324 17152
rect -14620 16448 -14572 17152
rect -15372 16400 -14572 16448
rect -13960 17152 -13160 17200
rect -13960 16448 -13912 17152
rect -13208 16448 -13160 17152
rect -13960 16400 -13160 16448
rect -12548 17152 -11748 17200
rect -12548 16448 -12500 17152
rect -11796 16448 -11748 17152
rect -12548 16400 -11748 16448
rect -11136 17152 -10336 17200
rect -11136 16448 -11088 17152
rect -10384 16448 -10336 17152
rect -11136 16400 -10336 16448
rect -9724 17152 -8924 17200
rect -9724 16448 -9676 17152
rect -8972 16448 -8924 17152
rect -9724 16400 -8924 16448
rect -8312 17152 -7512 17200
rect -8312 16448 -8264 17152
rect -7560 16448 -7512 17152
rect -8312 16400 -7512 16448
rect -6900 17152 -6100 17200
rect -6900 16448 -6852 17152
rect -6148 16448 -6100 17152
rect -6900 16400 -6100 16448
rect -5488 17152 -4688 17200
rect -5488 16448 -5440 17152
rect -4736 16448 -4688 17152
rect -5488 16400 -4688 16448
rect -4076 17152 -3276 17200
rect -4076 16448 -4028 17152
rect -3324 16448 -3276 17152
rect -4076 16400 -3276 16448
rect -2664 17152 -1864 17200
rect -2664 16448 -2616 17152
rect -1912 16448 -1864 17152
rect -2664 16400 -1864 16448
rect -1252 17152 -452 17200
rect -1252 16448 -1204 17152
rect -500 16448 -452 17152
rect -1252 16400 -452 16448
rect 160 17152 960 17200
rect 160 16448 208 17152
rect 912 16448 960 17152
rect 160 16400 960 16448
rect 1572 17152 2372 17200
rect 1572 16448 1620 17152
rect 2324 16448 2372 17152
rect 1572 16400 2372 16448
rect 2984 17152 3784 17200
rect 2984 16448 3032 17152
rect 3736 16448 3784 17152
rect 2984 16400 3784 16448
rect 4396 17152 5196 17200
rect 4396 16448 4444 17152
rect 5148 16448 5196 17152
rect 4396 16400 5196 16448
rect 5808 17152 6608 17200
rect 5808 16448 5856 17152
rect 6560 16448 6608 17152
rect 5808 16400 6608 16448
rect 7220 17152 8020 17200
rect 7220 16448 7268 17152
rect 7972 16448 8020 17152
rect 7220 16400 8020 16448
rect 8632 17152 9432 17200
rect 8632 16448 8680 17152
rect 9384 16448 9432 17152
rect 8632 16400 9432 16448
rect 10044 17152 10844 17200
rect 10044 16448 10092 17152
rect 10796 16448 10844 17152
rect 10044 16400 10844 16448
rect 11456 17152 12256 17200
rect 11456 16448 11504 17152
rect 12208 16448 12256 17152
rect 11456 16400 12256 16448
rect 12868 17152 13668 17200
rect 12868 16448 12916 17152
rect 13620 16448 13668 17152
rect 12868 16400 13668 16448
rect 14280 17152 15080 17200
rect 14280 16448 14328 17152
rect 15032 16448 15080 17152
rect 14280 16400 15080 16448
rect 15692 17152 16492 17200
rect 15692 16448 15740 17152
rect 16444 16448 16492 17152
rect 15692 16400 16492 16448
rect 17104 17152 17904 17200
rect 17104 16448 17152 17152
rect 17856 16448 17904 17152
rect 17104 16400 17904 16448
rect 18516 17152 19316 17200
rect 18516 16448 18564 17152
rect 19268 16448 19316 17152
rect 18516 16400 19316 16448
rect 19928 17152 20728 17200
rect 19928 16448 19976 17152
rect 20680 16448 20728 17152
rect 19928 16400 20728 16448
rect 21340 17152 22140 17200
rect 21340 16448 21388 17152
rect 22092 16448 22140 17152
rect 21340 16400 22140 16448
rect 22752 17152 23552 17200
rect 22752 16448 22800 17152
rect 23504 16448 23552 17152
rect 22752 16400 23552 16448
rect -23844 16032 -23044 16080
rect -23844 15328 -23796 16032
rect -23092 15328 -23044 16032
rect -23844 15280 -23044 15328
rect -22432 16032 -21632 16080
rect -22432 15328 -22384 16032
rect -21680 15328 -21632 16032
rect -22432 15280 -21632 15328
rect -21020 16032 -20220 16080
rect -21020 15328 -20972 16032
rect -20268 15328 -20220 16032
rect -21020 15280 -20220 15328
rect -19608 16032 -18808 16080
rect -19608 15328 -19560 16032
rect -18856 15328 -18808 16032
rect -19608 15280 -18808 15328
rect -18196 16032 -17396 16080
rect -18196 15328 -18148 16032
rect -17444 15328 -17396 16032
rect -18196 15280 -17396 15328
rect -16784 16032 -15984 16080
rect -16784 15328 -16736 16032
rect -16032 15328 -15984 16032
rect -16784 15280 -15984 15328
rect -15372 16032 -14572 16080
rect -15372 15328 -15324 16032
rect -14620 15328 -14572 16032
rect -15372 15280 -14572 15328
rect -13960 16032 -13160 16080
rect -13960 15328 -13912 16032
rect -13208 15328 -13160 16032
rect -13960 15280 -13160 15328
rect -12548 16032 -11748 16080
rect -12548 15328 -12500 16032
rect -11796 15328 -11748 16032
rect -12548 15280 -11748 15328
rect -11136 16032 -10336 16080
rect -11136 15328 -11088 16032
rect -10384 15328 -10336 16032
rect -11136 15280 -10336 15328
rect -9724 16032 -8924 16080
rect -9724 15328 -9676 16032
rect -8972 15328 -8924 16032
rect -9724 15280 -8924 15328
rect -8312 16032 -7512 16080
rect -8312 15328 -8264 16032
rect -7560 15328 -7512 16032
rect -8312 15280 -7512 15328
rect -6900 16032 -6100 16080
rect -6900 15328 -6852 16032
rect -6148 15328 -6100 16032
rect -6900 15280 -6100 15328
rect -5488 16032 -4688 16080
rect -5488 15328 -5440 16032
rect -4736 15328 -4688 16032
rect -5488 15280 -4688 15328
rect -4076 16032 -3276 16080
rect -4076 15328 -4028 16032
rect -3324 15328 -3276 16032
rect -4076 15280 -3276 15328
rect -2664 16032 -1864 16080
rect -2664 15328 -2616 16032
rect -1912 15328 -1864 16032
rect -2664 15280 -1864 15328
rect -1252 16032 -452 16080
rect -1252 15328 -1204 16032
rect -500 15328 -452 16032
rect -1252 15280 -452 15328
rect 160 16032 960 16080
rect 160 15328 208 16032
rect 912 15328 960 16032
rect 160 15280 960 15328
rect 1572 16032 2372 16080
rect 1572 15328 1620 16032
rect 2324 15328 2372 16032
rect 1572 15280 2372 15328
rect 2984 16032 3784 16080
rect 2984 15328 3032 16032
rect 3736 15328 3784 16032
rect 2984 15280 3784 15328
rect 4396 16032 5196 16080
rect 4396 15328 4444 16032
rect 5148 15328 5196 16032
rect 4396 15280 5196 15328
rect 5808 16032 6608 16080
rect 5808 15328 5856 16032
rect 6560 15328 6608 16032
rect 5808 15280 6608 15328
rect 7220 16032 8020 16080
rect 7220 15328 7268 16032
rect 7972 15328 8020 16032
rect 7220 15280 8020 15328
rect 8632 16032 9432 16080
rect 8632 15328 8680 16032
rect 9384 15328 9432 16032
rect 8632 15280 9432 15328
rect 10044 16032 10844 16080
rect 10044 15328 10092 16032
rect 10796 15328 10844 16032
rect 10044 15280 10844 15328
rect 11456 16032 12256 16080
rect 11456 15328 11504 16032
rect 12208 15328 12256 16032
rect 11456 15280 12256 15328
rect 12868 16032 13668 16080
rect 12868 15328 12916 16032
rect 13620 15328 13668 16032
rect 12868 15280 13668 15328
rect 14280 16032 15080 16080
rect 14280 15328 14328 16032
rect 15032 15328 15080 16032
rect 14280 15280 15080 15328
rect 15692 16032 16492 16080
rect 15692 15328 15740 16032
rect 16444 15328 16492 16032
rect 15692 15280 16492 15328
rect 17104 16032 17904 16080
rect 17104 15328 17152 16032
rect 17856 15328 17904 16032
rect 17104 15280 17904 15328
rect 18516 16032 19316 16080
rect 18516 15328 18564 16032
rect 19268 15328 19316 16032
rect 18516 15280 19316 15328
rect 19928 16032 20728 16080
rect 19928 15328 19976 16032
rect 20680 15328 20728 16032
rect 19928 15280 20728 15328
rect 21340 16032 22140 16080
rect 21340 15328 21388 16032
rect 22092 15328 22140 16032
rect 21340 15280 22140 15328
rect 22752 16032 23552 16080
rect 22752 15328 22800 16032
rect 23504 15328 23552 16032
rect 22752 15280 23552 15328
rect -23844 14912 -23044 14960
rect -23844 14208 -23796 14912
rect -23092 14208 -23044 14912
rect -23844 14160 -23044 14208
rect -22432 14912 -21632 14960
rect -22432 14208 -22384 14912
rect -21680 14208 -21632 14912
rect -22432 14160 -21632 14208
rect -21020 14912 -20220 14960
rect -21020 14208 -20972 14912
rect -20268 14208 -20220 14912
rect -21020 14160 -20220 14208
rect -19608 14912 -18808 14960
rect -19608 14208 -19560 14912
rect -18856 14208 -18808 14912
rect -19608 14160 -18808 14208
rect -18196 14912 -17396 14960
rect -18196 14208 -18148 14912
rect -17444 14208 -17396 14912
rect -18196 14160 -17396 14208
rect -16784 14912 -15984 14960
rect -16784 14208 -16736 14912
rect -16032 14208 -15984 14912
rect -16784 14160 -15984 14208
rect -15372 14912 -14572 14960
rect -15372 14208 -15324 14912
rect -14620 14208 -14572 14912
rect -15372 14160 -14572 14208
rect -13960 14912 -13160 14960
rect -13960 14208 -13912 14912
rect -13208 14208 -13160 14912
rect -13960 14160 -13160 14208
rect -12548 14912 -11748 14960
rect -12548 14208 -12500 14912
rect -11796 14208 -11748 14912
rect -12548 14160 -11748 14208
rect -11136 14912 -10336 14960
rect -11136 14208 -11088 14912
rect -10384 14208 -10336 14912
rect -11136 14160 -10336 14208
rect -9724 14912 -8924 14960
rect -9724 14208 -9676 14912
rect -8972 14208 -8924 14912
rect -9724 14160 -8924 14208
rect -8312 14912 -7512 14960
rect -8312 14208 -8264 14912
rect -7560 14208 -7512 14912
rect -8312 14160 -7512 14208
rect -6900 14912 -6100 14960
rect -6900 14208 -6852 14912
rect -6148 14208 -6100 14912
rect -6900 14160 -6100 14208
rect -5488 14912 -4688 14960
rect -5488 14208 -5440 14912
rect -4736 14208 -4688 14912
rect -5488 14160 -4688 14208
rect -4076 14912 -3276 14960
rect -4076 14208 -4028 14912
rect -3324 14208 -3276 14912
rect -4076 14160 -3276 14208
rect -2664 14912 -1864 14960
rect -2664 14208 -2616 14912
rect -1912 14208 -1864 14912
rect -2664 14160 -1864 14208
rect -1252 14912 -452 14960
rect -1252 14208 -1204 14912
rect -500 14208 -452 14912
rect -1252 14160 -452 14208
rect 160 14912 960 14960
rect 160 14208 208 14912
rect 912 14208 960 14912
rect 160 14160 960 14208
rect 1572 14912 2372 14960
rect 1572 14208 1620 14912
rect 2324 14208 2372 14912
rect 1572 14160 2372 14208
rect 2984 14912 3784 14960
rect 2984 14208 3032 14912
rect 3736 14208 3784 14912
rect 2984 14160 3784 14208
rect 4396 14912 5196 14960
rect 4396 14208 4444 14912
rect 5148 14208 5196 14912
rect 4396 14160 5196 14208
rect 5808 14912 6608 14960
rect 5808 14208 5856 14912
rect 6560 14208 6608 14912
rect 5808 14160 6608 14208
rect 7220 14912 8020 14960
rect 7220 14208 7268 14912
rect 7972 14208 8020 14912
rect 7220 14160 8020 14208
rect 8632 14912 9432 14960
rect 8632 14208 8680 14912
rect 9384 14208 9432 14912
rect 8632 14160 9432 14208
rect 10044 14912 10844 14960
rect 10044 14208 10092 14912
rect 10796 14208 10844 14912
rect 10044 14160 10844 14208
rect 11456 14912 12256 14960
rect 11456 14208 11504 14912
rect 12208 14208 12256 14912
rect 11456 14160 12256 14208
rect 12868 14912 13668 14960
rect 12868 14208 12916 14912
rect 13620 14208 13668 14912
rect 12868 14160 13668 14208
rect 14280 14912 15080 14960
rect 14280 14208 14328 14912
rect 15032 14208 15080 14912
rect 14280 14160 15080 14208
rect 15692 14912 16492 14960
rect 15692 14208 15740 14912
rect 16444 14208 16492 14912
rect 15692 14160 16492 14208
rect 17104 14912 17904 14960
rect 17104 14208 17152 14912
rect 17856 14208 17904 14912
rect 17104 14160 17904 14208
rect 18516 14912 19316 14960
rect 18516 14208 18564 14912
rect 19268 14208 19316 14912
rect 18516 14160 19316 14208
rect 19928 14912 20728 14960
rect 19928 14208 19976 14912
rect 20680 14208 20728 14912
rect 19928 14160 20728 14208
rect 21340 14912 22140 14960
rect 21340 14208 21388 14912
rect 22092 14208 22140 14912
rect 21340 14160 22140 14208
rect 22752 14912 23552 14960
rect 22752 14208 22800 14912
rect 23504 14208 23552 14912
rect 22752 14160 23552 14208
rect -23844 13792 -23044 13840
rect -23844 13088 -23796 13792
rect -23092 13088 -23044 13792
rect -23844 13040 -23044 13088
rect -22432 13792 -21632 13840
rect -22432 13088 -22384 13792
rect -21680 13088 -21632 13792
rect -22432 13040 -21632 13088
rect -21020 13792 -20220 13840
rect -21020 13088 -20972 13792
rect -20268 13088 -20220 13792
rect -21020 13040 -20220 13088
rect -19608 13792 -18808 13840
rect -19608 13088 -19560 13792
rect -18856 13088 -18808 13792
rect -19608 13040 -18808 13088
rect -18196 13792 -17396 13840
rect -18196 13088 -18148 13792
rect -17444 13088 -17396 13792
rect -18196 13040 -17396 13088
rect -16784 13792 -15984 13840
rect -16784 13088 -16736 13792
rect -16032 13088 -15984 13792
rect -16784 13040 -15984 13088
rect -15372 13792 -14572 13840
rect -15372 13088 -15324 13792
rect -14620 13088 -14572 13792
rect -15372 13040 -14572 13088
rect -13960 13792 -13160 13840
rect -13960 13088 -13912 13792
rect -13208 13088 -13160 13792
rect -13960 13040 -13160 13088
rect -12548 13792 -11748 13840
rect -12548 13088 -12500 13792
rect -11796 13088 -11748 13792
rect -12548 13040 -11748 13088
rect -11136 13792 -10336 13840
rect -11136 13088 -11088 13792
rect -10384 13088 -10336 13792
rect -11136 13040 -10336 13088
rect -9724 13792 -8924 13840
rect -9724 13088 -9676 13792
rect -8972 13088 -8924 13792
rect -9724 13040 -8924 13088
rect -8312 13792 -7512 13840
rect -8312 13088 -8264 13792
rect -7560 13088 -7512 13792
rect -8312 13040 -7512 13088
rect -6900 13792 -6100 13840
rect -6900 13088 -6852 13792
rect -6148 13088 -6100 13792
rect -6900 13040 -6100 13088
rect -5488 13792 -4688 13840
rect -5488 13088 -5440 13792
rect -4736 13088 -4688 13792
rect -5488 13040 -4688 13088
rect -4076 13792 -3276 13840
rect -4076 13088 -4028 13792
rect -3324 13088 -3276 13792
rect -4076 13040 -3276 13088
rect -2664 13792 -1864 13840
rect -2664 13088 -2616 13792
rect -1912 13088 -1864 13792
rect -2664 13040 -1864 13088
rect -1252 13792 -452 13840
rect -1252 13088 -1204 13792
rect -500 13088 -452 13792
rect -1252 13040 -452 13088
rect 160 13792 960 13840
rect 160 13088 208 13792
rect 912 13088 960 13792
rect 160 13040 960 13088
rect 1572 13792 2372 13840
rect 1572 13088 1620 13792
rect 2324 13088 2372 13792
rect 1572 13040 2372 13088
rect 2984 13792 3784 13840
rect 2984 13088 3032 13792
rect 3736 13088 3784 13792
rect 2984 13040 3784 13088
rect 4396 13792 5196 13840
rect 4396 13088 4444 13792
rect 5148 13088 5196 13792
rect 4396 13040 5196 13088
rect 5808 13792 6608 13840
rect 5808 13088 5856 13792
rect 6560 13088 6608 13792
rect 5808 13040 6608 13088
rect 7220 13792 8020 13840
rect 7220 13088 7268 13792
rect 7972 13088 8020 13792
rect 7220 13040 8020 13088
rect 8632 13792 9432 13840
rect 8632 13088 8680 13792
rect 9384 13088 9432 13792
rect 8632 13040 9432 13088
rect 10044 13792 10844 13840
rect 10044 13088 10092 13792
rect 10796 13088 10844 13792
rect 10044 13040 10844 13088
rect 11456 13792 12256 13840
rect 11456 13088 11504 13792
rect 12208 13088 12256 13792
rect 11456 13040 12256 13088
rect 12868 13792 13668 13840
rect 12868 13088 12916 13792
rect 13620 13088 13668 13792
rect 12868 13040 13668 13088
rect 14280 13792 15080 13840
rect 14280 13088 14328 13792
rect 15032 13088 15080 13792
rect 14280 13040 15080 13088
rect 15692 13792 16492 13840
rect 15692 13088 15740 13792
rect 16444 13088 16492 13792
rect 15692 13040 16492 13088
rect 17104 13792 17904 13840
rect 17104 13088 17152 13792
rect 17856 13088 17904 13792
rect 17104 13040 17904 13088
rect 18516 13792 19316 13840
rect 18516 13088 18564 13792
rect 19268 13088 19316 13792
rect 18516 13040 19316 13088
rect 19928 13792 20728 13840
rect 19928 13088 19976 13792
rect 20680 13088 20728 13792
rect 19928 13040 20728 13088
rect 21340 13792 22140 13840
rect 21340 13088 21388 13792
rect 22092 13088 22140 13792
rect 21340 13040 22140 13088
rect 22752 13792 23552 13840
rect 22752 13088 22800 13792
rect 23504 13088 23552 13792
rect 22752 13040 23552 13088
rect -23844 12672 -23044 12720
rect -23844 11968 -23796 12672
rect -23092 11968 -23044 12672
rect -23844 11920 -23044 11968
rect -22432 12672 -21632 12720
rect -22432 11968 -22384 12672
rect -21680 11968 -21632 12672
rect -22432 11920 -21632 11968
rect -21020 12672 -20220 12720
rect -21020 11968 -20972 12672
rect -20268 11968 -20220 12672
rect -21020 11920 -20220 11968
rect -19608 12672 -18808 12720
rect -19608 11968 -19560 12672
rect -18856 11968 -18808 12672
rect -19608 11920 -18808 11968
rect -18196 12672 -17396 12720
rect -18196 11968 -18148 12672
rect -17444 11968 -17396 12672
rect -18196 11920 -17396 11968
rect -16784 12672 -15984 12720
rect -16784 11968 -16736 12672
rect -16032 11968 -15984 12672
rect -16784 11920 -15984 11968
rect -15372 12672 -14572 12720
rect -15372 11968 -15324 12672
rect -14620 11968 -14572 12672
rect -15372 11920 -14572 11968
rect -13960 12672 -13160 12720
rect -13960 11968 -13912 12672
rect -13208 11968 -13160 12672
rect -13960 11920 -13160 11968
rect -12548 12672 -11748 12720
rect -12548 11968 -12500 12672
rect -11796 11968 -11748 12672
rect -12548 11920 -11748 11968
rect -11136 12672 -10336 12720
rect -11136 11968 -11088 12672
rect -10384 11968 -10336 12672
rect -11136 11920 -10336 11968
rect -9724 12672 -8924 12720
rect -9724 11968 -9676 12672
rect -8972 11968 -8924 12672
rect -9724 11920 -8924 11968
rect -8312 12672 -7512 12720
rect -8312 11968 -8264 12672
rect -7560 11968 -7512 12672
rect -8312 11920 -7512 11968
rect -6900 12672 -6100 12720
rect -6900 11968 -6852 12672
rect -6148 11968 -6100 12672
rect -6900 11920 -6100 11968
rect -5488 12672 -4688 12720
rect -5488 11968 -5440 12672
rect -4736 11968 -4688 12672
rect -5488 11920 -4688 11968
rect -4076 12672 -3276 12720
rect -4076 11968 -4028 12672
rect -3324 11968 -3276 12672
rect -4076 11920 -3276 11968
rect -2664 12672 -1864 12720
rect -2664 11968 -2616 12672
rect -1912 11968 -1864 12672
rect -2664 11920 -1864 11968
rect -1252 12672 -452 12720
rect -1252 11968 -1204 12672
rect -500 11968 -452 12672
rect -1252 11920 -452 11968
rect 160 12672 960 12720
rect 160 11968 208 12672
rect 912 11968 960 12672
rect 160 11920 960 11968
rect 1572 12672 2372 12720
rect 1572 11968 1620 12672
rect 2324 11968 2372 12672
rect 1572 11920 2372 11968
rect 2984 12672 3784 12720
rect 2984 11968 3032 12672
rect 3736 11968 3784 12672
rect 2984 11920 3784 11968
rect 4396 12672 5196 12720
rect 4396 11968 4444 12672
rect 5148 11968 5196 12672
rect 4396 11920 5196 11968
rect 5808 12672 6608 12720
rect 5808 11968 5856 12672
rect 6560 11968 6608 12672
rect 5808 11920 6608 11968
rect 7220 12672 8020 12720
rect 7220 11968 7268 12672
rect 7972 11968 8020 12672
rect 7220 11920 8020 11968
rect 8632 12672 9432 12720
rect 8632 11968 8680 12672
rect 9384 11968 9432 12672
rect 8632 11920 9432 11968
rect 10044 12672 10844 12720
rect 10044 11968 10092 12672
rect 10796 11968 10844 12672
rect 10044 11920 10844 11968
rect 11456 12672 12256 12720
rect 11456 11968 11504 12672
rect 12208 11968 12256 12672
rect 11456 11920 12256 11968
rect 12868 12672 13668 12720
rect 12868 11968 12916 12672
rect 13620 11968 13668 12672
rect 12868 11920 13668 11968
rect 14280 12672 15080 12720
rect 14280 11968 14328 12672
rect 15032 11968 15080 12672
rect 14280 11920 15080 11968
rect 15692 12672 16492 12720
rect 15692 11968 15740 12672
rect 16444 11968 16492 12672
rect 15692 11920 16492 11968
rect 17104 12672 17904 12720
rect 17104 11968 17152 12672
rect 17856 11968 17904 12672
rect 17104 11920 17904 11968
rect 18516 12672 19316 12720
rect 18516 11968 18564 12672
rect 19268 11968 19316 12672
rect 18516 11920 19316 11968
rect 19928 12672 20728 12720
rect 19928 11968 19976 12672
rect 20680 11968 20728 12672
rect 19928 11920 20728 11968
rect 21340 12672 22140 12720
rect 21340 11968 21388 12672
rect 22092 11968 22140 12672
rect 21340 11920 22140 11968
rect 22752 12672 23552 12720
rect 22752 11968 22800 12672
rect 23504 11968 23552 12672
rect 22752 11920 23552 11968
rect -23844 11552 -23044 11600
rect -23844 10848 -23796 11552
rect -23092 10848 -23044 11552
rect -23844 10800 -23044 10848
rect -22432 11552 -21632 11600
rect -22432 10848 -22384 11552
rect -21680 10848 -21632 11552
rect -22432 10800 -21632 10848
rect -21020 11552 -20220 11600
rect -21020 10848 -20972 11552
rect -20268 10848 -20220 11552
rect -21020 10800 -20220 10848
rect -19608 11552 -18808 11600
rect -19608 10848 -19560 11552
rect -18856 10848 -18808 11552
rect -19608 10800 -18808 10848
rect -18196 11552 -17396 11600
rect -18196 10848 -18148 11552
rect -17444 10848 -17396 11552
rect -18196 10800 -17396 10848
rect -16784 11552 -15984 11600
rect -16784 10848 -16736 11552
rect -16032 10848 -15984 11552
rect -16784 10800 -15984 10848
rect -15372 11552 -14572 11600
rect -15372 10848 -15324 11552
rect -14620 10848 -14572 11552
rect -15372 10800 -14572 10848
rect -13960 11552 -13160 11600
rect -13960 10848 -13912 11552
rect -13208 10848 -13160 11552
rect -13960 10800 -13160 10848
rect -12548 11552 -11748 11600
rect -12548 10848 -12500 11552
rect -11796 10848 -11748 11552
rect -12548 10800 -11748 10848
rect -11136 11552 -10336 11600
rect -11136 10848 -11088 11552
rect -10384 10848 -10336 11552
rect -11136 10800 -10336 10848
rect -9724 11552 -8924 11600
rect -9724 10848 -9676 11552
rect -8972 10848 -8924 11552
rect -9724 10800 -8924 10848
rect -8312 11552 -7512 11600
rect -8312 10848 -8264 11552
rect -7560 10848 -7512 11552
rect -8312 10800 -7512 10848
rect -6900 11552 -6100 11600
rect -6900 10848 -6852 11552
rect -6148 10848 -6100 11552
rect -6900 10800 -6100 10848
rect -5488 11552 -4688 11600
rect -5488 10848 -5440 11552
rect -4736 10848 -4688 11552
rect -5488 10800 -4688 10848
rect -4076 11552 -3276 11600
rect -4076 10848 -4028 11552
rect -3324 10848 -3276 11552
rect -4076 10800 -3276 10848
rect -2664 11552 -1864 11600
rect -2664 10848 -2616 11552
rect -1912 10848 -1864 11552
rect -2664 10800 -1864 10848
rect -1252 11552 -452 11600
rect -1252 10848 -1204 11552
rect -500 10848 -452 11552
rect -1252 10800 -452 10848
rect 160 11552 960 11600
rect 160 10848 208 11552
rect 912 10848 960 11552
rect 160 10800 960 10848
rect 1572 11552 2372 11600
rect 1572 10848 1620 11552
rect 2324 10848 2372 11552
rect 1572 10800 2372 10848
rect 2984 11552 3784 11600
rect 2984 10848 3032 11552
rect 3736 10848 3784 11552
rect 2984 10800 3784 10848
rect 4396 11552 5196 11600
rect 4396 10848 4444 11552
rect 5148 10848 5196 11552
rect 4396 10800 5196 10848
rect 5808 11552 6608 11600
rect 5808 10848 5856 11552
rect 6560 10848 6608 11552
rect 5808 10800 6608 10848
rect 7220 11552 8020 11600
rect 7220 10848 7268 11552
rect 7972 10848 8020 11552
rect 7220 10800 8020 10848
rect 8632 11552 9432 11600
rect 8632 10848 8680 11552
rect 9384 10848 9432 11552
rect 8632 10800 9432 10848
rect 10044 11552 10844 11600
rect 10044 10848 10092 11552
rect 10796 10848 10844 11552
rect 10044 10800 10844 10848
rect 11456 11552 12256 11600
rect 11456 10848 11504 11552
rect 12208 10848 12256 11552
rect 11456 10800 12256 10848
rect 12868 11552 13668 11600
rect 12868 10848 12916 11552
rect 13620 10848 13668 11552
rect 12868 10800 13668 10848
rect 14280 11552 15080 11600
rect 14280 10848 14328 11552
rect 15032 10848 15080 11552
rect 14280 10800 15080 10848
rect 15692 11552 16492 11600
rect 15692 10848 15740 11552
rect 16444 10848 16492 11552
rect 15692 10800 16492 10848
rect 17104 11552 17904 11600
rect 17104 10848 17152 11552
rect 17856 10848 17904 11552
rect 17104 10800 17904 10848
rect 18516 11552 19316 11600
rect 18516 10848 18564 11552
rect 19268 10848 19316 11552
rect 18516 10800 19316 10848
rect 19928 11552 20728 11600
rect 19928 10848 19976 11552
rect 20680 10848 20728 11552
rect 19928 10800 20728 10848
rect 21340 11552 22140 11600
rect 21340 10848 21388 11552
rect 22092 10848 22140 11552
rect 21340 10800 22140 10848
rect 22752 11552 23552 11600
rect 22752 10848 22800 11552
rect 23504 10848 23552 11552
rect 22752 10800 23552 10848
rect -23844 10432 -23044 10480
rect -23844 9728 -23796 10432
rect -23092 9728 -23044 10432
rect -23844 9680 -23044 9728
rect -22432 10432 -21632 10480
rect -22432 9728 -22384 10432
rect -21680 9728 -21632 10432
rect -22432 9680 -21632 9728
rect -21020 10432 -20220 10480
rect -21020 9728 -20972 10432
rect -20268 9728 -20220 10432
rect -21020 9680 -20220 9728
rect -19608 10432 -18808 10480
rect -19608 9728 -19560 10432
rect -18856 9728 -18808 10432
rect -19608 9680 -18808 9728
rect -18196 10432 -17396 10480
rect -18196 9728 -18148 10432
rect -17444 9728 -17396 10432
rect -18196 9680 -17396 9728
rect -16784 10432 -15984 10480
rect -16784 9728 -16736 10432
rect -16032 9728 -15984 10432
rect -16784 9680 -15984 9728
rect -15372 10432 -14572 10480
rect -15372 9728 -15324 10432
rect -14620 9728 -14572 10432
rect -15372 9680 -14572 9728
rect -13960 10432 -13160 10480
rect -13960 9728 -13912 10432
rect -13208 9728 -13160 10432
rect -13960 9680 -13160 9728
rect -12548 10432 -11748 10480
rect -12548 9728 -12500 10432
rect -11796 9728 -11748 10432
rect -12548 9680 -11748 9728
rect -11136 10432 -10336 10480
rect -11136 9728 -11088 10432
rect -10384 9728 -10336 10432
rect -11136 9680 -10336 9728
rect -9724 10432 -8924 10480
rect -9724 9728 -9676 10432
rect -8972 9728 -8924 10432
rect -9724 9680 -8924 9728
rect -8312 10432 -7512 10480
rect -8312 9728 -8264 10432
rect -7560 9728 -7512 10432
rect -8312 9680 -7512 9728
rect -6900 10432 -6100 10480
rect -6900 9728 -6852 10432
rect -6148 9728 -6100 10432
rect -6900 9680 -6100 9728
rect -5488 10432 -4688 10480
rect -5488 9728 -5440 10432
rect -4736 9728 -4688 10432
rect -5488 9680 -4688 9728
rect -4076 10432 -3276 10480
rect -4076 9728 -4028 10432
rect -3324 9728 -3276 10432
rect -4076 9680 -3276 9728
rect -2664 10432 -1864 10480
rect -2664 9728 -2616 10432
rect -1912 9728 -1864 10432
rect -2664 9680 -1864 9728
rect -1252 10432 -452 10480
rect -1252 9728 -1204 10432
rect -500 9728 -452 10432
rect -1252 9680 -452 9728
rect 160 10432 960 10480
rect 160 9728 208 10432
rect 912 9728 960 10432
rect 160 9680 960 9728
rect 1572 10432 2372 10480
rect 1572 9728 1620 10432
rect 2324 9728 2372 10432
rect 1572 9680 2372 9728
rect 2984 10432 3784 10480
rect 2984 9728 3032 10432
rect 3736 9728 3784 10432
rect 2984 9680 3784 9728
rect 4396 10432 5196 10480
rect 4396 9728 4444 10432
rect 5148 9728 5196 10432
rect 4396 9680 5196 9728
rect 5808 10432 6608 10480
rect 5808 9728 5856 10432
rect 6560 9728 6608 10432
rect 5808 9680 6608 9728
rect 7220 10432 8020 10480
rect 7220 9728 7268 10432
rect 7972 9728 8020 10432
rect 7220 9680 8020 9728
rect 8632 10432 9432 10480
rect 8632 9728 8680 10432
rect 9384 9728 9432 10432
rect 8632 9680 9432 9728
rect 10044 10432 10844 10480
rect 10044 9728 10092 10432
rect 10796 9728 10844 10432
rect 10044 9680 10844 9728
rect 11456 10432 12256 10480
rect 11456 9728 11504 10432
rect 12208 9728 12256 10432
rect 11456 9680 12256 9728
rect 12868 10432 13668 10480
rect 12868 9728 12916 10432
rect 13620 9728 13668 10432
rect 12868 9680 13668 9728
rect 14280 10432 15080 10480
rect 14280 9728 14328 10432
rect 15032 9728 15080 10432
rect 14280 9680 15080 9728
rect 15692 10432 16492 10480
rect 15692 9728 15740 10432
rect 16444 9728 16492 10432
rect 15692 9680 16492 9728
rect 17104 10432 17904 10480
rect 17104 9728 17152 10432
rect 17856 9728 17904 10432
rect 17104 9680 17904 9728
rect 18516 10432 19316 10480
rect 18516 9728 18564 10432
rect 19268 9728 19316 10432
rect 18516 9680 19316 9728
rect 19928 10432 20728 10480
rect 19928 9728 19976 10432
rect 20680 9728 20728 10432
rect 19928 9680 20728 9728
rect 21340 10432 22140 10480
rect 21340 9728 21388 10432
rect 22092 9728 22140 10432
rect 21340 9680 22140 9728
rect 22752 10432 23552 10480
rect 22752 9728 22800 10432
rect 23504 9728 23552 10432
rect 22752 9680 23552 9728
rect -23844 9312 -23044 9360
rect -23844 8608 -23796 9312
rect -23092 8608 -23044 9312
rect -23844 8560 -23044 8608
rect -22432 9312 -21632 9360
rect -22432 8608 -22384 9312
rect -21680 8608 -21632 9312
rect -22432 8560 -21632 8608
rect -21020 9312 -20220 9360
rect -21020 8608 -20972 9312
rect -20268 8608 -20220 9312
rect -21020 8560 -20220 8608
rect -19608 9312 -18808 9360
rect -19608 8608 -19560 9312
rect -18856 8608 -18808 9312
rect -19608 8560 -18808 8608
rect -18196 9312 -17396 9360
rect -18196 8608 -18148 9312
rect -17444 8608 -17396 9312
rect -18196 8560 -17396 8608
rect -16784 9312 -15984 9360
rect -16784 8608 -16736 9312
rect -16032 8608 -15984 9312
rect -16784 8560 -15984 8608
rect -15372 9312 -14572 9360
rect -15372 8608 -15324 9312
rect -14620 8608 -14572 9312
rect -15372 8560 -14572 8608
rect -13960 9312 -13160 9360
rect -13960 8608 -13912 9312
rect -13208 8608 -13160 9312
rect -13960 8560 -13160 8608
rect -12548 9312 -11748 9360
rect -12548 8608 -12500 9312
rect -11796 8608 -11748 9312
rect -12548 8560 -11748 8608
rect -11136 9312 -10336 9360
rect -11136 8608 -11088 9312
rect -10384 8608 -10336 9312
rect -11136 8560 -10336 8608
rect -9724 9312 -8924 9360
rect -9724 8608 -9676 9312
rect -8972 8608 -8924 9312
rect -9724 8560 -8924 8608
rect -8312 9312 -7512 9360
rect -8312 8608 -8264 9312
rect -7560 8608 -7512 9312
rect -8312 8560 -7512 8608
rect -6900 9312 -6100 9360
rect -6900 8608 -6852 9312
rect -6148 8608 -6100 9312
rect -6900 8560 -6100 8608
rect -5488 9312 -4688 9360
rect -5488 8608 -5440 9312
rect -4736 8608 -4688 9312
rect -5488 8560 -4688 8608
rect -4076 9312 -3276 9360
rect -4076 8608 -4028 9312
rect -3324 8608 -3276 9312
rect -4076 8560 -3276 8608
rect -2664 9312 -1864 9360
rect -2664 8608 -2616 9312
rect -1912 8608 -1864 9312
rect -2664 8560 -1864 8608
rect -1252 9312 -452 9360
rect -1252 8608 -1204 9312
rect -500 8608 -452 9312
rect -1252 8560 -452 8608
rect 160 9312 960 9360
rect 160 8608 208 9312
rect 912 8608 960 9312
rect 160 8560 960 8608
rect 1572 9312 2372 9360
rect 1572 8608 1620 9312
rect 2324 8608 2372 9312
rect 1572 8560 2372 8608
rect 2984 9312 3784 9360
rect 2984 8608 3032 9312
rect 3736 8608 3784 9312
rect 2984 8560 3784 8608
rect 4396 9312 5196 9360
rect 4396 8608 4444 9312
rect 5148 8608 5196 9312
rect 4396 8560 5196 8608
rect 5808 9312 6608 9360
rect 5808 8608 5856 9312
rect 6560 8608 6608 9312
rect 5808 8560 6608 8608
rect 7220 9312 8020 9360
rect 7220 8608 7268 9312
rect 7972 8608 8020 9312
rect 7220 8560 8020 8608
rect 8632 9312 9432 9360
rect 8632 8608 8680 9312
rect 9384 8608 9432 9312
rect 8632 8560 9432 8608
rect 10044 9312 10844 9360
rect 10044 8608 10092 9312
rect 10796 8608 10844 9312
rect 10044 8560 10844 8608
rect 11456 9312 12256 9360
rect 11456 8608 11504 9312
rect 12208 8608 12256 9312
rect 11456 8560 12256 8608
rect 12868 9312 13668 9360
rect 12868 8608 12916 9312
rect 13620 8608 13668 9312
rect 12868 8560 13668 8608
rect 14280 9312 15080 9360
rect 14280 8608 14328 9312
rect 15032 8608 15080 9312
rect 14280 8560 15080 8608
rect 15692 9312 16492 9360
rect 15692 8608 15740 9312
rect 16444 8608 16492 9312
rect 15692 8560 16492 8608
rect 17104 9312 17904 9360
rect 17104 8608 17152 9312
rect 17856 8608 17904 9312
rect 17104 8560 17904 8608
rect 18516 9312 19316 9360
rect 18516 8608 18564 9312
rect 19268 8608 19316 9312
rect 18516 8560 19316 8608
rect 19928 9312 20728 9360
rect 19928 8608 19976 9312
rect 20680 8608 20728 9312
rect 19928 8560 20728 8608
rect 21340 9312 22140 9360
rect 21340 8608 21388 9312
rect 22092 8608 22140 9312
rect 21340 8560 22140 8608
rect 22752 9312 23552 9360
rect 22752 8608 22800 9312
rect 23504 8608 23552 9312
rect 22752 8560 23552 8608
rect -23844 8192 -23044 8240
rect -23844 7488 -23796 8192
rect -23092 7488 -23044 8192
rect -23844 7440 -23044 7488
rect -22432 8192 -21632 8240
rect -22432 7488 -22384 8192
rect -21680 7488 -21632 8192
rect -22432 7440 -21632 7488
rect -21020 8192 -20220 8240
rect -21020 7488 -20972 8192
rect -20268 7488 -20220 8192
rect -21020 7440 -20220 7488
rect -19608 8192 -18808 8240
rect -19608 7488 -19560 8192
rect -18856 7488 -18808 8192
rect -19608 7440 -18808 7488
rect -18196 8192 -17396 8240
rect -18196 7488 -18148 8192
rect -17444 7488 -17396 8192
rect -18196 7440 -17396 7488
rect -16784 8192 -15984 8240
rect -16784 7488 -16736 8192
rect -16032 7488 -15984 8192
rect -16784 7440 -15984 7488
rect -15372 8192 -14572 8240
rect -15372 7488 -15324 8192
rect -14620 7488 -14572 8192
rect -15372 7440 -14572 7488
rect -13960 8192 -13160 8240
rect -13960 7488 -13912 8192
rect -13208 7488 -13160 8192
rect -13960 7440 -13160 7488
rect -12548 8192 -11748 8240
rect -12548 7488 -12500 8192
rect -11796 7488 -11748 8192
rect -12548 7440 -11748 7488
rect -11136 8192 -10336 8240
rect -11136 7488 -11088 8192
rect -10384 7488 -10336 8192
rect -11136 7440 -10336 7488
rect -9724 8192 -8924 8240
rect -9724 7488 -9676 8192
rect -8972 7488 -8924 8192
rect -9724 7440 -8924 7488
rect -8312 8192 -7512 8240
rect -8312 7488 -8264 8192
rect -7560 7488 -7512 8192
rect -8312 7440 -7512 7488
rect -6900 8192 -6100 8240
rect -6900 7488 -6852 8192
rect -6148 7488 -6100 8192
rect -6900 7440 -6100 7488
rect -5488 8192 -4688 8240
rect -5488 7488 -5440 8192
rect -4736 7488 -4688 8192
rect -5488 7440 -4688 7488
rect -4076 8192 -3276 8240
rect -4076 7488 -4028 8192
rect -3324 7488 -3276 8192
rect -4076 7440 -3276 7488
rect -2664 8192 -1864 8240
rect -2664 7488 -2616 8192
rect -1912 7488 -1864 8192
rect -2664 7440 -1864 7488
rect -1252 8192 -452 8240
rect -1252 7488 -1204 8192
rect -500 7488 -452 8192
rect -1252 7440 -452 7488
rect 160 8192 960 8240
rect 160 7488 208 8192
rect 912 7488 960 8192
rect 160 7440 960 7488
rect 1572 8192 2372 8240
rect 1572 7488 1620 8192
rect 2324 7488 2372 8192
rect 1572 7440 2372 7488
rect 2984 8192 3784 8240
rect 2984 7488 3032 8192
rect 3736 7488 3784 8192
rect 2984 7440 3784 7488
rect 4396 8192 5196 8240
rect 4396 7488 4444 8192
rect 5148 7488 5196 8192
rect 4396 7440 5196 7488
rect 5808 8192 6608 8240
rect 5808 7488 5856 8192
rect 6560 7488 6608 8192
rect 5808 7440 6608 7488
rect 7220 8192 8020 8240
rect 7220 7488 7268 8192
rect 7972 7488 8020 8192
rect 7220 7440 8020 7488
rect 8632 8192 9432 8240
rect 8632 7488 8680 8192
rect 9384 7488 9432 8192
rect 8632 7440 9432 7488
rect 10044 8192 10844 8240
rect 10044 7488 10092 8192
rect 10796 7488 10844 8192
rect 10044 7440 10844 7488
rect 11456 8192 12256 8240
rect 11456 7488 11504 8192
rect 12208 7488 12256 8192
rect 11456 7440 12256 7488
rect 12868 8192 13668 8240
rect 12868 7488 12916 8192
rect 13620 7488 13668 8192
rect 12868 7440 13668 7488
rect 14280 8192 15080 8240
rect 14280 7488 14328 8192
rect 15032 7488 15080 8192
rect 14280 7440 15080 7488
rect 15692 8192 16492 8240
rect 15692 7488 15740 8192
rect 16444 7488 16492 8192
rect 15692 7440 16492 7488
rect 17104 8192 17904 8240
rect 17104 7488 17152 8192
rect 17856 7488 17904 8192
rect 17104 7440 17904 7488
rect 18516 8192 19316 8240
rect 18516 7488 18564 8192
rect 19268 7488 19316 8192
rect 18516 7440 19316 7488
rect 19928 8192 20728 8240
rect 19928 7488 19976 8192
rect 20680 7488 20728 8192
rect 19928 7440 20728 7488
rect 21340 8192 22140 8240
rect 21340 7488 21388 8192
rect 22092 7488 22140 8192
rect 21340 7440 22140 7488
rect 22752 8192 23552 8240
rect 22752 7488 22800 8192
rect 23504 7488 23552 8192
rect 22752 7440 23552 7488
rect -23844 7072 -23044 7120
rect -23844 6368 -23796 7072
rect -23092 6368 -23044 7072
rect -23844 6320 -23044 6368
rect -22432 7072 -21632 7120
rect -22432 6368 -22384 7072
rect -21680 6368 -21632 7072
rect -22432 6320 -21632 6368
rect -21020 7072 -20220 7120
rect -21020 6368 -20972 7072
rect -20268 6368 -20220 7072
rect -21020 6320 -20220 6368
rect -19608 7072 -18808 7120
rect -19608 6368 -19560 7072
rect -18856 6368 -18808 7072
rect -19608 6320 -18808 6368
rect -18196 7072 -17396 7120
rect -18196 6368 -18148 7072
rect -17444 6368 -17396 7072
rect -18196 6320 -17396 6368
rect -16784 7072 -15984 7120
rect -16784 6368 -16736 7072
rect -16032 6368 -15984 7072
rect -16784 6320 -15984 6368
rect -15372 7072 -14572 7120
rect -15372 6368 -15324 7072
rect -14620 6368 -14572 7072
rect -15372 6320 -14572 6368
rect -13960 7072 -13160 7120
rect -13960 6368 -13912 7072
rect -13208 6368 -13160 7072
rect -13960 6320 -13160 6368
rect -12548 7072 -11748 7120
rect -12548 6368 -12500 7072
rect -11796 6368 -11748 7072
rect -12548 6320 -11748 6368
rect -11136 7072 -10336 7120
rect -11136 6368 -11088 7072
rect -10384 6368 -10336 7072
rect -11136 6320 -10336 6368
rect -9724 7072 -8924 7120
rect -9724 6368 -9676 7072
rect -8972 6368 -8924 7072
rect -9724 6320 -8924 6368
rect -8312 7072 -7512 7120
rect -8312 6368 -8264 7072
rect -7560 6368 -7512 7072
rect -8312 6320 -7512 6368
rect -6900 7072 -6100 7120
rect -6900 6368 -6852 7072
rect -6148 6368 -6100 7072
rect -6900 6320 -6100 6368
rect -5488 7072 -4688 7120
rect -5488 6368 -5440 7072
rect -4736 6368 -4688 7072
rect -5488 6320 -4688 6368
rect -4076 7072 -3276 7120
rect -4076 6368 -4028 7072
rect -3324 6368 -3276 7072
rect -4076 6320 -3276 6368
rect -2664 7072 -1864 7120
rect -2664 6368 -2616 7072
rect -1912 6368 -1864 7072
rect -2664 6320 -1864 6368
rect -1252 7072 -452 7120
rect -1252 6368 -1204 7072
rect -500 6368 -452 7072
rect -1252 6320 -452 6368
rect 160 7072 960 7120
rect 160 6368 208 7072
rect 912 6368 960 7072
rect 160 6320 960 6368
rect 1572 7072 2372 7120
rect 1572 6368 1620 7072
rect 2324 6368 2372 7072
rect 1572 6320 2372 6368
rect 2984 7072 3784 7120
rect 2984 6368 3032 7072
rect 3736 6368 3784 7072
rect 2984 6320 3784 6368
rect 4396 7072 5196 7120
rect 4396 6368 4444 7072
rect 5148 6368 5196 7072
rect 4396 6320 5196 6368
rect 5808 7072 6608 7120
rect 5808 6368 5856 7072
rect 6560 6368 6608 7072
rect 5808 6320 6608 6368
rect 7220 7072 8020 7120
rect 7220 6368 7268 7072
rect 7972 6368 8020 7072
rect 7220 6320 8020 6368
rect 8632 7072 9432 7120
rect 8632 6368 8680 7072
rect 9384 6368 9432 7072
rect 8632 6320 9432 6368
rect 10044 7072 10844 7120
rect 10044 6368 10092 7072
rect 10796 6368 10844 7072
rect 10044 6320 10844 6368
rect 11456 7072 12256 7120
rect 11456 6368 11504 7072
rect 12208 6368 12256 7072
rect 11456 6320 12256 6368
rect 12868 7072 13668 7120
rect 12868 6368 12916 7072
rect 13620 6368 13668 7072
rect 12868 6320 13668 6368
rect 14280 7072 15080 7120
rect 14280 6368 14328 7072
rect 15032 6368 15080 7072
rect 14280 6320 15080 6368
rect 15692 7072 16492 7120
rect 15692 6368 15740 7072
rect 16444 6368 16492 7072
rect 15692 6320 16492 6368
rect 17104 7072 17904 7120
rect 17104 6368 17152 7072
rect 17856 6368 17904 7072
rect 17104 6320 17904 6368
rect 18516 7072 19316 7120
rect 18516 6368 18564 7072
rect 19268 6368 19316 7072
rect 18516 6320 19316 6368
rect 19928 7072 20728 7120
rect 19928 6368 19976 7072
rect 20680 6368 20728 7072
rect 19928 6320 20728 6368
rect 21340 7072 22140 7120
rect 21340 6368 21388 7072
rect 22092 6368 22140 7072
rect 21340 6320 22140 6368
rect 22752 7072 23552 7120
rect 22752 6368 22800 7072
rect 23504 6368 23552 7072
rect 22752 6320 23552 6368
rect -23844 5952 -23044 6000
rect -23844 5248 -23796 5952
rect -23092 5248 -23044 5952
rect -23844 5200 -23044 5248
rect -22432 5952 -21632 6000
rect -22432 5248 -22384 5952
rect -21680 5248 -21632 5952
rect -22432 5200 -21632 5248
rect -21020 5952 -20220 6000
rect -21020 5248 -20972 5952
rect -20268 5248 -20220 5952
rect -21020 5200 -20220 5248
rect -19608 5952 -18808 6000
rect -19608 5248 -19560 5952
rect -18856 5248 -18808 5952
rect -19608 5200 -18808 5248
rect -18196 5952 -17396 6000
rect -18196 5248 -18148 5952
rect -17444 5248 -17396 5952
rect -18196 5200 -17396 5248
rect -16784 5952 -15984 6000
rect -16784 5248 -16736 5952
rect -16032 5248 -15984 5952
rect -16784 5200 -15984 5248
rect -15372 5952 -14572 6000
rect -15372 5248 -15324 5952
rect -14620 5248 -14572 5952
rect -15372 5200 -14572 5248
rect -13960 5952 -13160 6000
rect -13960 5248 -13912 5952
rect -13208 5248 -13160 5952
rect -13960 5200 -13160 5248
rect -12548 5952 -11748 6000
rect -12548 5248 -12500 5952
rect -11796 5248 -11748 5952
rect -12548 5200 -11748 5248
rect -11136 5952 -10336 6000
rect -11136 5248 -11088 5952
rect -10384 5248 -10336 5952
rect -11136 5200 -10336 5248
rect -9724 5952 -8924 6000
rect -9724 5248 -9676 5952
rect -8972 5248 -8924 5952
rect -9724 5200 -8924 5248
rect -8312 5952 -7512 6000
rect -8312 5248 -8264 5952
rect -7560 5248 -7512 5952
rect -8312 5200 -7512 5248
rect -6900 5952 -6100 6000
rect -6900 5248 -6852 5952
rect -6148 5248 -6100 5952
rect -6900 5200 -6100 5248
rect -5488 5952 -4688 6000
rect -5488 5248 -5440 5952
rect -4736 5248 -4688 5952
rect -5488 5200 -4688 5248
rect -4076 5952 -3276 6000
rect -4076 5248 -4028 5952
rect -3324 5248 -3276 5952
rect -4076 5200 -3276 5248
rect -2664 5952 -1864 6000
rect -2664 5248 -2616 5952
rect -1912 5248 -1864 5952
rect -2664 5200 -1864 5248
rect -1252 5952 -452 6000
rect -1252 5248 -1204 5952
rect -500 5248 -452 5952
rect -1252 5200 -452 5248
rect 160 5952 960 6000
rect 160 5248 208 5952
rect 912 5248 960 5952
rect 160 5200 960 5248
rect 1572 5952 2372 6000
rect 1572 5248 1620 5952
rect 2324 5248 2372 5952
rect 1572 5200 2372 5248
rect 2984 5952 3784 6000
rect 2984 5248 3032 5952
rect 3736 5248 3784 5952
rect 2984 5200 3784 5248
rect 4396 5952 5196 6000
rect 4396 5248 4444 5952
rect 5148 5248 5196 5952
rect 4396 5200 5196 5248
rect 5808 5952 6608 6000
rect 5808 5248 5856 5952
rect 6560 5248 6608 5952
rect 5808 5200 6608 5248
rect 7220 5952 8020 6000
rect 7220 5248 7268 5952
rect 7972 5248 8020 5952
rect 7220 5200 8020 5248
rect 8632 5952 9432 6000
rect 8632 5248 8680 5952
rect 9384 5248 9432 5952
rect 8632 5200 9432 5248
rect 10044 5952 10844 6000
rect 10044 5248 10092 5952
rect 10796 5248 10844 5952
rect 10044 5200 10844 5248
rect 11456 5952 12256 6000
rect 11456 5248 11504 5952
rect 12208 5248 12256 5952
rect 11456 5200 12256 5248
rect 12868 5952 13668 6000
rect 12868 5248 12916 5952
rect 13620 5248 13668 5952
rect 12868 5200 13668 5248
rect 14280 5952 15080 6000
rect 14280 5248 14328 5952
rect 15032 5248 15080 5952
rect 14280 5200 15080 5248
rect 15692 5952 16492 6000
rect 15692 5248 15740 5952
rect 16444 5248 16492 5952
rect 15692 5200 16492 5248
rect 17104 5952 17904 6000
rect 17104 5248 17152 5952
rect 17856 5248 17904 5952
rect 17104 5200 17904 5248
rect 18516 5952 19316 6000
rect 18516 5248 18564 5952
rect 19268 5248 19316 5952
rect 18516 5200 19316 5248
rect 19928 5952 20728 6000
rect 19928 5248 19976 5952
rect 20680 5248 20728 5952
rect 19928 5200 20728 5248
rect 21340 5952 22140 6000
rect 21340 5248 21388 5952
rect 22092 5248 22140 5952
rect 21340 5200 22140 5248
rect 22752 5952 23552 6000
rect 22752 5248 22800 5952
rect 23504 5248 23552 5952
rect 22752 5200 23552 5248
rect -23844 4832 -23044 4880
rect -23844 4128 -23796 4832
rect -23092 4128 -23044 4832
rect -23844 4080 -23044 4128
rect -22432 4832 -21632 4880
rect -22432 4128 -22384 4832
rect -21680 4128 -21632 4832
rect -22432 4080 -21632 4128
rect -21020 4832 -20220 4880
rect -21020 4128 -20972 4832
rect -20268 4128 -20220 4832
rect -21020 4080 -20220 4128
rect -19608 4832 -18808 4880
rect -19608 4128 -19560 4832
rect -18856 4128 -18808 4832
rect -19608 4080 -18808 4128
rect -18196 4832 -17396 4880
rect -18196 4128 -18148 4832
rect -17444 4128 -17396 4832
rect -18196 4080 -17396 4128
rect -16784 4832 -15984 4880
rect -16784 4128 -16736 4832
rect -16032 4128 -15984 4832
rect -16784 4080 -15984 4128
rect -15372 4832 -14572 4880
rect -15372 4128 -15324 4832
rect -14620 4128 -14572 4832
rect -15372 4080 -14572 4128
rect -13960 4832 -13160 4880
rect -13960 4128 -13912 4832
rect -13208 4128 -13160 4832
rect -13960 4080 -13160 4128
rect -12548 4832 -11748 4880
rect -12548 4128 -12500 4832
rect -11796 4128 -11748 4832
rect -12548 4080 -11748 4128
rect -11136 4832 -10336 4880
rect -11136 4128 -11088 4832
rect -10384 4128 -10336 4832
rect -11136 4080 -10336 4128
rect -9724 4832 -8924 4880
rect -9724 4128 -9676 4832
rect -8972 4128 -8924 4832
rect -9724 4080 -8924 4128
rect -8312 4832 -7512 4880
rect -8312 4128 -8264 4832
rect -7560 4128 -7512 4832
rect -8312 4080 -7512 4128
rect -6900 4832 -6100 4880
rect -6900 4128 -6852 4832
rect -6148 4128 -6100 4832
rect -6900 4080 -6100 4128
rect -5488 4832 -4688 4880
rect -5488 4128 -5440 4832
rect -4736 4128 -4688 4832
rect -5488 4080 -4688 4128
rect -4076 4832 -3276 4880
rect -4076 4128 -4028 4832
rect -3324 4128 -3276 4832
rect -4076 4080 -3276 4128
rect -2664 4832 -1864 4880
rect -2664 4128 -2616 4832
rect -1912 4128 -1864 4832
rect -2664 4080 -1864 4128
rect -1252 4832 -452 4880
rect -1252 4128 -1204 4832
rect -500 4128 -452 4832
rect -1252 4080 -452 4128
rect 160 4832 960 4880
rect 160 4128 208 4832
rect 912 4128 960 4832
rect 160 4080 960 4128
rect 1572 4832 2372 4880
rect 1572 4128 1620 4832
rect 2324 4128 2372 4832
rect 1572 4080 2372 4128
rect 2984 4832 3784 4880
rect 2984 4128 3032 4832
rect 3736 4128 3784 4832
rect 2984 4080 3784 4128
rect 4396 4832 5196 4880
rect 4396 4128 4444 4832
rect 5148 4128 5196 4832
rect 4396 4080 5196 4128
rect 5808 4832 6608 4880
rect 5808 4128 5856 4832
rect 6560 4128 6608 4832
rect 5808 4080 6608 4128
rect 7220 4832 8020 4880
rect 7220 4128 7268 4832
rect 7972 4128 8020 4832
rect 7220 4080 8020 4128
rect 8632 4832 9432 4880
rect 8632 4128 8680 4832
rect 9384 4128 9432 4832
rect 8632 4080 9432 4128
rect 10044 4832 10844 4880
rect 10044 4128 10092 4832
rect 10796 4128 10844 4832
rect 10044 4080 10844 4128
rect 11456 4832 12256 4880
rect 11456 4128 11504 4832
rect 12208 4128 12256 4832
rect 11456 4080 12256 4128
rect 12868 4832 13668 4880
rect 12868 4128 12916 4832
rect 13620 4128 13668 4832
rect 12868 4080 13668 4128
rect 14280 4832 15080 4880
rect 14280 4128 14328 4832
rect 15032 4128 15080 4832
rect 14280 4080 15080 4128
rect 15692 4832 16492 4880
rect 15692 4128 15740 4832
rect 16444 4128 16492 4832
rect 15692 4080 16492 4128
rect 17104 4832 17904 4880
rect 17104 4128 17152 4832
rect 17856 4128 17904 4832
rect 17104 4080 17904 4128
rect 18516 4832 19316 4880
rect 18516 4128 18564 4832
rect 19268 4128 19316 4832
rect 18516 4080 19316 4128
rect 19928 4832 20728 4880
rect 19928 4128 19976 4832
rect 20680 4128 20728 4832
rect 19928 4080 20728 4128
rect 21340 4832 22140 4880
rect 21340 4128 21388 4832
rect 22092 4128 22140 4832
rect 21340 4080 22140 4128
rect 22752 4832 23552 4880
rect 22752 4128 22800 4832
rect 23504 4128 23552 4832
rect 22752 4080 23552 4128
rect -23844 3712 -23044 3760
rect -23844 3008 -23796 3712
rect -23092 3008 -23044 3712
rect -23844 2960 -23044 3008
rect -22432 3712 -21632 3760
rect -22432 3008 -22384 3712
rect -21680 3008 -21632 3712
rect -22432 2960 -21632 3008
rect -21020 3712 -20220 3760
rect -21020 3008 -20972 3712
rect -20268 3008 -20220 3712
rect -21020 2960 -20220 3008
rect -19608 3712 -18808 3760
rect -19608 3008 -19560 3712
rect -18856 3008 -18808 3712
rect -19608 2960 -18808 3008
rect -18196 3712 -17396 3760
rect -18196 3008 -18148 3712
rect -17444 3008 -17396 3712
rect -18196 2960 -17396 3008
rect -16784 3712 -15984 3760
rect -16784 3008 -16736 3712
rect -16032 3008 -15984 3712
rect -16784 2960 -15984 3008
rect -15372 3712 -14572 3760
rect -15372 3008 -15324 3712
rect -14620 3008 -14572 3712
rect -15372 2960 -14572 3008
rect -13960 3712 -13160 3760
rect -13960 3008 -13912 3712
rect -13208 3008 -13160 3712
rect -13960 2960 -13160 3008
rect -12548 3712 -11748 3760
rect -12548 3008 -12500 3712
rect -11796 3008 -11748 3712
rect -12548 2960 -11748 3008
rect -11136 3712 -10336 3760
rect -11136 3008 -11088 3712
rect -10384 3008 -10336 3712
rect -11136 2960 -10336 3008
rect -9724 3712 -8924 3760
rect -9724 3008 -9676 3712
rect -8972 3008 -8924 3712
rect -9724 2960 -8924 3008
rect -8312 3712 -7512 3760
rect -8312 3008 -8264 3712
rect -7560 3008 -7512 3712
rect -8312 2960 -7512 3008
rect -6900 3712 -6100 3760
rect -6900 3008 -6852 3712
rect -6148 3008 -6100 3712
rect -6900 2960 -6100 3008
rect -5488 3712 -4688 3760
rect -5488 3008 -5440 3712
rect -4736 3008 -4688 3712
rect -5488 2960 -4688 3008
rect -4076 3712 -3276 3760
rect -4076 3008 -4028 3712
rect -3324 3008 -3276 3712
rect -4076 2960 -3276 3008
rect -2664 3712 -1864 3760
rect -2664 3008 -2616 3712
rect -1912 3008 -1864 3712
rect -2664 2960 -1864 3008
rect -1252 3712 -452 3760
rect -1252 3008 -1204 3712
rect -500 3008 -452 3712
rect -1252 2960 -452 3008
rect 160 3712 960 3760
rect 160 3008 208 3712
rect 912 3008 960 3712
rect 160 2960 960 3008
rect 1572 3712 2372 3760
rect 1572 3008 1620 3712
rect 2324 3008 2372 3712
rect 1572 2960 2372 3008
rect 2984 3712 3784 3760
rect 2984 3008 3032 3712
rect 3736 3008 3784 3712
rect 2984 2960 3784 3008
rect 4396 3712 5196 3760
rect 4396 3008 4444 3712
rect 5148 3008 5196 3712
rect 4396 2960 5196 3008
rect 5808 3712 6608 3760
rect 5808 3008 5856 3712
rect 6560 3008 6608 3712
rect 5808 2960 6608 3008
rect 7220 3712 8020 3760
rect 7220 3008 7268 3712
rect 7972 3008 8020 3712
rect 7220 2960 8020 3008
rect 8632 3712 9432 3760
rect 8632 3008 8680 3712
rect 9384 3008 9432 3712
rect 8632 2960 9432 3008
rect 10044 3712 10844 3760
rect 10044 3008 10092 3712
rect 10796 3008 10844 3712
rect 10044 2960 10844 3008
rect 11456 3712 12256 3760
rect 11456 3008 11504 3712
rect 12208 3008 12256 3712
rect 11456 2960 12256 3008
rect 12868 3712 13668 3760
rect 12868 3008 12916 3712
rect 13620 3008 13668 3712
rect 12868 2960 13668 3008
rect 14280 3712 15080 3760
rect 14280 3008 14328 3712
rect 15032 3008 15080 3712
rect 14280 2960 15080 3008
rect 15692 3712 16492 3760
rect 15692 3008 15740 3712
rect 16444 3008 16492 3712
rect 15692 2960 16492 3008
rect 17104 3712 17904 3760
rect 17104 3008 17152 3712
rect 17856 3008 17904 3712
rect 17104 2960 17904 3008
rect 18516 3712 19316 3760
rect 18516 3008 18564 3712
rect 19268 3008 19316 3712
rect 18516 2960 19316 3008
rect 19928 3712 20728 3760
rect 19928 3008 19976 3712
rect 20680 3008 20728 3712
rect 19928 2960 20728 3008
rect 21340 3712 22140 3760
rect 21340 3008 21388 3712
rect 22092 3008 22140 3712
rect 21340 2960 22140 3008
rect 22752 3712 23552 3760
rect 22752 3008 22800 3712
rect 23504 3008 23552 3712
rect 22752 2960 23552 3008
rect -23844 2592 -23044 2640
rect -23844 1888 -23796 2592
rect -23092 1888 -23044 2592
rect -23844 1840 -23044 1888
rect -22432 2592 -21632 2640
rect -22432 1888 -22384 2592
rect -21680 1888 -21632 2592
rect -22432 1840 -21632 1888
rect -21020 2592 -20220 2640
rect -21020 1888 -20972 2592
rect -20268 1888 -20220 2592
rect -21020 1840 -20220 1888
rect -19608 2592 -18808 2640
rect -19608 1888 -19560 2592
rect -18856 1888 -18808 2592
rect -19608 1840 -18808 1888
rect -18196 2592 -17396 2640
rect -18196 1888 -18148 2592
rect -17444 1888 -17396 2592
rect -18196 1840 -17396 1888
rect -16784 2592 -15984 2640
rect -16784 1888 -16736 2592
rect -16032 1888 -15984 2592
rect -16784 1840 -15984 1888
rect -15372 2592 -14572 2640
rect -15372 1888 -15324 2592
rect -14620 1888 -14572 2592
rect -15372 1840 -14572 1888
rect -13960 2592 -13160 2640
rect -13960 1888 -13912 2592
rect -13208 1888 -13160 2592
rect -13960 1840 -13160 1888
rect -12548 2592 -11748 2640
rect -12548 1888 -12500 2592
rect -11796 1888 -11748 2592
rect -12548 1840 -11748 1888
rect -11136 2592 -10336 2640
rect -11136 1888 -11088 2592
rect -10384 1888 -10336 2592
rect -11136 1840 -10336 1888
rect -9724 2592 -8924 2640
rect -9724 1888 -9676 2592
rect -8972 1888 -8924 2592
rect -9724 1840 -8924 1888
rect -8312 2592 -7512 2640
rect -8312 1888 -8264 2592
rect -7560 1888 -7512 2592
rect -8312 1840 -7512 1888
rect -6900 2592 -6100 2640
rect -6900 1888 -6852 2592
rect -6148 1888 -6100 2592
rect -6900 1840 -6100 1888
rect -5488 2592 -4688 2640
rect -5488 1888 -5440 2592
rect -4736 1888 -4688 2592
rect -5488 1840 -4688 1888
rect -4076 2592 -3276 2640
rect -4076 1888 -4028 2592
rect -3324 1888 -3276 2592
rect -4076 1840 -3276 1888
rect -2664 2592 -1864 2640
rect -2664 1888 -2616 2592
rect -1912 1888 -1864 2592
rect -2664 1840 -1864 1888
rect -1252 2592 -452 2640
rect -1252 1888 -1204 2592
rect -500 1888 -452 2592
rect -1252 1840 -452 1888
rect 160 2592 960 2640
rect 160 1888 208 2592
rect 912 1888 960 2592
rect 160 1840 960 1888
rect 1572 2592 2372 2640
rect 1572 1888 1620 2592
rect 2324 1888 2372 2592
rect 1572 1840 2372 1888
rect 2984 2592 3784 2640
rect 2984 1888 3032 2592
rect 3736 1888 3784 2592
rect 2984 1840 3784 1888
rect 4396 2592 5196 2640
rect 4396 1888 4444 2592
rect 5148 1888 5196 2592
rect 4396 1840 5196 1888
rect 5808 2592 6608 2640
rect 5808 1888 5856 2592
rect 6560 1888 6608 2592
rect 5808 1840 6608 1888
rect 7220 2592 8020 2640
rect 7220 1888 7268 2592
rect 7972 1888 8020 2592
rect 7220 1840 8020 1888
rect 8632 2592 9432 2640
rect 8632 1888 8680 2592
rect 9384 1888 9432 2592
rect 8632 1840 9432 1888
rect 10044 2592 10844 2640
rect 10044 1888 10092 2592
rect 10796 1888 10844 2592
rect 10044 1840 10844 1888
rect 11456 2592 12256 2640
rect 11456 1888 11504 2592
rect 12208 1888 12256 2592
rect 11456 1840 12256 1888
rect 12868 2592 13668 2640
rect 12868 1888 12916 2592
rect 13620 1888 13668 2592
rect 12868 1840 13668 1888
rect 14280 2592 15080 2640
rect 14280 1888 14328 2592
rect 15032 1888 15080 2592
rect 14280 1840 15080 1888
rect 15692 2592 16492 2640
rect 15692 1888 15740 2592
rect 16444 1888 16492 2592
rect 15692 1840 16492 1888
rect 17104 2592 17904 2640
rect 17104 1888 17152 2592
rect 17856 1888 17904 2592
rect 17104 1840 17904 1888
rect 18516 2592 19316 2640
rect 18516 1888 18564 2592
rect 19268 1888 19316 2592
rect 18516 1840 19316 1888
rect 19928 2592 20728 2640
rect 19928 1888 19976 2592
rect 20680 1888 20728 2592
rect 19928 1840 20728 1888
rect 21340 2592 22140 2640
rect 21340 1888 21388 2592
rect 22092 1888 22140 2592
rect 21340 1840 22140 1888
rect 22752 2592 23552 2640
rect 22752 1888 22800 2592
rect 23504 1888 23552 2592
rect 22752 1840 23552 1888
rect -23844 1472 -23044 1520
rect -23844 768 -23796 1472
rect -23092 768 -23044 1472
rect -23844 720 -23044 768
rect -22432 1472 -21632 1520
rect -22432 768 -22384 1472
rect -21680 768 -21632 1472
rect -22432 720 -21632 768
rect -21020 1472 -20220 1520
rect -21020 768 -20972 1472
rect -20268 768 -20220 1472
rect -21020 720 -20220 768
rect -19608 1472 -18808 1520
rect -19608 768 -19560 1472
rect -18856 768 -18808 1472
rect -19608 720 -18808 768
rect -18196 1472 -17396 1520
rect -18196 768 -18148 1472
rect -17444 768 -17396 1472
rect -18196 720 -17396 768
rect -16784 1472 -15984 1520
rect -16784 768 -16736 1472
rect -16032 768 -15984 1472
rect -16784 720 -15984 768
rect -15372 1472 -14572 1520
rect -15372 768 -15324 1472
rect -14620 768 -14572 1472
rect -15372 720 -14572 768
rect -13960 1472 -13160 1520
rect -13960 768 -13912 1472
rect -13208 768 -13160 1472
rect -13960 720 -13160 768
rect -12548 1472 -11748 1520
rect -12548 768 -12500 1472
rect -11796 768 -11748 1472
rect -12548 720 -11748 768
rect -11136 1472 -10336 1520
rect -11136 768 -11088 1472
rect -10384 768 -10336 1472
rect -11136 720 -10336 768
rect -9724 1472 -8924 1520
rect -9724 768 -9676 1472
rect -8972 768 -8924 1472
rect -9724 720 -8924 768
rect -8312 1472 -7512 1520
rect -8312 768 -8264 1472
rect -7560 768 -7512 1472
rect -8312 720 -7512 768
rect -6900 1472 -6100 1520
rect -6900 768 -6852 1472
rect -6148 768 -6100 1472
rect -6900 720 -6100 768
rect -5488 1472 -4688 1520
rect -5488 768 -5440 1472
rect -4736 768 -4688 1472
rect -5488 720 -4688 768
rect -4076 1472 -3276 1520
rect -4076 768 -4028 1472
rect -3324 768 -3276 1472
rect -4076 720 -3276 768
rect -2664 1472 -1864 1520
rect -2664 768 -2616 1472
rect -1912 768 -1864 1472
rect -2664 720 -1864 768
rect -1252 1472 -452 1520
rect -1252 768 -1204 1472
rect -500 768 -452 1472
rect -1252 720 -452 768
rect 160 1472 960 1520
rect 160 768 208 1472
rect 912 768 960 1472
rect 160 720 960 768
rect 1572 1472 2372 1520
rect 1572 768 1620 1472
rect 2324 768 2372 1472
rect 1572 720 2372 768
rect 2984 1472 3784 1520
rect 2984 768 3032 1472
rect 3736 768 3784 1472
rect 2984 720 3784 768
rect 4396 1472 5196 1520
rect 4396 768 4444 1472
rect 5148 768 5196 1472
rect 4396 720 5196 768
rect 5808 1472 6608 1520
rect 5808 768 5856 1472
rect 6560 768 6608 1472
rect 5808 720 6608 768
rect 7220 1472 8020 1520
rect 7220 768 7268 1472
rect 7972 768 8020 1472
rect 7220 720 8020 768
rect 8632 1472 9432 1520
rect 8632 768 8680 1472
rect 9384 768 9432 1472
rect 8632 720 9432 768
rect 10044 1472 10844 1520
rect 10044 768 10092 1472
rect 10796 768 10844 1472
rect 10044 720 10844 768
rect 11456 1472 12256 1520
rect 11456 768 11504 1472
rect 12208 768 12256 1472
rect 11456 720 12256 768
rect 12868 1472 13668 1520
rect 12868 768 12916 1472
rect 13620 768 13668 1472
rect 12868 720 13668 768
rect 14280 1472 15080 1520
rect 14280 768 14328 1472
rect 15032 768 15080 1472
rect 14280 720 15080 768
rect 15692 1472 16492 1520
rect 15692 768 15740 1472
rect 16444 768 16492 1472
rect 15692 720 16492 768
rect 17104 1472 17904 1520
rect 17104 768 17152 1472
rect 17856 768 17904 1472
rect 17104 720 17904 768
rect 18516 1472 19316 1520
rect 18516 768 18564 1472
rect 19268 768 19316 1472
rect 18516 720 19316 768
rect 19928 1472 20728 1520
rect 19928 768 19976 1472
rect 20680 768 20728 1472
rect 19928 720 20728 768
rect 21340 1472 22140 1520
rect 21340 768 21388 1472
rect 22092 768 22140 1472
rect 21340 720 22140 768
rect 22752 1472 23552 1520
rect 22752 768 22800 1472
rect 23504 768 23552 1472
rect 22752 720 23552 768
rect -23844 352 -23044 400
rect -23844 -352 -23796 352
rect -23092 -352 -23044 352
rect -23844 -400 -23044 -352
rect -22432 352 -21632 400
rect -22432 -352 -22384 352
rect -21680 -352 -21632 352
rect -22432 -400 -21632 -352
rect -21020 352 -20220 400
rect -21020 -352 -20972 352
rect -20268 -352 -20220 352
rect -21020 -400 -20220 -352
rect -19608 352 -18808 400
rect -19608 -352 -19560 352
rect -18856 -352 -18808 352
rect -19608 -400 -18808 -352
rect -18196 352 -17396 400
rect -18196 -352 -18148 352
rect -17444 -352 -17396 352
rect -18196 -400 -17396 -352
rect -16784 352 -15984 400
rect -16784 -352 -16736 352
rect -16032 -352 -15984 352
rect -16784 -400 -15984 -352
rect -15372 352 -14572 400
rect -15372 -352 -15324 352
rect -14620 -352 -14572 352
rect -15372 -400 -14572 -352
rect -13960 352 -13160 400
rect -13960 -352 -13912 352
rect -13208 -352 -13160 352
rect -13960 -400 -13160 -352
rect -12548 352 -11748 400
rect -12548 -352 -12500 352
rect -11796 -352 -11748 352
rect -12548 -400 -11748 -352
rect -11136 352 -10336 400
rect -11136 -352 -11088 352
rect -10384 -352 -10336 352
rect -11136 -400 -10336 -352
rect -9724 352 -8924 400
rect -9724 -352 -9676 352
rect -8972 -352 -8924 352
rect -9724 -400 -8924 -352
rect -8312 352 -7512 400
rect -8312 -352 -8264 352
rect -7560 -352 -7512 352
rect -8312 -400 -7512 -352
rect -6900 352 -6100 400
rect -6900 -352 -6852 352
rect -6148 -352 -6100 352
rect -6900 -400 -6100 -352
rect -5488 352 -4688 400
rect -5488 -352 -5440 352
rect -4736 -352 -4688 352
rect -5488 -400 -4688 -352
rect -4076 352 -3276 400
rect -4076 -352 -4028 352
rect -3324 -352 -3276 352
rect -4076 -400 -3276 -352
rect -2664 352 -1864 400
rect -2664 -352 -2616 352
rect -1912 -352 -1864 352
rect -2664 -400 -1864 -352
rect -1252 352 -452 400
rect -1252 -352 -1204 352
rect -500 -352 -452 352
rect -1252 -400 -452 -352
rect 160 352 960 400
rect 160 -352 208 352
rect 912 -352 960 352
rect 160 -400 960 -352
rect 1572 352 2372 400
rect 1572 -352 1620 352
rect 2324 -352 2372 352
rect 1572 -400 2372 -352
rect 2984 352 3784 400
rect 2984 -352 3032 352
rect 3736 -352 3784 352
rect 2984 -400 3784 -352
rect 4396 352 5196 400
rect 4396 -352 4444 352
rect 5148 -352 5196 352
rect 4396 -400 5196 -352
rect 5808 352 6608 400
rect 5808 -352 5856 352
rect 6560 -352 6608 352
rect 5808 -400 6608 -352
rect 7220 352 8020 400
rect 7220 -352 7268 352
rect 7972 -352 8020 352
rect 7220 -400 8020 -352
rect 8632 352 9432 400
rect 8632 -352 8680 352
rect 9384 -352 9432 352
rect 8632 -400 9432 -352
rect 10044 352 10844 400
rect 10044 -352 10092 352
rect 10796 -352 10844 352
rect 10044 -400 10844 -352
rect 11456 352 12256 400
rect 11456 -352 11504 352
rect 12208 -352 12256 352
rect 11456 -400 12256 -352
rect 12868 352 13668 400
rect 12868 -352 12916 352
rect 13620 -352 13668 352
rect 12868 -400 13668 -352
rect 14280 352 15080 400
rect 14280 -352 14328 352
rect 15032 -352 15080 352
rect 14280 -400 15080 -352
rect 15692 352 16492 400
rect 15692 -352 15740 352
rect 16444 -352 16492 352
rect 15692 -400 16492 -352
rect 17104 352 17904 400
rect 17104 -352 17152 352
rect 17856 -352 17904 352
rect 17104 -400 17904 -352
rect 18516 352 19316 400
rect 18516 -352 18564 352
rect 19268 -352 19316 352
rect 18516 -400 19316 -352
rect 19928 352 20728 400
rect 19928 -352 19976 352
rect 20680 -352 20728 352
rect 19928 -400 20728 -352
rect 21340 352 22140 400
rect 21340 -352 21388 352
rect 22092 -352 22140 352
rect 21340 -400 22140 -352
rect 22752 352 23552 400
rect 22752 -352 22800 352
rect 23504 -352 23552 352
rect 22752 -400 23552 -352
rect -23844 -768 -23044 -720
rect -23844 -1472 -23796 -768
rect -23092 -1472 -23044 -768
rect -23844 -1520 -23044 -1472
rect -22432 -768 -21632 -720
rect -22432 -1472 -22384 -768
rect -21680 -1472 -21632 -768
rect -22432 -1520 -21632 -1472
rect -21020 -768 -20220 -720
rect -21020 -1472 -20972 -768
rect -20268 -1472 -20220 -768
rect -21020 -1520 -20220 -1472
rect -19608 -768 -18808 -720
rect -19608 -1472 -19560 -768
rect -18856 -1472 -18808 -768
rect -19608 -1520 -18808 -1472
rect -18196 -768 -17396 -720
rect -18196 -1472 -18148 -768
rect -17444 -1472 -17396 -768
rect -18196 -1520 -17396 -1472
rect -16784 -768 -15984 -720
rect -16784 -1472 -16736 -768
rect -16032 -1472 -15984 -768
rect -16784 -1520 -15984 -1472
rect -15372 -768 -14572 -720
rect -15372 -1472 -15324 -768
rect -14620 -1472 -14572 -768
rect -15372 -1520 -14572 -1472
rect -13960 -768 -13160 -720
rect -13960 -1472 -13912 -768
rect -13208 -1472 -13160 -768
rect -13960 -1520 -13160 -1472
rect -12548 -768 -11748 -720
rect -12548 -1472 -12500 -768
rect -11796 -1472 -11748 -768
rect -12548 -1520 -11748 -1472
rect -11136 -768 -10336 -720
rect -11136 -1472 -11088 -768
rect -10384 -1472 -10336 -768
rect -11136 -1520 -10336 -1472
rect -9724 -768 -8924 -720
rect -9724 -1472 -9676 -768
rect -8972 -1472 -8924 -768
rect -9724 -1520 -8924 -1472
rect -8312 -768 -7512 -720
rect -8312 -1472 -8264 -768
rect -7560 -1472 -7512 -768
rect -8312 -1520 -7512 -1472
rect -6900 -768 -6100 -720
rect -6900 -1472 -6852 -768
rect -6148 -1472 -6100 -768
rect -6900 -1520 -6100 -1472
rect -5488 -768 -4688 -720
rect -5488 -1472 -5440 -768
rect -4736 -1472 -4688 -768
rect -5488 -1520 -4688 -1472
rect -4076 -768 -3276 -720
rect -4076 -1472 -4028 -768
rect -3324 -1472 -3276 -768
rect -4076 -1520 -3276 -1472
rect -2664 -768 -1864 -720
rect -2664 -1472 -2616 -768
rect -1912 -1472 -1864 -768
rect -2664 -1520 -1864 -1472
rect -1252 -768 -452 -720
rect -1252 -1472 -1204 -768
rect -500 -1472 -452 -768
rect -1252 -1520 -452 -1472
rect 160 -768 960 -720
rect 160 -1472 208 -768
rect 912 -1472 960 -768
rect 160 -1520 960 -1472
rect 1572 -768 2372 -720
rect 1572 -1472 1620 -768
rect 2324 -1472 2372 -768
rect 1572 -1520 2372 -1472
rect 2984 -768 3784 -720
rect 2984 -1472 3032 -768
rect 3736 -1472 3784 -768
rect 2984 -1520 3784 -1472
rect 4396 -768 5196 -720
rect 4396 -1472 4444 -768
rect 5148 -1472 5196 -768
rect 4396 -1520 5196 -1472
rect 5808 -768 6608 -720
rect 5808 -1472 5856 -768
rect 6560 -1472 6608 -768
rect 5808 -1520 6608 -1472
rect 7220 -768 8020 -720
rect 7220 -1472 7268 -768
rect 7972 -1472 8020 -768
rect 7220 -1520 8020 -1472
rect 8632 -768 9432 -720
rect 8632 -1472 8680 -768
rect 9384 -1472 9432 -768
rect 8632 -1520 9432 -1472
rect 10044 -768 10844 -720
rect 10044 -1472 10092 -768
rect 10796 -1472 10844 -768
rect 10044 -1520 10844 -1472
rect 11456 -768 12256 -720
rect 11456 -1472 11504 -768
rect 12208 -1472 12256 -768
rect 11456 -1520 12256 -1472
rect 12868 -768 13668 -720
rect 12868 -1472 12916 -768
rect 13620 -1472 13668 -768
rect 12868 -1520 13668 -1472
rect 14280 -768 15080 -720
rect 14280 -1472 14328 -768
rect 15032 -1472 15080 -768
rect 14280 -1520 15080 -1472
rect 15692 -768 16492 -720
rect 15692 -1472 15740 -768
rect 16444 -1472 16492 -768
rect 15692 -1520 16492 -1472
rect 17104 -768 17904 -720
rect 17104 -1472 17152 -768
rect 17856 -1472 17904 -768
rect 17104 -1520 17904 -1472
rect 18516 -768 19316 -720
rect 18516 -1472 18564 -768
rect 19268 -1472 19316 -768
rect 18516 -1520 19316 -1472
rect 19928 -768 20728 -720
rect 19928 -1472 19976 -768
rect 20680 -1472 20728 -768
rect 19928 -1520 20728 -1472
rect 21340 -768 22140 -720
rect 21340 -1472 21388 -768
rect 22092 -1472 22140 -768
rect 21340 -1520 22140 -1472
rect 22752 -768 23552 -720
rect 22752 -1472 22800 -768
rect 23504 -1472 23552 -768
rect 22752 -1520 23552 -1472
rect -23844 -1888 -23044 -1840
rect -23844 -2592 -23796 -1888
rect -23092 -2592 -23044 -1888
rect -23844 -2640 -23044 -2592
rect -22432 -1888 -21632 -1840
rect -22432 -2592 -22384 -1888
rect -21680 -2592 -21632 -1888
rect -22432 -2640 -21632 -2592
rect -21020 -1888 -20220 -1840
rect -21020 -2592 -20972 -1888
rect -20268 -2592 -20220 -1888
rect -21020 -2640 -20220 -2592
rect -19608 -1888 -18808 -1840
rect -19608 -2592 -19560 -1888
rect -18856 -2592 -18808 -1888
rect -19608 -2640 -18808 -2592
rect -18196 -1888 -17396 -1840
rect -18196 -2592 -18148 -1888
rect -17444 -2592 -17396 -1888
rect -18196 -2640 -17396 -2592
rect -16784 -1888 -15984 -1840
rect -16784 -2592 -16736 -1888
rect -16032 -2592 -15984 -1888
rect -16784 -2640 -15984 -2592
rect -15372 -1888 -14572 -1840
rect -15372 -2592 -15324 -1888
rect -14620 -2592 -14572 -1888
rect -15372 -2640 -14572 -2592
rect -13960 -1888 -13160 -1840
rect -13960 -2592 -13912 -1888
rect -13208 -2592 -13160 -1888
rect -13960 -2640 -13160 -2592
rect -12548 -1888 -11748 -1840
rect -12548 -2592 -12500 -1888
rect -11796 -2592 -11748 -1888
rect -12548 -2640 -11748 -2592
rect -11136 -1888 -10336 -1840
rect -11136 -2592 -11088 -1888
rect -10384 -2592 -10336 -1888
rect -11136 -2640 -10336 -2592
rect -9724 -1888 -8924 -1840
rect -9724 -2592 -9676 -1888
rect -8972 -2592 -8924 -1888
rect -9724 -2640 -8924 -2592
rect -8312 -1888 -7512 -1840
rect -8312 -2592 -8264 -1888
rect -7560 -2592 -7512 -1888
rect -8312 -2640 -7512 -2592
rect -6900 -1888 -6100 -1840
rect -6900 -2592 -6852 -1888
rect -6148 -2592 -6100 -1888
rect -6900 -2640 -6100 -2592
rect -5488 -1888 -4688 -1840
rect -5488 -2592 -5440 -1888
rect -4736 -2592 -4688 -1888
rect -5488 -2640 -4688 -2592
rect -4076 -1888 -3276 -1840
rect -4076 -2592 -4028 -1888
rect -3324 -2592 -3276 -1888
rect -4076 -2640 -3276 -2592
rect -2664 -1888 -1864 -1840
rect -2664 -2592 -2616 -1888
rect -1912 -2592 -1864 -1888
rect -2664 -2640 -1864 -2592
rect -1252 -1888 -452 -1840
rect -1252 -2592 -1204 -1888
rect -500 -2592 -452 -1888
rect -1252 -2640 -452 -2592
rect 160 -1888 960 -1840
rect 160 -2592 208 -1888
rect 912 -2592 960 -1888
rect 160 -2640 960 -2592
rect 1572 -1888 2372 -1840
rect 1572 -2592 1620 -1888
rect 2324 -2592 2372 -1888
rect 1572 -2640 2372 -2592
rect 2984 -1888 3784 -1840
rect 2984 -2592 3032 -1888
rect 3736 -2592 3784 -1888
rect 2984 -2640 3784 -2592
rect 4396 -1888 5196 -1840
rect 4396 -2592 4444 -1888
rect 5148 -2592 5196 -1888
rect 4396 -2640 5196 -2592
rect 5808 -1888 6608 -1840
rect 5808 -2592 5856 -1888
rect 6560 -2592 6608 -1888
rect 5808 -2640 6608 -2592
rect 7220 -1888 8020 -1840
rect 7220 -2592 7268 -1888
rect 7972 -2592 8020 -1888
rect 7220 -2640 8020 -2592
rect 8632 -1888 9432 -1840
rect 8632 -2592 8680 -1888
rect 9384 -2592 9432 -1888
rect 8632 -2640 9432 -2592
rect 10044 -1888 10844 -1840
rect 10044 -2592 10092 -1888
rect 10796 -2592 10844 -1888
rect 10044 -2640 10844 -2592
rect 11456 -1888 12256 -1840
rect 11456 -2592 11504 -1888
rect 12208 -2592 12256 -1888
rect 11456 -2640 12256 -2592
rect 12868 -1888 13668 -1840
rect 12868 -2592 12916 -1888
rect 13620 -2592 13668 -1888
rect 12868 -2640 13668 -2592
rect 14280 -1888 15080 -1840
rect 14280 -2592 14328 -1888
rect 15032 -2592 15080 -1888
rect 14280 -2640 15080 -2592
rect 15692 -1888 16492 -1840
rect 15692 -2592 15740 -1888
rect 16444 -2592 16492 -1888
rect 15692 -2640 16492 -2592
rect 17104 -1888 17904 -1840
rect 17104 -2592 17152 -1888
rect 17856 -2592 17904 -1888
rect 17104 -2640 17904 -2592
rect 18516 -1888 19316 -1840
rect 18516 -2592 18564 -1888
rect 19268 -2592 19316 -1888
rect 18516 -2640 19316 -2592
rect 19928 -1888 20728 -1840
rect 19928 -2592 19976 -1888
rect 20680 -2592 20728 -1888
rect 19928 -2640 20728 -2592
rect 21340 -1888 22140 -1840
rect 21340 -2592 21388 -1888
rect 22092 -2592 22140 -1888
rect 21340 -2640 22140 -2592
rect 22752 -1888 23552 -1840
rect 22752 -2592 22800 -1888
rect 23504 -2592 23552 -1888
rect 22752 -2640 23552 -2592
rect -23844 -3008 -23044 -2960
rect -23844 -3712 -23796 -3008
rect -23092 -3712 -23044 -3008
rect -23844 -3760 -23044 -3712
rect -22432 -3008 -21632 -2960
rect -22432 -3712 -22384 -3008
rect -21680 -3712 -21632 -3008
rect -22432 -3760 -21632 -3712
rect -21020 -3008 -20220 -2960
rect -21020 -3712 -20972 -3008
rect -20268 -3712 -20220 -3008
rect -21020 -3760 -20220 -3712
rect -19608 -3008 -18808 -2960
rect -19608 -3712 -19560 -3008
rect -18856 -3712 -18808 -3008
rect -19608 -3760 -18808 -3712
rect -18196 -3008 -17396 -2960
rect -18196 -3712 -18148 -3008
rect -17444 -3712 -17396 -3008
rect -18196 -3760 -17396 -3712
rect -16784 -3008 -15984 -2960
rect -16784 -3712 -16736 -3008
rect -16032 -3712 -15984 -3008
rect -16784 -3760 -15984 -3712
rect -15372 -3008 -14572 -2960
rect -15372 -3712 -15324 -3008
rect -14620 -3712 -14572 -3008
rect -15372 -3760 -14572 -3712
rect -13960 -3008 -13160 -2960
rect -13960 -3712 -13912 -3008
rect -13208 -3712 -13160 -3008
rect -13960 -3760 -13160 -3712
rect -12548 -3008 -11748 -2960
rect -12548 -3712 -12500 -3008
rect -11796 -3712 -11748 -3008
rect -12548 -3760 -11748 -3712
rect -11136 -3008 -10336 -2960
rect -11136 -3712 -11088 -3008
rect -10384 -3712 -10336 -3008
rect -11136 -3760 -10336 -3712
rect -9724 -3008 -8924 -2960
rect -9724 -3712 -9676 -3008
rect -8972 -3712 -8924 -3008
rect -9724 -3760 -8924 -3712
rect -8312 -3008 -7512 -2960
rect -8312 -3712 -8264 -3008
rect -7560 -3712 -7512 -3008
rect -8312 -3760 -7512 -3712
rect -6900 -3008 -6100 -2960
rect -6900 -3712 -6852 -3008
rect -6148 -3712 -6100 -3008
rect -6900 -3760 -6100 -3712
rect -5488 -3008 -4688 -2960
rect -5488 -3712 -5440 -3008
rect -4736 -3712 -4688 -3008
rect -5488 -3760 -4688 -3712
rect -4076 -3008 -3276 -2960
rect -4076 -3712 -4028 -3008
rect -3324 -3712 -3276 -3008
rect -4076 -3760 -3276 -3712
rect -2664 -3008 -1864 -2960
rect -2664 -3712 -2616 -3008
rect -1912 -3712 -1864 -3008
rect -2664 -3760 -1864 -3712
rect -1252 -3008 -452 -2960
rect -1252 -3712 -1204 -3008
rect -500 -3712 -452 -3008
rect -1252 -3760 -452 -3712
rect 160 -3008 960 -2960
rect 160 -3712 208 -3008
rect 912 -3712 960 -3008
rect 160 -3760 960 -3712
rect 1572 -3008 2372 -2960
rect 1572 -3712 1620 -3008
rect 2324 -3712 2372 -3008
rect 1572 -3760 2372 -3712
rect 2984 -3008 3784 -2960
rect 2984 -3712 3032 -3008
rect 3736 -3712 3784 -3008
rect 2984 -3760 3784 -3712
rect 4396 -3008 5196 -2960
rect 4396 -3712 4444 -3008
rect 5148 -3712 5196 -3008
rect 4396 -3760 5196 -3712
rect 5808 -3008 6608 -2960
rect 5808 -3712 5856 -3008
rect 6560 -3712 6608 -3008
rect 5808 -3760 6608 -3712
rect 7220 -3008 8020 -2960
rect 7220 -3712 7268 -3008
rect 7972 -3712 8020 -3008
rect 7220 -3760 8020 -3712
rect 8632 -3008 9432 -2960
rect 8632 -3712 8680 -3008
rect 9384 -3712 9432 -3008
rect 8632 -3760 9432 -3712
rect 10044 -3008 10844 -2960
rect 10044 -3712 10092 -3008
rect 10796 -3712 10844 -3008
rect 10044 -3760 10844 -3712
rect 11456 -3008 12256 -2960
rect 11456 -3712 11504 -3008
rect 12208 -3712 12256 -3008
rect 11456 -3760 12256 -3712
rect 12868 -3008 13668 -2960
rect 12868 -3712 12916 -3008
rect 13620 -3712 13668 -3008
rect 12868 -3760 13668 -3712
rect 14280 -3008 15080 -2960
rect 14280 -3712 14328 -3008
rect 15032 -3712 15080 -3008
rect 14280 -3760 15080 -3712
rect 15692 -3008 16492 -2960
rect 15692 -3712 15740 -3008
rect 16444 -3712 16492 -3008
rect 15692 -3760 16492 -3712
rect 17104 -3008 17904 -2960
rect 17104 -3712 17152 -3008
rect 17856 -3712 17904 -3008
rect 17104 -3760 17904 -3712
rect 18516 -3008 19316 -2960
rect 18516 -3712 18564 -3008
rect 19268 -3712 19316 -3008
rect 18516 -3760 19316 -3712
rect 19928 -3008 20728 -2960
rect 19928 -3712 19976 -3008
rect 20680 -3712 20728 -3008
rect 19928 -3760 20728 -3712
rect 21340 -3008 22140 -2960
rect 21340 -3712 21388 -3008
rect 22092 -3712 22140 -3008
rect 21340 -3760 22140 -3712
rect 22752 -3008 23552 -2960
rect 22752 -3712 22800 -3008
rect 23504 -3712 23552 -3008
rect 22752 -3760 23552 -3712
rect -23844 -4128 -23044 -4080
rect -23844 -4832 -23796 -4128
rect -23092 -4832 -23044 -4128
rect -23844 -4880 -23044 -4832
rect -22432 -4128 -21632 -4080
rect -22432 -4832 -22384 -4128
rect -21680 -4832 -21632 -4128
rect -22432 -4880 -21632 -4832
rect -21020 -4128 -20220 -4080
rect -21020 -4832 -20972 -4128
rect -20268 -4832 -20220 -4128
rect -21020 -4880 -20220 -4832
rect -19608 -4128 -18808 -4080
rect -19608 -4832 -19560 -4128
rect -18856 -4832 -18808 -4128
rect -19608 -4880 -18808 -4832
rect -18196 -4128 -17396 -4080
rect -18196 -4832 -18148 -4128
rect -17444 -4832 -17396 -4128
rect -18196 -4880 -17396 -4832
rect -16784 -4128 -15984 -4080
rect -16784 -4832 -16736 -4128
rect -16032 -4832 -15984 -4128
rect -16784 -4880 -15984 -4832
rect -15372 -4128 -14572 -4080
rect -15372 -4832 -15324 -4128
rect -14620 -4832 -14572 -4128
rect -15372 -4880 -14572 -4832
rect -13960 -4128 -13160 -4080
rect -13960 -4832 -13912 -4128
rect -13208 -4832 -13160 -4128
rect -13960 -4880 -13160 -4832
rect -12548 -4128 -11748 -4080
rect -12548 -4832 -12500 -4128
rect -11796 -4832 -11748 -4128
rect -12548 -4880 -11748 -4832
rect -11136 -4128 -10336 -4080
rect -11136 -4832 -11088 -4128
rect -10384 -4832 -10336 -4128
rect -11136 -4880 -10336 -4832
rect -9724 -4128 -8924 -4080
rect -9724 -4832 -9676 -4128
rect -8972 -4832 -8924 -4128
rect -9724 -4880 -8924 -4832
rect -8312 -4128 -7512 -4080
rect -8312 -4832 -8264 -4128
rect -7560 -4832 -7512 -4128
rect -8312 -4880 -7512 -4832
rect -6900 -4128 -6100 -4080
rect -6900 -4832 -6852 -4128
rect -6148 -4832 -6100 -4128
rect -6900 -4880 -6100 -4832
rect -5488 -4128 -4688 -4080
rect -5488 -4832 -5440 -4128
rect -4736 -4832 -4688 -4128
rect -5488 -4880 -4688 -4832
rect -4076 -4128 -3276 -4080
rect -4076 -4832 -4028 -4128
rect -3324 -4832 -3276 -4128
rect -4076 -4880 -3276 -4832
rect -2664 -4128 -1864 -4080
rect -2664 -4832 -2616 -4128
rect -1912 -4832 -1864 -4128
rect -2664 -4880 -1864 -4832
rect -1252 -4128 -452 -4080
rect -1252 -4832 -1204 -4128
rect -500 -4832 -452 -4128
rect -1252 -4880 -452 -4832
rect 160 -4128 960 -4080
rect 160 -4832 208 -4128
rect 912 -4832 960 -4128
rect 160 -4880 960 -4832
rect 1572 -4128 2372 -4080
rect 1572 -4832 1620 -4128
rect 2324 -4832 2372 -4128
rect 1572 -4880 2372 -4832
rect 2984 -4128 3784 -4080
rect 2984 -4832 3032 -4128
rect 3736 -4832 3784 -4128
rect 2984 -4880 3784 -4832
rect 4396 -4128 5196 -4080
rect 4396 -4832 4444 -4128
rect 5148 -4832 5196 -4128
rect 4396 -4880 5196 -4832
rect 5808 -4128 6608 -4080
rect 5808 -4832 5856 -4128
rect 6560 -4832 6608 -4128
rect 5808 -4880 6608 -4832
rect 7220 -4128 8020 -4080
rect 7220 -4832 7268 -4128
rect 7972 -4832 8020 -4128
rect 7220 -4880 8020 -4832
rect 8632 -4128 9432 -4080
rect 8632 -4832 8680 -4128
rect 9384 -4832 9432 -4128
rect 8632 -4880 9432 -4832
rect 10044 -4128 10844 -4080
rect 10044 -4832 10092 -4128
rect 10796 -4832 10844 -4128
rect 10044 -4880 10844 -4832
rect 11456 -4128 12256 -4080
rect 11456 -4832 11504 -4128
rect 12208 -4832 12256 -4128
rect 11456 -4880 12256 -4832
rect 12868 -4128 13668 -4080
rect 12868 -4832 12916 -4128
rect 13620 -4832 13668 -4128
rect 12868 -4880 13668 -4832
rect 14280 -4128 15080 -4080
rect 14280 -4832 14328 -4128
rect 15032 -4832 15080 -4128
rect 14280 -4880 15080 -4832
rect 15692 -4128 16492 -4080
rect 15692 -4832 15740 -4128
rect 16444 -4832 16492 -4128
rect 15692 -4880 16492 -4832
rect 17104 -4128 17904 -4080
rect 17104 -4832 17152 -4128
rect 17856 -4832 17904 -4128
rect 17104 -4880 17904 -4832
rect 18516 -4128 19316 -4080
rect 18516 -4832 18564 -4128
rect 19268 -4832 19316 -4128
rect 18516 -4880 19316 -4832
rect 19928 -4128 20728 -4080
rect 19928 -4832 19976 -4128
rect 20680 -4832 20728 -4128
rect 19928 -4880 20728 -4832
rect 21340 -4128 22140 -4080
rect 21340 -4832 21388 -4128
rect 22092 -4832 22140 -4128
rect 21340 -4880 22140 -4832
rect 22752 -4128 23552 -4080
rect 22752 -4832 22800 -4128
rect 23504 -4832 23552 -4128
rect 22752 -4880 23552 -4832
rect -23844 -5248 -23044 -5200
rect -23844 -5952 -23796 -5248
rect -23092 -5952 -23044 -5248
rect -23844 -6000 -23044 -5952
rect -22432 -5248 -21632 -5200
rect -22432 -5952 -22384 -5248
rect -21680 -5952 -21632 -5248
rect -22432 -6000 -21632 -5952
rect -21020 -5248 -20220 -5200
rect -21020 -5952 -20972 -5248
rect -20268 -5952 -20220 -5248
rect -21020 -6000 -20220 -5952
rect -19608 -5248 -18808 -5200
rect -19608 -5952 -19560 -5248
rect -18856 -5952 -18808 -5248
rect -19608 -6000 -18808 -5952
rect -18196 -5248 -17396 -5200
rect -18196 -5952 -18148 -5248
rect -17444 -5952 -17396 -5248
rect -18196 -6000 -17396 -5952
rect -16784 -5248 -15984 -5200
rect -16784 -5952 -16736 -5248
rect -16032 -5952 -15984 -5248
rect -16784 -6000 -15984 -5952
rect -15372 -5248 -14572 -5200
rect -15372 -5952 -15324 -5248
rect -14620 -5952 -14572 -5248
rect -15372 -6000 -14572 -5952
rect -13960 -5248 -13160 -5200
rect -13960 -5952 -13912 -5248
rect -13208 -5952 -13160 -5248
rect -13960 -6000 -13160 -5952
rect -12548 -5248 -11748 -5200
rect -12548 -5952 -12500 -5248
rect -11796 -5952 -11748 -5248
rect -12548 -6000 -11748 -5952
rect -11136 -5248 -10336 -5200
rect -11136 -5952 -11088 -5248
rect -10384 -5952 -10336 -5248
rect -11136 -6000 -10336 -5952
rect -9724 -5248 -8924 -5200
rect -9724 -5952 -9676 -5248
rect -8972 -5952 -8924 -5248
rect -9724 -6000 -8924 -5952
rect -8312 -5248 -7512 -5200
rect -8312 -5952 -8264 -5248
rect -7560 -5952 -7512 -5248
rect -8312 -6000 -7512 -5952
rect -6900 -5248 -6100 -5200
rect -6900 -5952 -6852 -5248
rect -6148 -5952 -6100 -5248
rect -6900 -6000 -6100 -5952
rect -5488 -5248 -4688 -5200
rect -5488 -5952 -5440 -5248
rect -4736 -5952 -4688 -5248
rect -5488 -6000 -4688 -5952
rect -4076 -5248 -3276 -5200
rect -4076 -5952 -4028 -5248
rect -3324 -5952 -3276 -5248
rect -4076 -6000 -3276 -5952
rect -2664 -5248 -1864 -5200
rect -2664 -5952 -2616 -5248
rect -1912 -5952 -1864 -5248
rect -2664 -6000 -1864 -5952
rect -1252 -5248 -452 -5200
rect -1252 -5952 -1204 -5248
rect -500 -5952 -452 -5248
rect -1252 -6000 -452 -5952
rect 160 -5248 960 -5200
rect 160 -5952 208 -5248
rect 912 -5952 960 -5248
rect 160 -6000 960 -5952
rect 1572 -5248 2372 -5200
rect 1572 -5952 1620 -5248
rect 2324 -5952 2372 -5248
rect 1572 -6000 2372 -5952
rect 2984 -5248 3784 -5200
rect 2984 -5952 3032 -5248
rect 3736 -5952 3784 -5248
rect 2984 -6000 3784 -5952
rect 4396 -5248 5196 -5200
rect 4396 -5952 4444 -5248
rect 5148 -5952 5196 -5248
rect 4396 -6000 5196 -5952
rect 5808 -5248 6608 -5200
rect 5808 -5952 5856 -5248
rect 6560 -5952 6608 -5248
rect 5808 -6000 6608 -5952
rect 7220 -5248 8020 -5200
rect 7220 -5952 7268 -5248
rect 7972 -5952 8020 -5248
rect 7220 -6000 8020 -5952
rect 8632 -5248 9432 -5200
rect 8632 -5952 8680 -5248
rect 9384 -5952 9432 -5248
rect 8632 -6000 9432 -5952
rect 10044 -5248 10844 -5200
rect 10044 -5952 10092 -5248
rect 10796 -5952 10844 -5248
rect 10044 -6000 10844 -5952
rect 11456 -5248 12256 -5200
rect 11456 -5952 11504 -5248
rect 12208 -5952 12256 -5248
rect 11456 -6000 12256 -5952
rect 12868 -5248 13668 -5200
rect 12868 -5952 12916 -5248
rect 13620 -5952 13668 -5248
rect 12868 -6000 13668 -5952
rect 14280 -5248 15080 -5200
rect 14280 -5952 14328 -5248
rect 15032 -5952 15080 -5248
rect 14280 -6000 15080 -5952
rect 15692 -5248 16492 -5200
rect 15692 -5952 15740 -5248
rect 16444 -5952 16492 -5248
rect 15692 -6000 16492 -5952
rect 17104 -5248 17904 -5200
rect 17104 -5952 17152 -5248
rect 17856 -5952 17904 -5248
rect 17104 -6000 17904 -5952
rect 18516 -5248 19316 -5200
rect 18516 -5952 18564 -5248
rect 19268 -5952 19316 -5248
rect 18516 -6000 19316 -5952
rect 19928 -5248 20728 -5200
rect 19928 -5952 19976 -5248
rect 20680 -5952 20728 -5248
rect 19928 -6000 20728 -5952
rect 21340 -5248 22140 -5200
rect 21340 -5952 21388 -5248
rect 22092 -5952 22140 -5248
rect 21340 -6000 22140 -5952
rect 22752 -5248 23552 -5200
rect 22752 -5952 22800 -5248
rect 23504 -5952 23552 -5248
rect 22752 -6000 23552 -5952
rect -23844 -6368 -23044 -6320
rect -23844 -7072 -23796 -6368
rect -23092 -7072 -23044 -6368
rect -23844 -7120 -23044 -7072
rect -22432 -6368 -21632 -6320
rect -22432 -7072 -22384 -6368
rect -21680 -7072 -21632 -6368
rect -22432 -7120 -21632 -7072
rect -21020 -6368 -20220 -6320
rect -21020 -7072 -20972 -6368
rect -20268 -7072 -20220 -6368
rect -21020 -7120 -20220 -7072
rect -19608 -6368 -18808 -6320
rect -19608 -7072 -19560 -6368
rect -18856 -7072 -18808 -6368
rect -19608 -7120 -18808 -7072
rect -18196 -6368 -17396 -6320
rect -18196 -7072 -18148 -6368
rect -17444 -7072 -17396 -6368
rect -18196 -7120 -17396 -7072
rect -16784 -6368 -15984 -6320
rect -16784 -7072 -16736 -6368
rect -16032 -7072 -15984 -6368
rect -16784 -7120 -15984 -7072
rect -15372 -6368 -14572 -6320
rect -15372 -7072 -15324 -6368
rect -14620 -7072 -14572 -6368
rect -15372 -7120 -14572 -7072
rect -13960 -6368 -13160 -6320
rect -13960 -7072 -13912 -6368
rect -13208 -7072 -13160 -6368
rect -13960 -7120 -13160 -7072
rect -12548 -6368 -11748 -6320
rect -12548 -7072 -12500 -6368
rect -11796 -7072 -11748 -6368
rect -12548 -7120 -11748 -7072
rect -11136 -6368 -10336 -6320
rect -11136 -7072 -11088 -6368
rect -10384 -7072 -10336 -6368
rect -11136 -7120 -10336 -7072
rect -9724 -6368 -8924 -6320
rect -9724 -7072 -9676 -6368
rect -8972 -7072 -8924 -6368
rect -9724 -7120 -8924 -7072
rect -8312 -6368 -7512 -6320
rect -8312 -7072 -8264 -6368
rect -7560 -7072 -7512 -6368
rect -8312 -7120 -7512 -7072
rect -6900 -6368 -6100 -6320
rect -6900 -7072 -6852 -6368
rect -6148 -7072 -6100 -6368
rect -6900 -7120 -6100 -7072
rect -5488 -6368 -4688 -6320
rect -5488 -7072 -5440 -6368
rect -4736 -7072 -4688 -6368
rect -5488 -7120 -4688 -7072
rect -4076 -6368 -3276 -6320
rect -4076 -7072 -4028 -6368
rect -3324 -7072 -3276 -6368
rect -4076 -7120 -3276 -7072
rect -2664 -6368 -1864 -6320
rect -2664 -7072 -2616 -6368
rect -1912 -7072 -1864 -6368
rect -2664 -7120 -1864 -7072
rect -1252 -6368 -452 -6320
rect -1252 -7072 -1204 -6368
rect -500 -7072 -452 -6368
rect -1252 -7120 -452 -7072
rect 160 -6368 960 -6320
rect 160 -7072 208 -6368
rect 912 -7072 960 -6368
rect 160 -7120 960 -7072
rect 1572 -6368 2372 -6320
rect 1572 -7072 1620 -6368
rect 2324 -7072 2372 -6368
rect 1572 -7120 2372 -7072
rect 2984 -6368 3784 -6320
rect 2984 -7072 3032 -6368
rect 3736 -7072 3784 -6368
rect 2984 -7120 3784 -7072
rect 4396 -6368 5196 -6320
rect 4396 -7072 4444 -6368
rect 5148 -7072 5196 -6368
rect 4396 -7120 5196 -7072
rect 5808 -6368 6608 -6320
rect 5808 -7072 5856 -6368
rect 6560 -7072 6608 -6368
rect 5808 -7120 6608 -7072
rect 7220 -6368 8020 -6320
rect 7220 -7072 7268 -6368
rect 7972 -7072 8020 -6368
rect 7220 -7120 8020 -7072
rect 8632 -6368 9432 -6320
rect 8632 -7072 8680 -6368
rect 9384 -7072 9432 -6368
rect 8632 -7120 9432 -7072
rect 10044 -6368 10844 -6320
rect 10044 -7072 10092 -6368
rect 10796 -7072 10844 -6368
rect 10044 -7120 10844 -7072
rect 11456 -6368 12256 -6320
rect 11456 -7072 11504 -6368
rect 12208 -7072 12256 -6368
rect 11456 -7120 12256 -7072
rect 12868 -6368 13668 -6320
rect 12868 -7072 12916 -6368
rect 13620 -7072 13668 -6368
rect 12868 -7120 13668 -7072
rect 14280 -6368 15080 -6320
rect 14280 -7072 14328 -6368
rect 15032 -7072 15080 -6368
rect 14280 -7120 15080 -7072
rect 15692 -6368 16492 -6320
rect 15692 -7072 15740 -6368
rect 16444 -7072 16492 -6368
rect 15692 -7120 16492 -7072
rect 17104 -6368 17904 -6320
rect 17104 -7072 17152 -6368
rect 17856 -7072 17904 -6368
rect 17104 -7120 17904 -7072
rect 18516 -6368 19316 -6320
rect 18516 -7072 18564 -6368
rect 19268 -7072 19316 -6368
rect 18516 -7120 19316 -7072
rect 19928 -6368 20728 -6320
rect 19928 -7072 19976 -6368
rect 20680 -7072 20728 -6368
rect 19928 -7120 20728 -7072
rect 21340 -6368 22140 -6320
rect 21340 -7072 21388 -6368
rect 22092 -7072 22140 -6368
rect 21340 -7120 22140 -7072
rect 22752 -6368 23552 -6320
rect 22752 -7072 22800 -6368
rect 23504 -7072 23552 -6368
rect 22752 -7120 23552 -7072
rect -23844 -7488 -23044 -7440
rect -23844 -8192 -23796 -7488
rect -23092 -8192 -23044 -7488
rect -23844 -8240 -23044 -8192
rect -22432 -7488 -21632 -7440
rect -22432 -8192 -22384 -7488
rect -21680 -8192 -21632 -7488
rect -22432 -8240 -21632 -8192
rect -21020 -7488 -20220 -7440
rect -21020 -8192 -20972 -7488
rect -20268 -8192 -20220 -7488
rect -21020 -8240 -20220 -8192
rect -19608 -7488 -18808 -7440
rect -19608 -8192 -19560 -7488
rect -18856 -8192 -18808 -7488
rect -19608 -8240 -18808 -8192
rect -18196 -7488 -17396 -7440
rect -18196 -8192 -18148 -7488
rect -17444 -8192 -17396 -7488
rect -18196 -8240 -17396 -8192
rect -16784 -7488 -15984 -7440
rect -16784 -8192 -16736 -7488
rect -16032 -8192 -15984 -7488
rect -16784 -8240 -15984 -8192
rect -15372 -7488 -14572 -7440
rect -15372 -8192 -15324 -7488
rect -14620 -8192 -14572 -7488
rect -15372 -8240 -14572 -8192
rect -13960 -7488 -13160 -7440
rect -13960 -8192 -13912 -7488
rect -13208 -8192 -13160 -7488
rect -13960 -8240 -13160 -8192
rect -12548 -7488 -11748 -7440
rect -12548 -8192 -12500 -7488
rect -11796 -8192 -11748 -7488
rect -12548 -8240 -11748 -8192
rect -11136 -7488 -10336 -7440
rect -11136 -8192 -11088 -7488
rect -10384 -8192 -10336 -7488
rect -11136 -8240 -10336 -8192
rect -9724 -7488 -8924 -7440
rect -9724 -8192 -9676 -7488
rect -8972 -8192 -8924 -7488
rect -9724 -8240 -8924 -8192
rect -8312 -7488 -7512 -7440
rect -8312 -8192 -8264 -7488
rect -7560 -8192 -7512 -7488
rect -8312 -8240 -7512 -8192
rect -6900 -7488 -6100 -7440
rect -6900 -8192 -6852 -7488
rect -6148 -8192 -6100 -7488
rect -6900 -8240 -6100 -8192
rect -5488 -7488 -4688 -7440
rect -5488 -8192 -5440 -7488
rect -4736 -8192 -4688 -7488
rect -5488 -8240 -4688 -8192
rect -4076 -7488 -3276 -7440
rect -4076 -8192 -4028 -7488
rect -3324 -8192 -3276 -7488
rect -4076 -8240 -3276 -8192
rect -2664 -7488 -1864 -7440
rect -2664 -8192 -2616 -7488
rect -1912 -8192 -1864 -7488
rect -2664 -8240 -1864 -8192
rect -1252 -7488 -452 -7440
rect -1252 -8192 -1204 -7488
rect -500 -8192 -452 -7488
rect -1252 -8240 -452 -8192
rect 160 -7488 960 -7440
rect 160 -8192 208 -7488
rect 912 -8192 960 -7488
rect 160 -8240 960 -8192
rect 1572 -7488 2372 -7440
rect 1572 -8192 1620 -7488
rect 2324 -8192 2372 -7488
rect 1572 -8240 2372 -8192
rect 2984 -7488 3784 -7440
rect 2984 -8192 3032 -7488
rect 3736 -8192 3784 -7488
rect 2984 -8240 3784 -8192
rect 4396 -7488 5196 -7440
rect 4396 -8192 4444 -7488
rect 5148 -8192 5196 -7488
rect 4396 -8240 5196 -8192
rect 5808 -7488 6608 -7440
rect 5808 -8192 5856 -7488
rect 6560 -8192 6608 -7488
rect 5808 -8240 6608 -8192
rect 7220 -7488 8020 -7440
rect 7220 -8192 7268 -7488
rect 7972 -8192 8020 -7488
rect 7220 -8240 8020 -8192
rect 8632 -7488 9432 -7440
rect 8632 -8192 8680 -7488
rect 9384 -8192 9432 -7488
rect 8632 -8240 9432 -8192
rect 10044 -7488 10844 -7440
rect 10044 -8192 10092 -7488
rect 10796 -8192 10844 -7488
rect 10044 -8240 10844 -8192
rect 11456 -7488 12256 -7440
rect 11456 -8192 11504 -7488
rect 12208 -8192 12256 -7488
rect 11456 -8240 12256 -8192
rect 12868 -7488 13668 -7440
rect 12868 -8192 12916 -7488
rect 13620 -8192 13668 -7488
rect 12868 -8240 13668 -8192
rect 14280 -7488 15080 -7440
rect 14280 -8192 14328 -7488
rect 15032 -8192 15080 -7488
rect 14280 -8240 15080 -8192
rect 15692 -7488 16492 -7440
rect 15692 -8192 15740 -7488
rect 16444 -8192 16492 -7488
rect 15692 -8240 16492 -8192
rect 17104 -7488 17904 -7440
rect 17104 -8192 17152 -7488
rect 17856 -8192 17904 -7488
rect 17104 -8240 17904 -8192
rect 18516 -7488 19316 -7440
rect 18516 -8192 18564 -7488
rect 19268 -8192 19316 -7488
rect 18516 -8240 19316 -8192
rect 19928 -7488 20728 -7440
rect 19928 -8192 19976 -7488
rect 20680 -8192 20728 -7488
rect 19928 -8240 20728 -8192
rect 21340 -7488 22140 -7440
rect 21340 -8192 21388 -7488
rect 22092 -8192 22140 -7488
rect 21340 -8240 22140 -8192
rect 22752 -7488 23552 -7440
rect 22752 -8192 22800 -7488
rect 23504 -8192 23552 -7488
rect 22752 -8240 23552 -8192
rect -23844 -8608 -23044 -8560
rect -23844 -9312 -23796 -8608
rect -23092 -9312 -23044 -8608
rect -23844 -9360 -23044 -9312
rect -22432 -8608 -21632 -8560
rect -22432 -9312 -22384 -8608
rect -21680 -9312 -21632 -8608
rect -22432 -9360 -21632 -9312
rect -21020 -8608 -20220 -8560
rect -21020 -9312 -20972 -8608
rect -20268 -9312 -20220 -8608
rect -21020 -9360 -20220 -9312
rect -19608 -8608 -18808 -8560
rect -19608 -9312 -19560 -8608
rect -18856 -9312 -18808 -8608
rect -19608 -9360 -18808 -9312
rect -18196 -8608 -17396 -8560
rect -18196 -9312 -18148 -8608
rect -17444 -9312 -17396 -8608
rect -18196 -9360 -17396 -9312
rect -16784 -8608 -15984 -8560
rect -16784 -9312 -16736 -8608
rect -16032 -9312 -15984 -8608
rect -16784 -9360 -15984 -9312
rect -15372 -8608 -14572 -8560
rect -15372 -9312 -15324 -8608
rect -14620 -9312 -14572 -8608
rect -15372 -9360 -14572 -9312
rect -13960 -8608 -13160 -8560
rect -13960 -9312 -13912 -8608
rect -13208 -9312 -13160 -8608
rect -13960 -9360 -13160 -9312
rect -12548 -8608 -11748 -8560
rect -12548 -9312 -12500 -8608
rect -11796 -9312 -11748 -8608
rect -12548 -9360 -11748 -9312
rect -11136 -8608 -10336 -8560
rect -11136 -9312 -11088 -8608
rect -10384 -9312 -10336 -8608
rect -11136 -9360 -10336 -9312
rect -9724 -8608 -8924 -8560
rect -9724 -9312 -9676 -8608
rect -8972 -9312 -8924 -8608
rect -9724 -9360 -8924 -9312
rect -8312 -8608 -7512 -8560
rect -8312 -9312 -8264 -8608
rect -7560 -9312 -7512 -8608
rect -8312 -9360 -7512 -9312
rect -6900 -8608 -6100 -8560
rect -6900 -9312 -6852 -8608
rect -6148 -9312 -6100 -8608
rect -6900 -9360 -6100 -9312
rect -5488 -8608 -4688 -8560
rect -5488 -9312 -5440 -8608
rect -4736 -9312 -4688 -8608
rect -5488 -9360 -4688 -9312
rect -4076 -8608 -3276 -8560
rect -4076 -9312 -4028 -8608
rect -3324 -9312 -3276 -8608
rect -4076 -9360 -3276 -9312
rect -2664 -8608 -1864 -8560
rect -2664 -9312 -2616 -8608
rect -1912 -9312 -1864 -8608
rect -2664 -9360 -1864 -9312
rect -1252 -8608 -452 -8560
rect -1252 -9312 -1204 -8608
rect -500 -9312 -452 -8608
rect -1252 -9360 -452 -9312
rect 160 -8608 960 -8560
rect 160 -9312 208 -8608
rect 912 -9312 960 -8608
rect 160 -9360 960 -9312
rect 1572 -8608 2372 -8560
rect 1572 -9312 1620 -8608
rect 2324 -9312 2372 -8608
rect 1572 -9360 2372 -9312
rect 2984 -8608 3784 -8560
rect 2984 -9312 3032 -8608
rect 3736 -9312 3784 -8608
rect 2984 -9360 3784 -9312
rect 4396 -8608 5196 -8560
rect 4396 -9312 4444 -8608
rect 5148 -9312 5196 -8608
rect 4396 -9360 5196 -9312
rect 5808 -8608 6608 -8560
rect 5808 -9312 5856 -8608
rect 6560 -9312 6608 -8608
rect 5808 -9360 6608 -9312
rect 7220 -8608 8020 -8560
rect 7220 -9312 7268 -8608
rect 7972 -9312 8020 -8608
rect 7220 -9360 8020 -9312
rect 8632 -8608 9432 -8560
rect 8632 -9312 8680 -8608
rect 9384 -9312 9432 -8608
rect 8632 -9360 9432 -9312
rect 10044 -8608 10844 -8560
rect 10044 -9312 10092 -8608
rect 10796 -9312 10844 -8608
rect 10044 -9360 10844 -9312
rect 11456 -8608 12256 -8560
rect 11456 -9312 11504 -8608
rect 12208 -9312 12256 -8608
rect 11456 -9360 12256 -9312
rect 12868 -8608 13668 -8560
rect 12868 -9312 12916 -8608
rect 13620 -9312 13668 -8608
rect 12868 -9360 13668 -9312
rect 14280 -8608 15080 -8560
rect 14280 -9312 14328 -8608
rect 15032 -9312 15080 -8608
rect 14280 -9360 15080 -9312
rect 15692 -8608 16492 -8560
rect 15692 -9312 15740 -8608
rect 16444 -9312 16492 -8608
rect 15692 -9360 16492 -9312
rect 17104 -8608 17904 -8560
rect 17104 -9312 17152 -8608
rect 17856 -9312 17904 -8608
rect 17104 -9360 17904 -9312
rect 18516 -8608 19316 -8560
rect 18516 -9312 18564 -8608
rect 19268 -9312 19316 -8608
rect 18516 -9360 19316 -9312
rect 19928 -8608 20728 -8560
rect 19928 -9312 19976 -8608
rect 20680 -9312 20728 -8608
rect 19928 -9360 20728 -9312
rect 21340 -8608 22140 -8560
rect 21340 -9312 21388 -8608
rect 22092 -9312 22140 -8608
rect 21340 -9360 22140 -9312
rect 22752 -8608 23552 -8560
rect 22752 -9312 22800 -8608
rect 23504 -9312 23552 -8608
rect 22752 -9360 23552 -9312
rect -23844 -9728 -23044 -9680
rect -23844 -10432 -23796 -9728
rect -23092 -10432 -23044 -9728
rect -23844 -10480 -23044 -10432
rect -22432 -9728 -21632 -9680
rect -22432 -10432 -22384 -9728
rect -21680 -10432 -21632 -9728
rect -22432 -10480 -21632 -10432
rect -21020 -9728 -20220 -9680
rect -21020 -10432 -20972 -9728
rect -20268 -10432 -20220 -9728
rect -21020 -10480 -20220 -10432
rect -19608 -9728 -18808 -9680
rect -19608 -10432 -19560 -9728
rect -18856 -10432 -18808 -9728
rect -19608 -10480 -18808 -10432
rect -18196 -9728 -17396 -9680
rect -18196 -10432 -18148 -9728
rect -17444 -10432 -17396 -9728
rect -18196 -10480 -17396 -10432
rect -16784 -9728 -15984 -9680
rect -16784 -10432 -16736 -9728
rect -16032 -10432 -15984 -9728
rect -16784 -10480 -15984 -10432
rect -15372 -9728 -14572 -9680
rect -15372 -10432 -15324 -9728
rect -14620 -10432 -14572 -9728
rect -15372 -10480 -14572 -10432
rect -13960 -9728 -13160 -9680
rect -13960 -10432 -13912 -9728
rect -13208 -10432 -13160 -9728
rect -13960 -10480 -13160 -10432
rect -12548 -9728 -11748 -9680
rect -12548 -10432 -12500 -9728
rect -11796 -10432 -11748 -9728
rect -12548 -10480 -11748 -10432
rect -11136 -9728 -10336 -9680
rect -11136 -10432 -11088 -9728
rect -10384 -10432 -10336 -9728
rect -11136 -10480 -10336 -10432
rect -9724 -9728 -8924 -9680
rect -9724 -10432 -9676 -9728
rect -8972 -10432 -8924 -9728
rect -9724 -10480 -8924 -10432
rect -8312 -9728 -7512 -9680
rect -8312 -10432 -8264 -9728
rect -7560 -10432 -7512 -9728
rect -8312 -10480 -7512 -10432
rect -6900 -9728 -6100 -9680
rect -6900 -10432 -6852 -9728
rect -6148 -10432 -6100 -9728
rect -6900 -10480 -6100 -10432
rect -5488 -9728 -4688 -9680
rect -5488 -10432 -5440 -9728
rect -4736 -10432 -4688 -9728
rect -5488 -10480 -4688 -10432
rect -4076 -9728 -3276 -9680
rect -4076 -10432 -4028 -9728
rect -3324 -10432 -3276 -9728
rect -4076 -10480 -3276 -10432
rect -2664 -9728 -1864 -9680
rect -2664 -10432 -2616 -9728
rect -1912 -10432 -1864 -9728
rect -2664 -10480 -1864 -10432
rect -1252 -9728 -452 -9680
rect -1252 -10432 -1204 -9728
rect -500 -10432 -452 -9728
rect -1252 -10480 -452 -10432
rect 160 -9728 960 -9680
rect 160 -10432 208 -9728
rect 912 -10432 960 -9728
rect 160 -10480 960 -10432
rect 1572 -9728 2372 -9680
rect 1572 -10432 1620 -9728
rect 2324 -10432 2372 -9728
rect 1572 -10480 2372 -10432
rect 2984 -9728 3784 -9680
rect 2984 -10432 3032 -9728
rect 3736 -10432 3784 -9728
rect 2984 -10480 3784 -10432
rect 4396 -9728 5196 -9680
rect 4396 -10432 4444 -9728
rect 5148 -10432 5196 -9728
rect 4396 -10480 5196 -10432
rect 5808 -9728 6608 -9680
rect 5808 -10432 5856 -9728
rect 6560 -10432 6608 -9728
rect 5808 -10480 6608 -10432
rect 7220 -9728 8020 -9680
rect 7220 -10432 7268 -9728
rect 7972 -10432 8020 -9728
rect 7220 -10480 8020 -10432
rect 8632 -9728 9432 -9680
rect 8632 -10432 8680 -9728
rect 9384 -10432 9432 -9728
rect 8632 -10480 9432 -10432
rect 10044 -9728 10844 -9680
rect 10044 -10432 10092 -9728
rect 10796 -10432 10844 -9728
rect 10044 -10480 10844 -10432
rect 11456 -9728 12256 -9680
rect 11456 -10432 11504 -9728
rect 12208 -10432 12256 -9728
rect 11456 -10480 12256 -10432
rect 12868 -9728 13668 -9680
rect 12868 -10432 12916 -9728
rect 13620 -10432 13668 -9728
rect 12868 -10480 13668 -10432
rect 14280 -9728 15080 -9680
rect 14280 -10432 14328 -9728
rect 15032 -10432 15080 -9728
rect 14280 -10480 15080 -10432
rect 15692 -9728 16492 -9680
rect 15692 -10432 15740 -9728
rect 16444 -10432 16492 -9728
rect 15692 -10480 16492 -10432
rect 17104 -9728 17904 -9680
rect 17104 -10432 17152 -9728
rect 17856 -10432 17904 -9728
rect 17104 -10480 17904 -10432
rect 18516 -9728 19316 -9680
rect 18516 -10432 18564 -9728
rect 19268 -10432 19316 -9728
rect 18516 -10480 19316 -10432
rect 19928 -9728 20728 -9680
rect 19928 -10432 19976 -9728
rect 20680 -10432 20728 -9728
rect 19928 -10480 20728 -10432
rect 21340 -9728 22140 -9680
rect 21340 -10432 21388 -9728
rect 22092 -10432 22140 -9728
rect 21340 -10480 22140 -10432
rect 22752 -9728 23552 -9680
rect 22752 -10432 22800 -9728
rect 23504 -10432 23552 -9728
rect 22752 -10480 23552 -10432
rect -23844 -10848 -23044 -10800
rect -23844 -11552 -23796 -10848
rect -23092 -11552 -23044 -10848
rect -23844 -11600 -23044 -11552
rect -22432 -10848 -21632 -10800
rect -22432 -11552 -22384 -10848
rect -21680 -11552 -21632 -10848
rect -22432 -11600 -21632 -11552
rect -21020 -10848 -20220 -10800
rect -21020 -11552 -20972 -10848
rect -20268 -11552 -20220 -10848
rect -21020 -11600 -20220 -11552
rect -19608 -10848 -18808 -10800
rect -19608 -11552 -19560 -10848
rect -18856 -11552 -18808 -10848
rect -19608 -11600 -18808 -11552
rect -18196 -10848 -17396 -10800
rect -18196 -11552 -18148 -10848
rect -17444 -11552 -17396 -10848
rect -18196 -11600 -17396 -11552
rect -16784 -10848 -15984 -10800
rect -16784 -11552 -16736 -10848
rect -16032 -11552 -15984 -10848
rect -16784 -11600 -15984 -11552
rect -15372 -10848 -14572 -10800
rect -15372 -11552 -15324 -10848
rect -14620 -11552 -14572 -10848
rect -15372 -11600 -14572 -11552
rect -13960 -10848 -13160 -10800
rect -13960 -11552 -13912 -10848
rect -13208 -11552 -13160 -10848
rect -13960 -11600 -13160 -11552
rect -12548 -10848 -11748 -10800
rect -12548 -11552 -12500 -10848
rect -11796 -11552 -11748 -10848
rect -12548 -11600 -11748 -11552
rect -11136 -10848 -10336 -10800
rect -11136 -11552 -11088 -10848
rect -10384 -11552 -10336 -10848
rect -11136 -11600 -10336 -11552
rect -9724 -10848 -8924 -10800
rect -9724 -11552 -9676 -10848
rect -8972 -11552 -8924 -10848
rect -9724 -11600 -8924 -11552
rect -8312 -10848 -7512 -10800
rect -8312 -11552 -8264 -10848
rect -7560 -11552 -7512 -10848
rect -8312 -11600 -7512 -11552
rect -6900 -10848 -6100 -10800
rect -6900 -11552 -6852 -10848
rect -6148 -11552 -6100 -10848
rect -6900 -11600 -6100 -11552
rect -5488 -10848 -4688 -10800
rect -5488 -11552 -5440 -10848
rect -4736 -11552 -4688 -10848
rect -5488 -11600 -4688 -11552
rect -4076 -10848 -3276 -10800
rect -4076 -11552 -4028 -10848
rect -3324 -11552 -3276 -10848
rect -4076 -11600 -3276 -11552
rect -2664 -10848 -1864 -10800
rect -2664 -11552 -2616 -10848
rect -1912 -11552 -1864 -10848
rect -2664 -11600 -1864 -11552
rect -1252 -10848 -452 -10800
rect -1252 -11552 -1204 -10848
rect -500 -11552 -452 -10848
rect -1252 -11600 -452 -11552
rect 160 -10848 960 -10800
rect 160 -11552 208 -10848
rect 912 -11552 960 -10848
rect 160 -11600 960 -11552
rect 1572 -10848 2372 -10800
rect 1572 -11552 1620 -10848
rect 2324 -11552 2372 -10848
rect 1572 -11600 2372 -11552
rect 2984 -10848 3784 -10800
rect 2984 -11552 3032 -10848
rect 3736 -11552 3784 -10848
rect 2984 -11600 3784 -11552
rect 4396 -10848 5196 -10800
rect 4396 -11552 4444 -10848
rect 5148 -11552 5196 -10848
rect 4396 -11600 5196 -11552
rect 5808 -10848 6608 -10800
rect 5808 -11552 5856 -10848
rect 6560 -11552 6608 -10848
rect 5808 -11600 6608 -11552
rect 7220 -10848 8020 -10800
rect 7220 -11552 7268 -10848
rect 7972 -11552 8020 -10848
rect 7220 -11600 8020 -11552
rect 8632 -10848 9432 -10800
rect 8632 -11552 8680 -10848
rect 9384 -11552 9432 -10848
rect 8632 -11600 9432 -11552
rect 10044 -10848 10844 -10800
rect 10044 -11552 10092 -10848
rect 10796 -11552 10844 -10848
rect 10044 -11600 10844 -11552
rect 11456 -10848 12256 -10800
rect 11456 -11552 11504 -10848
rect 12208 -11552 12256 -10848
rect 11456 -11600 12256 -11552
rect 12868 -10848 13668 -10800
rect 12868 -11552 12916 -10848
rect 13620 -11552 13668 -10848
rect 12868 -11600 13668 -11552
rect 14280 -10848 15080 -10800
rect 14280 -11552 14328 -10848
rect 15032 -11552 15080 -10848
rect 14280 -11600 15080 -11552
rect 15692 -10848 16492 -10800
rect 15692 -11552 15740 -10848
rect 16444 -11552 16492 -10848
rect 15692 -11600 16492 -11552
rect 17104 -10848 17904 -10800
rect 17104 -11552 17152 -10848
rect 17856 -11552 17904 -10848
rect 17104 -11600 17904 -11552
rect 18516 -10848 19316 -10800
rect 18516 -11552 18564 -10848
rect 19268 -11552 19316 -10848
rect 18516 -11600 19316 -11552
rect 19928 -10848 20728 -10800
rect 19928 -11552 19976 -10848
rect 20680 -11552 20728 -10848
rect 19928 -11600 20728 -11552
rect 21340 -10848 22140 -10800
rect 21340 -11552 21388 -10848
rect 22092 -11552 22140 -10848
rect 21340 -11600 22140 -11552
rect 22752 -10848 23552 -10800
rect 22752 -11552 22800 -10848
rect 23504 -11552 23552 -10848
rect 22752 -11600 23552 -11552
rect -23844 -11968 -23044 -11920
rect -23844 -12672 -23796 -11968
rect -23092 -12672 -23044 -11968
rect -23844 -12720 -23044 -12672
rect -22432 -11968 -21632 -11920
rect -22432 -12672 -22384 -11968
rect -21680 -12672 -21632 -11968
rect -22432 -12720 -21632 -12672
rect -21020 -11968 -20220 -11920
rect -21020 -12672 -20972 -11968
rect -20268 -12672 -20220 -11968
rect -21020 -12720 -20220 -12672
rect -19608 -11968 -18808 -11920
rect -19608 -12672 -19560 -11968
rect -18856 -12672 -18808 -11968
rect -19608 -12720 -18808 -12672
rect -18196 -11968 -17396 -11920
rect -18196 -12672 -18148 -11968
rect -17444 -12672 -17396 -11968
rect -18196 -12720 -17396 -12672
rect -16784 -11968 -15984 -11920
rect -16784 -12672 -16736 -11968
rect -16032 -12672 -15984 -11968
rect -16784 -12720 -15984 -12672
rect -15372 -11968 -14572 -11920
rect -15372 -12672 -15324 -11968
rect -14620 -12672 -14572 -11968
rect -15372 -12720 -14572 -12672
rect -13960 -11968 -13160 -11920
rect -13960 -12672 -13912 -11968
rect -13208 -12672 -13160 -11968
rect -13960 -12720 -13160 -12672
rect -12548 -11968 -11748 -11920
rect -12548 -12672 -12500 -11968
rect -11796 -12672 -11748 -11968
rect -12548 -12720 -11748 -12672
rect -11136 -11968 -10336 -11920
rect -11136 -12672 -11088 -11968
rect -10384 -12672 -10336 -11968
rect -11136 -12720 -10336 -12672
rect -9724 -11968 -8924 -11920
rect -9724 -12672 -9676 -11968
rect -8972 -12672 -8924 -11968
rect -9724 -12720 -8924 -12672
rect -8312 -11968 -7512 -11920
rect -8312 -12672 -8264 -11968
rect -7560 -12672 -7512 -11968
rect -8312 -12720 -7512 -12672
rect -6900 -11968 -6100 -11920
rect -6900 -12672 -6852 -11968
rect -6148 -12672 -6100 -11968
rect -6900 -12720 -6100 -12672
rect -5488 -11968 -4688 -11920
rect -5488 -12672 -5440 -11968
rect -4736 -12672 -4688 -11968
rect -5488 -12720 -4688 -12672
rect -4076 -11968 -3276 -11920
rect -4076 -12672 -4028 -11968
rect -3324 -12672 -3276 -11968
rect -4076 -12720 -3276 -12672
rect -2664 -11968 -1864 -11920
rect -2664 -12672 -2616 -11968
rect -1912 -12672 -1864 -11968
rect -2664 -12720 -1864 -12672
rect -1252 -11968 -452 -11920
rect -1252 -12672 -1204 -11968
rect -500 -12672 -452 -11968
rect -1252 -12720 -452 -12672
rect 160 -11968 960 -11920
rect 160 -12672 208 -11968
rect 912 -12672 960 -11968
rect 160 -12720 960 -12672
rect 1572 -11968 2372 -11920
rect 1572 -12672 1620 -11968
rect 2324 -12672 2372 -11968
rect 1572 -12720 2372 -12672
rect 2984 -11968 3784 -11920
rect 2984 -12672 3032 -11968
rect 3736 -12672 3784 -11968
rect 2984 -12720 3784 -12672
rect 4396 -11968 5196 -11920
rect 4396 -12672 4444 -11968
rect 5148 -12672 5196 -11968
rect 4396 -12720 5196 -12672
rect 5808 -11968 6608 -11920
rect 5808 -12672 5856 -11968
rect 6560 -12672 6608 -11968
rect 5808 -12720 6608 -12672
rect 7220 -11968 8020 -11920
rect 7220 -12672 7268 -11968
rect 7972 -12672 8020 -11968
rect 7220 -12720 8020 -12672
rect 8632 -11968 9432 -11920
rect 8632 -12672 8680 -11968
rect 9384 -12672 9432 -11968
rect 8632 -12720 9432 -12672
rect 10044 -11968 10844 -11920
rect 10044 -12672 10092 -11968
rect 10796 -12672 10844 -11968
rect 10044 -12720 10844 -12672
rect 11456 -11968 12256 -11920
rect 11456 -12672 11504 -11968
rect 12208 -12672 12256 -11968
rect 11456 -12720 12256 -12672
rect 12868 -11968 13668 -11920
rect 12868 -12672 12916 -11968
rect 13620 -12672 13668 -11968
rect 12868 -12720 13668 -12672
rect 14280 -11968 15080 -11920
rect 14280 -12672 14328 -11968
rect 15032 -12672 15080 -11968
rect 14280 -12720 15080 -12672
rect 15692 -11968 16492 -11920
rect 15692 -12672 15740 -11968
rect 16444 -12672 16492 -11968
rect 15692 -12720 16492 -12672
rect 17104 -11968 17904 -11920
rect 17104 -12672 17152 -11968
rect 17856 -12672 17904 -11968
rect 17104 -12720 17904 -12672
rect 18516 -11968 19316 -11920
rect 18516 -12672 18564 -11968
rect 19268 -12672 19316 -11968
rect 18516 -12720 19316 -12672
rect 19928 -11968 20728 -11920
rect 19928 -12672 19976 -11968
rect 20680 -12672 20728 -11968
rect 19928 -12720 20728 -12672
rect 21340 -11968 22140 -11920
rect 21340 -12672 21388 -11968
rect 22092 -12672 22140 -11968
rect 21340 -12720 22140 -12672
rect 22752 -11968 23552 -11920
rect 22752 -12672 22800 -11968
rect 23504 -12672 23552 -11968
rect 22752 -12720 23552 -12672
rect -23844 -13088 -23044 -13040
rect -23844 -13792 -23796 -13088
rect -23092 -13792 -23044 -13088
rect -23844 -13840 -23044 -13792
rect -22432 -13088 -21632 -13040
rect -22432 -13792 -22384 -13088
rect -21680 -13792 -21632 -13088
rect -22432 -13840 -21632 -13792
rect -21020 -13088 -20220 -13040
rect -21020 -13792 -20972 -13088
rect -20268 -13792 -20220 -13088
rect -21020 -13840 -20220 -13792
rect -19608 -13088 -18808 -13040
rect -19608 -13792 -19560 -13088
rect -18856 -13792 -18808 -13088
rect -19608 -13840 -18808 -13792
rect -18196 -13088 -17396 -13040
rect -18196 -13792 -18148 -13088
rect -17444 -13792 -17396 -13088
rect -18196 -13840 -17396 -13792
rect -16784 -13088 -15984 -13040
rect -16784 -13792 -16736 -13088
rect -16032 -13792 -15984 -13088
rect -16784 -13840 -15984 -13792
rect -15372 -13088 -14572 -13040
rect -15372 -13792 -15324 -13088
rect -14620 -13792 -14572 -13088
rect -15372 -13840 -14572 -13792
rect -13960 -13088 -13160 -13040
rect -13960 -13792 -13912 -13088
rect -13208 -13792 -13160 -13088
rect -13960 -13840 -13160 -13792
rect -12548 -13088 -11748 -13040
rect -12548 -13792 -12500 -13088
rect -11796 -13792 -11748 -13088
rect -12548 -13840 -11748 -13792
rect -11136 -13088 -10336 -13040
rect -11136 -13792 -11088 -13088
rect -10384 -13792 -10336 -13088
rect -11136 -13840 -10336 -13792
rect -9724 -13088 -8924 -13040
rect -9724 -13792 -9676 -13088
rect -8972 -13792 -8924 -13088
rect -9724 -13840 -8924 -13792
rect -8312 -13088 -7512 -13040
rect -8312 -13792 -8264 -13088
rect -7560 -13792 -7512 -13088
rect -8312 -13840 -7512 -13792
rect -6900 -13088 -6100 -13040
rect -6900 -13792 -6852 -13088
rect -6148 -13792 -6100 -13088
rect -6900 -13840 -6100 -13792
rect -5488 -13088 -4688 -13040
rect -5488 -13792 -5440 -13088
rect -4736 -13792 -4688 -13088
rect -5488 -13840 -4688 -13792
rect -4076 -13088 -3276 -13040
rect -4076 -13792 -4028 -13088
rect -3324 -13792 -3276 -13088
rect -4076 -13840 -3276 -13792
rect -2664 -13088 -1864 -13040
rect -2664 -13792 -2616 -13088
rect -1912 -13792 -1864 -13088
rect -2664 -13840 -1864 -13792
rect -1252 -13088 -452 -13040
rect -1252 -13792 -1204 -13088
rect -500 -13792 -452 -13088
rect -1252 -13840 -452 -13792
rect 160 -13088 960 -13040
rect 160 -13792 208 -13088
rect 912 -13792 960 -13088
rect 160 -13840 960 -13792
rect 1572 -13088 2372 -13040
rect 1572 -13792 1620 -13088
rect 2324 -13792 2372 -13088
rect 1572 -13840 2372 -13792
rect 2984 -13088 3784 -13040
rect 2984 -13792 3032 -13088
rect 3736 -13792 3784 -13088
rect 2984 -13840 3784 -13792
rect 4396 -13088 5196 -13040
rect 4396 -13792 4444 -13088
rect 5148 -13792 5196 -13088
rect 4396 -13840 5196 -13792
rect 5808 -13088 6608 -13040
rect 5808 -13792 5856 -13088
rect 6560 -13792 6608 -13088
rect 5808 -13840 6608 -13792
rect 7220 -13088 8020 -13040
rect 7220 -13792 7268 -13088
rect 7972 -13792 8020 -13088
rect 7220 -13840 8020 -13792
rect 8632 -13088 9432 -13040
rect 8632 -13792 8680 -13088
rect 9384 -13792 9432 -13088
rect 8632 -13840 9432 -13792
rect 10044 -13088 10844 -13040
rect 10044 -13792 10092 -13088
rect 10796 -13792 10844 -13088
rect 10044 -13840 10844 -13792
rect 11456 -13088 12256 -13040
rect 11456 -13792 11504 -13088
rect 12208 -13792 12256 -13088
rect 11456 -13840 12256 -13792
rect 12868 -13088 13668 -13040
rect 12868 -13792 12916 -13088
rect 13620 -13792 13668 -13088
rect 12868 -13840 13668 -13792
rect 14280 -13088 15080 -13040
rect 14280 -13792 14328 -13088
rect 15032 -13792 15080 -13088
rect 14280 -13840 15080 -13792
rect 15692 -13088 16492 -13040
rect 15692 -13792 15740 -13088
rect 16444 -13792 16492 -13088
rect 15692 -13840 16492 -13792
rect 17104 -13088 17904 -13040
rect 17104 -13792 17152 -13088
rect 17856 -13792 17904 -13088
rect 17104 -13840 17904 -13792
rect 18516 -13088 19316 -13040
rect 18516 -13792 18564 -13088
rect 19268 -13792 19316 -13088
rect 18516 -13840 19316 -13792
rect 19928 -13088 20728 -13040
rect 19928 -13792 19976 -13088
rect 20680 -13792 20728 -13088
rect 19928 -13840 20728 -13792
rect 21340 -13088 22140 -13040
rect 21340 -13792 21388 -13088
rect 22092 -13792 22140 -13088
rect 21340 -13840 22140 -13792
rect 22752 -13088 23552 -13040
rect 22752 -13792 22800 -13088
rect 23504 -13792 23552 -13088
rect 22752 -13840 23552 -13792
rect -23844 -14208 -23044 -14160
rect -23844 -14912 -23796 -14208
rect -23092 -14912 -23044 -14208
rect -23844 -14960 -23044 -14912
rect -22432 -14208 -21632 -14160
rect -22432 -14912 -22384 -14208
rect -21680 -14912 -21632 -14208
rect -22432 -14960 -21632 -14912
rect -21020 -14208 -20220 -14160
rect -21020 -14912 -20972 -14208
rect -20268 -14912 -20220 -14208
rect -21020 -14960 -20220 -14912
rect -19608 -14208 -18808 -14160
rect -19608 -14912 -19560 -14208
rect -18856 -14912 -18808 -14208
rect -19608 -14960 -18808 -14912
rect -18196 -14208 -17396 -14160
rect -18196 -14912 -18148 -14208
rect -17444 -14912 -17396 -14208
rect -18196 -14960 -17396 -14912
rect -16784 -14208 -15984 -14160
rect -16784 -14912 -16736 -14208
rect -16032 -14912 -15984 -14208
rect -16784 -14960 -15984 -14912
rect -15372 -14208 -14572 -14160
rect -15372 -14912 -15324 -14208
rect -14620 -14912 -14572 -14208
rect -15372 -14960 -14572 -14912
rect -13960 -14208 -13160 -14160
rect -13960 -14912 -13912 -14208
rect -13208 -14912 -13160 -14208
rect -13960 -14960 -13160 -14912
rect -12548 -14208 -11748 -14160
rect -12548 -14912 -12500 -14208
rect -11796 -14912 -11748 -14208
rect -12548 -14960 -11748 -14912
rect -11136 -14208 -10336 -14160
rect -11136 -14912 -11088 -14208
rect -10384 -14912 -10336 -14208
rect -11136 -14960 -10336 -14912
rect -9724 -14208 -8924 -14160
rect -9724 -14912 -9676 -14208
rect -8972 -14912 -8924 -14208
rect -9724 -14960 -8924 -14912
rect -8312 -14208 -7512 -14160
rect -8312 -14912 -8264 -14208
rect -7560 -14912 -7512 -14208
rect -8312 -14960 -7512 -14912
rect -6900 -14208 -6100 -14160
rect -6900 -14912 -6852 -14208
rect -6148 -14912 -6100 -14208
rect -6900 -14960 -6100 -14912
rect -5488 -14208 -4688 -14160
rect -5488 -14912 -5440 -14208
rect -4736 -14912 -4688 -14208
rect -5488 -14960 -4688 -14912
rect -4076 -14208 -3276 -14160
rect -4076 -14912 -4028 -14208
rect -3324 -14912 -3276 -14208
rect -4076 -14960 -3276 -14912
rect -2664 -14208 -1864 -14160
rect -2664 -14912 -2616 -14208
rect -1912 -14912 -1864 -14208
rect -2664 -14960 -1864 -14912
rect -1252 -14208 -452 -14160
rect -1252 -14912 -1204 -14208
rect -500 -14912 -452 -14208
rect -1252 -14960 -452 -14912
rect 160 -14208 960 -14160
rect 160 -14912 208 -14208
rect 912 -14912 960 -14208
rect 160 -14960 960 -14912
rect 1572 -14208 2372 -14160
rect 1572 -14912 1620 -14208
rect 2324 -14912 2372 -14208
rect 1572 -14960 2372 -14912
rect 2984 -14208 3784 -14160
rect 2984 -14912 3032 -14208
rect 3736 -14912 3784 -14208
rect 2984 -14960 3784 -14912
rect 4396 -14208 5196 -14160
rect 4396 -14912 4444 -14208
rect 5148 -14912 5196 -14208
rect 4396 -14960 5196 -14912
rect 5808 -14208 6608 -14160
rect 5808 -14912 5856 -14208
rect 6560 -14912 6608 -14208
rect 5808 -14960 6608 -14912
rect 7220 -14208 8020 -14160
rect 7220 -14912 7268 -14208
rect 7972 -14912 8020 -14208
rect 7220 -14960 8020 -14912
rect 8632 -14208 9432 -14160
rect 8632 -14912 8680 -14208
rect 9384 -14912 9432 -14208
rect 8632 -14960 9432 -14912
rect 10044 -14208 10844 -14160
rect 10044 -14912 10092 -14208
rect 10796 -14912 10844 -14208
rect 10044 -14960 10844 -14912
rect 11456 -14208 12256 -14160
rect 11456 -14912 11504 -14208
rect 12208 -14912 12256 -14208
rect 11456 -14960 12256 -14912
rect 12868 -14208 13668 -14160
rect 12868 -14912 12916 -14208
rect 13620 -14912 13668 -14208
rect 12868 -14960 13668 -14912
rect 14280 -14208 15080 -14160
rect 14280 -14912 14328 -14208
rect 15032 -14912 15080 -14208
rect 14280 -14960 15080 -14912
rect 15692 -14208 16492 -14160
rect 15692 -14912 15740 -14208
rect 16444 -14912 16492 -14208
rect 15692 -14960 16492 -14912
rect 17104 -14208 17904 -14160
rect 17104 -14912 17152 -14208
rect 17856 -14912 17904 -14208
rect 17104 -14960 17904 -14912
rect 18516 -14208 19316 -14160
rect 18516 -14912 18564 -14208
rect 19268 -14912 19316 -14208
rect 18516 -14960 19316 -14912
rect 19928 -14208 20728 -14160
rect 19928 -14912 19976 -14208
rect 20680 -14912 20728 -14208
rect 19928 -14960 20728 -14912
rect 21340 -14208 22140 -14160
rect 21340 -14912 21388 -14208
rect 22092 -14912 22140 -14208
rect 21340 -14960 22140 -14912
rect 22752 -14208 23552 -14160
rect 22752 -14912 22800 -14208
rect 23504 -14912 23552 -14208
rect 22752 -14960 23552 -14912
rect -23844 -15328 -23044 -15280
rect -23844 -16032 -23796 -15328
rect -23092 -16032 -23044 -15328
rect -23844 -16080 -23044 -16032
rect -22432 -15328 -21632 -15280
rect -22432 -16032 -22384 -15328
rect -21680 -16032 -21632 -15328
rect -22432 -16080 -21632 -16032
rect -21020 -15328 -20220 -15280
rect -21020 -16032 -20972 -15328
rect -20268 -16032 -20220 -15328
rect -21020 -16080 -20220 -16032
rect -19608 -15328 -18808 -15280
rect -19608 -16032 -19560 -15328
rect -18856 -16032 -18808 -15328
rect -19608 -16080 -18808 -16032
rect -18196 -15328 -17396 -15280
rect -18196 -16032 -18148 -15328
rect -17444 -16032 -17396 -15328
rect -18196 -16080 -17396 -16032
rect -16784 -15328 -15984 -15280
rect -16784 -16032 -16736 -15328
rect -16032 -16032 -15984 -15328
rect -16784 -16080 -15984 -16032
rect -15372 -15328 -14572 -15280
rect -15372 -16032 -15324 -15328
rect -14620 -16032 -14572 -15328
rect -15372 -16080 -14572 -16032
rect -13960 -15328 -13160 -15280
rect -13960 -16032 -13912 -15328
rect -13208 -16032 -13160 -15328
rect -13960 -16080 -13160 -16032
rect -12548 -15328 -11748 -15280
rect -12548 -16032 -12500 -15328
rect -11796 -16032 -11748 -15328
rect -12548 -16080 -11748 -16032
rect -11136 -15328 -10336 -15280
rect -11136 -16032 -11088 -15328
rect -10384 -16032 -10336 -15328
rect -11136 -16080 -10336 -16032
rect -9724 -15328 -8924 -15280
rect -9724 -16032 -9676 -15328
rect -8972 -16032 -8924 -15328
rect -9724 -16080 -8924 -16032
rect -8312 -15328 -7512 -15280
rect -8312 -16032 -8264 -15328
rect -7560 -16032 -7512 -15328
rect -8312 -16080 -7512 -16032
rect -6900 -15328 -6100 -15280
rect -6900 -16032 -6852 -15328
rect -6148 -16032 -6100 -15328
rect -6900 -16080 -6100 -16032
rect -5488 -15328 -4688 -15280
rect -5488 -16032 -5440 -15328
rect -4736 -16032 -4688 -15328
rect -5488 -16080 -4688 -16032
rect -4076 -15328 -3276 -15280
rect -4076 -16032 -4028 -15328
rect -3324 -16032 -3276 -15328
rect -4076 -16080 -3276 -16032
rect -2664 -15328 -1864 -15280
rect -2664 -16032 -2616 -15328
rect -1912 -16032 -1864 -15328
rect -2664 -16080 -1864 -16032
rect -1252 -15328 -452 -15280
rect -1252 -16032 -1204 -15328
rect -500 -16032 -452 -15328
rect -1252 -16080 -452 -16032
rect 160 -15328 960 -15280
rect 160 -16032 208 -15328
rect 912 -16032 960 -15328
rect 160 -16080 960 -16032
rect 1572 -15328 2372 -15280
rect 1572 -16032 1620 -15328
rect 2324 -16032 2372 -15328
rect 1572 -16080 2372 -16032
rect 2984 -15328 3784 -15280
rect 2984 -16032 3032 -15328
rect 3736 -16032 3784 -15328
rect 2984 -16080 3784 -16032
rect 4396 -15328 5196 -15280
rect 4396 -16032 4444 -15328
rect 5148 -16032 5196 -15328
rect 4396 -16080 5196 -16032
rect 5808 -15328 6608 -15280
rect 5808 -16032 5856 -15328
rect 6560 -16032 6608 -15328
rect 5808 -16080 6608 -16032
rect 7220 -15328 8020 -15280
rect 7220 -16032 7268 -15328
rect 7972 -16032 8020 -15328
rect 7220 -16080 8020 -16032
rect 8632 -15328 9432 -15280
rect 8632 -16032 8680 -15328
rect 9384 -16032 9432 -15328
rect 8632 -16080 9432 -16032
rect 10044 -15328 10844 -15280
rect 10044 -16032 10092 -15328
rect 10796 -16032 10844 -15328
rect 10044 -16080 10844 -16032
rect 11456 -15328 12256 -15280
rect 11456 -16032 11504 -15328
rect 12208 -16032 12256 -15328
rect 11456 -16080 12256 -16032
rect 12868 -15328 13668 -15280
rect 12868 -16032 12916 -15328
rect 13620 -16032 13668 -15328
rect 12868 -16080 13668 -16032
rect 14280 -15328 15080 -15280
rect 14280 -16032 14328 -15328
rect 15032 -16032 15080 -15328
rect 14280 -16080 15080 -16032
rect 15692 -15328 16492 -15280
rect 15692 -16032 15740 -15328
rect 16444 -16032 16492 -15328
rect 15692 -16080 16492 -16032
rect 17104 -15328 17904 -15280
rect 17104 -16032 17152 -15328
rect 17856 -16032 17904 -15328
rect 17104 -16080 17904 -16032
rect 18516 -15328 19316 -15280
rect 18516 -16032 18564 -15328
rect 19268 -16032 19316 -15328
rect 18516 -16080 19316 -16032
rect 19928 -15328 20728 -15280
rect 19928 -16032 19976 -15328
rect 20680 -16032 20728 -15328
rect 19928 -16080 20728 -16032
rect 21340 -15328 22140 -15280
rect 21340 -16032 21388 -15328
rect 22092 -16032 22140 -15328
rect 21340 -16080 22140 -16032
rect 22752 -15328 23552 -15280
rect 22752 -16032 22800 -15328
rect 23504 -16032 23552 -15328
rect 22752 -16080 23552 -16032
rect -23844 -16448 -23044 -16400
rect -23844 -17152 -23796 -16448
rect -23092 -17152 -23044 -16448
rect -23844 -17200 -23044 -17152
rect -22432 -16448 -21632 -16400
rect -22432 -17152 -22384 -16448
rect -21680 -17152 -21632 -16448
rect -22432 -17200 -21632 -17152
rect -21020 -16448 -20220 -16400
rect -21020 -17152 -20972 -16448
rect -20268 -17152 -20220 -16448
rect -21020 -17200 -20220 -17152
rect -19608 -16448 -18808 -16400
rect -19608 -17152 -19560 -16448
rect -18856 -17152 -18808 -16448
rect -19608 -17200 -18808 -17152
rect -18196 -16448 -17396 -16400
rect -18196 -17152 -18148 -16448
rect -17444 -17152 -17396 -16448
rect -18196 -17200 -17396 -17152
rect -16784 -16448 -15984 -16400
rect -16784 -17152 -16736 -16448
rect -16032 -17152 -15984 -16448
rect -16784 -17200 -15984 -17152
rect -15372 -16448 -14572 -16400
rect -15372 -17152 -15324 -16448
rect -14620 -17152 -14572 -16448
rect -15372 -17200 -14572 -17152
rect -13960 -16448 -13160 -16400
rect -13960 -17152 -13912 -16448
rect -13208 -17152 -13160 -16448
rect -13960 -17200 -13160 -17152
rect -12548 -16448 -11748 -16400
rect -12548 -17152 -12500 -16448
rect -11796 -17152 -11748 -16448
rect -12548 -17200 -11748 -17152
rect -11136 -16448 -10336 -16400
rect -11136 -17152 -11088 -16448
rect -10384 -17152 -10336 -16448
rect -11136 -17200 -10336 -17152
rect -9724 -16448 -8924 -16400
rect -9724 -17152 -9676 -16448
rect -8972 -17152 -8924 -16448
rect -9724 -17200 -8924 -17152
rect -8312 -16448 -7512 -16400
rect -8312 -17152 -8264 -16448
rect -7560 -17152 -7512 -16448
rect -8312 -17200 -7512 -17152
rect -6900 -16448 -6100 -16400
rect -6900 -17152 -6852 -16448
rect -6148 -17152 -6100 -16448
rect -6900 -17200 -6100 -17152
rect -5488 -16448 -4688 -16400
rect -5488 -17152 -5440 -16448
rect -4736 -17152 -4688 -16448
rect -5488 -17200 -4688 -17152
rect -4076 -16448 -3276 -16400
rect -4076 -17152 -4028 -16448
rect -3324 -17152 -3276 -16448
rect -4076 -17200 -3276 -17152
rect -2664 -16448 -1864 -16400
rect -2664 -17152 -2616 -16448
rect -1912 -17152 -1864 -16448
rect -2664 -17200 -1864 -17152
rect -1252 -16448 -452 -16400
rect -1252 -17152 -1204 -16448
rect -500 -17152 -452 -16448
rect -1252 -17200 -452 -17152
rect 160 -16448 960 -16400
rect 160 -17152 208 -16448
rect 912 -17152 960 -16448
rect 160 -17200 960 -17152
rect 1572 -16448 2372 -16400
rect 1572 -17152 1620 -16448
rect 2324 -17152 2372 -16448
rect 1572 -17200 2372 -17152
rect 2984 -16448 3784 -16400
rect 2984 -17152 3032 -16448
rect 3736 -17152 3784 -16448
rect 2984 -17200 3784 -17152
rect 4396 -16448 5196 -16400
rect 4396 -17152 4444 -16448
rect 5148 -17152 5196 -16448
rect 4396 -17200 5196 -17152
rect 5808 -16448 6608 -16400
rect 5808 -17152 5856 -16448
rect 6560 -17152 6608 -16448
rect 5808 -17200 6608 -17152
rect 7220 -16448 8020 -16400
rect 7220 -17152 7268 -16448
rect 7972 -17152 8020 -16448
rect 7220 -17200 8020 -17152
rect 8632 -16448 9432 -16400
rect 8632 -17152 8680 -16448
rect 9384 -17152 9432 -16448
rect 8632 -17200 9432 -17152
rect 10044 -16448 10844 -16400
rect 10044 -17152 10092 -16448
rect 10796 -17152 10844 -16448
rect 10044 -17200 10844 -17152
rect 11456 -16448 12256 -16400
rect 11456 -17152 11504 -16448
rect 12208 -17152 12256 -16448
rect 11456 -17200 12256 -17152
rect 12868 -16448 13668 -16400
rect 12868 -17152 12916 -16448
rect 13620 -17152 13668 -16448
rect 12868 -17200 13668 -17152
rect 14280 -16448 15080 -16400
rect 14280 -17152 14328 -16448
rect 15032 -17152 15080 -16448
rect 14280 -17200 15080 -17152
rect 15692 -16448 16492 -16400
rect 15692 -17152 15740 -16448
rect 16444 -17152 16492 -16448
rect 15692 -17200 16492 -17152
rect 17104 -16448 17904 -16400
rect 17104 -17152 17152 -16448
rect 17856 -17152 17904 -16448
rect 17104 -17200 17904 -17152
rect 18516 -16448 19316 -16400
rect 18516 -17152 18564 -16448
rect 19268 -17152 19316 -16448
rect 18516 -17200 19316 -17152
rect 19928 -16448 20728 -16400
rect 19928 -17152 19976 -16448
rect 20680 -17152 20728 -16448
rect 19928 -17200 20728 -17152
rect 21340 -16448 22140 -16400
rect 21340 -17152 21388 -16448
rect 22092 -17152 22140 -16448
rect 21340 -17200 22140 -17152
rect 22752 -16448 23552 -16400
rect 22752 -17152 22800 -16448
rect 23504 -17152 23552 -16448
rect 22752 -17200 23552 -17152
rect -23844 -17568 -23044 -17520
rect -23844 -18272 -23796 -17568
rect -23092 -18272 -23044 -17568
rect -23844 -18320 -23044 -18272
rect -22432 -17568 -21632 -17520
rect -22432 -18272 -22384 -17568
rect -21680 -18272 -21632 -17568
rect -22432 -18320 -21632 -18272
rect -21020 -17568 -20220 -17520
rect -21020 -18272 -20972 -17568
rect -20268 -18272 -20220 -17568
rect -21020 -18320 -20220 -18272
rect -19608 -17568 -18808 -17520
rect -19608 -18272 -19560 -17568
rect -18856 -18272 -18808 -17568
rect -19608 -18320 -18808 -18272
rect -18196 -17568 -17396 -17520
rect -18196 -18272 -18148 -17568
rect -17444 -18272 -17396 -17568
rect -18196 -18320 -17396 -18272
rect -16784 -17568 -15984 -17520
rect -16784 -18272 -16736 -17568
rect -16032 -18272 -15984 -17568
rect -16784 -18320 -15984 -18272
rect -15372 -17568 -14572 -17520
rect -15372 -18272 -15324 -17568
rect -14620 -18272 -14572 -17568
rect -15372 -18320 -14572 -18272
rect -13960 -17568 -13160 -17520
rect -13960 -18272 -13912 -17568
rect -13208 -18272 -13160 -17568
rect -13960 -18320 -13160 -18272
rect -12548 -17568 -11748 -17520
rect -12548 -18272 -12500 -17568
rect -11796 -18272 -11748 -17568
rect -12548 -18320 -11748 -18272
rect -11136 -17568 -10336 -17520
rect -11136 -18272 -11088 -17568
rect -10384 -18272 -10336 -17568
rect -11136 -18320 -10336 -18272
rect -9724 -17568 -8924 -17520
rect -9724 -18272 -9676 -17568
rect -8972 -18272 -8924 -17568
rect -9724 -18320 -8924 -18272
rect -8312 -17568 -7512 -17520
rect -8312 -18272 -8264 -17568
rect -7560 -18272 -7512 -17568
rect -8312 -18320 -7512 -18272
rect -6900 -17568 -6100 -17520
rect -6900 -18272 -6852 -17568
rect -6148 -18272 -6100 -17568
rect -6900 -18320 -6100 -18272
rect -5488 -17568 -4688 -17520
rect -5488 -18272 -5440 -17568
rect -4736 -18272 -4688 -17568
rect -5488 -18320 -4688 -18272
rect -4076 -17568 -3276 -17520
rect -4076 -18272 -4028 -17568
rect -3324 -18272 -3276 -17568
rect -4076 -18320 -3276 -18272
rect -2664 -17568 -1864 -17520
rect -2664 -18272 -2616 -17568
rect -1912 -18272 -1864 -17568
rect -2664 -18320 -1864 -18272
rect -1252 -17568 -452 -17520
rect -1252 -18272 -1204 -17568
rect -500 -18272 -452 -17568
rect -1252 -18320 -452 -18272
rect 160 -17568 960 -17520
rect 160 -18272 208 -17568
rect 912 -18272 960 -17568
rect 160 -18320 960 -18272
rect 1572 -17568 2372 -17520
rect 1572 -18272 1620 -17568
rect 2324 -18272 2372 -17568
rect 1572 -18320 2372 -18272
rect 2984 -17568 3784 -17520
rect 2984 -18272 3032 -17568
rect 3736 -18272 3784 -17568
rect 2984 -18320 3784 -18272
rect 4396 -17568 5196 -17520
rect 4396 -18272 4444 -17568
rect 5148 -18272 5196 -17568
rect 4396 -18320 5196 -18272
rect 5808 -17568 6608 -17520
rect 5808 -18272 5856 -17568
rect 6560 -18272 6608 -17568
rect 5808 -18320 6608 -18272
rect 7220 -17568 8020 -17520
rect 7220 -18272 7268 -17568
rect 7972 -18272 8020 -17568
rect 7220 -18320 8020 -18272
rect 8632 -17568 9432 -17520
rect 8632 -18272 8680 -17568
rect 9384 -18272 9432 -17568
rect 8632 -18320 9432 -18272
rect 10044 -17568 10844 -17520
rect 10044 -18272 10092 -17568
rect 10796 -18272 10844 -17568
rect 10044 -18320 10844 -18272
rect 11456 -17568 12256 -17520
rect 11456 -18272 11504 -17568
rect 12208 -18272 12256 -17568
rect 11456 -18320 12256 -18272
rect 12868 -17568 13668 -17520
rect 12868 -18272 12916 -17568
rect 13620 -18272 13668 -17568
rect 12868 -18320 13668 -18272
rect 14280 -17568 15080 -17520
rect 14280 -18272 14328 -17568
rect 15032 -18272 15080 -17568
rect 14280 -18320 15080 -18272
rect 15692 -17568 16492 -17520
rect 15692 -18272 15740 -17568
rect 16444 -18272 16492 -17568
rect 15692 -18320 16492 -18272
rect 17104 -17568 17904 -17520
rect 17104 -18272 17152 -17568
rect 17856 -18272 17904 -17568
rect 17104 -18320 17904 -18272
rect 18516 -17568 19316 -17520
rect 18516 -18272 18564 -17568
rect 19268 -18272 19316 -17568
rect 18516 -18320 19316 -18272
rect 19928 -17568 20728 -17520
rect 19928 -18272 19976 -17568
rect 20680 -18272 20728 -17568
rect 19928 -18320 20728 -18272
rect 21340 -17568 22140 -17520
rect 21340 -18272 21388 -17568
rect 22092 -18272 22140 -17568
rect 21340 -18320 22140 -18272
rect 22752 -17568 23552 -17520
rect 22752 -18272 22800 -17568
rect 23504 -18272 23552 -17568
rect 22752 -18320 23552 -18272
<< mimcapcontact >>
rect -23796 17568 -23092 18272
rect -22384 17568 -21680 18272
rect -20972 17568 -20268 18272
rect -19560 17568 -18856 18272
rect -18148 17568 -17444 18272
rect -16736 17568 -16032 18272
rect -15324 17568 -14620 18272
rect -13912 17568 -13208 18272
rect -12500 17568 -11796 18272
rect -11088 17568 -10384 18272
rect -9676 17568 -8972 18272
rect -8264 17568 -7560 18272
rect -6852 17568 -6148 18272
rect -5440 17568 -4736 18272
rect -4028 17568 -3324 18272
rect -2616 17568 -1912 18272
rect -1204 17568 -500 18272
rect 208 17568 912 18272
rect 1620 17568 2324 18272
rect 3032 17568 3736 18272
rect 4444 17568 5148 18272
rect 5856 17568 6560 18272
rect 7268 17568 7972 18272
rect 8680 17568 9384 18272
rect 10092 17568 10796 18272
rect 11504 17568 12208 18272
rect 12916 17568 13620 18272
rect 14328 17568 15032 18272
rect 15740 17568 16444 18272
rect 17152 17568 17856 18272
rect 18564 17568 19268 18272
rect 19976 17568 20680 18272
rect 21388 17568 22092 18272
rect 22800 17568 23504 18272
rect -23796 16448 -23092 17152
rect -22384 16448 -21680 17152
rect -20972 16448 -20268 17152
rect -19560 16448 -18856 17152
rect -18148 16448 -17444 17152
rect -16736 16448 -16032 17152
rect -15324 16448 -14620 17152
rect -13912 16448 -13208 17152
rect -12500 16448 -11796 17152
rect -11088 16448 -10384 17152
rect -9676 16448 -8972 17152
rect -8264 16448 -7560 17152
rect -6852 16448 -6148 17152
rect -5440 16448 -4736 17152
rect -4028 16448 -3324 17152
rect -2616 16448 -1912 17152
rect -1204 16448 -500 17152
rect 208 16448 912 17152
rect 1620 16448 2324 17152
rect 3032 16448 3736 17152
rect 4444 16448 5148 17152
rect 5856 16448 6560 17152
rect 7268 16448 7972 17152
rect 8680 16448 9384 17152
rect 10092 16448 10796 17152
rect 11504 16448 12208 17152
rect 12916 16448 13620 17152
rect 14328 16448 15032 17152
rect 15740 16448 16444 17152
rect 17152 16448 17856 17152
rect 18564 16448 19268 17152
rect 19976 16448 20680 17152
rect 21388 16448 22092 17152
rect 22800 16448 23504 17152
rect -23796 15328 -23092 16032
rect -22384 15328 -21680 16032
rect -20972 15328 -20268 16032
rect -19560 15328 -18856 16032
rect -18148 15328 -17444 16032
rect -16736 15328 -16032 16032
rect -15324 15328 -14620 16032
rect -13912 15328 -13208 16032
rect -12500 15328 -11796 16032
rect -11088 15328 -10384 16032
rect -9676 15328 -8972 16032
rect -8264 15328 -7560 16032
rect -6852 15328 -6148 16032
rect -5440 15328 -4736 16032
rect -4028 15328 -3324 16032
rect -2616 15328 -1912 16032
rect -1204 15328 -500 16032
rect 208 15328 912 16032
rect 1620 15328 2324 16032
rect 3032 15328 3736 16032
rect 4444 15328 5148 16032
rect 5856 15328 6560 16032
rect 7268 15328 7972 16032
rect 8680 15328 9384 16032
rect 10092 15328 10796 16032
rect 11504 15328 12208 16032
rect 12916 15328 13620 16032
rect 14328 15328 15032 16032
rect 15740 15328 16444 16032
rect 17152 15328 17856 16032
rect 18564 15328 19268 16032
rect 19976 15328 20680 16032
rect 21388 15328 22092 16032
rect 22800 15328 23504 16032
rect -23796 14208 -23092 14912
rect -22384 14208 -21680 14912
rect -20972 14208 -20268 14912
rect -19560 14208 -18856 14912
rect -18148 14208 -17444 14912
rect -16736 14208 -16032 14912
rect -15324 14208 -14620 14912
rect -13912 14208 -13208 14912
rect -12500 14208 -11796 14912
rect -11088 14208 -10384 14912
rect -9676 14208 -8972 14912
rect -8264 14208 -7560 14912
rect -6852 14208 -6148 14912
rect -5440 14208 -4736 14912
rect -4028 14208 -3324 14912
rect -2616 14208 -1912 14912
rect -1204 14208 -500 14912
rect 208 14208 912 14912
rect 1620 14208 2324 14912
rect 3032 14208 3736 14912
rect 4444 14208 5148 14912
rect 5856 14208 6560 14912
rect 7268 14208 7972 14912
rect 8680 14208 9384 14912
rect 10092 14208 10796 14912
rect 11504 14208 12208 14912
rect 12916 14208 13620 14912
rect 14328 14208 15032 14912
rect 15740 14208 16444 14912
rect 17152 14208 17856 14912
rect 18564 14208 19268 14912
rect 19976 14208 20680 14912
rect 21388 14208 22092 14912
rect 22800 14208 23504 14912
rect -23796 13088 -23092 13792
rect -22384 13088 -21680 13792
rect -20972 13088 -20268 13792
rect -19560 13088 -18856 13792
rect -18148 13088 -17444 13792
rect -16736 13088 -16032 13792
rect -15324 13088 -14620 13792
rect -13912 13088 -13208 13792
rect -12500 13088 -11796 13792
rect -11088 13088 -10384 13792
rect -9676 13088 -8972 13792
rect -8264 13088 -7560 13792
rect -6852 13088 -6148 13792
rect -5440 13088 -4736 13792
rect -4028 13088 -3324 13792
rect -2616 13088 -1912 13792
rect -1204 13088 -500 13792
rect 208 13088 912 13792
rect 1620 13088 2324 13792
rect 3032 13088 3736 13792
rect 4444 13088 5148 13792
rect 5856 13088 6560 13792
rect 7268 13088 7972 13792
rect 8680 13088 9384 13792
rect 10092 13088 10796 13792
rect 11504 13088 12208 13792
rect 12916 13088 13620 13792
rect 14328 13088 15032 13792
rect 15740 13088 16444 13792
rect 17152 13088 17856 13792
rect 18564 13088 19268 13792
rect 19976 13088 20680 13792
rect 21388 13088 22092 13792
rect 22800 13088 23504 13792
rect -23796 11968 -23092 12672
rect -22384 11968 -21680 12672
rect -20972 11968 -20268 12672
rect -19560 11968 -18856 12672
rect -18148 11968 -17444 12672
rect -16736 11968 -16032 12672
rect -15324 11968 -14620 12672
rect -13912 11968 -13208 12672
rect -12500 11968 -11796 12672
rect -11088 11968 -10384 12672
rect -9676 11968 -8972 12672
rect -8264 11968 -7560 12672
rect -6852 11968 -6148 12672
rect -5440 11968 -4736 12672
rect -4028 11968 -3324 12672
rect -2616 11968 -1912 12672
rect -1204 11968 -500 12672
rect 208 11968 912 12672
rect 1620 11968 2324 12672
rect 3032 11968 3736 12672
rect 4444 11968 5148 12672
rect 5856 11968 6560 12672
rect 7268 11968 7972 12672
rect 8680 11968 9384 12672
rect 10092 11968 10796 12672
rect 11504 11968 12208 12672
rect 12916 11968 13620 12672
rect 14328 11968 15032 12672
rect 15740 11968 16444 12672
rect 17152 11968 17856 12672
rect 18564 11968 19268 12672
rect 19976 11968 20680 12672
rect 21388 11968 22092 12672
rect 22800 11968 23504 12672
rect -23796 10848 -23092 11552
rect -22384 10848 -21680 11552
rect -20972 10848 -20268 11552
rect -19560 10848 -18856 11552
rect -18148 10848 -17444 11552
rect -16736 10848 -16032 11552
rect -15324 10848 -14620 11552
rect -13912 10848 -13208 11552
rect -12500 10848 -11796 11552
rect -11088 10848 -10384 11552
rect -9676 10848 -8972 11552
rect -8264 10848 -7560 11552
rect -6852 10848 -6148 11552
rect -5440 10848 -4736 11552
rect -4028 10848 -3324 11552
rect -2616 10848 -1912 11552
rect -1204 10848 -500 11552
rect 208 10848 912 11552
rect 1620 10848 2324 11552
rect 3032 10848 3736 11552
rect 4444 10848 5148 11552
rect 5856 10848 6560 11552
rect 7268 10848 7972 11552
rect 8680 10848 9384 11552
rect 10092 10848 10796 11552
rect 11504 10848 12208 11552
rect 12916 10848 13620 11552
rect 14328 10848 15032 11552
rect 15740 10848 16444 11552
rect 17152 10848 17856 11552
rect 18564 10848 19268 11552
rect 19976 10848 20680 11552
rect 21388 10848 22092 11552
rect 22800 10848 23504 11552
rect -23796 9728 -23092 10432
rect -22384 9728 -21680 10432
rect -20972 9728 -20268 10432
rect -19560 9728 -18856 10432
rect -18148 9728 -17444 10432
rect -16736 9728 -16032 10432
rect -15324 9728 -14620 10432
rect -13912 9728 -13208 10432
rect -12500 9728 -11796 10432
rect -11088 9728 -10384 10432
rect -9676 9728 -8972 10432
rect -8264 9728 -7560 10432
rect -6852 9728 -6148 10432
rect -5440 9728 -4736 10432
rect -4028 9728 -3324 10432
rect -2616 9728 -1912 10432
rect -1204 9728 -500 10432
rect 208 9728 912 10432
rect 1620 9728 2324 10432
rect 3032 9728 3736 10432
rect 4444 9728 5148 10432
rect 5856 9728 6560 10432
rect 7268 9728 7972 10432
rect 8680 9728 9384 10432
rect 10092 9728 10796 10432
rect 11504 9728 12208 10432
rect 12916 9728 13620 10432
rect 14328 9728 15032 10432
rect 15740 9728 16444 10432
rect 17152 9728 17856 10432
rect 18564 9728 19268 10432
rect 19976 9728 20680 10432
rect 21388 9728 22092 10432
rect 22800 9728 23504 10432
rect -23796 8608 -23092 9312
rect -22384 8608 -21680 9312
rect -20972 8608 -20268 9312
rect -19560 8608 -18856 9312
rect -18148 8608 -17444 9312
rect -16736 8608 -16032 9312
rect -15324 8608 -14620 9312
rect -13912 8608 -13208 9312
rect -12500 8608 -11796 9312
rect -11088 8608 -10384 9312
rect -9676 8608 -8972 9312
rect -8264 8608 -7560 9312
rect -6852 8608 -6148 9312
rect -5440 8608 -4736 9312
rect -4028 8608 -3324 9312
rect -2616 8608 -1912 9312
rect -1204 8608 -500 9312
rect 208 8608 912 9312
rect 1620 8608 2324 9312
rect 3032 8608 3736 9312
rect 4444 8608 5148 9312
rect 5856 8608 6560 9312
rect 7268 8608 7972 9312
rect 8680 8608 9384 9312
rect 10092 8608 10796 9312
rect 11504 8608 12208 9312
rect 12916 8608 13620 9312
rect 14328 8608 15032 9312
rect 15740 8608 16444 9312
rect 17152 8608 17856 9312
rect 18564 8608 19268 9312
rect 19976 8608 20680 9312
rect 21388 8608 22092 9312
rect 22800 8608 23504 9312
rect -23796 7488 -23092 8192
rect -22384 7488 -21680 8192
rect -20972 7488 -20268 8192
rect -19560 7488 -18856 8192
rect -18148 7488 -17444 8192
rect -16736 7488 -16032 8192
rect -15324 7488 -14620 8192
rect -13912 7488 -13208 8192
rect -12500 7488 -11796 8192
rect -11088 7488 -10384 8192
rect -9676 7488 -8972 8192
rect -8264 7488 -7560 8192
rect -6852 7488 -6148 8192
rect -5440 7488 -4736 8192
rect -4028 7488 -3324 8192
rect -2616 7488 -1912 8192
rect -1204 7488 -500 8192
rect 208 7488 912 8192
rect 1620 7488 2324 8192
rect 3032 7488 3736 8192
rect 4444 7488 5148 8192
rect 5856 7488 6560 8192
rect 7268 7488 7972 8192
rect 8680 7488 9384 8192
rect 10092 7488 10796 8192
rect 11504 7488 12208 8192
rect 12916 7488 13620 8192
rect 14328 7488 15032 8192
rect 15740 7488 16444 8192
rect 17152 7488 17856 8192
rect 18564 7488 19268 8192
rect 19976 7488 20680 8192
rect 21388 7488 22092 8192
rect 22800 7488 23504 8192
rect -23796 6368 -23092 7072
rect -22384 6368 -21680 7072
rect -20972 6368 -20268 7072
rect -19560 6368 -18856 7072
rect -18148 6368 -17444 7072
rect -16736 6368 -16032 7072
rect -15324 6368 -14620 7072
rect -13912 6368 -13208 7072
rect -12500 6368 -11796 7072
rect -11088 6368 -10384 7072
rect -9676 6368 -8972 7072
rect -8264 6368 -7560 7072
rect -6852 6368 -6148 7072
rect -5440 6368 -4736 7072
rect -4028 6368 -3324 7072
rect -2616 6368 -1912 7072
rect -1204 6368 -500 7072
rect 208 6368 912 7072
rect 1620 6368 2324 7072
rect 3032 6368 3736 7072
rect 4444 6368 5148 7072
rect 5856 6368 6560 7072
rect 7268 6368 7972 7072
rect 8680 6368 9384 7072
rect 10092 6368 10796 7072
rect 11504 6368 12208 7072
rect 12916 6368 13620 7072
rect 14328 6368 15032 7072
rect 15740 6368 16444 7072
rect 17152 6368 17856 7072
rect 18564 6368 19268 7072
rect 19976 6368 20680 7072
rect 21388 6368 22092 7072
rect 22800 6368 23504 7072
rect -23796 5248 -23092 5952
rect -22384 5248 -21680 5952
rect -20972 5248 -20268 5952
rect -19560 5248 -18856 5952
rect -18148 5248 -17444 5952
rect -16736 5248 -16032 5952
rect -15324 5248 -14620 5952
rect -13912 5248 -13208 5952
rect -12500 5248 -11796 5952
rect -11088 5248 -10384 5952
rect -9676 5248 -8972 5952
rect -8264 5248 -7560 5952
rect -6852 5248 -6148 5952
rect -5440 5248 -4736 5952
rect -4028 5248 -3324 5952
rect -2616 5248 -1912 5952
rect -1204 5248 -500 5952
rect 208 5248 912 5952
rect 1620 5248 2324 5952
rect 3032 5248 3736 5952
rect 4444 5248 5148 5952
rect 5856 5248 6560 5952
rect 7268 5248 7972 5952
rect 8680 5248 9384 5952
rect 10092 5248 10796 5952
rect 11504 5248 12208 5952
rect 12916 5248 13620 5952
rect 14328 5248 15032 5952
rect 15740 5248 16444 5952
rect 17152 5248 17856 5952
rect 18564 5248 19268 5952
rect 19976 5248 20680 5952
rect 21388 5248 22092 5952
rect 22800 5248 23504 5952
rect -23796 4128 -23092 4832
rect -22384 4128 -21680 4832
rect -20972 4128 -20268 4832
rect -19560 4128 -18856 4832
rect -18148 4128 -17444 4832
rect -16736 4128 -16032 4832
rect -15324 4128 -14620 4832
rect -13912 4128 -13208 4832
rect -12500 4128 -11796 4832
rect -11088 4128 -10384 4832
rect -9676 4128 -8972 4832
rect -8264 4128 -7560 4832
rect -6852 4128 -6148 4832
rect -5440 4128 -4736 4832
rect -4028 4128 -3324 4832
rect -2616 4128 -1912 4832
rect -1204 4128 -500 4832
rect 208 4128 912 4832
rect 1620 4128 2324 4832
rect 3032 4128 3736 4832
rect 4444 4128 5148 4832
rect 5856 4128 6560 4832
rect 7268 4128 7972 4832
rect 8680 4128 9384 4832
rect 10092 4128 10796 4832
rect 11504 4128 12208 4832
rect 12916 4128 13620 4832
rect 14328 4128 15032 4832
rect 15740 4128 16444 4832
rect 17152 4128 17856 4832
rect 18564 4128 19268 4832
rect 19976 4128 20680 4832
rect 21388 4128 22092 4832
rect 22800 4128 23504 4832
rect -23796 3008 -23092 3712
rect -22384 3008 -21680 3712
rect -20972 3008 -20268 3712
rect -19560 3008 -18856 3712
rect -18148 3008 -17444 3712
rect -16736 3008 -16032 3712
rect -15324 3008 -14620 3712
rect -13912 3008 -13208 3712
rect -12500 3008 -11796 3712
rect -11088 3008 -10384 3712
rect -9676 3008 -8972 3712
rect -8264 3008 -7560 3712
rect -6852 3008 -6148 3712
rect -5440 3008 -4736 3712
rect -4028 3008 -3324 3712
rect -2616 3008 -1912 3712
rect -1204 3008 -500 3712
rect 208 3008 912 3712
rect 1620 3008 2324 3712
rect 3032 3008 3736 3712
rect 4444 3008 5148 3712
rect 5856 3008 6560 3712
rect 7268 3008 7972 3712
rect 8680 3008 9384 3712
rect 10092 3008 10796 3712
rect 11504 3008 12208 3712
rect 12916 3008 13620 3712
rect 14328 3008 15032 3712
rect 15740 3008 16444 3712
rect 17152 3008 17856 3712
rect 18564 3008 19268 3712
rect 19976 3008 20680 3712
rect 21388 3008 22092 3712
rect 22800 3008 23504 3712
rect -23796 1888 -23092 2592
rect -22384 1888 -21680 2592
rect -20972 1888 -20268 2592
rect -19560 1888 -18856 2592
rect -18148 1888 -17444 2592
rect -16736 1888 -16032 2592
rect -15324 1888 -14620 2592
rect -13912 1888 -13208 2592
rect -12500 1888 -11796 2592
rect -11088 1888 -10384 2592
rect -9676 1888 -8972 2592
rect -8264 1888 -7560 2592
rect -6852 1888 -6148 2592
rect -5440 1888 -4736 2592
rect -4028 1888 -3324 2592
rect -2616 1888 -1912 2592
rect -1204 1888 -500 2592
rect 208 1888 912 2592
rect 1620 1888 2324 2592
rect 3032 1888 3736 2592
rect 4444 1888 5148 2592
rect 5856 1888 6560 2592
rect 7268 1888 7972 2592
rect 8680 1888 9384 2592
rect 10092 1888 10796 2592
rect 11504 1888 12208 2592
rect 12916 1888 13620 2592
rect 14328 1888 15032 2592
rect 15740 1888 16444 2592
rect 17152 1888 17856 2592
rect 18564 1888 19268 2592
rect 19976 1888 20680 2592
rect 21388 1888 22092 2592
rect 22800 1888 23504 2592
rect -23796 768 -23092 1472
rect -22384 768 -21680 1472
rect -20972 768 -20268 1472
rect -19560 768 -18856 1472
rect -18148 768 -17444 1472
rect -16736 768 -16032 1472
rect -15324 768 -14620 1472
rect -13912 768 -13208 1472
rect -12500 768 -11796 1472
rect -11088 768 -10384 1472
rect -9676 768 -8972 1472
rect -8264 768 -7560 1472
rect -6852 768 -6148 1472
rect -5440 768 -4736 1472
rect -4028 768 -3324 1472
rect -2616 768 -1912 1472
rect -1204 768 -500 1472
rect 208 768 912 1472
rect 1620 768 2324 1472
rect 3032 768 3736 1472
rect 4444 768 5148 1472
rect 5856 768 6560 1472
rect 7268 768 7972 1472
rect 8680 768 9384 1472
rect 10092 768 10796 1472
rect 11504 768 12208 1472
rect 12916 768 13620 1472
rect 14328 768 15032 1472
rect 15740 768 16444 1472
rect 17152 768 17856 1472
rect 18564 768 19268 1472
rect 19976 768 20680 1472
rect 21388 768 22092 1472
rect 22800 768 23504 1472
rect -23796 -352 -23092 352
rect -22384 -352 -21680 352
rect -20972 -352 -20268 352
rect -19560 -352 -18856 352
rect -18148 -352 -17444 352
rect -16736 -352 -16032 352
rect -15324 -352 -14620 352
rect -13912 -352 -13208 352
rect -12500 -352 -11796 352
rect -11088 -352 -10384 352
rect -9676 -352 -8972 352
rect -8264 -352 -7560 352
rect -6852 -352 -6148 352
rect -5440 -352 -4736 352
rect -4028 -352 -3324 352
rect -2616 -352 -1912 352
rect -1204 -352 -500 352
rect 208 -352 912 352
rect 1620 -352 2324 352
rect 3032 -352 3736 352
rect 4444 -352 5148 352
rect 5856 -352 6560 352
rect 7268 -352 7972 352
rect 8680 -352 9384 352
rect 10092 -352 10796 352
rect 11504 -352 12208 352
rect 12916 -352 13620 352
rect 14328 -352 15032 352
rect 15740 -352 16444 352
rect 17152 -352 17856 352
rect 18564 -352 19268 352
rect 19976 -352 20680 352
rect 21388 -352 22092 352
rect 22800 -352 23504 352
rect -23796 -1472 -23092 -768
rect -22384 -1472 -21680 -768
rect -20972 -1472 -20268 -768
rect -19560 -1472 -18856 -768
rect -18148 -1472 -17444 -768
rect -16736 -1472 -16032 -768
rect -15324 -1472 -14620 -768
rect -13912 -1472 -13208 -768
rect -12500 -1472 -11796 -768
rect -11088 -1472 -10384 -768
rect -9676 -1472 -8972 -768
rect -8264 -1472 -7560 -768
rect -6852 -1472 -6148 -768
rect -5440 -1472 -4736 -768
rect -4028 -1472 -3324 -768
rect -2616 -1472 -1912 -768
rect -1204 -1472 -500 -768
rect 208 -1472 912 -768
rect 1620 -1472 2324 -768
rect 3032 -1472 3736 -768
rect 4444 -1472 5148 -768
rect 5856 -1472 6560 -768
rect 7268 -1472 7972 -768
rect 8680 -1472 9384 -768
rect 10092 -1472 10796 -768
rect 11504 -1472 12208 -768
rect 12916 -1472 13620 -768
rect 14328 -1472 15032 -768
rect 15740 -1472 16444 -768
rect 17152 -1472 17856 -768
rect 18564 -1472 19268 -768
rect 19976 -1472 20680 -768
rect 21388 -1472 22092 -768
rect 22800 -1472 23504 -768
rect -23796 -2592 -23092 -1888
rect -22384 -2592 -21680 -1888
rect -20972 -2592 -20268 -1888
rect -19560 -2592 -18856 -1888
rect -18148 -2592 -17444 -1888
rect -16736 -2592 -16032 -1888
rect -15324 -2592 -14620 -1888
rect -13912 -2592 -13208 -1888
rect -12500 -2592 -11796 -1888
rect -11088 -2592 -10384 -1888
rect -9676 -2592 -8972 -1888
rect -8264 -2592 -7560 -1888
rect -6852 -2592 -6148 -1888
rect -5440 -2592 -4736 -1888
rect -4028 -2592 -3324 -1888
rect -2616 -2592 -1912 -1888
rect -1204 -2592 -500 -1888
rect 208 -2592 912 -1888
rect 1620 -2592 2324 -1888
rect 3032 -2592 3736 -1888
rect 4444 -2592 5148 -1888
rect 5856 -2592 6560 -1888
rect 7268 -2592 7972 -1888
rect 8680 -2592 9384 -1888
rect 10092 -2592 10796 -1888
rect 11504 -2592 12208 -1888
rect 12916 -2592 13620 -1888
rect 14328 -2592 15032 -1888
rect 15740 -2592 16444 -1888
rect 17152 -2592 17856 -1888
rect 18564 -2592 19268 -1888
rect 19976 -2592 20680 -1888
rect 21388 -2592 22092 -1888
rect 22800 -2592 23504 -1888
rect -23796 -3712 -23092 -3008
rect -22384 -3712 -21680 -3008
rect -20972 -3712 -20268 -3008
rect -19560 -3712 -18856 -3008
rect -18148 -3712 -17444 -3008
rect -16736 -3712 -16032 -3008
rect -15324 -3712 -14620 -3008
rect -13912 -3712 -13208 -3008
rect -12500 -3712 -11796 -3008
rect -11088 -3712 -10384 -3008
rect -9676 -3712 -8972 -3008
rect -8264 -3712 -7560 -3008
rect -6852 -3712 -6148 -3008
rect -5440 -3712 -4736 -3008
rect -4028 -3712 -3324 -3008
rect -2616 -3712 -1912 -3008
rect -1204 -3712 -500 -3008
rect 208 -3712 912 -3008
rect 1620 -3712 2324 -3008
rect 3032 -3712 3736 -3008
rect 4444 -3712 5148 -3008
rect 5856 -3712 6560 -3008
rect 7268 -3712 7972 -3008
rect 8680 -3712 9384 -3008
rect 10092 -3712 10796 -3008
rect 11504 -3712 12208 -3008
rect 12916 -3712 13620 -3008
rect 14328 -3712 15032 -3008
rect 15740 -3712 16444 -3008
rect 17152 -3712 17856 -3008
rect 18564 -3712 19268 -3008
rect 19976 -3712 20680 -3008
rect 21388 -3712 22092 -3008
rect 22800 -3712 23504 -3008
rect -23796 -4832 -23092 -4128
rect -22384 -4832 -21680 -4128
rect -20972 -4832 -20268 -4128
rect -19560 -4832 -18856 -4128
rect -18148 -4832 -17444 -4128
rect -16736 -4832 -16032 -4128
rect -15324 -4832 -14620 -4128
rect -13912 -4832 -13208 -4128
rect -12500 -4832 -11796 -4128
rect -11088 -4832 -10384 -4128
rect -9676 -4832 -8972 -4128
rect -8264 -4832 -7560 -4128
rect -6852 -4832 -6148 -4128
rect -5440 -4832 -4736 -4128
rect -4028 -4832 -3324 -4128
rect -2616 -4832 -1912 -4128
rect -1204 -4832 -500 -4128
rect 208 -4832 912 -4128
rect 1620 -4832 2324 -4128
rect 3032 -4832 3736 -4128
rect 4444 -4832 5148 -4128
rect 5856 -4832 6560 -4128
rect 7268 -4832 7972 -4128
rect 8680 -4832 9384 -4128
rect 10092 -4832 10796 -4128
rect 11504 -4832 12208 -4128
rect 12916 -4832 13620 -4128
rect 14328 -4832 15032 -4128
rect 15740 -4832 16444 -4128
rect 17152 -4832 17856 -4128
rect 18564 -4832 19268 -4128
rect 19976 -4832 20680 -4128
rect 21388 -4832 22092 -4128
rect 22800 -4832 23504 -4128
rect -23796 -5952 -23092 -5248
rect -22384 -5952 -21680 -5248
rect -20972 -5952 -20268 -5248
rect -19560 -5952 -18856 -5248
rect -18148 -5952 -17444 -5248
rect -16736 -5952 -16032 -5248
rect -15324 -5952 -14620 -5248
rect -13912 -5952 -13208 -5248
rect -12500 -5952 -11796 -5248
rect -11088 -5952 -10384 -5248
rect -9676 -5952 -8972 -5248
rect -8264 -5952 -7560 -5248
rect -6852 -5952 -6148 -5248
rect -5440 -5952 -4736 -5248
rect -4028 -5952 -3324 -5248
rect -2616 -5952 -1912 -5248
rect -1204 -5952 -500 -5248
rect 208 -5952 912 -5248
rect 1620 -5952 2324 -5248
rect 3032 -5952 3736 -5248
rect 4444 -5952 5148 -5248
rect 5856 -5952 6560 -5248
rect 7268 -5952 7972 -5248
rect 8680 -5952 9384 -5248
rect 10092 -5952 10796 -5248
rect 11504 -5952 12208 -5248
rect 12916 -5952 13620 -5248
rect 14328 -5952 15032 -5248
rect 15740 -5952 16444 -5248
rect 17152 -5952 17856 -5248
rect 18564 -5952 19268 -5248
rect 19976 -5952 20680 -5248
rect 21388 -5952 22092 -5248
rect 22800 -5952 23504 -5248
rect -23796 -7072 -23092 -6368
rect -22384 -7072 -21680 -6368
rect -20972 -7072 -20268 -6368
rect -19560 -7072 -18856 -6368
rect -18148 -7072 -17444 -6368
rect -16736 -7072 -16032 -6368
rect -15324 -7072 -14620 -6368
rect -13912 -7072 -13208 -6368
rect -12500 -7072 -11796 -6368
rect -11088 -7072 -10384 -6368
rect -9676 -7072 -8972 -6368
rect -8264 -7072 -7560 -6368
rect -6852 -7072 -6148 -6368
rect -5440 -7072 -4736 -6368
rect -4028 -7072 -3324 -6368
rect -2616 -7072 -1912 -6368
rect -1204 -7072 -500 -6368
rect 208 -7072 912 -6368
rect 1620 -7072 2324 -6368
rect 3032 -7072 3736 -6368
rect 4444 -7072 5148 -6368
rect 5856 -7072 6560 -6368
rect 7268 -7072 7972 -6368
rect 8680 -7072 9384 -6368
rect 10092 -7072 10796 -6368
rect 11504 -7072 12208 -6368
rect 12916 -7072 13620 -6368
rect 14328 -7072 15032 -6368
rect 15740 -7072 16444 -6368
rect 17152 -7072 17856 -6368
rect 18564 -7072 19268 -6368
rect 19976 -7072 20680 -6368
rect 21388 -7072 22092 -6368
rect 22800 -7072 23504 -6368
rect -23796 -8192 -23092 -7488
rect -22384 -8192 -21680 -7488
rect -20972 -8192 -20268 -7488
rect -19560 -8192 -18856 -7488
rect -18148 -8192 -17444 -7488
rect -16736 -8192 -16032 -7488
rect -15324 -8192 -14620 -7488
rect -13912 -8192 -13208 -7488
rect -12500 -8192 -11796 -7488
rect -11088 -8192 -10384 -7488
rect -9676 -8192 -8972 -7488
rect -8264 -8192 -7560 -7488
rect -6852 -8192 -6148 -7488
rect -5440 -8192 -4736 -7488
rect -4028 -8192 -3324 -7488
rect -2616 -8192 -1912 -7488
rect -1204 -8192 -500 -7488
rect 208 -8192 912 -7488
rect 1620 -8192 2324 -7488
rect 3032 -8192 3736 -7488
rect 4444 -8192 5148 -7488
rect 5856 -8192 6560 -7488
rect 7268 -8192 7972 -7488
rect 8680 -8192 9384 -7488
rect 10092 -8192 10796 -7488
rect 11504 -8192 12208 -7488
rect 12916 -8192 13620 -7488
rect 14328 -8192 15032 -7488
rect 15740 -8192 16444 -7488
rect 17152 -8192 17856 -7488
rect 18564 -8192 19268 -7488
rect 19976 -8192 20680 -7488
rect 21388 -8192 22092 -7488
rect 22800 -8192 23504 -7488
rect -23796 -9312 -23092 -8608
rect -22384 -9312 -21680 -8608
rect -20972 -9312 -20268 -8608
rect -19560 -9312 -18856 -8608
rect -18148 -9312 -17444 -8608
rect -16736 -9312 -16032 -8608
rect -15324 -9312 -14620 -8608
rect -13912 -9312 -13208 -8608
rect -12500 -9312 -11796 -8608
rect -11088 -9312 -10384 -8608
rect -9676 -9312 -8972 -8608
rect -8264 -9312 -7560 -8608
rect -6852 -9312 -6148 -8608
rect -5440 -9312 -4736 -8608
rect -4028 -9312 -3324 -8608
rect -2616 -9312 -1912 -8608
rect -1204 -9312 -500 -8608
rect 208 -9312 912 -8608
rect 1620 -9312 2324 -8608
rect 3032 -9312 3736 -8608
rect 4444 -9312 5148 -8608
rect 5856 -9312 6560 -8608
rect 7268 -9312 7972 -8608
rect 8680 -9312 9384 -8608
rect 10092 -9312 10796 -8608
rect 11504 -9312 12208 -8608
rect 12916 -9312 13620 -8608
rect 14328 -9312 15032 -8608
rect 15740 -9312 16444 -8608
rect 17152 -9312 17856 -8608
rect 18564 -9312 19268 -8608
rect 19976 -9312 20680 -8608
rect 21388 -9312 22092 -8608
rect 22800 -9312 23504 -8608
rect -23796 -10432 -23092 -9728
rect -22384 -10432 -21680 -9728
rect -20972 -10432 -20268 -9728
rect -19560 -10432 -18856 -9728
rect -18148 -10432 -17444 -9728
rect -16736 -10432 -16032 -9728
rect -15324 -10432 -14620 -9728
rect -13912 -10432 -13208 -9728
rect -12500 -10432 -11796 -9728
rect -11088 -10432 -10384 -9728
rect -9676 -10432 -8972 -9728
rect -8264 -10432 -7560 -9728
rect -6852 -10432 -6148 -9728
rect -5440 -10432 -4736 -9728
rect -4028 -10432 -3324 -9728
rect -2616 -10432 -1912 -9728
rect -1204 -10432 -500 -9728
rect 208 -10432 912 -9728
rect 1620 -10432 2324 -9728
rect 3032 -10432 3736 -9728
rect 4444 -10432 5148 -9728
rect 5856 -10432 6560 -9728
rect 7268 -10432 7972 -9728
rect 8680 -10432 9384 -9728
rect 10092 -10432 10796 -9728
rect 11504 -10432 12208 -9728
rect 12916 -10432 13620 -9728
rect 14328 -10432 15032 -9728
rect 15740 -10432 16444 -9728
rect 17152 -10432 17856 -9728
rect 18564 -10432 19268 -9728
rect 19976 -10432 20680 -9728
rect 21388 -10432 22092 -9728
rect 22800 -10432 23504 -9728
rect -23796 -11552 -23092 -10848
rect -22384 -11552 -21680 -10848
rect -20972 -11552 -20268 -10848
rect -19560 -11552 -18856 -10848
rect -18148 -11552 -17444 -10848
rect -16736 -11552 -16032 -10848
rect -15324 -11552 -14620 -10848
rect -13912 -11552 -13208 -10848
rect -12500 -11552 -11796 -10848
rect -11088 -11552 -10384 -10848
rect -9676 -11552 -8972 -10848
rect -8264 -11552 -7560 -10848
rect -6852 -11552 -6148 -10848
rect -5440 -11552 -4736 -10848
rect -4028 -11552 -3324 -10848
rect -2616 -11552 -1912 -10848
rect -1204 -11552 -500 -10848
rect 208 -11552 912 -10848
rect 1620 -11552 2324 -10848
rect 3032 -11552 3736 -10848
rect 4444 -11552 5148 -10848
rect 5856 -11552 6560 -10848
rect 7268 -11552 7972 -10848
rect 8680 -11552 9384 -10848
rect 10092 -11552 10796 -10848
rect 11504 -11552 12208 -10848
rect 12916 -11552 13620 -10848
rect 14328 -11552 15032 -10848
rect 15740 -11552 16444 -10848
rect 17152 -11552 17856 -10848
rect 18564 -11552 19268 -10848
rect 19976 -11552 20680 -10848
rect 21388 -11552 22092 -10848
rect 22800 -11552 23504 -10848
rect -23796 -12672 -23092 -11968
rect -22384 -12672 -21680 -11968
rect -20972 -12672 -20268 -11968
rect -19560 -12672 -18856 -11968
rect -18148 -12672 -17444 -11968
rect -16736 -12672 -16032 -11968
rect -15324 -12672 -14620 -11968
rect -13912 -12672 -13208 -11968
rect -12500 -12672 -11796 -11968
rect -11088 -12672 -10384 -11968
rect -9676 -12672 -8972 -11968
rect -8264 -12672 -7560 -11968
rect -6852 -12672 -6148 -11968
rect -5440 -12672 -4736 -11968
rect -4028 -12672 -3324 -11968
rect -2616 -12672 -1912 -11968
rect -1204 -12672 -500 -11968
rect 208 -12672 912 -11968
rect 1620 -12672 2324 -11968
rect 3032 -12672 3736 -11968
rect 4444 -12672 5148 -11968
rect 5856 -12672 6560 -11968
rect 7268 -12672 7972 -11968
rect 8680 -12672 9384 -11968
rect 10092 -12672 10796 -11968
rect 11504 -12672 12208 -11968
rect 12916 -12672 13620 -11968
rect 14328 -12672 15032 -11968
rect 15740 -12672 16444 -11968
rect 17152 -12672 17856 -11968
rect 18564 -12672 19268 -11968
rect 19976 -12672 20680 -11968
rect 21388 -12672 22092 -11968
rect 22800 -12672 23504 -11968
rect -23796 -13792 -23092 -13088
rect -22384 -13792 -21680 -13088
rect -20972 -13792 -20268 -13088
rect -19560 -13792 -18856 -13088
rect -18148 -13792 -17444 -13088
rect -16736 -13792 -16032 -13088
rect -15324 -13792 -14620 -13088
rect -13912 -13792 -13208 -13088
rect -12500 -13792 -11796 -13088
rect -11088 -13792 -10384 -13088
rect -9676 -13792 -8972 -13088
rect -8264 -13792 -7560 -13088
rect -6852 -13792 -6148 -13088
rect -5440 -13792 -4736 -13088
rect -4028 -13792 -3324 -13088
rect -2616 -13792 -1912 -13088
rect -1204 -13792 -500 -13088
rect 208 -13792 912 -13088
rect 1620 -13792 2324 -13088
rect 3032 -13792 3736 -13088
rect 4444 -13792 5148 -13088
rect 5856 -13792 6560 -13088
rect 7268 -13792 7972 -13088
rect 8680 -13792 9384 -13088
rect 10092 -13792 10796 -13088
rect 11504 -13792 12208 -13088
rect 12916 -13792 13620 -13088
rect 14328 -13792 15032 -13088
rect 15740 -13792 16444 -13088
rect 17152 -13792 17856 -13088
rect 18564 -13792 19268 -13088
rect 19976 -13792 20680 -13088
rect 21388 -13792 22092 -13088
rect 22800 -13792 23504 -13088
rect -23796 -14912 -23092 -14208
rect -22384 -14912 -21680 -14208
rect -20972 -14912 -20268 -14208
rect -19560 -14912 -18856 -14208
rect -18148 -14912 -17444 -14208
rect -16736 -14912 -16032 -14208
rect -15324 -14912 -14620 -14208
rect -13912 -14912 -13208 -14208
rect -12500 -14912 -11796 -14208
rect -11088 -14912 -10384 -14208
rect -9676 -14912 -8972 -14208
rect -8264 -14912 -7560 -14208
rect -6852 -14912 -6148 -14208
rect -5440 -14912 -4736 -14208
rect -4028 -14912 -3324 -14208
rect -2616 -14912 -1912 -14208
rect -1204 -14912 -500 -14208
rect 208 -14912 912 -14208
rect 1620 -14912 2324 -14208
rect 3032 -14912 3736 -14208
rect 4444 -14912 5148 -14208
rect 5856 -14912 6560 -14208
rect 7268 -14912 7972 -14208
rect 8680 -14912 9384 -14208
rect 10092 -14912 10796 -14208
rect 11504 -14912 12208 -14208
rect 12916 -14912 13620 -14208
rect 14328 -14912 15032 -14208
rect 15740 -14912 16444 -14208
rect 17152 -14912 17856 -14208
rect 18564 -14912 19268 -14208
rect 19976 -14912 20680 -14208
rect 21388 -14912 22092 -14208
rect 22800 -14912 23504 -14208
rect -23796 -16032 -23092 -15328
rect -22384 -16032 -21680 -15328
rect -20972 -16032 -20268 -15328
rect -19560 -16032 -18856 -15328
rect -18148 -16032 -17444 -15328
rect -16736 -16032 -16032 -15328
rect -15324 -16032 -14620 -15328
rect -13912 -16032 -13208 -15328
rect -12500 -16032 -11796 -15328
rect -11088 -16032 -10384 -15328
rect -9676 -16032 -8972 -15328
rect -8264 -16032 -7560 -15328
rect -6852 -16032 -6148 -15328
rect -5440 -16032 -4736 -15328
rect -4028 -16032 -3324 -15328
rect -2616 -16032 -1912 -15328
rect -1204 -16032 -500 -15328
rect 208 -16032 912 -15328
rect 1620 -16032 2324 -15328
rect 3032 -16032 3736 -15328
rect 4444 -16032 5148 -15328
rect 5856 -16032 6560 -15328
rect 7268 -16032 7972 -15328
rect 8680 -16032 9384 -15328
rect 10092 -16032 10796 -15328
rect 11504 -16032 12208 -15328
rect 12916 -16032 13620 -15328
rect 14328 -16032 15032 -15328
rect 15740 -16032 16444 -15328
rect 17152 -16032 17856 -15328
rect 18564 -16032 19268 -15328
rect 19976 -16032 20680 -15328
rect 21388 -16032 22092 -15328
rect 22800 -16032 23504 -15328
rect -23796 -17152 -23092 -16448
rect -22384 -17152 -21680 -16448
rect -20972 -17152 -20268 -16448
rect -19560 -17152 -18856 -16448
rect -18148 -17152 -17444 -16448
rect -16736 -17152 -16032 -16448
rect -15324 -17152 -14620 -16448
rect -13912 -17152 -13208 -16448
rect -12500 -17152 -11796 -16448
rect -11088 -17152 -10384 -16448
rect -9676 -17152 -8972 -16448
rect -8264 -17152 -7560 -16448
rect -6852 -17152 -6148 -16448
rect -5440 -17152 -4736 -16448
rect -4028 -17152 -3324 -16448
rect -2616 -17152 -1912 -16448
rect -1204 -17152 -500 -16448
rect 208 -17152 912 -16448
rect 1620 -17152 2324 -16448
rect 3032 -17152 3736 -16448
rect 4444 -17152 5148 -16448
rect 5856 -17152 6560 -16448
rect 7268 -17152 7972 -16448
rect 8680 -17152 9384 -16448
rect 10092 -17152 10796 -16448
rect 11504 -17152 12208 -16448
rect 12916 -17152 13620 -16448
rect 14328 -17152 15032 -16448
rect 15740 -17152 16444 -16448
rect 17152 -17152 17856 -16448
rect 18564 -17152 19268 -16448
rect 19976 -17152 20680 -16448
rect 21388 -17152 22092 -16448
rect 22800 -17152 23504 -16448
rect -23796 -18272 -23092 -17568
rect -22384 -18272 -21680 -17568
rect -20972 -18272 -20268 -17568
rect -19560 -18272 -18856 -17568
rect -18148 -18272 -17444 -17568
rect -16736 -18272 -16032 -17568
rect -15324 -18272 -14620 -17568
rect -13912 -18272 -13208 -17568
rect -12500 -18272 -11796 -17568
rect -11088 -18272 -10384 -17568
rect -9676 -18272 -8972 -17568
rect -8264 -18272 -7560 -17568
rect -6852 -18272 -6148 -17568
rect -5440 -18272 -4736 -17568
rect -4028 -18272 -3324 -17568
rect -2616 -18272 -1912 -17568
rect -1204 -18272 -500 -17568
rect 208 -18272 912 -17568
rect 1620 -18272 2324 -17568
rect 3032 -18272 3736 -17568
rect 4444 -18272 5148 -17568
rect 5856 -18272 6560 -17568
rect 7268 -18272 7972 -17568
rect 8680 -18272 9384 -17568
rect 10092 -18272 10796 -17568
rect 11504 -18272 12208 -17568
rect 12916 -18272 13620 -17568
rect 14328 -18272 15032 -17568
rect 15740 -18272 16444 -17568
rect 17152 -18272 17856 -17568
rect 18564 -18272 19268 -17568
rect 19976 -18272 20680 -17568
rect 21388 -18272 22092 -17568
rect 22800 -18272 23504 -17568
<< metal4 >>
rect -22812 18312 -22716 18348
rect -23805 18272 -23083 18281
rect -23805 17568 -23796 18272
rect -23092 17568 -23083 18272
rect -23805 17559 -23083 17568
rect -22812 18248 -22796 18312
rect -22732 18248 -22716 18312
rect -21400 18312 -21304 18348
rect -22812 18232 -22716 18248
rect -22812 18168 -22796 18232
rect -22732 18168 -22716 18232
rect -22812 18152 -22716 18168
rect -22812 18088 -22796 18152
rect -22732 18088 -22716 18152
rect -22812 18072 -22716 18088
rect -22812 18008 -22796 18072
rect -22732 18008 -22716 18072
rect -22812 17992 -22716 18008
rect -22812 17928 -22796 17992
rect -22732 17928 -22716 17992
rect -22812 17912 -22716 17928
rect -22812 17848 -22796 17912
rect -22732 17848 -22716 17912
rect -22812 17832 -22716 17848
rect -22812 17768 -22796 17832
rect -22732 17768 -22716 17832
rect -22812 17752 -22716 17768
rect -22812 17688 -22796 17752
rect -22732 17688 -22716 17752
rect -22812 17672 -22716 17688
rect -22812 17608 -22796 17672
rect -22732 17608 -22716 17672
rect -22812 17592 -22716 17608
rect -22812 17528 -22796 17592
rect -22732 17528 -22716 17592
rect -22393 18272 -21671 18281
rect -22393 17568 -22384 18272
rect -21680 17568 -21671 18272
rect -22393 17559 -21671 17568
rect -21400 18248 -21384 18312
rect -21320 18248 -21304 18312
rect -19988 18312 -19892 18348
rect -21400 18232 -21304 18248
rect -21400 18168 -21384 18232
rect -21320 18168 -21304 18232
rect -21400 18152 -21304 18168
rect -21400 18088 -21384 18152
rect -21320 18088 -21304 18152
rect -21400 18072 -21304 18088
rect -21400 18008 -21384 18072
rect -21320 18008 -21304 18072
rect -21400 17992 -21304 18008
rect -21400 17928 -21384 17992
rect -21320 17928 -21304 17992
rect -21400 17912 -21304 17928
rect -21400 17848 -21384 17912
rect -21320 17848 -21304 17912
rect -21400 17832 -21304 17848
rect -21400 17768 -21384 17832
rect -21320 17768 -21304 17832
rect -21400 17752 -21304 17768
rect -21400 17688 -21384 17752
rect -21320 17688 -21304 17752
rect -21400 17672 -21304 17688
rect -21400 17608 -21384 17672
rect -21320 17608 -21304 17672
rect -21400 17592 -21304 17608
rect -22812 17492 -22716 17528
rect -21400 17528 -21384 17592
rect -21320 17528 -21304 17592
rect -20981 18272 -20259 18281
rect -20981 17568 -20972 18272
rect -20268 17568 -20259 18272
rect -20981 17559 -20259 17568
rect -19988 18248 -19972 18312
rect -19908 18248 -19892 18312
rect -18576 18312 -18480 18348
rect -19988 18232 -19892 18248
rect -19988 18168 -19972 18232
rect -19908 18168 -19892 18232
rect -19988 18152 -19892 18168
rect -19988 18088 -19972 18152
rect -19908 18088 -19892 18152
rect -19988 18072 -19892 18088
rect -19988 18008 -19972 18072
rect -19908 18008 -19892 18072
rect -19988 17992 -19892 18008
rect -19988 17928 -19972 17992
rect -19908 17928 -19892 17992
rect -19988 17912 -19892 17928
rect -19988 17848 -19972 17912
rect -19908 17848 -19892 17912
rect -19988 17832 -19892 17848
rect -19988 17768 -19972 17832
rect -19908 17768 -19892 17832
rect -19988 17752 -19892 17768
rect -19988 17688 -19972 17752
rect -19908 17688 -19892 17752
rect -19988 17672 -19892 17688
rect -19988 17608 -19972 17672
rect -19908 17608 -19892 17672
rect -19988 17592 -19892 17608
rect -21400 17492 -21304 17528
rect -19988 17528 -19972 17592
rect -19908 17528 -19892 17592
rect -19569 18272 -18847 18281
rect -19569 17568 -19560 18272
rect -18856 17568 -18847 18272
rect -19569 17559 -18847 17568
rect -18576 18248 -18560 18312
rect -18496 18248 -18480 18312
rect -17164 18312 -17068 18348
rect -18576 18232 -18480 18248
rect -18576 18168 -18560 18232
rect -18496 18168 -18480 18232
rect -18576 18152 -18480 18168
rect -18576 18088 -18560 18152
rect -18496 18088 -18480 18152
rect -18576 18072 -18480 18088
rect -18576 18008 -18560 18072
rect -18496 18008 -18480 18072
rect -18576 17992 -18480 18008
rect -18576 17928 -18560 17992
rect -18496 17928 -18480 17992
rect -18576 17912 -18480 17928
rect -18576 17848 -18560 17912
rect -18496 17848 -18480 17912
rect -18576 17832 -18480 17848
rect -18576 17768 -18560 17832
rect -18496 17768 -18480 17832
rect -18576 17752 -18480 17768
rect -18576 17688 -18560 17752
rect -18496 17688 -18480 17752
rect -18576 17672 -18480 17688
rect -18576 17608 -18560 17672
rect -18496 17608 -18480 17672
rect -18576 17592 -18480 17608
rect -19988 17492 -19892 17528
rect -18576 17528 -18560 17592
rect -18496 17528 -18480 17592
rect -18157 18272 -17435 18281
rect -18157 17568 -18148 18272
rect -17444 17568 -17435 18272
rect -18157 17559 -17435 17568
rect -17164 18248 -17148 18312
rect -17084 18248 -17068 18312
rect -15752 18312 -15656 18348
rect -17164 18232 -17068 18248
rect -17164 18168 -17148 18232
rect -17084 18168 -17068 18232
rect -17164 18152 -17068 18168
rect -17164 18088 -17148 18152
rect -17084 18088 -17068 18152
rect -17164 18072 -17068 18088
rect -17164 18008 -17148 18072
rect -17084 18008 -17068 18072
rect -17164 17992 -17068 18008
rect -17164 17928 -17148 17992
rect -17084 17928 -17068 17992
rect -17164 17912 -17068 17928
rect -17164 17848 -17148 17912
rect -17084 17848 -17068 17912
rect -17164 17832 -17068 17848
rect -17164 17768 -17148 17832
rect -17084 17768 -17068 17832
rect -17164 17752 -17068 17768
rect -17164 17688 -17148 17752
rect -17084 17688 -17068 17752
rect -17164 17672 -17068 17688
rect -17164 17608 -17148 17672
rect -17084 17608 -17068 17672
rect -17164 17592 -17068 17608
rect -18576 17492 -18480 17528
rect -17164 17528 -17148 17592
rect -17084 17528 -17068 17592
rect -16745 18272 -16023 18281
rect -16745 17568 -16736 18272
rect -16032 17568 -16023 18272
rect -16745 17559 -16023 17568
rect -15752 18248 -15736 18312
rect -15672 18248 -15656 18312
rect -14340 18312 -14244 18348
rect -15752 18232 -15656 18248
rect -15752 18168 -15736 18232
rect -15672 18168 -15656 18232
rect -15752 18152 -15656 18168
rect -15752 18088 -15736 18152
rect -15672 18088 -15656 18152
rect -15752 18072 -15656 18088
rect -15752 18008 -15736 18072
rect -15672 18008 -15656 18072
rect -15752 17992 -15656 18008
rect -15752 17928 -15736 17992
rect -15672 17928 -15656 17992
rect -15752 17912 -15656 17928
rect -15752 17848 -15736 17912
rect -15672 17848 -15656 17912
rect -15752 17832 -15656 17848
rect -15752 17768 -15736 17832
rect -15672 17768 -15656 17832
rect -15752 17752 -15656 17768
rect -15752 17688 -15736 17752
rect -15672 17688 -15656 17752
rect -15752 17672 -15656 17688
rect -15752 17608 -15736 17672
rect -15672 17608 -15656 17672
rect -15752 17592 -15656 17608
rect -17164 17492 -17068 17528
rect -15752 17528 -15736 17592
rect -15672 17528 -15656 17592
rect -15333 18272 -14611 18281
rect -15333 17568 -15324 18272
rect -14620 17568 -14611 18272
rect -15333 17559 -14611 17568
rect -14340 18248 -14324 18312
rect -14260 18248 -14244 18312
rect -12928 18312 -12832 18348
rect -14340 18232 -14244 18248
rect -14340 18168 -14324 18232
rect -14260 18168 -14244 18232
rect -14340 18152 -14244 18168
rect -14340 18088 -14324 18152
rect -14260 18088 -14244 18152
rect -14340 18072 -14244 18088
rect -14340 18008 -14324 18072
rect -14260 18008 -14244 18072
rect -14340 17992 -14244 18008
rect -14340 17928 -14324 17992
rect -14260 17928 -14244 17992
rect -14340 17912 -14244 17928
rect -14340 17848 -14324 17912
rect -14260 17848 -14244 17912
rect -14340 17832 -14244 17848
rect -14340 17768 -14324 17832
rect -14260 17768 -14244 17832
rect -14340 17752 -14244 17768
rect -14340 17688 -14324 17752
rect -14260 17688 -14244 17752
rect -14340 17672 -14244 17688
rect -14340 17608 -14324 17672
rect -14260 17608 -14244 17672
rect -14340 17592 -14244 17608
rect -15752 17492 -15656 17528
rect -14340 17528 -14324 17592
rect -14260 17528 -14244 17592
rect -13921 18272 -13199 18281
rect -13921 17568 -13912 18272
rect -13208 17568 -13199 18272
rect -13921 17559 -13199 17568
rect -12928 18248 -12912 18312
rect -12848 18248 -12832 18312
rect -11516 18312 -11420 18348
rect -12928 18232 -12832 18248
rect -12928 18168 -12912 18232
rect -12848 18168 -12832 18232
rect -12928 18152 -12832 18168
rect -12928 18088 -12912 18152
rect -12848 18088 -12832 18152
rect -12928 18072 -12832 18088
rect -12928 18008 -12912 18072
rect -12848 18008 -12832 18072
rect -12928 17992 -12832 18008
rect -12928 17928 -12912 17992
rect -12848 17928 -12832 17992
rect -12928 17912 -12832 17928
rect -12928 17848 -12912 17912
rect -12848 17848 -12832 17912
rect -12928 17832 -12832 17848
rect -12928 17768 -12912 17832
rect -12848 17768 -12832 17832
rect -12928 17752 -12832 17768
rect -12928 17688 -12912 17752
rect -12848 17688 -12832 17752
rect -12928 17672 -12832 17688
rect -12928 17608 -12912 17672
rect -12848 17608 -12832 17672
rect -12928 17592 -12832 17608
rect -14340 17492 -14244 17528
rect -12928 17528 -12912 17592
rect -12848 17528 -12832 17592
rect -12509 18272 -11787 18281
rect -12509 17568 -12500 18272
rect -11796 17568 -11787 18272
rect -12509 17559 -11787 17568
rect -11516 18248 -11500 18312
rect -11436 18248 -11420 18312
rect -10104 18312 -10008 18348
rect -11516 18232 -11420 18248
rect -11516 18168 -11500 18232
rect -11436 18168 -11420 18232
rect -11516 18152 -11420 18168
rect -11516 18088 -11500 18152
rect -11436 18088 -11420 18152
rect -11516 18072 -11420 18088
rect -11516 18008 -11500 18072
rect -11436 18008 -11420 18072
rect -11516 17992 -11420 18008
rect -11516 17928 -11500 17992
rect -11436 17928 -11420 17992
rect -11516 17912 -11420 17928
rect -11516 17848 -11500 17912
rect -11436 17848 -11420 17912
rect -11516 17832 -11420 17848
rect -11516 17768 -11500 17832
rect -11436 17768 -11420 17832
rect -11516 17752 -11420 17768
rect -11516 17688 -11500 17752
rect -11436 17688 -11420 17752
rect -11516 17672 -11420 17688
rect -11516 17608 -11500 17672
rect -11436 17608 -11420 17672
rect -11516 17592 -11420 17608
rect -12928 17492 -12832 17528
rect -11516 17528 -11500 17592
rect -11436 17528 -11420 17592
rect -11097 18272 -10375 18281
rect -11097 17568 -11088 18272
rect -10384 17568 -10375 18272
rect -11097 17559 -10375 17568
rect -10104 18248 -10088 18312
rect -10024 18248 -10008 18312
rect -8692 18312 -8596 18348
rect -10104 18232 -10008 18248
rect -10104 18168 -10088 18232
rect -10024 18168 -10008 18232
rect -10104 18152 -10008 18168
rect -10104 18088 -10088 18152
rect -10024 18088 -10008 18152
rect -10104 18072 -10008 18088
rect -10104 18008 -10088 18072
rect -10024 18008 -10008 18072
rect -10104 17992 -10008 18008
rect -10104 17928 -10088 17992
rect -10024 17928 -10008 17992
rect -10104 17912 -10008 17928
rect -10104 17848 -10088 17912
rect -10024 17848 -10008 17912
rect -10104 17832 -10008 17848
rect -10104 17768 -10088 17832
rect -10024 17768 -10008 17832
rect -10104 17752 -10008 17768
rect -10104 17688 -10088 17752
rect -10024 17688 -10008 17752
rect -10104 17672 -10008 17688
rect -10104 17608 -10088 17672
rect -10024 17608 -10008 17672
rect -10104 17592 -10008 17608
rect -11516 17492 -11420 17528
rect -10104 17528 -10088 17592
rect -10024 17528 -10008 17592
rect -9685 18272 -8963 18281
rect -9685 17568 -9676 18272
rect -8972 17568 -8963 18272
rect -9685 17559 -8963 17568
rect -8692 18248 -8676 18312
rect -8612 18248 -8596 18312
rect -7280 18312 -7184 18348
rect -8692 18232 -8596 18248
rect -8692 18168 -8676 18232
rect -8612 18168 -8596 18232
rect -8692 18152 -8596 18168
rect -8692 18088 -8676 18152
rect -8612 18088 -8596 18152
rect -8692 18072 -8596 18088
rect -8692 18008 -8676 18072
rect -8612 18008 -8596 18072
rect -8692 17992 -8596 18008
rect -8692 17928 -8676 17992
rect -8612 17928 -8596 17992
rect -8692 17912 -8596 17928
rect -8692 17848 -8676 17912
rect -8612 17848 -8596 17912
rect -8692 17832 -8596 17848
rect -8692 17768 -8676 17832
rect -8612 17768 -8596 17832
rect -8692 17752 -8596 17768
rect -8692 17688 -8676 17752
rect -8612 17688 -8596 17752
rect -8692 17672 -8596 17688
rect -8692 17608 -8676 17672
rect -8612 17608 -8596 17672
rect -8692 17592 -8596 17608
rect -10104 17492 -10008 17528
rect -8692 17528 -8676 17592
rect -8612 17528 -8596 17592
rect -8273 18272 -7551 18281
rect -8273 17568 -8264 18272
rect -7560 17568 -7551 18272
rect -8273 17559 -7551 17568
rect -7280 18248 -7264 18312
rect -7200 18248 -7184 18312
rect -5868 18312 -5772 18348
rect -7280 18232 -7184 18248
rect -7280 18168 -7264 18232
rect -7200 18168 -7184 18232
rect -7280 18152 -7184 18168
rect -7280 18088 -7264 18152
rect -7200 18088 -7184 18152
rect -7280 18072 -7184 18088
rect -7280 18008 -7264 18072
rect -7200 18008 -7184 18072
rect -7280 17992 -7184 18008
rect -7280 17928 -7264 17992
rect -7200 17928 -7184 17992
rect -7280 17912 -7184 17928
rect -7280 17848 -7264 17912
rect -7200 17848 -7184 17912
rect -7280 17832 -7184 17848
rect -7280 17768 -7264 17832
rect -7200 17768 -7184 17832
rect -7280 17752 -7184 17768
rect -7280 17688 -7264 17752
rect -7200 17688 -7184 17752
rect -7280 17672 -7184 17688
rect -7280 17608 -7264 17672
rect -7200 17608 -7184 17672
rect -7280 17592 -7184 17608
rect -8692 17492 -8596 17528
rect -7280 17528 -7264 17592
rect -7200 17528 -7184 17592
rect -6861 18272 -6139 18281
rect -6861 17568 -6852 18272
rect -6148 17568 -6139 18272
rect -6861 17559 -6139 17568
rect -5868 18248 -5852 18312
rect -5788 18248 -5772 18312
rect -4456 18312 -4360 18348
rect -5868 18232 -5772 18248
rect -5868 18168 -5852 18232
rect -5788 18168 -5772 18232
rect -5868 18152 -5772 18168
rect -5868 18088 -5852 18152
rect -5788 18088 -5772 18152
rect -5868 18072 -5772 18088
rect -5868 18008 -5852 18072
rect -5788 18008 -5772 18072
rect -5868 17992 -5772 18008
rect -5868 17928 -5852 17992
rect -5788 17928 -5772 17992
rect -5868 17912 -5772 17928
rect -5868 17848 -5852 17912
rect -5788 17848 -5772 17912
rect -5868 17832 -5772 17848
rect -5868 17768 -5852 17832
rect -5788 17768 -5772 17832
rect -5868 17752 -5772 17768
rect -5868 17688 -5852 17752
rect -5788 17688 -5772 17752
rect -5868 17672 -5772 17688
rect -5868 17608 -5852 17672
rect -5788 17608 -5772 17672
rect -5868 17592 -5772 17608
rect -7280 17492 -7184 17528
rect -5868 17528 -5852 17592
rect -5788 17528 -5772 17592
rect -5449 18272 -4727 18281
rect -5449 17568 -5440 18272
rect -4736 17568 -4727 18272
rect -5449 17559 -4727 17568
rect -4456 18248 -4440 18312
rect -4376 18248 -4360 18312
rect -3044 18312 -2948 18348
rect -4456 18232 -4360 18248
rect -4456 18168 -4440 18232
rect -4376 18168 -4360 18232
rect -4456 18152 -4360 18168
rect -4456 18088 -4440 18152
rect -4376 18088 -4360 18152
rect -4456 18072 -4360 18088
rect -4456 18008 -4440 18072
rect -4376 18008 -4360 18072
rect -4456 17992 -4360 18008
rect -4456 17928 -4440 17992
rect -4376 17928 -4360 17992
rect -4456 17912 -4360 17928
rect -4456 17848 -4440 17912
rect -4376 17848 -4360 17912
rect -4456 17832 -4360 17848
rect -4456 17768 -4440 17832
rect -4376 17768 -4360 17832
rect -4456 17752 -4360 17768
rect -4456 17688 -4440 17752
rect -4376 17688 -4360 17752
rect -4456 17672 -4360 17688
rect -4456 17608 -4440 17672
rect -4376 17608 -4360 17672
rect -4456 17592 -4360 17608
rect -5868 17492 -5772 17528
rect -4456 17528 -4440 17592
rect -4376 17528 -4360 17592
rect -4037 18272 -3315 18281
rect -4037 17568 -4028 18272
rect -3324 17568 -3315 18272
rect -4037 17559 -3315 17568
rect -3044 18248 -3028 18312
rect -2964 18248 -2948 18312
rect -1632 18312 -1536 18348
rect -3044 18232 -2948 18248
rect -3044 18168 -3028 18232
rect -2964 18168 -2948 18232
rect -3044 18152 -2948 18168
rect -3044 18088 -3028 18152
rect -2964 18088 -2948 18152
rect -3044 18072 -2948 18088
rect -3044 18008 -3028 18072
rect -2964 18008 -2948 18072
rect -3044 17992 -2948 18008
rect -3044 17928 -3028 17992
rect -2964 17928 -2948 17992
rect -3044 17912 -2948 17928
rect -3044 17848 -3028 17912
rect -2964 17848 -2948 17912
rect -3044 17832 -2948 17848
rect -3044 17768 -3028 17832
rect -2964 17768 -2948 17832
rect -3044 17752 -2948 17768
rect -3044 17688 -3028 17752
rect -2964 17688 -2948 17752
rect -3044 17672 -2948 17688
rect -3044 17608 -3028 17672
rect -2964 17608 -2948 17672
rect -3044 17592 -2948 17608
rect -4456 17492 -4360 17528
rect -3044 17528 -3028 17592
rect -2964 17528 -2948 17592
rect -2625 18272 -1903 18281
rect -2625 17568 -2616 18272
rect -1912 17568 -1903 18272
rect -2625 17559 -1903 17568
rect -1632 18248 -1616 18312
rect -1552 18248 -1536 18312
rect -220 18312 -124 18348
rect -1632 18232 -1536 18248
rect -1632 18168 -1616 18232
rect -1552 18168 -1536 18232
rect -1632 18152 -1536 18168
rect -1632 18088 -1616 18152
rect -1552 18088 -1536 18152
rect -1632 18072 -1536 18088
rect -1632 18008 -1616 18072
rect -1552 18008 -1536 18072
rect -1632 17992 -1536 18008
rect -1632 17928 -1616 17992
rect -1552 17928 -1536 17992
rect -1632 17912 -1536 17928
rect -1632 17848 -1616 17912
rect -1552 17848 -1536 17912
rect -1632 17832 -1536 17848
rect -1632 17768 -1616 17832
rect -1552 17768 -1536 17832
rect -1632 17752 -1536 17768
rect -1632 17688 -1616 17752
rect -1552 17688 -1536 17752
rect -1632 17672 -1536 17688
rect -1632 17608 -1616 17672
rect -1552 17608 -1536 17672
rect -1632 17592 -1536 17608
rect -3044 17492 -2948 17528
rect -1632 17528 -1616 17592
rect -1552 17528 -1536 17592
rect -1213 18272 -491 18281
rect -1213 17568 -1204 18272
rect -500 17568 -491 18272
rect -1213 17559 -491 17568
rect -220 18248 -204 18312
rect -140 18248 -124 18312
rect 1192 18312 1288 18348
rect -220 18232 -124 18248
rect -220 18168 -204 18232
rect -140 18168 -124 18232
rect -220 18152 -124 18168
rect -220 18088 -204 18152
rect -140 18088 -124 18152
rect -220 18072 -124 18088
rect -220 18008 -204 18072
rect -140 18008 -124 18072
rect -220 17992 -124 18008
rect -220 17928 -204 17992
rect -140 17928 -124 17992
rect -220 17912 -124 17928
rect -220 17848 -204 17912
rect -140 17848 -124 17912
rect -220 17832 -124 17848
rect -220 17768 -204 17832
rect -140 17768 -124 17832
rect -220 17752 -124 17768
rect -220 17688 -204 17752
rect -140 17688 -124 17752
rect -220 17672 -124 17688
rect -220 17608 -204 17672
rect -140 17608 -124 17672
rect -220 17592 -124 17608
rect -1632 17492 -1536 17528
rect -220 17528 -204 17592
rect -140 17528 -124 17592
rect 199 18272 921 18281
rect 199 17568 208 18272
rect 912 17568 921 18272
rect 199 17559 921 17568
rect 1192 18248 1208 18312
rect 1272 18248 1288 18312
rect 2604 18312 2700 18348
rect 1192 18232 1288 18248
rect 1192 18168 1208 18232
rect 1272 18168 1288 18232
rect 1192 18152 1288 18168
rect 1192 18088 1208 18152
rect 1272 18088 1288 18152
rect 1192 18072 1288 18088
rect 1192 18008 1208 18072
rect 1272 18008 1288 18072
rect 1192 17992 1288 18008
rect 1192 17928 1208 17992
rect 1272 17928 1288 17992
rect 1192 17912 1288 17928
rect 1192 17848 1208 17912
rect 1272 17848 1288 17912
rect 1192 17832 1288 17848
rect 1192 17768 1208 17832
rect 1272 17768 1288 17832
rect 1192 17752 1288 17768
rect 1192 17688 1208 17752
rect 1272 17688 1288 17752
rect 1192 17672 1288 17688
rect 1192 17608 1208 17672
rect 1272 17608 1288 17672
rect 1192 17592 1288 17608
rect -220 17492 -124 17528
rect 1192 17528 1208 17592
rect 1272 17528 1288 17592
rect 1611 18272 2333 18281
rect 1611 17568 1620 18272
rect 2324 17568 2333 18272
rect 1611 17559 2333 17568
rect 2604 18248 2620 18312
rect 2684 18248 2700 18312
rect 4016 18312 4112 18348
rect 2604 18232 2700 18248
rect 2604 18168 2620 18232
rect 2684 18168 2700 18232
rect 2604 18152 2700 18168
rect 2604 18088 2620 18152
rect 2684 18088 2700 18152
rect 2604 18072 2700 18088
rect 2604 18008 2620 18072
rect 2684 18008 2700 18072
rect 2604 17992 2700 18008
rect 2604 17928 2620 17992
rect 2684 17928 2700 17992
rect 2604 17912 2700 17928
rect 2604 17848 2620 17912
rect 2684 17848 2700 17912
rect 2604 17832 2700 17848
rect 2604 17768 2620 17832
rect 2684 17768 2700 17832
rect 2604 17752 2700 17768
rect 2604 17688 2620 17752
rect 2684 17688 2700 17752
rect 2604 17672 2700 17688
rect 2604 17608 2620 17672
rect 2684 17608 2700 17672
rect 2604 17592 2700 17608
rect 1192 17492 1288 17528
rect 2604 17528 2620 17592
rect 2684 17528 2700 17592
rect 3023 18272 3745 18281
rect 3023 17568 3032 18272
rect 3736 17568 3745 18272
rect 3023 17559 3745 17568
rect 4016 18248 4032 18312
rect 4096 18248 4112 18312
rect 5428 18312 5524 18348
rect 4016 18232 4112 18248
rect 4016 18168 4032 18232
rect 4096 18168 4112 18232
rect 4016 18152 4112 18168
rect 4016 18088 4032 18152
rect 4096 18088 4112 18152
rect 4016 18072 4112 18088
rect 4016 18008 4032 18072
rect 4096 18008 4112 18072
rect 4016 17992 4112 18008
rect 4016 17928 4032 17992
rect 4096 17928 4112 17992
rect 4016 17912 4112 17928
rect 4016 17848 4032 17912
rect 4096 17848 4112 17912
rect 4016 17832 4112 17848
rect 4016 17768 4032 17832
rect 4096 17768 4112 17832
rect 4016 17752 4112 17768
rect 4016 17688 4032 17752
rect 4096 17688 4112 17752
rect 4016 17672 4112 17688
rect 4016 17608 4032 17672
rect 4096 17608 4112 17672
rect 4016 17592 4112 17608
rect 2604 17492 2700 17528
rect 4016 17528 4032 17592
rect 4096 17528 4112 17592
rect 4435 18272 5157 18281
rect 4435 17568 4444 18272
rect 5148 17568 5157 18272
rect 4435 17559 5157 17568
rect 5428 18248 5444 18312
rect 5508 18248 5524 18312
rect 6840 18312 6936 18348
rect 5428 18232 5524 18248
rect 5428 18168 5444 18232
rect 5508 18168 5524 18232
rect 5428 18152 5524 18168
rect 5428 18088 5444 18152
rect 5508 18088 5524 18152
rect 5428 18072 5524 18088
rect 5428 18008 5444 18072
rect 5508 18008 5524 18072
rect 5428 17992 5524 18008
rect 5428 17928 5444 17992
rect 5508 17928 5524 17992
rect 5428 17912 5524 17928
rect 5428 17848 5444 17912
rect 5508 17848 5524 17912
rect 5428 17832 5524 17848
rect 5428 17768 5444 17832
rect 5508 17768 5524 17832
rect 5428 17752 5524 17768
rect 5428 17688 5444 17752
rect 5508 17688 5524 17752
rect 5428 17672 5524 17688
rect 5428 17608 5444 17672
rect 5508 17608 5524 17672
rect 5428 17592 5524 17608
rect 4016 17492 4112 17528
rect 5428 17528 5444 17592
rect 5508 17528 5524 17592
rect 5847 18272 6569 18281
rect 5847 17568 5856 18272
rect 6560 17568 6569 18272
rect 5847 17559 6569 17568
rect 6840 18248 6856 18312
rect 6920 18248 6936 18312
rect 8252 18312 8348 18348
rect 6840 18232 6936 18248
rect 6840 18168 6856 18232
rect 6920 18168 6936 18232
rect 6840 18152 6936 18168
rect 6840 18088 6856 18152
rect 6920 18088 6936 18152
rect 6840 18072 6936 18088
rect 6840 18008 6856 18072
rect 6920 18008 6936 18072
rect 6840 17992 6936 18008
rect 6840 17928 6856 17992
rect 6920 17928 6936 17992
rect 6840 17912 6936 17928
rect 6840 17848 6856 17912
rect 6920 17848 6936 17912
rect 6840 17832 6936 17848
rect 6840 17768 6856 17832
rect 6920 17768 6936 17832
rect 6840 17752 6936 17768
rect 6840 17688 6856 17752
rect 6920 17688 6936 17752
rect 6840 17672 6936 17688
rect 6840 17608 6856 17672
rect 6920 17608 6936 17672
rect 6840 17592 6936 17608
rect 5428 17492 5524 17528
rect 6840 17528 6856 17592
rect 6920 17528 6936 17592
rect 7259 18272 7981 18281
rect 7259 17568 7268 18272
rect 7972 17568 7981 18272
rect 7259 17559 7981 17568
rect 8252 18248 8268 18312
rect 8332 18248 8348 18312
rect 9664 18312 9760 18348
rect 8252 18232 8348 18248
rect 8252 18168 8268 18232
rect 8332 18168 8348 18232
rect 8252 18152 8348 18168
rect 8252 18088 8268 18152
rect 8332 18088 8348 18152
rect 8252 18072 8348 18088
rect 8252 18008 8268 18072
rect 8332 18008 8348 18072
rect 8252 17992 8348 18008
rect 8252 17928 8268 17992
rect 8332 17928 8348 17992
rect 8252 17912 8348 17928
rect 8252 17848 8268 17912
rect 8332 17848 8348 17912
rect 8252 17832 8348 17848
rect 8252 17768 8268 17832
rect 8332 17768 8348 17832
rect 8252 17752 8348 17768
rect 8252 17688 8268 17752
rect 8332 17688 8348 17752
rect 8252 17672 8348 17688
rect 8252 17608 8268 17672
rect 8332 17608 8348 17672
rect 8252 17592 8348 17608
rect 6840 17492 6936 17528
rect 8252 17528 8268 17592
rect 8332 17528 8348 17592
rect 8671 18272 9393 18281
rect 8671 17568 8680 18272
rect 9384 17568 9393 18272
rect 8671 17559 9393 17568
rect 9664 18248 9680 18312
rect 9744 18248 9760 18312
rect 11076 18312 11172 18348
rect 9664 18232 9760 18248
rect 9664 18168 9680 18232
rect 9744 18168 9760 18232
rect 9664 18152 9760 18168
rect 9664 18088 9680 18152
rect 9744 18088 9760 18152
rect 9664 18072 9760 18088
rect 9664 18008 9680 18072
rect 9744 18008 9760 18072
rect 9664 17992 9760 18008
rect 9664 17928 9680 17992
rect 9744 17928 9760 17992
rect 9664 17912 9760 17928
rect 9664 17848 9680 17912
rect 9744 17848 9760 17912
rect 9664 17832 9760 17848
rect 9664 17768 9680 17832
rect 9744 17768 9760 17832
rect 9664 17752 9760 17768
rect 9664 17688 9680 17752
rect 9744 17688 9760 17752
rect 9664 17672 9760 17688
rect 9664 17608 9680 17672
rect 9744 17608 9760 17672
rect 9664 17592 9760 17608
rect 8252 17492 8348 17528
rect 9664 17528 9680 17592
rect 9744 17528 9760 17592
rect 10083 18272 10805 18281
rect 10083 17568 10092 18272
rect 10796 17568 10805 18272
rect 10083 17559 10805 17568
rect 11076 18248 11092 18312
rect 11156 18248 11172 18312
rect 12488 18312 12584 18348
rect 11076 18232 11172 18248
rect 11076 18168 11092 18232
rect 11156 18168 11172 18232
rect 11076 18152 11172 18168
rect 11076 18088 11092 18152
rect 11156 18088 11172 18152
rect 11076 18072 11172 18088
rect 11076 18008 11092 18072
rect 11156 18008 11172 18072
rect 11076 17992 11172 18008
rect 11076 17928 11092 17992
rect 11156 17928 11172 17992
rect 11076 17912 11172 17928
rect 11076 17848 11092 17912
rect 11156 17848 11172 17912
rect 11076 17832 11172 17848
rect 11076 17768 11092 17832
rect 11156 17768 11172 17832
rect 11076 17752 11172 17768
rect 11076 17688 11092 17752
rect 11156 17688 11172 17752
rect 11076 17672 11172 17688
rect 11076 17608 11092 17672
rect 11156 17608 11172 17672
rect 11076 17592 11172 17608
rect 9664 17492 9760 17528
rect 11076 17528 11092 17592
rect 11156 17528 11172 17592
rect 11495 18272 12217 18281
rect 11495 17568 11504 18272
rect 12208 17568 12217 18272
rect 11495 17559 12217 17568
rect 12488 18248 12504 18312
rect 12568 18248 12584 18312
rect 13900 18312 13996 18348
rect 12488 18232 12584 18248
rect 12488 18168 12504 18232
rect 12568 18168 12584 18232
rect 12488 18152 12584 18168
rect 12488 18088 12504 18152
rect 12568 18088 12584 18152
rect 12488 18072 12584 18088
rect 12488 18008 12504 18072
rect 12568 18008 12584 18072
rect 12488 17992 12584 18008
rect 12488 17928 12504 17992
rect 12568 17928 12584 17992
rect 12488 17912 12584 17928
rect 12488 17848 12504 17912
rect 12568 17848 12584 17912
rect 12488 17832 12584 17848
rect 12488 17768 12504 17832
rect 12568 17768 12584 17832
rect 12488 17752 12584 17768
rect 12488 17688 12504 17752
rect 12568 17688 12584 17752
rect 12488 17672 12584 17688
rect 12488 17608 12504 17672
rect 12568 17608 12584 17672
rect 12488 17592 12584 17608
rect 11076 17492 11172 17528
rect 12488 17528 12504 17592
rect 12568 17528 12584 17592
rect 12907 18272 13629 18281
rect 12907 17568 12916 18272
rect 13620 17568 13629 18272
rect 12907 17559 13629 17568
rect 13900 18248 13916 18312
rect 13980 18248 13996 18312
rect 15312 18312 15408 18348
rect 13900 18232 13996 18248
rect 13900 18168 13916 18232
rect 13980 18168 13996 18232
rect 13900 18152 13996 18168
rect 13900 18088 13916 18152
rect 13980 18088 13996 18152
rect 13900 18072 13996 18088
rect 13900 18008 13916 18072
rect 13980 18008 13996 18072
rect 13900 17992 13996 18008
rect 13900 17928 13916 17992
rect 13980 17928 13996 17992
rect 13900 17912 13996 17928
rect 13900 17848 13916 17912
rect 13980 17848 13996 17912
rect 13900 17832 13996 17848
rect 13900 17768 13916 17832
rect 13980 17768 13996 17832
rect 13900 17752 13996 17768
rect 13900 17688 13916 17752
rect 13980 17688 13996 17752
rect 13900 17672 13996 17688
rect 13900 17608 13916 17672
rect 13980 17608 13996 17672
rect 13900 17592 13996 17608
rect 12488 17492 12584 17528
rect 13900 17528 13916 17592
rect 13980 17528 13996 17592
rect 14319 18272 15041 18281
rect 14319 17568 14328 18272
rect 15032 17568 15041 18272
rect 14319 17559 15041 17568
rect 15312 18248 15328 18312
rect 15392 18248 15408 18312
rect 16724 18312 16820 18348
rect 15312 18232 15408 18248
rect 15312 18168 15328 18232
rect 15392 18168 15408 18232
rect 15312 18152 15408 18168
rect 15312 18088 15328 18152
rect 15392 18088 15408 18152
rect 15312 18072 15408 18088
rect 15312 18008 15328 18072
rect 15392 18008 15408 18072
rect 15312 17992 15408 18008
rect 15312 17928 15328 17992
rect 15392 17928 15408 17992
rect 15312 17912 15408 17928
rect 15312 17848 15328 17912
rect 15392 17848 15408 17912
rect 15312 17832 15408 17848
rect 15312 17768 15328 17832
rect 15392 17768 15408 17832
rect 15312 17752 15408 17768
rect 15312 17688 15328 17752
rect 15392 17688 15408 17752
rect 15312 17672 15408 17688
rect 15312 17608 15328 17672
rect 15392 17608 15408 17672
rect 15312 17592 15408 17608
rect 13900 17492 13996 17528
rect 15312 17528 15328 17592
rect 15392 17528 15408 17592
rect 15731 18272 16453 18281
rect 15731 17568 15740 18272
rect 16444 17568 16453 18272
rect 15731 17559 16453 17568
rect 16724 18248 16740 18312
rect 16804 18248 16820 18312
rect 18136 18312 18232 18348
rect 16724 18232 16820 18248
rect 16724 18168 16740 18232
rect 16804 18168 16820 18232
rect 16724 18152 16820 18168
rect 16724 18088 16740 18152
rect 16804 18088 16820 18152
rect 16724 18072 16820 18088
rect 16724 18008 16740 18072
rect 16804 18008 16820 18072
rect 16724 17992 16820 18008
rect 16724 17928 16740 17992
rect 16804 17928 16820 17992
rect 16724 17912 16820 17928
rect 16724 17848 16740 17912
rect 16804 17848 16820 17912
rect 16724 17832 16820 17848
rect 16724 17768 16740 17832
rect 16804 17768 16820 17832
rect 16724 17752 16820 17768
rect 16724 17688 16740 17752
rect 16804 17688 16820 17752
rect 16724 17672 16820 17688
rect 16724 17608 16740 17672
rect 16804 17608 16820 17672
rect 16724 17592 16820 17608
rect 15312 17492 15408 17528
rect 16724 17528 16740 17592
rect 16804 17528 16820 17592
rect 17143 18272 17865 18281
rect 17143 17568 17152 18272
rect 17856 17568 17865 18272
rect 17143 17559 17865 17568
rect 18136 18248 18152 18312
rect 18216 18248 18232 18312
rect 19548 18312 19644 18348
rect 18136 18232 18232 18248
rect 18136 18168 18152 18232
rect 18216 18168 18232 18232
rect 18136 18152 18232 18168
rect 18136 18088 18152 18152
rect 18216 18088 18232 18152
rect 18136 18072 18232 18088
rect 18136 18008 18152 18072
rect 18216 18008 18232 18072
rect 18136 17992 18232 18008
rect 18136 17928 18152 17992
rect 18216 17928 18232 17992
rect 18136 17912 18232 17928
rect 18136 17848 18152 17912
rect 18216 17848 18232 17912
rect 18136 17832 18232 17848
rect 18136 17768 18152 17832
rect 18216 17768 18232 17832
rect 18136 17752 18232 17768
rect 18136 17688 18152 17752
rect 18216 17688 18232 17752
rect 18136 17672 18232 17688
rect 18136 17608 18152 17672
rect 18216 17608 18232 17672
rect 18136 17592 18232 17608
rect 16724 17492 16820 17528
rect 18136 17528 18152 17592
rect 18216 17528 18232 17592
rect 18555 18272 19277 18281
rect 18555 17568 18564 18272
rect 19268 17568 19277 18272
rect 18555 17559 19277 17568
rect 19548 18248 19564 18312
rect 19628 18248 19644 18312
rect 20960 18312 21056 18348
rect 19548 18232 19644 18248
rect 19548 18168 19564 18232
rect 19628 18168 19644 18232
rect 19548 18152 19644 18168
rect 19548 18088 19564 18152
rect 19628 18088 19644 18152
rect 19548 18072 19644 18088
rect 19548 18008 19564 18072
rect 19628 18008 19644 18072
rect 19548 17992 19644 18008
rect 19548 17928 19564 17992
rect 19628 17928 19644 17992
rect 19548 17912 19644 17928
rect 19548 17848 19564 17912
rect 19628 17848 19644 17912
rect 19548 17832 19644 17848
rect 19548 17768 19564 17832
rect 19628 17768 19644 17832
rect 19548 17752 19644 17768
rect 19548 17688 19564 17752
rect 19628 17688 19644 17752
rect 19548 17672 19644 17688
rect 19548 17608 19564 17672
rect 19628 17608 19644 17672
rect 19548 17592 19644 17608
rect 18136 17492 18232 17528
rect 19548 17528 19564 17592
rect 19628 17528 19644 17592
rect 19967 18272 20689 18281
rect 19967 17568 19976 18272
rect 20680 17568 20689 18272
rect 19967 17559 20689 17568
rect 20960 18248 20976 18312
rect 21040 18248 21056 18312
rect 22372 18312 22468 18348
rect 20960 18232 21056 18248
rect 20960 18168 20976 18232
rect 21040 18168 21056 18232
rect 20960 18152 21056 18168
rect 20960 18088 20976 18152
rect 21040 18088 21056 18152
rect 20960 18072 21056 18088
rect 20960 18008 20976 18072
rect 21040 18008 21056 18072
rect 20960 17992 21056 18008
rect 20960 17928 20976 17992
rect 21040 17928 21056 17992
rect 20960 17912 21056 17928
rect 20960 17848 20976 17912
rect 21040 17848 21056 17912
rect 20960 17832 21056 17848
rect 20960 17768 20976 17832
rect 21040 17768 21056 17832
rect 20960 17752 21056 17768
rect 20960 17688 20976 17752
rect 21040 17688 21056 17752
rect 20960 17672 21056 17688
rect 20960 17608 20976 17672
rect 21040 17608 21056 17672
rect 20960 17592 21056 17608
rect 19548 17492 19644 17528
rect 20960 17528 20976 17592
rect 21040 17528 21056 17592
rect 21379 18272 22101 18281
rect 21379 17568 21388 18272
rect 22092 17568 22101 18272
rect 21379 17559 22101 17568
rect 22372 18248 22388 18312
rect 22452 18248 22468 18312
rect 23784 18312 23880 18348
rect 22372 18232 22468 18248
rect 22372 18168 22388 18232
rect 22452 18168 22468 18232
rect 22372 18152 22468 18168
rect 22372 18088 22388 18152
rect 22452 18088 22468 18152
rect 22372 18072 22468 18088
rect 22372 18008 22388 18072
rect 22452 18008 22468 18072
rect 22372 17992 22468 18008
rect 22372 17928 22388 17992
rect 22452 17928 22468 17992
rect 22372 17912 22468 17928
rect 22372 17848 22388 17912
rect 22452 17848 22468 17912
rect 22372 17832 22468 17848
rect 22372 17768 22388 17832
rect 22452 17768 22468 17832
rect 22372 17752 22468 17768
rect 22372 17688 22388 17752
rect 22452 17688 22468 17752
rect 22372 17672 22468 17688
rect 22372 17608 22388 17672
rect 22452 17608 22468 17672
rect 22372 17592 22468 17608
rect 20960 17492 21056 17528
rect 22372 17528 22388 17592
rect 22452 17528 22468 17592
rect 22791 18272 23513 18281
rect 22791 17568 22800 18272
rect 23504 17568 23513 18272
rect 22791 17559 23513 17568
rect 23784 18248 23800 18312
rect 23864 18248 23880 18312
rect 23784 18232 23880 18248
rect 23784 18168 23800 18232
rect 23864 18168 23880 18232
rect 23784 18152 23880 18168
rect 23784 18088 23800 18152
rect 23864 18088 23880 18152
rect 23784 18072 23880 18088
rect 23784 18008 23800 18072
rect 23864 18008 23880 18072
rect 23784 17992 23880 18008
rect 23784 17928 23800 17992
rect 23864 17928 23880 17992
rect 23784 17912 23880 17928
rect 23784 17848 23800 17912
rect 23864 17848 23880 17912
rect 23784 17832 23880 17848
rect 23784 17768 23800 17832
rect 23864 17768 23880 17832
rect 23784 17752 23880 17768
rect 23784 17688 23800 17752
rect 23864 17688 23880 17752
rect 23784 17672 23880 17688
rect 23784 17608 23800 17672
rect 23864 17608 23880 17672
rect 23784 17592 23880 17608
rect 22372 17492 22468 17528
rect 23784 17528 23800 17592
rect 23864 17528 23880 17592
rect 23784 17492 23880 17528
rect -22812 17192 -22716 17228
rect -23805 17152 -23083 17161
rect -23805 16448 -23796 17152
rect -23092 16448 -23083 17152
rect -23805 16439 -23083 16448
rect -22812 17128 -22796 17192
rect -22732 17128 -22716 17192
rect -21400 17192 -21304 17228
rect -22812 17112 -22716 17128
rect -22812 17048 -22796 17112
rect -22732 17048 -22716 17112
rect -22812 17032 -22716 17048
rect -22812 16968 -22796 17032
rect -22732 16968 -22716 17032
rect -22812 16952 -22716 16968
rect -22812 16888 -22796 16952
rect -22732 16888 -22716 16952
rect -22812 16872 -22716 16888
rect -22812 16808 -22796 16872
rect -22732 16808 -22716 16872
rect -22812 16792 -22716 16808
rect -22812 16728 -22796 16792
rect -22732 16728 -22716 16792
rect -22812 16712 -22716 16728
rect -22812 16648 -22796 16712
rect -22732 16648 -22716 16712
rect -22812 16632 -22716 16648
rect -22812 16568 -22796 16632
rect -22732 16568 -22716 16632
rect -22812 16552 -22716 16568
rect -22812 16488 -22796 16552
rect -22732 16488 -22716 16552
rect -22812 16472 -22716 16488
rect -22812 16408 -22796 16472
rect -22732 16408 -22716 16472
rect -22393 17152 -21671 17161
rect -22393 16448 -22384 17152
rect -21680 16448 -21671 17152
rect -22393 16439 -21671 16448
rect -21400 17128 -21384 17192
rect -21320 17128 -21304 17192
rect -19988 17192 -19892 17228
rect -21400 17112 -21304 17128
rect -21400 17048 -21384 17112
rect -21320 17048 -21304 17112
rect -21400 17032 -21304 17048
rect -21400 16968 -21384 17032
rect -21320 16968 -21304 17032
rect -21400 16952 -21304 16968
rect -21400 16888 -21384 16952
rect -21320 16888 -21304 16952
rect -21400 16872 -21304 16888
rect -21400 16808 -21384 16872
rect -21320 16808 -21304 16872
rect -21400 16792 -21304 16808
rect -21400 16728 -21384 16792
rect -21320 16728 -21304 16792
rect -21400 16712 -21304 16728
rect -21400 16648 -21384 16712
rect -21320 16648 -21304 16712
rect -21400 16632 -21304 16648
rect -21400 16568 -21384 16632
rect -21320 16568 -21304 16632
rect -21400 16552 -21304 16568
rect -21400 16488 -21384 16552
rect -21320 16488 -21304 16552
rect -21400 16472 -21304 16488
rect -22812 16372 -22716 16408
rect -21400 16408 -21384 16472
rect -21320 16408 -21304 16472
rect -20981 17152 -20259 17161
rect -20981 16448 -20972 17152
rect -20268 16448 -20259 17152
rect -20981 16439 -20259 16448
rect -19988 17128 -19972 17192
rect -19908 17128 -19892 17192
rect -18576 17192 -18480 17228
rect -19988 17112 -19892 17128
rect -19988 17048 -19972 17112
rect -19908 17048 -19892 17112
rect -19988 17032 -19892 17048
rect -19988 16968 -19972 17032
rect -19908 16968 -19892 17032
rect -19988 16952 -19892 16968
rect -19988 16888 -19972 16952
rect -19908 16888 -19892 16952
rect -19988 16872 -19892 16888
rect -19988 16808 -19972 16872
rect -19908 16808 -19892 16872
rect -19988 16792 -19892 16808
rect -19988 16728 -19972 16792
rect -19908 16728 -19892 16792
rect -19988 16712 -19892 16728
rect -19988 16648 -19972 16712
rect -19908 16648 -19892 16712
rect -19988 16632 -19892 16648
rect -19988 16568 -19972 16632
rect -19908 16568 -19892 16632
rect -19988 16552 -19892 16568
rect -19988 16488 -19972 16552
rect -19908 16488 -19892 16552
rect -19988 16472 -19892 16488
rect -21400 16372 -21304 16408
rect -19988 16408 -19972 16472
rect -19908 16408 -19892 16472
rect -19569 17152 -18847 17161
rect -19569 16448 -19560 17152
rect -18856 16448 -18847 17152
rect -19569 16439 -18847 16448
rect -18576 17128 -18560 17192
rect -18496 17128 -18480 17192
rect -17164 17192 -17068 17228
rect -18576 17112 -18480 17128
rect -18576 17048 -18560 17112
rect -18496 17048 -18480 17112
rect -18576 17032 -18480 17048
rect -18576 16968 -18560 17032
rect -18496 16968 -18480 17032
rect -18576 16952 -18480 16968
rect -18576 16888 -18560 16952
rect -18496 16888 -18480 16952
rect -18576 16872 -18480 16888
rect -18576 16808 -18560 16872
rect -18496 16808 -18480 16872
rect -18576 16792 -18480 16808
rect -18576 16728 -18560 16792
rect -18496 16728 -18480 16792
rect -18576 16712 -18480 16728
rect -18576 16648 -18560 16712
rect -18496 16648 -18480 16712
rect -18576 16632 -18480 16648
rect -18576 16568 -18560 16632
rect -18496 16568 -18480 16632
rect -18576 16552 -18480 16568
rect -18576 16488 -18560 16552
rect -18496 16488 -18480 16552
rect -18576 16472 -18480 16488
rect -19988 16372 -19892 16408
rect -18576 16408 -18560 16472
rect -18496 16408 -18480 16472
rect -18157 17152 -17435 17161
rect -18157 16448 -18148 17152
rect -17444 16448 -17435 17152
rect -18157 16439 -17435 16448
rect -17164 17128 -17148 17192
rect -17084 17128 -17068 17192
rect -15752 17192 -15656 17228
rect -17164 17112 -17068 17128
rect -17164 17048 -17148 17112
rect -17084 17048 -17068 17112
rect -17164 17032 -17068 17048
rect -17164 16968 -17148 17032
rect -17084 16968 -17068 17032
rect -17164 16952 -17068 16968
rect -17164 16888 -17148 16952
rect -17084 16888 -17068 16952
rect -17164 16872 -17068 16888
rect -17164 16808 -17148 16872
rect -17084 16808 -17068 16872
rect -17164 16792 -17068 16808
rect -17164 16728 -17148 16792
rect -17084 16728 -17068 16792
rect -17164 16712 -17068 16728
rect -17164 16648 -17148 16712
rect -17084 16648 -17068 16712
rect -17164 16632 -17068 16648
rect -17164 16568 -17148 16632
rect -17084 16568 -17068 16632
rect -17164 16552 -17068 16568
rect -17164 16488 -17148 16552
rect -17084 16488 -17068 16552
rect -17164 16472 -17068 16488
rect -18576 16372 -18480 16408
rect -17164 16408 -17148 16472
rect -17084 16408 -17068 16472
rect -16745 17152 -16023 17161
rect -16745 16448 -16736 17152
rect -16032 16448 -16023 17152
rect -16745 16439 -16023 16448
rect -15752 17128 -15736 17192
rect -15672 17128 -15656 17192
rect -14340 17192 -14244 17228
rect -15752 17112 -15656 17128
rect -15752 17048 -15736 17112
rect -15672 17048 -15656 17112
rect -15752 17032 -15656 17048
rect -15752 16968 -15736 17032
rect -15672 16968 -15656 17032
rect -15752 16952 -15656 16968
rect -15752 16888 -15736 16952
rect -15672 16888 -15656 16952
rect -15752 16872 -15656 16888
rect -15752 16808 -15736 16872
rect -15672 16808 -15656 16872
rect -15752 16792 -15656 16808
rect -15752 16728 -15736 16792
rect -15672 16728 -15656 16792
rect -15752 16712 -15656 16728
rect -15752 16648 -15736 16712
rect -15672 16648 -15656 16712
rect -15752 16632 -15656 16648
rect -15752 16568 -15736 16632
rect -15672 16568 -15656 16632
rect -15752 16552 -15656 16568
rect -15752 16488 -15736 16552
rect -15672 16488 -15656 16552
rect -15752 16472 -15656 16488
rect -17164 16372 -17068 16408
rect -15752 16408 -15736 16472
rect -15672 16408 -15656 16472
rect -15333 17152 -14611 17161
rect -15333 16448 -15324 17152
rect -14620 16448 -14611 17152
rect -15333 16439 -14611 16448
rect -14340 17128 -14324 17192
rect -14260 17128 -14244 17192
rect -12928 17192 -12832 17228
rect -14340 17112 -14244 17128
rect -14340 17048 -14324 17112
rect -14260 17048 -14244 17112
rect -14340 17032 -14244 17048
rect -14340 16968 -14324 17032
rect -14260 16968 -14244 17032
rect -14340 16952 -14244 16968
rect -14340 16888 -14324 16952
rect -14260 16888 -14244 16952
rect -14340 16872 -14244 16888
rect -14340 16808 -14324 16872
rect -14260 16808 -14244 16872
rect -14340 16792 -14244 16808
rect -14340 16728 -14324 16792
rect -14260 16728 -14244 16792
rect -14340 16712 -14244 16728
rect -14340 16648 -14324 16712
rect -14260 16648 -14244 16712
rect -14340 16632 -14244 16648
rect -14340 16568 -14324 16632
rect -14260 16568 -14244 16632
rect -14340 16552 -14244 16568
rect -14340 16488 -14324 16552
rect -14260 16488 -14244 16552
rect -14340 16472 -14244 16488
rect -15752 16372 -15656 16408
rect -14340 16408 -14324 16472
rect -14260 16408 -14244 16472
rect -13921 17152 -13199 17161
rect -13921 16448 -13912 17152
rect -13208 16448 -13199 17152
rect -13921 16439 -13199 16448
rect -12928 17128 -12912 17192
rect -12848 17128 -12832 17192
rect -11516 17192 -11420 17228
rect -12928 17112 -12832 17128
rect -12928 17048 -12912 17112
rect -12848 17048 -12832 17112
rect -12928 17032 -12832 17048
rect -12928 16968 -12912 17032
rect -12848 16968 -12832 17032
rect -12928 16952 -12832 16968
rect -12928 16888 -12912 16952
rect -12848 16888 -12832 16952
rect -12928 16872 -12832 16888
rect -12928 16808 -12912 16872
rect -12848 16808 -12832 16872
rect -12928 16792 -12832 16808
rect -12928 16728 -12912 16792
rect -12848 16728 -12832 16792
rect -12928 16712 -12832 16728
rect -12928 16648 -12912 16712
rect -12848 16648 -12832 16712
rect -12928 16632 -12832 16648
rect -12928 16568 -12912 16632
rect -12848 16568 -12832 16632
rect -12928 16552 -12832 16568
rect -12928 16488 -12912 16552
rect -12848 16488 -12832 16552
rect -12928 16472 -12832 16488
rect -14340 16372 -14244 16408
rect -12928 16408 -12912 16472
rect -12848 16408 -12832 16472
rect -12509 17152 -11787 17161
rect -12509 16448 -12500 17152
rect -11796 16448 -11787 17152
rect -12509 16439 -11787 16448
rect -11516 17128 -11500 17192
rect -11436 17128 -11420 17192
rect -10104 17192 -10008 17228
rect -11516 17112 -11420 17128
rect -11516 17048 -11500 17112
rect -11436 17048 -11420 17112
rect -11516 17032 -11420 17048
rect -11516 16968 -11500 17032
rect -11436 16968 -11420 17032
rect -11516 16952 -11420 16968
rect -11516 16888 -11500 16952
rect -11436 16888 -11420 16952
rect -11516 16872 -11420 16888
rect -11516 16808 -11500 16872
rect -11436 16808 -11420 16872
rect -11516 16792 -11420 16808
rect -11516 16728 -11500 16792
rect -11436 16728 -11420 16792
rect -11516 16712 -11420 16728
rect -11516 16648 -11500 16712
rect -11436 16648 -11420 16712
rect -11516 16632 -11420 16648
rect -11516 16568 -11500 16632
rect -11436 16568 -11420 16632
rect -11516 16552 -11420 16568
rect -11516 16488 -11500 16552
rect -11436 16488 -11420 16552
rect -11516 16472 -11420 16488
rect -12928 16372 -12832 16408
rect -11516 16408 -11500 16472
rect -11436 16408 -11420 16472
rect -11097 17152 -10375 17161
rect -11097 16448 -11088 17152
rect -10384 16448 -10375 17152
rect -11097 16439 -10375 16448
rect -10104 17128 -10088 17192
rect -10024 17128 -10008 17192
rect -8692 17192 -8596 17228
rect -10104 17112 -10008 17128
rect -10104 17048 -10088 17112
rect -10024 17048 -10008 17112
rect -10104 17032 -10008 17048
rect -10104 16968 -10088 17032
rect -10024 16968 -10008 17032
rect -10104 16952 -10008 16968
rect -10104 16888 -10088 16952
rect -10024 16888 -10008 16952
rect -10104 16872 -10008 16888
rect -10104 16808 -10088 16872
rect -10024 16808 -10008 16872
rect -10104 16792 -10008 16808
rect -10104 16728 -10088 16792
rect -10024 16728 -10008 16792
rect -10104 16712 -10008 16728
rect -10104 16648 -10088 16712
rect -10024 16648 -10008 16712
rect -10104 16632 -10008 16648
rect -10104 16568 -10088 16632
rect -10024 16568 -10008 16632
rect -10104 16552 -10008 16568
rect -10104 16488 -10088 16552
rect -10024 16488 -10008 16552
rect -10104 16472 -10008 16488
rect -11516 16372 -11420 16408
rect -10104 16408 -10088 16472
rect -10024 16408 -10008 16472
rect -9685 17152 -8963 17161
rect -9685 16448 -9676 17152
rect -8972 16448 -8963 17152
rect -9685 16439 -8963 16448
rect -8692 17128 -8676 17192
rect -8612 17128 -8596 17192
rect -7280 17192 -7184 17228
rect -8692 17112 -8596 17128
rect -8692 17048 -8676 17112
rect -8612 17048 -8596 17112
rect -8692 17032 -8596 17048
rect -8692 16968 -8676 17032
rect -8612 16968 -8596 17032
rect -8692 16952 -8596 16968
rect -8692 16888 -8676 16952
rect -8612 16888 -8596 16952
rect -8692 16872 -8596 16888
rect -8692 16808 -8676 16872
rect -8612 16808 -8596 16872
rect -8692 16792 -8596 16808
rect -8692 16728 -8676 16792
rect -8612 16728 -8596 16792
rect -8692 16712 -8596 16728
rect -8692 16648 -8676 16712
rect -8612 16648 -8596 16712
rect -8692 16632 -8596 16648
rect -8692 16568 -8676 16632
rect -8612 16568 -8596 16632
rect -8692 16552 -8596 16568
rect -8692 16488 -8676 16552
rect -8612 16488 -8596 16552
rect -8692 16472 -8596 16488
rect -10104 16372 -10008 16408
rect -8692 16408 -8676 16472
rect -8612 16408 -8596 16472
rect -8273 17152 -7551 17161
rect -8273 16448 -8264 17152
rect -7560 16448 -7551 17152
rect -8273 16439 -7551 16448
rect -7280 17128 -7264 17192
rect -7200 17128 -7184 17192
rect -5868 17192 -5772 17228
rect -7280 17112 -7184 17128
rect -7280 17048 -7264 17112
rect -7200 17048 -7184 17112
rect -7280 17032 -7184 17048
rect -7280 16968 -7264 17032
rect -7200 16968 -7184 17032
rect -7280 16952 -7184 16968
rect -7280 16888 -7264 16952
rect -7200 16888 -7184 16952
rect -7280 16872 -7184 16888
rect -7280 16808 -7264 16872
rect -7200 16808 -7184 16872
rect -7280 16792 -7184 16808
rect -7280 16728 -7264 16792
rect -7200 16728 -7184 16792
rect -7280 16712 -7184 16728
rect -7280 16648 -7264 16712
rect -7200 16648 -7184 16712
rect -7280 16632 -7184 16648
rect -7280 16568 -7264 16632
rect -7200 16568 -7184 16632
rect -7280 16552 -7184 16568
rect -7280 16488 -7264 16552
rect -7200 16488 -7184 16552
rect -7280 16472 -7184 16488
rect -8692 16372 -8596 16408
rect -7280 16408 -7264 16472
rect -7200 16408 -7184 16472
rect -6861 17152 -6139 17161
rect -6861 16448 -6852 17152
rect -6148 16448 -6139 17152
rect -6861 16439 -6139 16448
rect -5868 17128 -5852 17192
rect -5788 17128 -5772 17192
rect -4456 17192 -4360 17228
rect -5868 17112 -5772 17128
rect -5868 17048 -5852 17112
rect -5788 17048 -5772 17112
rect -5868 17032 -5772 17048
rect -5868 16968 -5852 17032
rect -5788 16968 -5772 17032
rect -5868 16952 -5772 16968
rect -5868 16888 -5852 16952
rect -5788 16888 -5772 16952
rect -5868 16872 -5772 16888
rect -5868 16808 -5852 16872
rect -5788 16808 -5772 16872
rect -5868 16792 -5772 16808
rect -5868 16728 -5852 16792
rect -5788 16728 -5772 16792
rect -5868 16712 -5772 16728
rect -5868 16648 -5852 16712
rect -5788 16648 -5772 16712
rect -5868 16632 -5772 16648
rect -5868 16568 -5852 16632
rect -5788 16568 -5772 16632
rect -5868 16552 -5772 16568
rect -5868 16488 -5852 16552
rect -5788 16488 -5772 16552
rect -5868 16472 -5772 16488
rect -7280 16372 -7184 16408
rect -5868 16408 -5852 16472
rect -5788 16408 -5772 16472
rect -5449 17152 -4727 17161
rect -5449 16448 -5440 17152
rect -4736 16448 -4727 17152
rect -5449 16439 -4727 16448
rect -4456 17128 -4440 17192
rect -4376 17128 -4360 17192
rect -3044 17192 -2948 17228
rect -4456 17112 -4360 17128
rect -4456 17048 -4440 17112
rect -4376 17048 -4360 17112
rect -4456 17032 -4360 17048
rect -4456 16968 -4440 17032
rect -4376 16968 -4360 17032
rect -4456 16952 -4360 16968
rect -4456 16888 -4440 16952
rect -4376 16888 -4360 16952
rect -4456 16872 -4360 16888
rect -4456 16808 -4440 16872
rect -4376 16808 -4360 16872
rect -4456 16792 -4360 16808
rect -4456 16728 -4440 16792
rect -4376 16728 -4360 16792
rect -4456 16712 -4360 16728
rect -4456 16648 -4440 16712
rect -4376 16648 -4360 16712
rect -4456 16632 -4360 16648
rect -4456 16568 -4440 16632
rect -4376 16568 -4360 16632
rect -4456 16552 -4360 16568
rect -4456 16488 -4440 16552
rect -4376 16488 -4360 16552
rect -4456 16472 -4360 16488
rect -5868 16372 -5772 16408
rect -4456 16408 -4440 16472
rect -4376 16408 -4360 16472
rect -4037 17152 -3315 17161
rect -4037 16448 -4028 17152
rect -3324 16448 -3315 17152
rect -4037 16439 -3315 16448
rect -3044 17128 -3028 17192
rect -2964 17128 -2948 17192
rect -1632 17192 -1536 17228
rect -3044 17112 -2948 17128
rect -3044 17048 -3028 17112
rect -2964 17048 -2948 17112
rect -3044 17032 -2948 17048
rect -3044 16968 -3028 17032
rect -2964 16968 -2948 17032
rect -3044 16952 -2948 16968
rect -3044 16888 -3028 16952
rect -2964 16888 -2948 16952
rect -3044 16872 -2948 16888
rect -3044 16808 -3028 16872
rect -2964 16808 -2948 16872
rect -3044 16792 -2948 16808
rect -3044 16728 -3028 16792
rect -2964 16728 -2948 16792
rect -3044 16712 -2948 16728
rect -3044 16648 -3028 16712
rect -2964 16648 -2948 16712
rect -3044 16632 -2948 16648
rect -3044 16568 -3028 16632
rect -2964 16568 -2948 16632
rect -3044 16552 -2948 16568
rect -3044 16488 -3028 16552
rect -2964 16488 -2948 16552
rect -3044 16472 -2948 16488
rect -4456 16372 -4360 16408
rect -3044 16408 -3028 16472
rect -2964 16408 -2948 16472
rect -2625 17152 -1903 17161
rect -2625 16448 -2616 17152
rect -1912 16448 -1903 17152
rect -2625 16439 -1903 16448
rect -1632 17128 -1616 17192
rect -1552 17128 -1536 17192
rect -220 17192 -124 17228
rect -1632 17112 -1536 17128
rect -1632 17048 -1616 17112
rect -1552 17048 -1536 17112
rect -1632 17032 -1536 17048
rect -1632 16968 -1616 17032
rect -1552 16968 -1536 17032
rect -1632 16952 -1536 16968
rect -1632 16888 -1616 16952
rect -1552 16888 -1536 16952
rect -1632 16872 -1536 16888
rect -1632 16808 -1616 16872
rect -1552 16808 -1536 16872
rect -1632 16792 -1536 16808
rect -1632 16728 -1616 16792
rect -1552 16728 -1536 16792
rect -1632 16712 -1536 16728
rect -1632 16648 -1616 16712
rect -1552 16648 -1536 16712
rect -1632 16632 -1536 16648
rect -1632 16568 -1616 16632
rect -1552 16568 -1536 16632
rect -1632 16552 -1536 16568
rect -1632 16488 -1616 16552
rect -1552 16488 -1536 16552
rect -1632 16472 -1536 16488
rect -3044 16372 -2948 16408
rect -1632 16408 -1616 16472
rect -1552 16408 -1536 16472
rect -1213 17152 -491 17161
rect -1213 16448 -1204 17152
rect -500 16448 -491 17152
rect -1213 16439 -491 16448
rect -220 17128 -204 17192
rect -140 17128 -124 17192
rect 1192 17192 1288 17228
rect -220 17112 -124 17128
rect -220 17048 -204 17112
rect -140 17048 -124 17112
rect -220 17032 -124 17048
rect -220 16968 -204 17032
rect -140 16968 -124 17032
rect -220 16952 -124 16968
rect -220 16888 -204 16952
rect -140 16888 -124 16952
rect -220 16872 -124 16888
rect -220 16808 -204 16872
rect -140 16808 -124 16872
rect -220 16792 -124 16808
rect -220 16728 -204 16792
rect -140 16728 -124 16792
rect -220 16712 -124 16728
rect -220 16648 -204 16712
rect -140 16648 -124 16712
rect -220 16632 -124 16648
rect -220 16568 -204 16632
rect -140 16568 -124 16632
rect -220 16552 -124 16568
rect -220 16488 -204 16552
rect -140 16488 -124 16552
rect -220 16472 -124 16488
rect -1632 16372 -1536 16408
rect -220 16408 -204 16472
rect -140 16408 -124 16472
rect 199 17152 921 17161
rect 199 16448 208 17152
rect 912 16448 921 17152
rect 199 16439 921 16448
rect 1192 17128 1208 17192
rect 1272 17128 1288 17192
rect 2604 17192 2700 17228
rect 1192 17112 1288 17128
rect 1192 17048 1208 17112
rect 1272 17048 1288 17112
rect 1192 17032 1288 17048
rect 1192 16968 1208 17032
rect 1272 16968 1288 17032
rect 1192 16952 1288 16968
rect 1192 16888 1208 16952
rect 1272 16888 1288 16952
rect 1192 16872 1288 16888
rect 1192 16808 1208 16872
rect 1272 16808 1288 16872
rect 1192 16792 1288 16808
rect 1192 16728 1208 16792
rect 1272 16728 1288 16792
rect 1192 16712 1288 16728
rect 1192 16648 1208 16712
rect 1272 16648 1288 16712
rect 1192 16632 1288 16648
rect 1192 16568 1208 16632
rect 1272 16568 1288 16632
rect 1192 16552 1288 16568
rect 1192 16488 1208 16552
rect 1272 16488 1288 16552
rect 1192 16472 1288 16488
rect -220 16372 -124 16408
rect 1192 16408 1208 16472
rect 1272 16408 1288 16472
rect 1611 17152 2333 17161
rect 1611 16448 1620 17152
rect 2324 16448 2333 17152
rect 1611 16439 2333 16448
rect 2604 17128 2620 17192
rect 2684 17128 2700 17192
rect 4016 17192 4112 17228
rect 2604 17112 2700 17128
rect 2604 17048 2620 17112
rect 2684 17048 2700 17112
rect 2604 17032 2700 17048
rect 2604 16968 2620 17032
rect 2684 16968 2700 17032
rect 2604 16952 2700 16968
rect 2604 16888 2620 16952
rect 2684 16888 2700 16952
rect 2604 16872 2700 16888
rect 2604 16808 2620 16872
rect 2684 16808 2700 16872
rect 2604 16792 2700 16808
rect 2604 16728 2620 16792
rect 2684 16728 2700 16792
rect 2604 16712 2700 16728
rect 2604 16648 2620 16712
rect 2684 16648 2700 16712
rect 2604 16632 2700 16648
rect 2604 16568 2620 16632
rect 2684 16568 2700 16632
rect 2604 16552 2700 16568
rect 2604 16488 2620 16552
rect 2684 16488 2700 16552
rect 2604 16472 2700 16488
rect 1192 16372 1288 16408
rect 2604 16408 2620 16472
rect 2684 16408 2700 16472
rect 3023 17152 3745 17161
rect 3023 16448 3032 17152
rect 3736 16448 3745 17152
rect 3023 16439 3745 16448
rect 4016 17128 4032 17192
rect 4096 17128 4112 17192
rect 5428 17192 5524 17228
rect 4016 17112 4112 17128
rect 4016 17048 4032 17112
rect 4096 17048 4112 17112
rect 4016 17032 4112 17048
rect 4016 16968 4032 17032
rect 4096 16968 4112 17032
rect 4016 16952 4112 16968
rect 4016 16888 4032 16952
rect 4096 16888 4112 16952
rect 4016 16872 4112 16888
rect 4016 16808 4032 16872
rect 4096 16808 4112 16872
rect 4016 16792 4112 16808
rect 4016 16728 4032 16792
rect 4096 16728 4112 16792
rect 4016 16712 4112 16728
rect 4016 16648 4032 16712
rect 4096 16648 4112 16712
rect 4016 16632 4112 16648
rect 4016 16568 4032 16632
rect 4096 16568 4112 16632
rect 4016 16552 4112 16568
rect 4016 16488 4032 16552
rect 4096 16488 4112 16552
rect 4016 16472 4112 16488
rect 2604 16372 2700 16408
rect 4016 16408 4032 16472
rect 4096 16408 4112 16472
rect 4435 17152 5157 17161
rect 4435 16448 4444 17152
rect 5148 16448 5157 17152
rect 4435 16439 5157 16448
rect 5428 17128 5444 17192
rect 5508 17128 5524 17192
rect 6840 17192 6936 17228
rect 5428 17112 5524 17128
rect 5428 17048 5444 17112
rect 5508 17048 5524 17112
rect 5428 17032 5524 17048
rect 5428 16968 5444 17032
rect 5508 16968 5524 17032
rect 5428 16952 5524 16968
rect 5428 16888 5444 16952
rect 5508 16888 5524 16952
rect 5428 16872 5524 16888
rect 5428 16808 5444 16872
rect 5508 16808 5524 16872
rect 5428 16792 5524 16808
rect 5428 16728 5444 16792
rect 5508 16728 5524 16792
rect 5428 16712 5524 16728
rect 5428 16648 5444 16712
rect 5508 16648 5524 16712
rect 5428 16632 5524 16648
rect 5428 16568 5444 16632
rect 5508 16568 5524 16632
rect 5428 16552 5524 16568
rect 5428 16488 5444 16552
rect 5508 16488 5524 16552
rect 5428 16472 5524 16488
rect 4016 16372 4112 16408
rect 5428 16408 5444 16472
rect 5508 16408 5524 16472
rect 5847 17152 6569 17161
rect 5847 16448 5856 17152
rect 6560 16448 6569 17152
rect 5847 16439 6569 16448
rect 6840 17128 6856 17192
rect 6920 17128 6936 17192
rect 8252 17192 8348 17228
rect 6840 17112 6936 17128
rect 6840 17048 6856 17112
rect 6920 17048 6936 17112
rect 6840 17032 6936 17048
rect 6840 16968 6856 17032
rect 6920 16968 6936 17032
rect 6840 16952 6936 16968
rect 6840 16888 6856 16952
rect 6920 16888 6936 16952
rect 6840 16872 6936 16888
rect 6840 16808 6856 16872
rect 6920 16808 6936 16872
rect 6840 16792 6936 16808
rect 6840 16728 6856 16792
rect 6920 16728 6936 16792
rect 6840 16712 6936 16728
rect 6840 16648 6856 16712
rect 6920 16648 6936 16712
rect 6840 16632 6936 16648
rect 6840 16568 6856 16632
rect 6920 16568 6936 16632
rect 6840 16552 6936 16568
rect 6840 16488 6856 16552
rect 6920 16488 6936 16552
rect 6840 16472 6936 16488
rect 5428 16372 5524 16408
rect 6840 16408 6856 16472
rect 6920 16408 6936 16472
rect 7259 17152 7981 17161
rect 7259 16448 7268 17152
rect 7972 16448 7981 17152
rect 7259 16439 7981 16448
rect 8252 17128 8268 17192
rect 8332 17128 8348 17192
rect 9664 17192 9760 17228
rect 8252 17112 8348 17128
rect 8252 17048 8268 17112
rect 8332 17048 8348 17112
rect 8252 17032 8348 17048
rect 8252 16968 8268 17032
rect 8332 16968 8348 17032
rect 8252 16952 8348 16968
rect 8252 16888 8268 16952
rect 8332 16888 8348 16952
rect 8252 16872 8348 16888
rect 8252 16808 8268 16872
rect 8332 16808 8348 16872
rect 8252 16792 8348 16808
rect 8252 16728 8268 16792
rect 8332 16728 8348 16792
rect 8252 16712 8348 16728
rect 8252 16648 8268 16712
rect 8332 16648 8348 16712
rect 8252 16632 8348 16648
rect 8252 16568 8268 16632
rect 8332 16568 8348 16632
rect 8252 16552 8348 16568
rect 8252 16488 8268 16552
rect 8332 16488 8348 16552
rect 8252 16472 8348 16488
rect 6840 16372 6936 16408
rect 8252 16408 8268 16472
rect 8332 16408 8348 16472
rect 8671 17152 9393 17161
rect 8671 16448 8680 17152
rect 9384 16448 9393 17152
rect 8671 16439 9393 16448
rect 9664 17128 9680 17192
rect 9744 17128 9760 17192
rect 11076 17192 11172 17228
rect 9664 17112 9760 17128
rect 9664 17048 9680 17112
rect 9744 17048 9760 17112
rect 9664 17032 9760 17048
rect 9664 16968 9680 17032
rect 9744 16968 9760 17032
rect 9664 16952 9760 16968
rect 9664 16888 9680 16952
rect 9744 16888 9760 16952
rect 9664 16872 9760 16888
rect 9664 16808 9680 16872
rect 9744 16808 9760 16872
rect 9664 16792 9760 16808
rect 9664 16728 9680 16792
rect 9744 16728 9760 16792
rect 9664 16712 9760 16728
rect 9664 16648 9680 16712
rect 9744 16648 9760 16712
rect 9664 16632 9760 16648
rect 9664 16568 9680 16632
rect 9744 16568 9760 16632
rect 9664 16552 9760 16568
rect 9664 16488 9680 16552
rect 9744 16488 9760 16552
rect 9664 16472 9760 16488
rect 8252 16372 8348 16408
rect 9664 16408 9680 16472
rect 9744 16408 9760 16472
rect 10083 17152 10805 17161
rect 10083 16448 10092 17152
rect 10796 16448 10805 17152
rect 10083 16439 10805 16448
rect 11076 17128 11092 17192
rect 11156 17128 11172 17192
rect 12488 17192 12584 17228
rect 11076 17112 11172 17128
rect 11076 17048 11092 17112
rect 11156 17048 11172 17112
rect 11076 17032 11172 17048
rect 11076 16968 11092 17032
rect 11156 16968 11172 17032
rect 11076 16952 11172 16968
rect 11076 16888 11092 16952
rect 11156 16888 11172 16952
rect 11076 16872 11172 16888
rect 11076 16808 11092 16872
rect 11156 16808 11172 16872
rect 11076 16792 11172 16808
rect 11076 16728 11092 16792
rect 11156 16728 11172 16792
rect 11076 16712 11172 16728
rect 11076 16648 11092 16712
rect 11156 16648 11172 16712
rect 11076 16632 11172 16648
rect 11076 16568 11092 16632
rect 11156 16568 11172 16632
rect 11076 16552 11172 16568
rect 11076 16488 11092 16552
rect 11156 16488 11172 16552
rect 11076 16472 11172 16488
rect 9664 16372 9760 16408
rect 11076 16408 11092 16472
rect 11156 16408 11172 16472
rect 11495 17152 12217 17161
rect 11495 16448 11504 17152
rect 12208 16448 12217 17152
rect 11495 16439 12217 16448
rect 12488 17128 12504 17192
rect 12568 17128 12584 17192
rect 13900 17192 13996 17228
rect 12488 17112 12584 17128
rect 12488 17048 12504 17112
rect 12568 17048 12584 17112
rect 12488 17032 12584 17048
rect 12488 16968 12504 17032
rect 12568 16968 12584 17032
rect 12488 16952 12584 16968
rect 12488 16888 12504 16952
rect 12568 16888 12584 16952
rect 12488 16872 12584 16888
rect 12488 16808 12504 16872
rect 12568 16808 12584 16872
rect 12488 16792 12584 16808
rect 12488 16728 12504 16792
rect 12568 16728 12584 16792
rect 12488 16712 12584 16728
rect 12488 16648 12504 16712
rect 12568 16648 12584 16712
rect 12488 16632 12584 16648
rect 12488 16568 12504 16632
rect 12568 16568 12584 16632
rect 12488 16552 12584 16568
rect 12488 16488 12504 16552
rect 12568 16488 12584 16552
rect 12488 16472 12584 16488
rect 11076 16372 11172 16408
rect 12488 16408 12504 16472
rect 12568 16408 12584 16472
rect 12907 17152 13629 17161
rect 12907 16448 12916 17152
rect 13620 16448 13629 17152
rect 12907 16439 13629 16448
rect 13900 17128 13916 17192
rect 13980 17128 13996 17192
rect 15312 17192 15408 17228
rect 13900 17112 13996 17128
rect 13900 17048 13916 17112
rect 13980 17048 13996 17112
rect 13900 17032 13996 17048
rect 13900 16968 13916 17032
rect 13980 16968 13996 17032
rect 13900 16952 13996 16968
rect 13900 16888 13916 16952
rect 13980 16888 13996 16952
rect 13900 16872 13996 16888
rect 13900 16808 13916 16872
rect 13980 16808 13996 16872
rect 13900 16792 13996 16808
rect 13900 16728 13916 16792
rect 13980 16728 13996 16792
rect 13900 16712 13996 16728
rect 13900 16648 13916 16712
rect 13980 16648 13996 16712
rect 13900 16632 13996 16648
rect 13900 16568 13916 16632
rect 13980 16568 13996 16632
rect 13900 16552 13996 16568
rect 13900 16488 13916 16552
rect 13980 16488 13996 16552
rect 13900 16472 13996 16488
rect 12488 16372 12584 16408
rect 13900 16408 13916 16472
rect 13980 16408 13996 16472
rect 14319 17152 15041 17161
rect 14319 16448 14328 17152
rect 15032 16448 15041 17152
rect 14319 16439 15041 16448
rect 15312 17128 15328 17192
rect 15392 17128 15408 17192
rect 16724 17192 16820 17228
rect 15312 17112 15408 17128
rect 15312 17048 15328 17112
rect 15392 17048 15408 17112
rect 15312 17032 15408 17048
rect 15312 16968 15328 17032
rect 15392 16968 15408 17032
rect 15312 16952 15408 16968
rect 15312 16888 15328 16952
rect 15392 16888 15408 16952
rect 15312 16872 15408 16888
rect 15312 16808 15328 16872
rect 15392 16808 15408 16872
rect 15312 16792 15408 16808
rect 15312 16728 15328 16792
rect 15392 16728 15408 16792
rect 15312 16712 15408 16728
rect 15312 16648 15328 16712
rect 15392 16648 15408 16712
rect 15312 16632 15408 16648
rect 15312 16568 15328 16632
rect 15392 16568 15408 16632
rect 15312 16552 15408 16568
rect 15312 16488 15328 16552
rect 15392 16488 15408 16552
rect 15312 16472 15408 16488
rect 13900 16372 13996 16408
rect 15312 16408 15328 16472
rect 15392 16408 15408 16472
rect 15731 17152 16453 17161
rect 15731 16448 15740 17152
rect 16444 16448 16453 17152
rect 15731 16439 16453 16448
rect 16724 17128 16740 17192
rect 16804 17128 16820 17192
rect 18136 17192 18232 17228
rect 16724 17112 16820 17128
rect 16724 17048 16740 17112
rect 16804 17048 16820 17112
rect 16724 17032 16820 17048
rect 16724 16968 16740 17032
rect 16804 16968 16820 17032
rect 16724 16952 16820 16968
rect 16724 16888 16740 16952
rect 16804 16888 16820 16952
rect 16724 16872 16820 16888
rect 16724 16808 16740 16872
rect 16804 16808 16820 16872
rect 16724 16792 16820 16808
rect 16724 16728 16740 16792
rect 16804 16728 16820 16792
rect 16724 16712 16820 16728
rect 16724 16648 16740 16712
rect 16804 16648 16820 16712
rect 16724 16632 16820 16648
rect 16724 16568 16740 16632
rect 16804 16568 16820 16632
rect 16724 16552 16820 16568
rect 16724 16488 16740 16552
rect 16804 16488 16820 16552
rect 16724 16472 16820 16488
rect 15312 16372 15408 16408
rect 16724 16408 16740 16472
rect 16804 16408 16820 16472
rect 17143 17152 17865 17161
rect 17143 16448 17152 17152
rect 17856 16448 17865 17152
rect 17143 16439 17865 16448
rect 18136 17128 18152 17192
rect 18216 17128 18232 17192
rect 19548 17192 19644 17228
rect 18136 17112 18232 17128
rect 18136 17048 18152 17112
rect 18216 17048 18232 17112
rect 18136 17032 18232 17048
rect 18136 16968 18152 17032
rect 18216 16968 18232 17032
rect 18136 16952 18232 16968
rect 18136 16888 18152 16952
rect 18216 16888 18232 16952
rect 18136 16872 18232 16888
rect 18136 16808 18152 16872
rect 18216 16808 18232 16872
rect 18136 16792 18232 16808
rect 18136 16728 18152 16792
rect 18216 16728 18232 16792
rect 18136 16712 18232 16728
rect 18136 16648 18152 16712
rect 18216 16648 18232 16712
rect 18136 16632 18232 16648
rect 18136 16568 18152 16632
rect 18216 16568 18232 16632
rect 18136 16552 18232 16568
rect 18136 16488 18152 16552
rect 18216 16488 18232 16552
rect 18136 16472 18232 16488
rect 16724 16372 16820 16408
rect 18136 16408 18152 16472
rect 18216 16408 18232 16472
rect 18555 17152 19277 17161
rect 18555 16448 18564 17152
rect 19268 16448 19277 17152
rect 18555 16439 19277 16448
rect 19548 17128 19564 17192
rect 19628 17128 19644 17192
rect 20960 17192 21056 17228
rect 19548 17112 19644 17128
rect 19548 17048 19564 17112
rect 19628 17048 19644 17112
rect 19548 17032 19644 17048
rect 19548 16968 19564 17032
rect 19628 16968 19644 17032
rect 19548 16952 19644 16968
rect 19548 16888 19564 16952
rect 19628 16888 19644 16952
rect 19548 16872 19644 16888
rect 19548 16808 19564 16872
rect 19628 16808 19644 16872
rect 19548 16792 19644 16808
rect 19548 16728 19564 16792
rect 19628 16728 19644 16792
rect 19548 16712 19644 16728
rect 19548 16648 19564 16712
rect 19628 16648 19644 16712
rect 19548 16632 19644 16648
rect 19548 16568 19564 16632
rect 19628 16568 19644 16632
rect 19548 16552 19644 16568
rect 19548 16488 19564 16552
rect 19628 16488 19644 16552
rect 19548 16472 19644 16488
rect 18136 16372 18232 16408
rect 19548 16408 19564 16472
rect 19628 16408 19644 16472
rect 19967 17152 20689 17161
rect 19967 16448 19976 17152
rect 20680 16448 20689 17152
rect 19967 16439 20689 16448
rect 20960 17128 20976 17192
rect 21040 17128 21056 17192
rect 22372 17192 22468 17228
rect 20960 17112 21056 17128
rect 20960 17048 20976 17112
rect 21040 17048 21056 17112
rect 20960 17032 21056 17048
rect 20960 16968 20976 17032
rect 21040 16968 21056 17032
rect 20960 16952 21056 16968
rect 20960 16888 20976 16952
rect 21040 16888 21056 16952
rect 20960 16872 21056 16888
rect 20960 16808 20976 16872
rect 21040 16808 21056 16872
rect 20960 16792 21056 16808
rect 20960 16728 20976 16792
rect 21040 16728 21056 16792
rect 20960 16712 21056 16728
rect 20960 16648 20976 16712
rect 21040 16648 21056 16712
rect 20960 16632 21056 16648
rect 20960 16568 20976 16632
rect 21040 16568 21056 16632
rect 20960 16552 21056 16568
rect 20960 16488 20976 16552
rect 21040 16488 21056 16552
rect 20960 16472 21056 16488
rect 19548 16372 19644 16408
rect 20960 16408 20976 16472
rect 21040 16408 21056 16472
rect 21379 17152 22101 17161
rect 21379 16448 21388 17152
rect 22092 16448 22101 17152
rect 21379 16439 22101 16448
rect 22372 17128 22388 17192
rect 22452 17128 22468 17192
rect 23784 17192 23880 17228
rect 22372 17112 22468 17128
rect 22372 17048 22388 17112
rect 22452 17048 22468 17112
rect 22372 17032 22468 17048
rect 22372 16968 22388 17032
rect 22452 16968 22468 17032
rect 22372 16952 22468 16968
rect 22372 16888 22388 16952
rect 22452 16888 22468 16952
rect 22372 16872 22468 16888
rect 22372 16808 22388 16872
rect 22452 16808 22468 16872
rect 22372 16792 22468 16808
rect 22372 16728 22388 16792
rect 22452 16728 22468 16792
rect 22372 16712 22468 16728
rect 22372 16648 22388 16712
rect 22452 16648 22468 16712
rect 22372 16632 22468 16648
rect 22372 16568 22388 16632
rect 22452 16568 22468 16632
rect 22372 16552 22468 16568
rect 22372 16488 22388 16552
rect 22452 16488 22468 16552
rect 22372 16472 22468 16488
rect 20960 16372 21056 16408
rect 22372 16408 22388 16472
rect 22452 16408 22468 16472
rect 22791 17152 23513 17161
rect 22791 16448 22800 17152
rect 23504 16448 23513 17152
rect 22791 16439 23513 16448
rect 23784 17128 23800 17192
rect 23864 17128 23880 17192
rect 23784 17112 23880 17128
rect 23784 17048 23800 17112
rect 23864 17048 23880 17112
rect 23784 17032 23880 17048
rect 23784 16968 23800 17032
rect 23864 16968 23880 17032
rect 23784 16952 23880 16968
rect 23784 16888 23800 16952
rect 23864 16888 23880 16952
rect 23784 16872 23880 16888
rect 23784 16808 23800 16872
rect 23864 16808 23880 16872
rect 23784 16792 23880 16808
rect 23784 16728 23800 16792
rect 23864 16728 23880 16792
rect 23784 16712 23880 16728
rect 23784 16648 23800 16712
rect 23864 16648 23880 16712
rect 23784 16632 23880 16648
rect 23784 16568 23800 16632
rect 23864 16568 23880 16632
rect 23784 16552 23880 16568
rect 23784 16488 23800 16552
rect 23864 16488 23880 16552
rect 23784 16472 23880 16488
rect 22372 16372 22468 16408
rect 23784 16408 23800 16472
rect 23864 16408 23880 16472
rect 23784 16372 23880 16408
rect -22812 16072 -22716 16108
rect -23805 16032 -23083 16041
rect -23805 15328 -23796 16032
rect -23092 15328 -23083 16032
rect -23805 15319 -23083 15328
rect -22812 16008 -22796 16072
rect -22732 16008 -22716 16072
rect -21400 16072 -21304 16108
rect -22812 15992 -22716 16008
rect -22812 15928 -22796 15992
rect -22732 15928 -22716 15992
rect -22812 15912 -22716 15928
rect -22812 15848 -22796 15912
rect -22732 15848 -22716 15912
rect -22812 15832 -22716 15848
rect -22812 15768 -22796 15832
rect -22732 15768 -22716 15832
rect -22812 15752 -22716 15768
rect -22812 15688 -22796 15752
rect -22732 15688 -22716 15752
rect -22812 15672 -22716 15688
rect -22812 15608 -22796 15672
rect -22732 15608 -22716 15672
rect -22812 15592 -22716 15608
rect -22812 15528 -22796 15592
rect -22732 15528 -22716 15592
rect -22812 15512 -22716 15528
rect -22812 15448 -22796 15512
rect -22732 15448 -22716 15512
rect -22812 15432 -22716 15448
rect -22812 15368 -22796 15432
rect -22732 15368 -22716 15432
rect -22812 15352 -22716 15368
rect -22812 15288 -22796 15352
rect -22732 15288 -22716 15352
rect -22393 16032 -21671 16041
rect -22393 15328 -22384 16032
rect -21680 15328 -21671 16032
rect -22393 15319 -21671 15328
rect -21400 16008 -21384 16072
rect -21320 16008 -21304 16072
rect -19988 16072 -19892 16108
rect -21400 15992 -21304 16008
rect -21400 15928 -21384 15992
rect -21320 15928 -21304 15992
rect -21400 15912 -21304 15928
rect -21400 15848 -21384 15912
rect -21320 15848 -21304 15912
rect -21400 15832 -21304 15848
rect -21400 15768 -21384 15832
rect -21320 15768 -21304 15832
rect -21400 15752 -21304 15768
rect -21400 15688 -21384 15752
rect -21320 15688 -21304 15752
rect -21400 15672 -21304 15688
rect -21400 15608 -21384 15672
rect -21320 15608 -21304 15672
rect -21400 15592 -21304 15608
rect -21400 15528 -21384 15592
rect -21320 15528 -21304 15592
rect -21400 15512 -21304 15528
rect -21400 15448 -21384 15512
rect -21320 15448 -21304 15512
rect -21400 15432 -21304 15448
rect -21400 15368 -21384 15432
rect -21320 15368 -21304 15432
rect -21400 15352 -21304 15368
rect -22812 15252 -22716 15288
rect -21400 15288 -21384 15352
rect -21320 15288 -21304 15352
rect -20981 16032 -20259 16041
rect -20981 15328 -20972 16032
rect -20268 15328 -20259 16032
rect -20981 15319 -20259 15328
rect -19988 16008 -19972 16072
rect -19908 16008 -19892 16072
rect -18576 16072 -18480 16108
rect -19988 15992 -19892 16008
rect -19988 15928 -19972 15992
rect -19908 15928 -19892 15992
rect -19988 15912 -19892 15928
rect -19988 15848 -19972 15912
rect -19908 15848 -19892 15912
rect -19988 15832 -19892 15848
rect -19988 15768 -19972 15832
rect -19908 15768 -19892 15832
rect -19988 15752 -19892 15768
rect -19988 15688 -19972 15752
rect -19908 15688 -19892 15752
rect -19988 15672 -19892 15688
rect -19988 15608 -19972 15672
rect -19908 15608 -19892 15672
rect -19988 15592 -19892 15608
rect -19988 15528 -19972 15592
rect -19908 15528 -19892 15592
rect -19988 15512 -19892 15528
rect -19988 15448 -19972 15512
rect -19908 15448 -19892 15512
rect -19988 15432 -19892 15448
rect -19988 15368 -19972 15432
rect -19908 15368 -19892 15432
rect -19988 15352 -19892 15368
rect -21400 15252 -21304 15288
rect -19988 15288 -19972 15352
rect -19908 15288 -19892 15352
rect -19569 16032 -18847 16041
rect -19569 15328 -19560 16032
rect -18856 15328 -18847 16032
rect -19569 15319 -18847 15328
rect -18576 16008 -18560 16072
rect -18496 16008 -18480 16072
rect -17164 16072 -17068 16108
rect -18576 15992 -18480 16008
rect -18576 15928 -18560 15992
rect -18496 15928 -18480 15992
rect -18576 15912 -18480 15928
rect -18576 15848 -18560 15912
rect -18496 15848 -18480 15912
rect -18576 15832 -18480 15848
rect -18576 15768 -18560 15832
rect -18496 15768 -18480 15832
rect -18576 15752 -18480 15768
rect -18576 15688 -18560 15752
rect -18496 15688 -18480 15752
rect -18576 15672 -18480 15688
rect -18576 15608 -18560 15672
rect -18496 15608 -18480 15672
rect -18576 15592 -18480 15608
rect -18576 15528 -18560 15592
rect -18496 15528 -18480 15592
rect -18576 15512 -18480 15528
rect -18576 15448 -18560 15512
rect -18496 15448 -18480 15512
rect -18576 15432 -18480 15448
rect -18576 15368 -18560 15432
rect -18496 15368 -18480 15432
rect -18576 15352 -18480 15368
rect -19988 15252 -19892 15288
rect -18576 15288 -18560 15352
rect -18496 15288 -18480 15352
rect -18157 16032 -17435 16041
rect -18157 15328 -18148 16032
rect -17444 15328 -17435 16032
rect -18157 15319 -17435 15328
rect -17164 16008 -17148 16072
rect -17084 16008 -17068 16072
rect -15752 16072 -15656 16108
rect -17164 15992 -17068 16008
rect -17164 15928 -17148 15992
rect -17084 15928 -17068 15992
rect -17164 15912 -17068 15928
rect -17164 15848 -17148 15912
rect -17084 15848 -17068 15912
rect -17164 15832 -17068 15848
rect -17164 15768 -17148 15832
rect -17084 15768 -17068 15832
rect -17164 15752 -17068 15768
rect -17164 15688 -17148 15752
rect -17084 15688 -17068 15752
rect -17164 15672 -17068 15688
rect -17164 15608 -17148 15672
rect -17084 15608 -17068 15672
rect -17164 15592 -17068 15608
rect -17164 15528 -17148 15592
rect -17084 15528 -17068 15592
rect -17164 15512 -17068 15528
rect -17164 15448 -17148 15512
rect -17084 15448 -17068 15512
rect -17164 15432 -17068 15448
rect -17164 15368 -17148 15432
rect -17084 15368 -17068 15432
rect -17164 15352 -17068 15368
rect -18576 15252 -18480 15288
rect -17164 15288 -17148 15352
rect -17084 15288 -17068 15352
rect -16745 16032 -16023 16041
rect -16745 15328 -16736 16032
rect -16032 15328 -16023 16032
rect -16745 15319 -16023 15328
rect -15752 16008 -15736 16072
rect -15672 16008 -15656 16072
rect -14340 16072 -14244 16108
rect -15752 15992 -15656 16008
rect -15752 15928 -15736 15992
rect -15672 15928 -15656 15992
rect -15752 15912 -15656 15928
rect -15752 15848 -15736 15912
rect -15672 15848 -15656 15912
rect -15752 15832 -15656 15848
rect -15752 15768 -15736 15832
rect -15672 15768 -15656 15832
rect -15752 15752 -15656 15768
rect -15752 15688 -15736 15752
rect -15672 15688 -15656 15752
rect -15752 15672 -15656 15688
rect -15752 15608 -15736 15672
rect -15672 15608 -15656 15672
rect -15752 15592 -15656 15608
rect -15752 15528 -15736 15592
rect -15672 15528 -15656 15592
rect -15752 15512 -15656 15528
rect -15752 15448 -15736 15512
rect -15672 15448 -15656 15512
rect -15752 15432 -15656 15448
rect -15752 15368 -15736 15432
rect -15672 15368 -15656 15432
rect -15752 15352 -15656 15368
rect -17164 15252 -17068 15288
rect -15752 15288 -15736 15352
rect -15672 15288 -15656 15352
rect -15333 16032 -14611 16041
rect -15333 15328 -15324 16032
rect -14620 15328 -14611 16032
rect -15333 15319 -14611 15328
rect -14340 16008 -14324 16072
rect -14260 16008 -14244 16072
rect -12928 16072 -12832 16108
rect -14340 15992 -14244 16008
rect -14340 15928 -14324 15992
rect -14260 15928 -14244 15992
rect -14340 15912 -14244 15928
rect -14340 15848 -14324 15912
rect -14260 15848 -14244 15912
rect -14340 15832 -14244 15848
rect -14340 15768 -14324 15832
rect -14260 15768 -14244 15832
rect -14340 15752 -14244 15768
rect -14340 15688 -14324 15752
rect -14260 15688 -14244 15752
rect -14340 15672 -14244 15688
rect -14340 15608 -14324 15672
rect -14260 15608 -14244 15672
rect -14340 15592 -14244 15608
rect -14340 15528 -14324 15592
rect -14260 15528 -14244 15592
rect -14340 15512 -14244 15528
rect -14340 15448 -14324 15512
rect -14260 15448 -14244 15512
rect -14340 15432 -14244 15448
rect -14340 15368 -14324 15432
rect -14260 15368 -14244 15432
rect -14340 15352 -14244 15368
rect -15752 15252 -15656 15288
rect -14340 15288 -14324 15352
rect -14260 15288 -14244 15352
rect -13921 16032 -13199 16041
rect -13921 15328 -13912 16032
rect -13208 15328 -13199 16032
rect -13921 15319 -13199 15328
rect -12928 16008 -12912 16072
rect -12848 16008 -12832 16072
rect -11516 16072 -11420 16108
rect -12928 15992 -12832 16008
rect -12928 15928 -12912 15992
rect -12848 15928 -12832 15992
rect -12928 15912 -12832 15928
rect -12928 15848 -12912 15912
rect -12848 15848 -12832 15912
rect -12928 15832 -12832 15848
rect -12928 15768 -12912 15832
rect -12848 15768 -12832 15832
rect -12928 15752 -12832 15768
rect -12928 15688 -12912 15752
rect -12848 15688 -12832 15752
rect -12928 15672 -12832 15688
rect -12928 15608 -12912 15672
rect -12848 15608 -12832 15672
rect -12928 15592 -12832 15608
rect -12928 15528 -12912 15592
rect -12848 15528 -12832 15592
rect -12928 15512 -12832 15528
rect -12928 15448 -12912 15512
rect -12848 15448 -12832 15512
rect -12928 15432 -12832 15448
rect -12928 15368 -12912 15432
rect -12848 15368 -12832 15432
rect -12928 15352 -12832 15368
rect -14340 15252 -14244 15288
rect -12928 15288 -12912 15352
rect -12848 15288 -12832 15352
rect -12509 16032 -11787 16041
rect -12509 15328 -12500 16032
rect -11796 15328 -11787 16032
rect -12509 15319 -11787 15328
rect -11516 16008 -11500 16072
rect -11436 16008 -11420 16072
rect -10104 16072 -10008 16108
rect -11516 15992 -11420 16008
rect -11516 15928 -11500 15992
rect -11436 15928 -11420 15992
rect -11516 15912 -11420 15928
rect -11516 15848 -11500 15912
rect -11436 15848 -11420 15912
rect -11516 15832 -11420 15848
rect -11516 15768 -11500 15832
rect -11436 15768 -11420 15832
rect -11516 15752 -11420 15768
rect -11516 15688 -11500 15752
rect -11436 15688 -11420 15752
rect -11516 15672 -11420 15688
rect -11516 15608 -11500 15672
rect -11436 15608 -11420 15672
rect -11516 15592 -11420 15608
rect -11516 15528 -11500 15592
rect -11436 15528 -11420 15592
rect -11516 15512 -11420 15528
rect -11516 15448 -11500 15512
rect -11436 15448 -11420 15512
rect -11516 15432 -11420 15448
rect -11516 15368 -11500 15432
rect -11436 15368 -11420 15432
rect -11516 15352 -11420 15368
rect -12928 15252 -12832 15288
rect -11516 15288 -11500 15352
rect -11436 15288 -11420 15352
rect -11097 16032 -10375 16041
rect -11097 15328 -11088 16032
rect -10384 15328 -10375 16032
rect -11097 15319 -10375 15328
rect -10104 16008 -10088 16072
rect -10024 16008 -10008 16072
rect -8692 16072 -8596 16108
rect -10104 15992 -10008 16008
rect -10104 15928 -10088 15992
rect -10024 15928 -10008 15992
rect -10104 15912 -10008 15928
rect -10104 15848 -10088 15912
rect -10024 15848 -10008 15912
rect -10104 15832 -10008 15848
rect -10104 15768 -10088 15832
rect -10024 15768 -10008 15832
rect -10104 15752 -10008 15768
rect -10104 15688 -10088 15752
rect -10024 15688 -10008 15752
rect -10104 15672 -10008 15688
rect -10104 15608 -10088 15672
rect -10024 15608 -10008 15672
rect -10104 15592 -10008 15608
rect -10104 15528 -10088 15592
rect -10024 15528 -10008 15592
rect -10104 15512 -10008 15528
rect -10104 15448 -10088 15512
rect -10024 15448 -10008 15512
rect -10104 15432 -10008 15448
rect -10104 15368 -10088 15432
rect -10024 15368 -10008 15432
rect -10104 15352 -10008 15368
rect -11516 15252 -11420 15288
rect -10104 15288 -10088 15352
rect -10024 15288 -10008 15352
rect -9685 16032 -8963 16041
rect -9685 15328 -9676 16032
rect -8972 15328 -8963 16032
rect -9685 15319 -8963 15328
rect -8692 16008 -8676 16072
rect -8612 16008 -8596 16072
rect -7280 16072 -7184 16108
rect -8692 15992 -8596 16008
rect -8692 15928 -8676 15992
rect -8612 15928 -8596 15992
rect -8692 15912 -8596 15928
rect -8692 15848 -8676 15912
rect -8612 15848 -8596 15912
rect -8692 15832 -8596 15848
rect -8692 15768 -8676 15832
rect -8612 15768 -8596 15832
rect -8692 15752 -8596 15768
rect -8692 15688 -8676 15752
rect -8612 15688 -8596 15752
rect -8692 15672 -8596 15688
rect -8692 15608 -8676 15672
rect -8612 15608 -8596 15672
rect -8692 15592 -8596 15608
rect -8692 15528 -8676 15592
rect -8612 15528 -8596 15592
rect -8692 15512 -8596 15528
rect -8692 15448 -8676 15512
rect -8612 15448 -8596 15512
rect -8692 15432 -8596 15448
rect -8692 15368 -8676 15432
rect -8612 15368 -8596 15432
rect -8692 15352 -8596 15368
rect -10104 15252 -10008 15288
rect -8692 15288 -8676 15352
rect -8612 15288 -8596 15352
rect -8273 16032 -7551 16041
rect -8273 15328 -8264 16032
rect -7560 15328 -7551 16032
rect -8273 15319 -7551 15328
rect -7280 16008 -7264 16072
rect -7200 16008 -7184 16072
rect -5868 16072 -5772 16108
rect -7280 15992 -7184 16008
rect -7280 15928 -7264 15992
rect -7200 15928 -7184 15992
rect -7280 15912 -7184 15928
rect -7280 15848 -7264 15912
rect -7200 15848 -7184 15912
rect -7280 15832 -7184 15848
rect -7280 15768 -7264 15832
rect -7200 15768 -7184 15832
rect -7280 15752 -7184 15768
rect -7280 15688 -7264 15752
rect -7200 15688 -7184 15752
rect -7280 15672 -7184 15688
rect -7280 15608 -7264 15672
rect -7200 15608 -7184 15672
rect -7280 15592 -7184 15608
rect -7280 15528 -7264 15592
rect -7200 15528 -7184 15592
rect -7280 15512 -7184 15528
rect -7280 15448 -7264 15512
rect -7200 15448 -7184 15512
rect -7280 15432 -7184 15448
rect -7280 15368 -7264 15432
rect -7200 15368 -7184 15432
rect -7280 15352 -7184 15368
rect -8692 15252 -8596 15288
rect -7280 15288 -7264 15352
rect -7200 15288 -7184 15352
rect -6861 16032 -6139 16041
rect -6861 15328 -6852 16032
rect -6148 15328 -6139 16032
rect -6861 15319 -6139 15328
rect -5868 16008 -5852 16072
rect -5788 16008 -5772 16072
rect -4456 16072 -4360 16108
rect -5868 15992 -5772 16008
rect -5868 15928 -5852 15992
rect -5788 15928 -5772 15992
rect -5868 15912 -5772 15928
rect -5868 15848 -5852 15912
rect -5788 15848 -5772 15912
rect -5868 15832 -5772 15848
rect -5868 15768 -5852 15832
rect -5788 15768 -5772 15832
rect -5868 15752 -5772 15768
rect -5868 15688 -5852 15752
rect -5788 15688 -5772 15752
rect -5868 15672 -5772 15688
rect -5868 15608 -5852 15672
rect -5788 15608 -5772 15672
rect -5868 15592 -5772 15608
rect -5868 15528 -5852 15592
rect -5788 15528 -5772 15592
rect -5868 15512 -5772 15528
rect -5868 15448 -5852 15512
rect -5788 15448 -5772 15512
rect -5868 15432 -5772 15448
rect -5868 15368 -5852 15432
rect -5788 15368 -5772 15432
rect -5868 15352 -5772 15368
rect -7280 15252 -7184 15288
rect -5868 15288 -5852 15352
rect -5788 15288 -5772 15352
rect -5449 16032 -4727 16041
rect -5449 15328 -5440 16032
rect -4736 15328 -4727 16032
rect -5449 15319 -4727 15328
rect -4456 16008 -4440 16072
rect -4376 16008 -4360 16072
rect -3044 16072 -2948 16108
rect -4456 15992 -4360 16008
rect -4456 15928 -4440 15992
rect -4376 15928 -4360 15992
rect -4456 15912 -4360 15928
rect -4456 15848 -4440 15912
rect -4376 15848 -4360 15912
rect -4456 15832 -4360 15848
rect -4456 15768 -4440 15832
rect -4376 15768 -4360 15832
rect -4456 15752 -4360 15768
rect -4456 15688 -4440 15752
rect -4376 15688 -4360 15752
rect -4456 15672 -4360 15688
rect -4456 15608 -4440 15672
rect -4376 15608 -4360 15672
rect -4456 15592 -4360 15608
rect -4456 15528 -4440 15592
rect -4376 15528 -4360 15592
rect -4456 15512 -4360 15528
rect -4456 15448 -4440 15512
rect -4376 15448 -4360 15512
rect -4456 15432 -4360 15448
rect -4456 15368 -4440 15432
rect -4376 15368 -4360 15432
rect -4456 15352 -4360 15368
rect -5868 15252 -5772 15288
rect -4456 15288 -4440 15352
rect -4376 15288 -4360 15352
rect -4037 16032 -3315 16041
rect -4037 15328 -4028 16032
rect -3324 15328 -3315 16032
rect -4037 15319 -3315 15328
rect -3044 16008 -3028 16072
rect -2964 16008 -2948 16072
rect -1632 16072 -1536 16108
rect -3044 15992 -2948 16008
rect -3044 15928 -3028 15992
rect -2964 15928 -2948 15992
rect -3044 15912 -2948 15928
rect -3044 15848 -3028 15912
rect -2964 15848 -2948 15912
rect -3044 15832 -2948 15848
rect -3044 15768 -3028 15832
rect -2964 15768 -2948 15832
rect -3044 15752 -2948 15768
rect -3044 15688 -3028 15752
rect -2964 15688 -2948 15752
rect -3044 15672 -2948 15688
rect -3044 15608 -3028 15672
rect -2964 15608 -2948 15672
rect -3044 15592 -2948 15608
rect -3044 15528 -3028 15592
rect -2964 15528 -2948 15592
rect -3044 15512 -2948 15528
rect -3044 15448 -3028 15512
rect -2964 15448 -2948 15512
rect -3044 15432 -2948 15448
rect -3044 15368 -3028 15432
rect -2964 15368 -2948 15432
rect -3044 15352 -2948 15368
rect -4456 15252 -4360 15288
rect -3044 15288 -3028 15352
rect -2964 15288 -2948 15352
rect -2625 16032 -1903 16041
rect -2625 15328 -2616 16032
rect -1912 15328 -1903 16032
rect -2625 15319 -1903 15328
rect -1632 16008 -1616 16072
rect -1552 16008 -1536 16072
rect -220 16072 -124 16108
rect -1632 15992 -1536 16008
rect -1632 15928 -1616 15992
rect -1552 15928 -1536 15992
rect -1632 15912 -1536 15928
rect -1632 15848 -1616 15912
rect -1552 15848 -1536 15912
rect -1632 15832 -1536 15848
rect -1632 15768 -1616 15832
rect -1552 15768 -1536 15832
rect -1632 15752 -1536 15768
rect -1632 15688 -1616 15752
rect -1552 15688 -1536 15752
rect -1632 15672 -1536 15688
rect -1632 15608 -1616 15672
rect -1552 15608 -1536 15672
rect -1632 15592 -1536 15608
rect -1632 15528 -1616 15592
rect -1552 15528 -1536 15592
rect -1632 15512 -1536 15528
rect -1632 15448 -1616 15512
rect -1552 15448 -1536 15512
rect -1632 15432 -1536 15448
rect -1632 15368 -1616 15432
rect -1552 15368 -1536 15432
rect -1632 15352 -1536 15368
rect -3044 15252 -2948 15288
rect -1632 15288 -1616 15352
rect -1552 15288 -1536 15352
rect -1213 16032 -491 16041
rect -1213 15328 -1204 16032
rect -500 15328 -491 16032
rect -1213 15319 -491 15328
rect -220 16008 -204 16072
rect -140 16008 -124 16072
rect 1192 16072 1288 16108
rect -220 15992 -124 16008
rect -220 15928 -204 15992
rect -140 15928 -124 15992
rect -220 15912 -124 15928
rect -220 15848 -204 15912
rect -140 15848 -124 15912
rect -220 15832 -124 15848
rect -220 15768 -204 15832
rect -140 15768 -124 15832
rect -220 15752 -124 15768
rect -220 15688 -204 15752
rect -140 15688 -124 15752
rect -220 15672 -124 15688
rect -220 15608 -204 15672
rect -140 15608 -124 15672
rect -220 15592 -124 15608
rect -220 15528 -204 15592
rect -140 15528 -124 15592
rect -220 15512 -124 15528
rect -220 15448 -204 15512
rect -140 15448 -124 15512
rect -220 15432 -124 15448
rect -220 15368 -204 15432
rect -140 15368 -124 15432
rect -220 15352 -124 15368
rect -1632 15252 -1536 15288
rect -220 15288 -204 15352
rect -140 15288 -124 15352
rect 199 16032 921 16041
rect 199 15328 208 16032
rect 912 15328 921 16032
rect 199 15319 921 15328
rect 1192 16008 1208 16072
rect 1272 16008 1288 16072
rect 2604 16072 2700 16108
rect 1192 15992 1288 16008
rect 1192 15928 1208 15992
rect 1272 15928 1288 15992
rect 1192 15912 1288 15928
rect 1192 15848 1208 15912
rect 1272 15848 1288 15912
rect 1192 15832 1288 15848
rect 1192 15768 1208 15832
rect 1272 15768 1288 15832
rect 1192 15752 1288 15768
rect 1192 15688 1208 15752
rect 1272 15688 1288 15752
rect 1192 15672 1288 15688
rect 1192 15608 1208 15672
rect 1272 15608 1288 15672
rect 1192 15592 1288 15608
rect 1192 15528 1208 15592
rect 1272 15528 1288 15592
rect 1192 15512 1288 15528
rect 1192 15448 1208 15512
rect 1272 15448 1288 15512
rect 1192 15432 1288 15448
rect 1192 15368 1208 15432
rect 1272 15368 1288 15432
rect 1192 15352 1288 15368
rect -220 15252 -124 15288
rect 1192 15288 1208 15352
rect 1272 15288 1288 15352
rect 1611 16032 2333 16041
rect 1611 15328 1620 16032
rect 2324 15328 2333 16032
rect 1611 15319 2333 15328
rect 2604 16008 2620 16072
rect 2684 16008 2700 16072
rect 4016 16072 4112 16108
rect 2604 15992 2700 16008
rect 2604 15928 2620 15992
rect 2684 15928 2700 15992
rect 2604 15912 2700 15928
rect 2604 15848 2620 15912
rect 2684 15848 2700 15912
rect 2604 15832 2700 15848
rect 2604 15768 2620 15832
rect 2684 15768 2700 15832
rect 2604 15752 2700 15768
rect 2604 15688 2620 15752
rect 2684 15688 2700 15752
rect 2604 15672 2700 15688
rect 2604 15608 2620 15672
rect 2684 15608 2700 15672
rect 2604 15592 2700 15608
rect 2604 15528 2620 15592
rect 2684 15528 2700 15592
rect 2604 15512 2700 15528
rect 2604 15448 2620 15512
rect 2684 15448 2700 15512
rect 2604 15432 2700 15448
rect 2604 15368 2620 15432
rect 2684 15368 2700 15432
rect 2604 15352 2700 15368
rect 1192 15252 1288 15288
rect 2604 15288 2620 15352
rect 2684 15288 2700 15352
rect 3023 16032 3745 16041
rect 3023 15328 3032 16032
rect 3736 15328 3745 16032
rect 3023 15319 3745 15328
rect 4016 16008 4032 16072
rect 4096 16008 4112 16072
rect 5428 16072 5524 16108
rect 4016 15992 4112 16008
rect 4016 15928 4032 15992
rect 4096 15928 4112 15992
rect 4016 15912 4112 15928
rect 4016 15848 4032 15912
rect 4096 15848 4112 15912
rect 4016 15832 4112 15848
rect 4016 15768 4032 15832
rect 4096 15768 4112 15832
rect 4016 15752 4112 15768
rect 4016 15688 4032 15752
rect 4096 15688 4112 15752
rect 4016 15672 4112 15688
rect 4016 15608 4032 15672
rect 4096 15608 4112 15672
rect 4016 15592 4112 15608
rect 4016 15528 4032 15592
rect 4096 15528 4112 15592
rect 4016 15512 4112 15528
rect 4016 15448 4032 15512
rect 4096 15448 4112 15512
rect 4016 15432 4112 15448
rect 4016 15368 4032 15432
rect 4096 15368 4112 15432
rect 4016 15352 4112 15368
rect 2604 15252 2700 15288
rect 4016 15288 4032 15352
rect 4096 15288 4112 15352
rect 4435 16032 5157 16041
rect 4435 15328 4444 16032
rect 5148 15328 5157 16032
rect 4435 15319 5157 15328
rect 5428 16008 5444 16072
rect 5508 16008 5524 16072
rect 6840 16072 6936 16108
rect 5428 15992 5524 16008
rect 5428 15928 5444 15992
rect 5508 15928 5524 15992
rect 5428 15912 5524 15928
rect 5428 15848 5444 15912
rect 5508 15848 5524 15912
rect 5428 15832 5524 15848
rect 5428 15768 5444 15832
rect 5508 15768 5524 15832
rect 5428 15752 5524 15768
rect 5428 15688 5444 15752
rect 5508 15688 5524 15752
rect 5428 15672 5524 15688
rect 5428 15608 5444 15672
rect 5508 15608 5524 15672
rect 5428 15592 5524 15608
rect 5428 15528 5444 15592
rect 5508 15528 5524 15592
rect 5428 15512 5524 15528
rect 5428 15448 5444 15512
rect 5508 15448 5524 15512
rect 5428 15432 5524 15448
rect 5428 15368 5444 15432
rect 5508 15368 5524 15432
rect 5428 15352 5524 15368
rect 4016 15252 4112 15288
rect 5428 15288 5444 15352
rect 5508 15288 5524 15352
rect 5847 16032 6569 16041
rect 5847 15328 5856 16032
rect 6560 15328 6569 16032
rect 5847 15319 6569 15328
rect 6840 16008 6856 16072
rect 6920 16008 6936 16072
rect 8252 16072 8348 16108
rect 6840 15992 6936 16008
rect 6840 15928 6856 15992
rect 6920 15928 6936 15992
rect 6840 15912 6936 15928
rect 6840 15848 6856 15912
rect 6920 15848 6936 15912
rect 6840 15832 6936 15848
rect 6840 15768 6856 15832
rect 6920 15768 6936 15832
rect 6840 15752 6936 15768
rect 6840 15688 6856 15752
rect 6920 15688 6936 15752
rect 6840 15672 6936 15688
rect 6840 15608 6856 15672
rect 6920 15608 6936 15672
rect 6840 15592 6936 15608
rect 6840 15528 6856 15592
rect 6920 15528 6936 15592
rect 6840 15512 6936 15528
rect 6840 15448 6856 15512
rect 6920 15448 6936 15512
rect 6840 15432 6936 15448
rect 6840 15368 6856 15432
rect 6920 15368 6936 15432
rect 6840 15352 6936 15368
rect 5428 15252 5524 15288
rect 6840 15288 6856 15352
rect 6920 15288 6936 15352
rect 7259 16032 7981 16041
rect 7259 15328 7268 16032
rect 7972 15328 7981 16032
rect 7259 15319 7981 15328
rect 8252 16008 8268 16072
rect 8332 16008 8348 16072
rect 9664 16072 9760 16108
rect 8252 15992 8348 16008
rect 8252 15928 8268 15992
rect 8332 15928 8348 15992
rect 8252 15912 8348 15928
rect 8252 15848 8268 15912
rect 8332 15848 8348 15912
rect 8252 15832 8348 15848
rect 8252 15768 8268 15832
rect 8332 15768 8348 15832
rect 8252 15752 8348 15768
rect 8252 15688 8268 15752
rect 8332 15688 8348 15752
rect 8252 15672 8348 15688
rect 8252 15608 8268 15672
rect 8332 15608 8348 15672
rect 8252 15592 8348 15608
rect 8252 15528 8268 15592
rect 8332 15528 8348 15592
rect 8252 15512 8348 15528
rect 8252 15448 8268 15512
rect 8332 15448 8348 15512
rect 8252 15432 8348 15448
rect 8252 15368 8268 15432
rect 8332 15368 8348 15432
rect 8252 15352 8348 15368
rect 6840 15252 6936 15288
rect 8252 15288 8268 15352
rect 8332 15288 8348 15352
rect 8671 16032 9393 16041
rect 8671 15328 8680 16032
rect 9384 15328 9393 16032
rect 8671 15319 9393 15328
rect 9664 16008 9680 16072
rect 9744 16008 9760 16072
rect 11076 16072 11172 16108
rect 9664 15992 9760 16008
rect 9664 15928 9680 15992
rect 9744 15928 9760 15992
rect 9664 15912 9760 15928
rect 9664 15848 9680 15912
rect 9744 15848 9760 15912
rect 9664 15832 9760 15848
rect 9664 15768 9680 15832
rect 9744 15768 9760 15832
rect 9664 15752 9760 15768
rect 9664 15688 9680 15752
rect 9744 15688 9760 15752
rect 9664 15672 9760 15688
rect 9664 15608 9680 15672
rect 9744 15608 9760 15672
rect 9664 15592 9760 15608
rect 9664 15528 9680 15592
rect 9744 15528 9760 15592
rect 9664 15512 9760 15528
rect 9664 15448 9680 15512
rect 9744 15448 9760 15512
rect 9664 15432 9760 15448
rect 9664 15368 9680 15432
rect 9744 15368 9760 15432
rect 9664 15352 9760 15368
rect 8252 15252 8348 15288
rect 9664 15288 9680 15352
rect 9744 15288 9760 15352
rect 10083 16032 10805 16041
rect 10083 15328 10092 16032
rect 10796 15328 10805 16032
rect 10083 15319 10805 15328
rect 11076 16008 11092 16072
rect 11156 16008 11172 16072
rect 12488 16072 12584 16108
rect 11076 15992 11172 16008
rect 11076 15928 11092 15992
rect 11156 15928 11172 15992
rect 11076 15912 11172 15928
rect 11076 15848 11092 15912
rect 11156 15848 11172 15912
rect 11076 15832 11172 15848
rect 11076 15768 11092 15832
rect 11156 15768 11172 15832
rect 11076 15752 11172 15768
rect 11076 15688 11092 15752
rect 11156 15688 11172 15752
rect 11076 15672 11172 15688
rect 11076 15608 11092 15672
rect 11156 15608 11172 15672
rect 11076 15592 11172 15608
rect 11076 15528 11092 15592
rect 11156 15528 11172 15592
rect 11076 15512 11172 15528
rect 11076 15448 11092 15512
rect 11156 15448 11172 15512
rect 11076 15432 11172 15448
rect 11076 15368 11092 15432
rect 11156 15368 11172 15432
rect 11076 15352 11172 15368
rect 9664 15252 9760 15288
rect 11076 15288 11092 15352
rect 11156 15288 11172 15352
rect 11495 16032 12217 16041
rect 11495 15328 11504 16032
rect 12208 15328 12217 16032
rect 11495 15319 12217 15328
rect 12488 16008 12504 16072
rect 12568 16008 12584 16072
rect 13900 16072 13996 16108
rect 12488 15992 12584 16008
rect 12488 15928 12504 15992
rect 12568 15928 12584 15992
rect 12488 15912 12584 15928
rect 12488 15848 12504 15912
rect 12568 15848 12584 15912
rect 12488 15832 12584 15848
rect 12488 15768 12504 15832
rect 12568 15768 12584 15832
rect 12488 15752 12584 15768
rect 12488 15688 12504 15752
rect 12568 15688 12584 15752
rect 12488 15672 12584 15688
rect 12488 15608 12504 15672
rect 12568 15608 12584 15672
rect 12488 15592 12584 15608
rect 12488 15528 12504 15592
rect 12568 15528 12584 15592
rect 12488 15512 12584 15528
rect 12488 15448 12504 15512
rect 12568 15448 12584 15512
rect 12488 15432 12584 15448
rect 12488 15368 12504 15432
rect 12568 15368 12584 15432
rect 12488 15352 12584 15368
rect 11076 15252 11172 15288
rect 12488 15288 12504 15352
rect 12568 15288 12584 15352
rect 12907 16032 13629 16041
rect 12907 15328 12916 16032
rect 13620 15328 13629 16032
rect 12907 15319 13629 15328
rect 13900 16008 13916 16072
rect 13980 16008 13996 16072
rect 15312 16072 15408 16108
rect 13900 15992 13996 16008
rect 13900 15928 13916 15992
rect 13980 15928 13996 15992
rect 13900 15912 13996 15928
rect 13900 15848 13916 15912
rect 13980 15848 13996 15912
rect 13900 15832 13996 15848
rect 13900 15768 13916 15832
rect 13980 15768 13996 15832
rect 13900 15752 13996 15768
rect 13900 15688 13916 15752
rect 13980 15688 13996 15752
rect 13900 15672 13996 15688
rect 13900 15608 13916 15672
rect 13980 15608 13996 15672
rect 13900 15592 13996 15608
rect 13900 15528 13916 15592
rect 13980 15528 13996 15592
rect 13900 15512 13996 15528
rect 13900 15448 13916 15512
rect 13980 15448 13996 15512
rect 13900 15432 13996 15448
rect 13900 15368 13916 15432
rect 13980 15368 13996 15432
rect 13900 15352 13996 15368
rect 12488 15252 12584 15288
rect 13900 15288 13916 15352
rect 13980 15288 13996 15352
rect 14319 16032 15041 16041
rect 14319 15328 14328 16032
rect 15032 15328 15041 16032
rect 14319 15319 15041 15328
rect 15312 16008 15328 16072
rect 15392 16008 15408 16072
rect 16724 16072 16820 16108
rect 15312 15992 15408 16008
rect 15312 15928 15328 15992
rect 15392 15928 15408 15992
rect 15312 15912 15408 15928
rect 15312 15848 15328 15912
rect 15392 15848 15408 15912
rect 15312 15832 15408 15848
rect 15312 15768 15328 15832
rect 15392 15768 15408 15832
rect 15312 15752 15408 15768
rect 15312 15688 15328 15752
rect 15392 15688 15408 15752
rect 15312 15672 15408 15688
rect 15312 15608 15328 15672
rect 15392 15608 15408 15672
rect 15312 15592 15408 15608
rect 15312 15528 15328 15592
rect 15392 15528 15408 15592
rect 15312 15512 15408 15528
rect 15312 15448 15328 15512
rect 15392 15448 15408 15512
rect 15312 15432 15408 15448
rect 15312 15368 15328 15432
rect 15392 15368 15408 15432
rect 15312 15352 15408 15368
rect 13900 15252 13996 15288
rect 15312 15288 15328 15352
rect 15392 15288 15408 15352
rect 15731 16032 16453 16041
rect 15731 15328 15740 16032
rect 16444 15328 16453 16032
rect 15731 15319 16453 15328
rect 16724 16008 16740 16072
rect 16804 16008 16820 16072
rect 18136 16072 18232 16108
rect 16724 15992 16820 16008
rect 16724 15928 16740 15992
rect 16804 15928 16820 15992
rect 16724 15912 16820 15928
rect 16724 15848 16740 15912
rect 16804 15848 16820 15912
rect 16724 15832 16820 15848
rect 16724 15768 16740 15832
rect 16804 15768 16820 15832
rect 16724 15752 16820 15768
rect 16724 15688 16740 15752
rect 16804 15688 16820 15752
rect 16724 15672 16820 15688
rect 16724 15608 16740 15672
rect 16804 15608 16820 15672
rect 16724 15592 16820 15608
rect 16724 15528 16740 15592
rect 16804 15528 16820 15592
rect 16724 15512 16820 15528
rect 16724 15448 16740 15512
rect 16804 15448 16820 15512
rect 16724 15432 16820 15448
rect 16724 15368 16740 15432
rect 16804 15368 16820 15432
rect 16724 15352 16820 15368
rect 15312 15252 15408 15288
rect 16724 15288 16740 15352
rect 16804 15288 16820 15352
rect 17143 16032 17865 16041
rect 17143 15328 17152 16032
rect 17856 15328 17865 16032
rect 17143 15319 17865 15328
rect 18136 16008 18152 16072
rect 18216 16008 18232 16072
rect 19548 16072 19644 16108
rect 18136 15992 18232 16008
rect 18136 15928 18152 15992
rect 18216 15928 18232 15992
rect 18136 15912 18232 15928
rect 18136 15848 18152 15912
rect 18216 15848 18232 15912
rect 18136 15832 18232 15848
rect 18136 15768 18152 15832
rect 18216 15768 18232 15832
rect 18136 15752 18232 15768
rect 18136 15688 18152 15752
rect 18216 15688 18232 15752
rect 18136 15672 18232 15688
rect 18136 15608 18152 15672
rect 18216 15608 18232 15672
rect 18136 15592 18232 15608
rect 18136 15528 18152 15592
rect 18216 15528 18232 15592
rect 18136 15512 18232 15528
rect 18136 15448 18152 15512
rect 18216 15448 18232 15512
rect 18136 15432 18232 15448
rect 18136 15368 18152 15432
rect 18216 15368 18232 15432
rect 18136 15352 18232 15368
rect 16724 15252 16820 15288
rect 18136 15288 18152 15352
rect 18216 15288 18232 15352
rect 18555 16032 19277 16041
rect 18555 15328 18564 16032
rect 19268 15328 19277 16032
rect 18555 15319 19277 15328
rect 19548 16008 19564 16072
rect 19628 16008 19644 16072
rect 20960 16072 21056 16108
rect 19548 15992 19644 16008
rect 19548 15928 19564 15992
rect 19628 15928 19644 15992
rect 19548 15912 19644 15928
rect 19548 15848 19564 15912
rect 19628 15848 19644 15912
rect 19548 15832 19644 15848
rect 19548 15768 19564 15832
rect 19628 15768 19644 15832
rect 19548 15752 19644 15768
rect 19548 15688 19564 15752
rect 19628 15688 19644 15752
rect 19548 15672 19644 15688
rect 19548 15608 19564 15672
rect 19628 15608 19644 15672
rect 19548 15592 19644 15608
rect 19548 15528 19564 15592
rect 19628 15528 19644 15592
rect 19548 15512 19644 15528
rect 19548 15448 19564 15512
rect 19628 15448 19644 15512
rect 19548 15432 19644 15448
rect 19548 15368 19564 15432
rect 19628 15368 19644 15432
rect 19548 15352 19644 15368
rect 18136 15252 18232 15288
rect 19548 15288 19564 15352
rect 19628 15288 19644 15352
rect 19967 16032 20689 16041
rect 19967 15328 19976 16032
rect 20680 15328 20689 16032
rect 19967 15319 20689 15328
rect 20960 16008 20976 16072
rect 21040 16008 21056 16072
rect 22372 16072 22468 16108
rect 20960 15992 21056 16008
rect 20960 15928 20976 15992
rect 21040 15928 21056 15992
rect 20960 15912 21056 15928
rect 20960 15848 20976 15912
rect 21040 15848 21056 15912
rect 20960 15832 21056 15848
rect 20960 15768 20976 15832
rect 21040 15768 21056 15832
rect 20960 15752 21056 15768
rect 20960 15688 20976 15752
rect 21040 15688 21056 15752
rect 20960 15672 21056 15688
rect 20960 15608 20976 15672
rect 21040 15608 21056 15672
rect 20960 15592 21056 15608
rect 20960 15528 20976 15592
rect 21040 15528 21056 15592
rect 20960 15512 21056 15528
rect 20960 15448 20976 15512
rect 21040 15448 21056 15512
rect 20960 15432 21056 15448
rect 20960 15368 20976 15432
rect 21040 15368 21056 15432
rect 20960 15352 21056 15368
rect 19548 15252 19644 15288
rect 20960 15288 20976 15352
rect 21040 15288 21056 15352
rect 21379 16032 22101 16041
rect 21379 15328 21388 16032
rect 22092 15328 22101 16032
rect 21379 15319 22101 15328
rect 22372 16008 22388 16072
rect 22452 16008 22468 16072
rect 23784 16072 23880 16108
rect 22372 15992 22468 16008
rect 22372 15928 22388 15992
rect 22452 15928 22468 15992
rect 22372 15912 22468 15928
rect 22372 15848 22388 15912
rect 22452 15848 22468 15912
rect 22372 15832 22468 15848
rect 22372 15768 22388 15832
rect 22452 15768 22468 15832
rect 22372 15752 22468 15768
rect 22372 15688 22388 15752
rect 22452 15688 22468 15752
rect 22372 15672 22468 15688
rect 22372 15608 22388 15672
rect 22452 15608 22468 15672
rect 22372 15592 22468 15608
rect 22372 15528 22388 15592
rect 22452 15528 22468 15592
rect 22372 15512 22468 15528
rect 22372 15448 22388 15512
rect 22452 15448 22468 15512
rect 22372 15432 22468 15448
rect 22372 15368 22388 15432
rect 22452 15368 22468 15432
rect 22372 15352 22468 15368
rect 20960 15252 21056 15288
rect 22372 15288 22388 15352
rect 22452 15288 22468 15352
rect 22791 16032 23513 16041
rect 22791 15328 22800 16032
rect 23504 15328 23513 16032
rect 22791 15319 23513 15328
rect 23784 16008 23800 16072
rect 23864 16008 23880 16072
rect 23784 15992 23880 16008
rect 23784 15928 23800 15992
rect 23864 15928 23880 15992
rect 23784 15912 23880 15928
rect 23784 15848 23800 15912
rect 23864 15848 23880 15912
rect 23784 15832 23880 15848
rect 23784 15768 23800 15832
rect 23864 15768 23880 15832
rect 23784 15752 23880 15768
rect 23784 15688 23800 15752
rect 23864 15688 23880 15752
rect 23784 15672 23880 15688
rect 23784 15608 23800 15672
rect 23864 15608 23880 15672
rect 23784 15592 23880 15608
rect 23784 15528 23800 15592
rect 23864 15528 23880 15592
rect 23784 15512 23880 15528
rect 23784 15448 23800 15512
rect 23864 15448 23880 15512
rect 23784 15432 23880 15448
rect 23784 15368 23800 15432
rect 23864 15368 23880 15432
rect 23784 15352 23880 15368
rect 22372 15252 22468 15288
rect 23784 15288 23800 15352
rect 23864 15288 23880 15352
rect 23784 15252 23880 15288
rect -22812 14952 -22716 14988
rect -23805 14912 -23083 14921
rect -23805 14208 -23796 14912
rect -23092 14208 -23083 14912
rect -23805 14199 -23083 14208
rect -22812 14888 -22796 14952
rect -22732 14888 -22716 14952
rect -21400 14952 -21304 14988
rect -22812 14872 -22716 14888
rect -22812 14808 -22796 14872
rect -22732 14808 -22716 14872
rect -22812 14792 -22716 14808
rect -22812 14728 -22796 14792
rect -22732 14728 -22716 14792
rect -22812 14712 -22716 14728
rect -22812 14648 -22796 14712
rect -22732 14648 -22716 14712
rect -22812 14632 -22716 14648
rect -22812 14568 -22796 14632
rect -22732 14568 -22716 14632
rect -22812 14552 -22716 14568
rect -22812 14488 -22796 14552
rect -22732 14488 -22716 14552
rect -22812 14472 -22716 14488
rect -22812 14408 -22796 14472
rect -22732 14408 -22716 14472
rect -22812 14392 -22716 14408
rect -22812 14328 -22796 14392
rect -22732 14328 -22716 14392
rect -22812 14312 -22716 14328
rect -22812 14248 -22796 14312
rect -22732 14248 -22716 14312
rect -22812 14232 -22716 14248
rect -22812 14168 -22796 14232
rect -22732 14168 -22716 14232
rect -22393 14912 -21671 14921
rect -22393 14208 -22384 14912
rect -21680 14208 -21671 14912
rect -22393 14199 -21671 14208
rect -21400 14888 -21384 14952
rect -21320 14888 -21304 14952
rect -19988 14952 -19892 14988
rect -21400 14872 -21304 14888
rect -21400 14808 -21384 14872
rect -21320 14808 -21304 14872
rect -21400 14792 -21304 14808
rect -21400 14728 -21384 14792
rect -21320 14728 -21304 14792
rect -21400 14712 -21304 14728
rect -21400 14648 -21384 14712
rect -21320 14648 -21304 14712
rect -21400 14632 -21304 14648
rect -21400 14568 -21384 14632
rect -21320 14568 -21304 14632
rect -21400 14552 -21304 14568
rect -21400 14488 -21384 14552
rect -21320 14488 -21304 14552
rect -21400 14472 -21304 14488
rect -21400 14408 -21384 14472
rect -21320 14408 -21304 14472
rect -21400 14392 -21304 14408
rect -21400 14328 -21384 14392
rect -21320 14328 -21304 14392
rect -21400 14312 -21304 14328
rect -21400 14248 -21384 14312
rect -21320 14248 -21304 14312
rect -21400 14232 -21304 14248
rect -22812 14132 -22716 14168
rect -21400 14168 -21384 14232
rect -21320 14168 -21304 14232
rect -20981 14912 -20259 14921
rect -20981 14208 -20972 14912
rect -20268 14208 -20259 14912
rect -20981 14199 -20259 14208
rect -19988 14888 -19972 14952
rect -19908 14888 -19892 14952
rect -18576 14952 -18480 14988
rect -19988 14872 -19892 14888
rect -19988 14808 -19972 14872
rect -19908 14808 -19892 14872
rect -19988 14792 -19892 14808
rect -19988 14728 -19972 14792
rect -19908 14728 -19892 14792
rect -19988 14712 -19892 14728
rect -19988 14648 -19972 14712
rect -19908 14648 -19892 14712
rect -19988 14632 -19892 14648
rect -19988 14568 -19972 14632
rect -19908 14568 -19892 14632
rect -19988 14552 -19892 14568
rect -19988 14488 -19972 14552
rect -19908 14488 -19892 14552
rect -19988 14472 -19892 14488
rect -19988 14408 -19972 14472
rect -19908 14408 -19892 14472
rect -19988 14392 -19892 14408
rect -19988 14328 -19972 14392
rect -19908 14328 -19892 14392
rect -19988 14312 -19892 14328
rect -19988 14248 -19972 14312
rect -19908 14248 -19892 14312
rect -19988 14232 -19892 14248
rect -21400 14132 -21304 14168
rect -19988 14168 -19972 14232
rect -19908 14168 -19892 14232
rect -19569 14912 -18847 14921
rect -19569 14208 -19560 14912
rect -18856 14208 -18847 14912
rect -19569 14199 -18847 14208
rect -18576 14888 -18560 14952
rect -18496 14888 -18480 14952
rect -17164 14952 -17068 14988
rect -18576 14872 -18480 14888
rect -18576 14808 -18560 14872
rect -18496 14808 -18480 14872
rect -18576 14792 -18480 14808
rect -18576 14728 -18560 14792
rect -18496 14728 -18480 14792
rect -18576 14712 -18480 14728
rect -18576 14648 -18560 14712
rect -18496 14648 -18480 14712
rect -18576 14632 -18480 14648
rect -18576 14568 -18560 14632
rect -18496 14568 -18480 14632
rect -18576 14552 -18480 14568
rect -18576 14488 -18560 14552
rect -18496 14488 -18480 14552
rect -18576 14472 -18480 14488
rect -18576 14408 -18560 14472
rect -18496 14408 -18480 14472
rect -18576 14392 -18480 14408
rect -18576 14328 -18560 14392
rect -18496 14328 -18480 14392
rect -18576 14312 -18480 14328
rect -18576 14248 -18560 14312
rect -18496 14248 -18480 14312
rect -18576 14232 -18480 14248
rect -19988 14132 -19892 14168
rect -18576 14168 -18560 14232
rect -18496 14168 -18480 14232
rect -18157 14912 -17435 14921
rect -18157 14208 -18148 14912
rect -17444 14208 -17435 14912
rect -18157 14199 -17435 14208
rect -17164 14888 -17148 14952
rect -17084 14888 -17068 14952
rect -15752 14952 -15656 14988
rect -17164 14872 -17068 14888
rect -17164 14808 -17148 14872
rect -17084 14808 -17068 14872
rect -17164 14792 -17068 14808
rect -17164 14728 -17148 14792
rect -17084 14728 -17068 14792
rect -17164 14712 -17068 14728
rect -17164 14648 -17148 14712
rect -17084 14648 -17068 14712
rect -17164 14632 -17068 14648
rect -17164 14568 -17148 14632
rect -17084 14568 -17068 14632
rect -17164 14552 -17068 14568
rect -17164 14488 -17148 14552
rect -17084 14488 -17068 14552
rect -17164 14472 -17068 14488
rect -17164 14408 -17148 14472
rect -17084 14408 -17068 14472
rect -17164 14392 -17068 14408
rect -17164 14328 -17148 14392
rect -17084 14328 -17068 14392
rect -17164 14312 -17068 14328
rect -17164 14248 -17148 14312
rect -17084 14248 -17068 14312
rect -17164 14232 -17068 14248
rect -18576 14132 -18480 14168
rect -17164 14168 -17148 14232
rect -17084 14168 -17068 14232
rect -16745 14912 -16023 14921
rect -16745 14208 -16736 14912
rect -16032 14208 -16023 14912
rect -16745 14199 -16023 14208
rect -15752 14888 -15736 14952
rect -15672 14888 -15656 14952
rect -14340 14952 -14244 14988
rect -15752 14872 -15656 14888
rect -15752 14808 -15736 14872
rect -15672 14808 -15656 14872
rect -15752 14792 -15656 14808
rect -15752 14728 -15736 14792
rect -15672 14728 -15656 14792
rect -15752 14712 -15656 14728
rect -15752 14648 -15736 14712
rect -15672 14648 -15656 14712
rect -15752 14632 -15656 14648
rect -15752 14568 -15736 14632
rect -15672 14568 -15656 14632
rect -15752 14552 -15656 14568
rect -15752 14488 -15736 14552
rect -15672 14488 -15656 14552
rect -15752 14472 -15656 14488
rect -15752 14408 -15736 14472
rect -15672 14408 -15656 14472
rect -15752 14392 -15656 14408
rect -15752 14328 -15736 14392
rect -15672 14328 -15656 14392
rect -15752 14312 -15656 14328
rect -15752 14248 -15736 14312
rect -15672 14248 -15656 14312
rect -15752 14232 -15656 14248
rect -17164 14132 -17068 14168
rect -15752 14168 -15736 14232
rect -15672 14168 -15656 14232
rect -15333 14912 -14611 14921
rect -15333 14208 -15324 14912
rect -14620 14208 -14611 14912
rect -15333 14199 -14611 14208
rect -14340 14888 -14324 14952
rect -14260 14888 -14244 14952
rect -12928 14952 -12832 14988
rect -14340 14872 -14244 14888
rect -14340 14808 -14324 14872
rect -14260 14808 -14244 14872
rect -14340 14792 -14244 14808
rect -14340 14728 -14324 14792
rect -14260 14728 -14244 14792
rect -14340 14712 -14244 14728
rect -14340 14648 -14324 14712
rect -14260 14648 -14244 14712
rect -14340 14632 -14244 14648
rect -14340 14568 -14324 14632
rect -14260 14568 -14244 14632
rect -14340 14552 -14244 14568
rect -14340 14488 -14324 14552
rect -14260 14488 -14244 14552
rect -14340 14472 -14244 14488
rect -14340 14408 -14324 14472
rect -14260 14408 -14244 14472
rect -14340 14392 -14244 14408
rect -14340 14328 -14324 14392
rect -14260 14328 -14244 14392
rect -14340 14312 -14244 14328
rect -14340 14248 -14324 14312
rect -14260 14248 -14244 14312
rect -14340 14232 -14244 14248
rect -15752 14132 -15656 14168
rect -14340 14168 -14324 14232
rect -14260 14168 -14244 14232
rect -13921 14912 -13199 14921
rect -13921 14208 -13912 14912
rect -13208 14208 -13199 14912
rect -13921 14199 -13199 14208
rect -12928 14888 -12912 14952
rect -12848 14888 -12832 14952
rect -11516 14952 -11420 14988
rect -12928 14872 -12832 14888
rect -12928 14808 -12912 14872
rect -12848 14808 -12832 14872
rect -12928 14792 -12832 14808
rect -12928 14728 -12912 14792
rect -12848 14728 -12832 14792
rect -12928 14712 -12832 14728
rect -12928 14648 -12912 14712
rect -12848 14648 -12832 14712
rect -12928 14632 -12832 14648
rect -12928 14568 -12912 14632
rect -12848 14568 -12832 14632
rect -12928 14552 -12832 14568
rect -12928 14488 -12912 14552
rect -12848 14488 -12832 14552
rect -12928 14472 -12832 14488
rect -12928 14408 -12912 14472
rect -12848 14408 -12832 14472
rect -12928 14392 -12832 14408
rect -12928 14328 -12912 14392
rect -12848 14328 -12832 14392
rect -12928 14312 -12832 14328
rect -12928 14248 -12912 14312
rect -12848 14248 -12832 14312
rect -12928 14232 -12832 14248
rect -14340 14132 -14244 14168
rect -12928 14168 -12912 14232
rect -12848 14168 -12832 14232
rect -12509 14912 -11787 14921
rect -12509 14208 -12500 14912
rect -11796 14208 -11787 14912
rect -12509 14199 -11787 14208
rect -11516 14888 -11500 14952
rect -11436 14888 -11420 14952
rect -10104 14952 -10008 14988
rect -11516 14872 -11420 14888
rect -11516 14808 -11500 14872
rect -11436 14808 -11420 14872
rect -11516 14792 -11420 14808
rect -11516 14728 -11500 14792
rect -11436 14728 -11420 14792
rect -11516 14712 -11420 14728
rect -11516 14648 -11500 14712
rect -11436 14648 -11420 14712
rect -11516 14632 -11420 14648
rect -11516 14568 -11500 14632
rect -11436 14568 -11420 14632
rect -11516 14552 -11420 14568
rect -11516 14488 -11500 14552
rect -11436 14488 -11420 14552
rect -11516 14472 -11420 14488
rect -11516 14408 -11500 14472
rect -11436 14408 -11420 14472
rect -11516 14392 -11420 14408
rect -11516 14328 -11500 14392
rect -11436 14328 -11420 14392
rect -11516 14312 -11420 14328
rect -11516 14248 -11500 14312
rect -11436 14248 -11420 14312
rect -11516 14232 -11420 14248
rect -12928 14132 -12832 14168
rect -11516 14168 -11500 14232
rect -11436 14168 -11420 14232
rect -11097 14912 -10375 14921
rect -11097 14208 -11088 14912
rect -10384 14208 -10375 14912
rect -11097 14199 -10375 14208
rect -10104 14888 -10088 14952
rect -10024 14888 -10008 14952
rect -8692 14952 -8596 14988
rect -10104 14872 -10008 14888
rect -10104 14808 -10088 14872
rect -10024 14808 -10008 14872
rect -10104 14792 -10008 14808
rect -10104 14728 -10088 14792
rect -10024 14728 -10008 14792
rect -10104 14712 -10008 14728
rect -10104 14648 -10088 14712
rect -10024 14648 -10008 14712
rect -10104 14632 -10008 14648
rect -10104 14568 -10088 14632
rect -10024 14568 -10008 14632
rect -10104 14552 -10008 14568
rect -10104 14488 -10088 14552
rect -10024 14488 -10008 14552
rect -10104 14472 -10008 14488
rect -10104 14408 -10088 14472
rect -10024 14408 -10008 14472
rect -10104 14392 -10008 14408
rect -10104 14328 -10088 14392
rect -10024 14328 -10008 14392
rect -10104 14312 -10008 14328
rect -10104 14248 -10088 14312
rect -10024 14248 -10008 14312
rect -10104 14232 -10008 14248
rect -11516 14132 -11420 14168
rect -10104 14168 -10088 14232
rect -10024 14168 -10008 14232
rect -9685 14912 -8963 14921
rect -9685 14208 -9676 14912
rect -8972 14208 -8963 14912
rect -9685 14199 -8963 14208
rect -8692 14888 -8676 14952
rect -8612 14888 -8596 14952
rect -7280 14952 -7184 14988
rect -8692 14872 -8596 14888
rect -8692 14808 -8676 14872
rect -8612 14808 -8596 14872
rect -8692 14792 -8596 14808
rect -8692 14728 -8676 14792
rect -8612 14728 -8596 14792
rect -8692 14712 -8596 14728
rect -8692 14648 -8676 14712
rect -8612 14648 -8596 14712
rect -8692 14632 -8596 14648
rect -8692 14568 -8676 14632
rect -8612 14568 -8596 14632
rect -8692 14552 -8596 14568
rect -8692 14488 -8676 14552
rect -8612 14488 -8596 14552
rect -8692 14472 -8596 14488
rect -8692 14408 -8676 14472
rect -8612 14408 -8596 14472
rect -8692 14392 -8596 14408
rect -8692 14328 -8676 14392
rect -8612 14328 -8596 14392
rect -8692 14312 -8596 14328
rect -8692 14248 -8676 14312
rect -8612 14248 -8596 14312
rect -8692 14232 -8596 14248
rect -10104 14132 -10008 14168
rect -8692 14168 -8676 14232
rect -8612 14168 -8596 14232
rect -8273 14912 -7551 14921
rect -8273 14208 -8264 14912
rect -7560 14208 -7551 14912
rect -8273 14199 -7551 14208
rect -7280 14888 -7264 14952
rect -7200 14888 -7184 14952
rect -5868 14952 -5772 14988
rect -7280 14872 -7184 14888
rect -7280 14808 -7264 14872
rect -7200 14808 -7184 14872
rect -7280 14792 -7184 14808
rect -7280 14728 -7264 14792
rect -7200 14728 -7184 14792
rect -7280 14712 -7184 14728
rect -7280 14648 -7264 14712
rect -7200 14648 -7184 14712
rect -7280 14632 -7184 14648
rect -7280 14568 -7264 14632
rect -7200 14568 -7184 14632
rect -7280 14552 -7184 14568
rect -7280 14488 -7264 14552
rect -7200 14488 -7184 14552
rect -7280 14472 -7184 14488
rect -7280 14408 -7264 14472
rect -7200 14408 -7184 14472
rect -7280 14392 -7184 14408
rect -7280 14328 -7264 14392
rect -7200 14328 -7184 14392
rect -7280 14312 -7184 14328
rect -7280 14248 -7264 14312
rect -7200 14248 -7184 14312
rect -7280 14232 -7184 14248
rect -8692 14132 -8596 14168
rect -7280 14168 -7264 14232
rect -7200 14168 -7184 14232
rect -6861 14912 -6139 14921
rect -6861 14208 -6852 14912
rect -6148 14208 -6139 14912
rect -6861 14199 -6139 14208
rect -5868 14888 -5852 14952
rect -5788 14888 -5772 14952
rect -4456 14952 -4360 14988
rect -5868 14872 -5772 14888
rect -5868 14808 -5852 14872
rect -5788 14808 -5772 14872
rect -5868 14792 -5772 14808
rect -5868 14728 -5852 14792
rect -5788 14728 -5772 14792
rect -5868 14712 -5772 14728
rect -5868 14648 -5852 14712
rect -5788 14648 -5772 14712
rect -5868 14632 -5772 14648
rect -5868 14568 -5852 14632
rect -5788 14568 -5772 14632
rect -5868 14552 -5772 14568
rect -5868 14488 -5852 14552
rect -5788 14488 -5772 14552
rect -5868 14472 -5772 14488
rect -5868 14408 -5852 14472
rect -5788 14408 -5772 14472
rect -5868 14392 -5772 14408
rect -5868 14328 -5852 14392
rect -5788 14328 -5772 14392
rect -5868 14312 -5772 14328
rect -5868 14248 -5852 14312
rect -5788 14248 -5772 14312
rect -5868 14232 -5772 14248
rect -7280 14132 -7184 14168
rect -5868 14168 -5852 14232
rect -5788 14168 -5772 14232
rect -5449 14912 -4727 14921
rect -5449 14208 -5440 14912
rect -4736 14208 -4727 14912
rect -5449 14199 -4727 14208
rect -4456 14888 -4440 14952
rect -4376 14888 -4360 14952
rect -3044 14952 -2948 14988
rect -4456 14872 -4360 14888
rect -4456 14808 -4440 14872
rect -4376 14808 -4360 14872
rect -4456 14792 -4360 14808
rect -4456 14728 -4440 14792
rect -4376 14728 -4360 14792
rect -4456 14712 -4360 14728
rect -4456 14648 -4440 14712
rect -4376 14648 -4360 14712
rect -4456 14632 -4360 14648
rect -4456 14568 -4440 14632
rect -4376 14568 -4360 14632
rect -4456 14552 -4360 14568
rect -4456 14488 -4440 14552
rect -4376 14488 -4360 14552
rect -4456 14472 -4360 14488
rect -4456 14408 -4440 14472
rect -4376 14408 -4360 14472
rect -4456 14392 -4360 14408
rect -4456 14328 -4440 14392
rect -4376 14328 -4360 14392
rect -4456 14312 -4360 14328
rect -4456 14248 -4440 14312
rect -4376 14248 -4360 14312
rect -4456 14232 -4360 14248
rect -5868 14132 -5772 14168
rect -4456 14168 -4440 14232
rect -4376 14168 -4360 14232
rect -4037 14912 -3315 14921
rect -4037 14208 -4028 14912
rect -3324 14208 -3315 14912
rect -4037 14199 -3315 14208
rect -3044 14888 -3028 14952
rect -2964 14888 -2948 14952
rect -1632 14952 -1536 14988
rect -3044 14872 -2948 14888
rect -3044 14808 -3028 14872
rect -2964 14808 -2948 14872
rect -3044 14792 -2948 14808
rect -3044 14728 -3028 14792
rect -2964 14728 -2948 14792
rect -3044 14712 -2948 14728
rect -3044 14648 -3028 14712
rect -2964 14648 -2948 14712
rect -3044 14632 -2948 14648
rect -3044 14568 -3028 14632
rect -2964 14568 -2948 14632
rect -3044 14552 -2948 14568
rect -3044 14488 -3028 14552
rect -2964 14488 -2948 14552
rect -3044 14472 -2948 14488
rect -3044 14408 -3028 14472
rect -2964 14408 -2948 14472
rect -3044 14392 -2948 14408
rect -3044 14328 -3028 14392
rect -2964 14328 -2948 14392
rect -3044 14312 -2948 14328
rect -3044 14248 -3028 14312
rect -2964 14248 -2948 14312
rect -3044 14232 -2948 14248
rect -4456 14132 -4360 14168
rect -3044 14168 -3028 14232
rect -2964 14168 -2948 14232
rect -2625 14912 -1903 14921
rect -2625 14208 -2616 14912
rect -1912 14208 -1903 14912
rect -2625 14199 -1903 14208
rect -1632 14888 -1616 14952
rect -1552 14888 -1536 14952
rect -220 14952 -124 14988
rect -1632 14872 -1536 14888
rect -1632 14808 -1616 14872
rect -1552 14808 -1536 14872
rect -1632 14792 -1536 14808
rect -1632 14728 -1616 14792
rect -1552 14728 -1536 14792
rect -1632 14712 -1536 14728
rect -1632 14648 -1616 14712
rect -1552 14648 -1536 14712
rect -1632 14632 -1536 14648
rect -1632 14568 -1616 14632
rect -1552 14568 -1536 14632
rect -1632 14552 -1536 14568
rect -1632 14488 -1616 14552
rect -1552 14488 -1536 14552
rect -1632 14472 -1536 14488
rect -1632 14408 -1616 14472
rect -1552 14408 -1536 14472
rect -1632 14392 -1536 14408
rect -1632 14328 -1616 14392
rect -1552 14328 -1536 14392
rect -1632 14312 -1536 14328
rect -1632 14248 -1616 14312
rect -1552 14248 -1536 14312
rect -1632 14232 -1536 14248
rect -3044 14132 -2948 14168
rect -1632 14168 -1616 14232
rect -1552 14168 -1536 14232
rect -1213 14912 -491 14921
rect -1213 14208 -1204 14912
rect -500 14208 -491 14912
rect -1213 14199 -491 14208
rect -220 14888 -204 14952
rect -140 14888 -124 14952
rect 1192 14952 1288 14988
rect -220 14872 -124 14888
rect -220 14808 -204 14872
rect -140 14808 -124 14872
rect -220 14792 -124 14808
rect -220 14728 -204 14792
rect -140 14728 -124 14792
rect -220 14712 -124 14728
rect -220 14648 -204 14712
rect -140 14648 -124 14712
rect -220 14632 -124 14648
rect -220 14568 -204 14632
rect -140 14568 -124 14632
rect -220 14552 -124 14568
rect -220 14488 -204 14552
rect -140 14488 -124 14552
rect -220 14472 -124 14488
rect -220 14408 -204 14472
rect -140 14408 -124 14472
rect -220 14392 -124 14408
rect -220 14328 -204 14392
rect -140 14328 -124 14392
rect -220 14312 -124 14328
rect -220 14248 -204 14312
rect -140 14248 -124 14312
rect -220 14232 -124 14248
rect -1632 14132 -1536 14168
rect -220 14168 -204 14232
rect -140 14168 -124 14232
rect 199 14912 921 14921
rect 199 14208 208 14912
rect 912 14208 921 14912
rect 199 14199 921 14208
rect 1192 14888 1208 14952
rect 1272 14888 1288 14952
rect 2604 14952 2700 14988
rect 1192 14872 1288 14888
rect 1192 14808 1208 14872
rect 1272 14808 1288 14872
rect 1192 14792 1288 14808
rect 1192 14728 1208 14792
rect 1272 14728 1288 14792
rect 1192 14712 1288 14728
rect 1192 14648 1208 14712
rect 1272 14648 1288 14712
rect 1192 14632 1288 14648
rect 1192 14568 1208 14632
rect 1272 14568 1288 14632
rect 1192 14552 1288 14568
rect 1192 14488 1208 14552
rect 1272 14488 1288 14552
rect 1192 14472 1288 14488
rect 1192 14408 1208 14472
rect 1272 14408 1288 14472
rect 1192 14392 1288 14408
rect 1192 14328 1208 14392
rect 1272 14328 1288 14392
rect 1192 14312 1288 14328
rect 1192 14248 1208 14312
rect 1272 14248 1288 14312
rect 1192 14232 1288 14248
rect -220 14132 -124 14168
rect 1192 14168 1208 14232
rect 1272 14168 1288 14232
rect 1611 14912 2333 14921
rect 1611 14208 1620 14912
rect 2324 14208 2333 14912
rect 1611 14199 2333 14208
rect 2604 14888 2620 14952
rect 2684 14888 2700 14952
rect 4016 14952 4112 14988
rect 2604 14872 2700 14888
rect 2604 14808 2620 14872
rect 2684 14808 2700 14872
rect 2604 14792 2700 14808
rect 2604 14728 2620 14792
rect 2684 14728 2700 14792
rect 2604 14712 2700 14728
rect 2604 14648 2620 14712
rect 2684 14648 2700 14712
rect 2604 14632 2700 14648
rect 2604 14568 2620 14632
rect 2684 14568 2700 14632
rect 2604 14552 2700 14568
rect 2604 14488 2620 14552
rect 2684 14488 2700 14552
rect 2604 14472 2700 14488
rect 2604 14408 2620 14472
rect 2684 14408 2700 14472
rect 2604 14392 2700 14408
rect 2604 14328 2620 14392
rect 2684 14328 2700 14392
rect 2604 14312 2700 14328
rect 2604 14248 2620 14312
rect 2684 14248 2700 14312
rect 2604 14232 2700 14248
rect 1192 14132 1288 14168
rect 2604 14168 2620 14232
rect 2684 14168 2700 14232
rect 3023 14912 3745 14921
rect 3023 14208 3032 14912
rect 3736 14208 3745 14912
rect 3023 14199 3745 14208
rect 4016 14888 4032 14952
rect 4096 14888 4112 14952
rect 5428 14952 5524 14988
rect 4016 14872 4112 14888
rect 4016 14808 4032 14872
rect 4096 14808 4112 14872
rect 4016 14792 4112 14808
rect 4016 14728 4032 14792
rect 4096 14728 4112 14792
rect 4016 14712 4112 14728
rect 4016 14648 4032 14712
rect 4096 14648 4112 14712
rect 4016 14632 4112 14648
rect 4016 14568 4032 14632
rect 4096 14568 4112 14632
rect 4016 14552 4112 14568
rect 4016 14488 4032 14552
rect 4096 14488 4112 14552
rect 4016 14472 4112 14488
rect 4016 14408 4032 14472
rect 4096 14408 4112 14472
rect 4016 14392 4112 14408
rect 4016 14328 4032 14392
rect 4096 14328 4112 14392
rect 4016 14312 4112 14328
rect 4016 14248 4032 14312
rect 4096 14248 4112 14312
rect 4016 14232 4112 14248
rect 2604 14132 2700 14168
rect 4016 14168 4032 14232
rect 4096 14168 4112 14232
rect 4435 14912 5157 14921
rect 4435 14208 4444 14912
rect 5148 14208 5157 14912
rect 4435 14199 5157 14208
rect 5428 14888 5444 14952
rect 5508 14888 5524 14952
rect 6840 14952 6936 14988
rect 5428 14872 5524 14888
rect 5428 14808 5444 14872
rect 5508 14808 5524 14872
rect 5428 14792 5524 14808
rect 5428 14728 5444 14792
rect 5508 14728 5524 14792
rect 5428 14712 5524 14728
rect 5428 14648 5444 14712
rect 5508 14648 5524 14712
rect 5428 14632 5524 14648
rect 5428 14568 5444 14632
rect 5508 14568 5524 14632
rect 5428 14552 5524 14568
rect 5428 14488 5444 14552
rect 5508 14488 5524 14552
rect 5428 14472 5524 14488
rect 5428 14408 5444 14472
rect 5508 14408 5524 14472
rect 5428 14392 5524 14408
rect 5428 14328 5444 14392
rect 5508 14328 5524 14392
rect 5428 14312 5524 14328
rect 5428 14248 5444 14312
rect 5508 14248 5524 14312
rect 5428 14232 5524 14248
rect 4016 14132 4112 14168
rect 5428 14168 5444 14232
rect 5508 14168 5524 14232
rect 5847 14912 6569 14921
rect 5847 14208 5856 14912
rect 6560 14208 6569 14912
rect 5847 14199 6569 14208
rect 6840 14888 6856 14952
rect 6920 14888 6936 14952
rect 8252 14952 8348 14988
rect 6840 14872 6936 14888
rect 6840 14808 6856 14872
rect 6920 14808 6936 14872
rect 6840 14792 6936 14808
rect 6840 14728 6856 14792
rect 6920 14728 6936 14792
rect 6840 14712 6936 14728
rect 6840 14648 6856 14712
rect 6920 14648 6936 14712
rect 6840 14632 6936 14648
rect 6840 14568 6856 14632
rect 6920 14568 6936 14632
rect 6840 14552 6936 14568
rect 6840 14488 6856 14552
rect 6920 14488 6936 14552
rect 6840 14472 6936 14488
rect 6840 14408 6856 14472
rect 6920 14408 6936 14472
rect 6840 14392 6936 14408
rect 6840 14328 6856 14392
rect 6920 14328 6936 14392
rect 6840 14312 6936 14328
rect 6840 14248 6856 14312
rect 6920 14248 6936 14312
rect 6840 14232 6936 14248
rect 5428 14132 5524 14168
rect 6840 14168 6856 14232
rect 6920 14168 6936 14232
rect 7259 14912 7981 14921
rect 7259 14208 7268 14912
rect 7972 14208 7981 14912
rect 7259 14199 7981 14208
rect 8252 14888 8268 14952
rect 8332 14888 8348 14952
rect 9664 14952 9760 14988
rect 8252 14872 8348 14888
rect 8252 14808 8268 14872
rect 8332 14808 8348 14872
rect 8252 14792 8348 14808
rect 8252 14728 8268 14792
rect 8332 14728 8348 14792
rect 8252 14712 8348 14728
rect 8252 14648 8268 14712
rect 8332 14648 8348 14712
rect 8252 14632 8348 14648
rect 8252 14568 8268 14632
rect 8332 14568 8348 14632
rect 8252 14552 8348 14568
rect 8252 14488 8268 14552
rect 8332 14488 8348 14552
rect 8252 14472 8348 14488
rect 8252 14408 8268 14472
rect 8332 14408 8348 14472
rect 8252 14392 8348 14408
rect 8252 14328 8268 14392
rect 8332 14328 8348 14392
rect 8252 14312 8348 14328
rect 8252 14248 8268 14312
rect 8332 14248 8348 14312
rect 8252 14232 8348 14248
rect 6840 14132 6936 14168
rect 8252 14168 8268 14232
rect 8332 14168 8348 14232
rect 8671 14912 9393 14921
rect 8671 14208 8680 14912
rect 9384 14208 9393 14912
rect 8671 14199 9393 14208
rect 9664 14888 9680 14952
rect 9744 14888 9760 14952
rect 11076 14952 11172 14988
rect 9664 14872 9760 14888
rect 9664 14808 9680 14872
rect 9744 14808 9760 14872
rect 9664 14792 9760 14808
rect 9664 14728 9680 14792
rect 9744 14728 9760 14792
rect 9664 14712 9760 14728
rect 9664 14648 9680 14712
rect 9744 14648 9760 14712
rect 9664 14632 9760 14648
rect 9664 14568 9680 14632
rect 9744 14568 9760 14632
rect 9664 14552 9760 14568
rect 9664 14488 9680 14552
rect 9744 14488 9760 14552
rect 9664 14472 9760 14488
rect 9664 14408 9680 14472
rect 9744 14408 9760 14472
rect 9664 14392 9760 14408
rect 9664 14328 9680 14392
rect 9744 14328 9760 14392
rect 9664 14312 9760 14328
rect 9664 14248 9680 14312
rect 9744 14248 9760 14312
rect 9664 14232 9760 14248
rect 8252 14132 8348 14168
rect 9664 14168 9680 14232
rect 9744 14168 9760 14232
rect 10083 14912 10805 14921
rect 10083 14208 10092 14912
rect 10796 14208 10805 14912
rect 10083 14199 10805 14208
rect 11076 14888 11092 14952
rect 11156 14888 11172 14952
rect 12488 14952 12584 14988
rect 11076 14872 11172 14888
rect 11076 14808 11092 14872
rect 11156 14808 11172 14872
rect 11076 14792 11172 14808
rect 11076 14728 11092 14792
rect 11156 14728 11172 14792
rect 11076 14712 11172 14728
rect 11076 14648 11092 14712
rect 11156 14648 11172 14712
rect 11076 14632 11172 14648
rect 11076 14568 11092 14632
rect 11156 14568 11172 14632
rect 11076 14552 11172 14568
rect 11076 14488 11092 14552
rect 11156 14488 11172 14552
rect 11076 14472 11172 14488
rect 11076 14408 11092 14472
rect 11156 14408 11172 14472
rect 11076 14392 11172 14408
rect 11076 14328 11092 14392
rect 11156 14328 11172 14392
rect 11076 14312 11172 14328
rect 11076 14248 11092 14312
rect 11156 14248 11172 14312
rect 11076 14232 11172 14248
rect 9664 14132 9760 14168
rect 11076 14168 11092 14232
rect 11156 14168 11172 14232
rect 11495 14912 12217 14921
rect 11495 14208 11504 14912
rect 12208 14208 12217 14912
rect 11495 14199 12217 14208
rect 12488 14888 12504 14952
rect 12568 14888 12584 14952
rect 13900 14952 13996 14988
rect 12488 14872 12584 14888
rect 12488 14808 12504 14872
rect 12568 14808 12584 14872
rect 12488 14792 12584 14808
rect 12488 14728 12504 14792
rect 12568 14728 12584 14792
rect 12488 14712 12584 14728
rect 12488 14648 12504 14712
rect 12568 14648 12584 14712
rect 12488 14632 12584 14648
rect 12488 14568 12504 14632
rect 12568 14568 12584 14632
rect 12488 14552 12584 14568
rect 12488 14488 12504 14552
rect 12568 14488 12584 14552
rect 12488 14472 12584 14488
rect 12488 14408 12504 14472
rect 12568 14408 12584 14472
rect 12488 14392 12584 14408
rect 12488 14328 12504 14392
rect 12568 14328 12584 14392
rect 12488 14312 12584 14328
rect 12488 14248 12504 14312
rect 12568 14248 12584 14312
rect 12488 14232 12584 14248
rect 11076 14132 11172 14168
rect 12488 14168 12504 14232
rect 12568 14168 12584 14232
rect 12907 14912 13629 14921
rect 12907 14208 12916 14912
rect 13620 14208 13629 14912
rect 12907 14199 13629 14208
rect 13900 14888 13916 14952
rect 13980 14888 13996 14952
rect 15312 14952 15408 14988
rect 13900 14872 13996 14888
rect 13900 14808 13916 14872
rect 13980 14808 13996 14872
rect 13900 14792 13996 14808
rect 13900 14728 13916 14792
rect 13980 14728 13996 14792
rect 13900 14712 13996 14728
rect 13900 14648 13916 14712
rect 13980 14648 13996 14712
rect 13900 14632 13996 14648
rect 13900 14568 13916 14632
rect 13980 14568 13996 14632
rect 13900 14552 13996 14568
rect 13900 14488 13916 14552
rect 13980 14488 13996 14552
rect 13900 14472 13996 14488
rect 13900 14408 13916 14472
rect 13980 14408 13996 14472
rect 13900 14392 13996 14408
rect 13900 14328 13916 14392
rect 13980 14328 13996 14392
rect 13900 14312 13996 14328
rect 13900 14248 13916 14312
rect 13980 14248 13996 14312
rect 13900 14232 13996 14248
rect 12488 14132 12584 14168
rect 13900 14168 13916 14232
rect 13980 14168 13996 14232
rect 14319 14912 15041 14921
rect 14319 14208 14328 14912
rect 15032 14208 15041 14912
rect 14319 14199 15041 14208
rect 15312 14888 15328 14952
rect 15392 14888 15408 14952
rect 16724 14952 16820 14988
rect 15312 14872 15408 14888
rect 15312 14808 15328 14872
rect 15392 14808 15408 14872
rect 15312 14792 15408 14808
rect 15312 14728 15328 14792
rect 15392 14728 15408 14792
rect 15312 14712 15408 14728
rect 15312 14648 15328 14712
rect 15392 14648 15408 14712
rect 15312 14632 15408 14648
rect 15312 14568 15328 14632
rect 15392 14568 15408 14632
rect 15312 14552 15408 14568
rect 15312 14488 15328 14552
rect 15392 14488 15408 14552
rect 15312 14472 15408 14488
rect 15312 14408 15328 14472
rect 15392 14408 15408 14472
rect 15312 14392 15408 14408
rect 15312 14328 15328 14392
rect 15392 14328 15408 14392
rect 15312 14312 15408 14328
rect 15312 14248 15328 14312
rect 15392 14248 15408 14312
rect 15312 14232 15408 14248
rect 13900 14132 13996 14168
rect 15312 14168 15328 14232
rect 15392 14168 15408 14232
rect 15731 14912 16453 14921
rect 15731 14208 15740 14912
rect 16444 14208 16453 14912
rect 15731 14199 16453 14208
rect 16724 14888 16740 14952
rect 16804 14888 16820 14952
rect 18136 14952 18232 14988
rect 16724 14872 16820 14888
rect 16724 14808 16740 14872
rect 16804 14808 16820 14872
rect 16724 14792 16820 14808
rect 16724 14728 16740 14792
rect 16804 14728 16820 14792
rect 16724 14712 16820 14728
rect 16724 14648 16740 14712
rect 16804 14648 16820 14712
rect 16724 14632 16820 14648
rect 16724 14568 16740 14632
rect 16804 14568 16820 14632
rect 16724 14552 16820 14568
rect 16724 14488 16740 14552
rect 16804 14488 16820 14552
rect 16724 14472 16820 14488
rect 16724 14408 16740 14472
rect 16804 14408 16820 14472
rect 16724 14392 16820 14408
rect 16724 14328 16740 14392
rect 16804 14328 16820 14392
rect 16724 14312 16820 14328
rect 16724 14248 16740 14312
rect 16804 14248 16820 14312
rect 16724 14232 16820 14248
rect 15312 14132 15408 14168
rect 16724 14168 16740 14232
rect 16804 14168 16820 14232
rect 17143 14912 17865 14921
rect 17143 14208 17152 14912
rect 17856 14208 17865 14912
rect 17143 14199 17865 14208
rect 18136 14888 18152 14952
rect 18216 14888 18232 14952
rect 19548 14952 19644 14988
rect 18136 14872 18232 14888
rect 18136 14808 18152 14872
rect 18216 14808 18232 14872
rect 18136 14792 18232 14808
rect 18136 14728 18152 14792
rect 18216 14728 18232 14792
rect 18136 14712 18232 14728
rect 18136 14648 18152 14712
rect 18216 14648 18232 14712
rect 18136 14632 18232 14648
rect 18136 14568 18152 14632
rect 18216 14568 18232 14632
rect 18136 14552 18232 14568
rect 18136 14488 18152 14552
rect 18216 14488 18232 14552
rect 18136 14472 18232 14488
rect 18136 14408 18152 14472
rect 18216 14408 18232 14472
rect 18136 14392 18232 14408
rect 18136 14328 18152 14392
rect 18216 14328 18232 14392
rect 18136 14312 18232 14328
rect 18136 14248 18152 14312
rect 18216 14248 18232 14312
rect 18136 14232 18232 14248
rect 16724 14132 16820 14168
rect 18136 14168 18152 14232
rect 18216 14168 18232 14232
rect 18555 14912 19277 14921
rect 18555 14208 18564 14912
rect 19268 14208 19277 14912
rect 18555 14199 19277 14208
rect 19548 14888 19564 14952
rect 19628 14888 19644 14952
rect 20960 14952 21056 14988
rect 19548 14872 19644 14888
rect 19548 14808 19564 14872
rect 19628 14808 19644 14872
rect 19548 14792 19644 14808
rect 19548 14728 19564 14792
rect 19628 14728 19644 14792
rect 19548 14712 19644 14728
rect 19548 14648 19564 14712
rect 19628 14648 19644 14712
rect 19548 14632 19644 14648
rect 19548 14568 19564 14632
rect 19628 14568 19644 14632
rect 19548 14552 19644 14568
rect 19548 14488 19564 14552
rect 19628 14488 19644 14552
rect 19548 14472 19644 14488
rect 19548 14408 19564 14472
rect 19628 14408 19644 14472
rect 19548 14392 19644 14408
rect 19548 14328 19564 14392
rect 19628 14328 19644 14392
rect 19548 14312 19644 14328
rect 19548 14248 19564 14312
rect 19628 14248 19644 14312
rect 19548 14232 19644 14248
rect 18136 14132 18232 14168
rect 19548 14168 19564 14232
rect 19628 14168 19644 14232
rect 19967 14912 20689 14921
rect 19967 14208 19976 14912
rect 20680 14208 20689 14912
rect 19967 14199 20689 14208
rect 20960 14888 20976 14952
rect 21040 14888 21056 14952
rect 22372 14952 22468 14988
rect 20960 14872 21056 14888
rect 20960 14808 20976 14872
rect 21040 14808 21056 14872
rect 20960 14792 21056 14808
rect 20960 14728 20976 14792
rect 21040 14728 21056 14792
rect 20960 14712 21056 14728
rect 20960 14648 20976 14712
rect 21040 14648 21056 14712
rect 20960 14632 21056 14648
rect 20960 14568 20976 14632
rect 21040 14568 21056 14632
rect 20960 14552 21056 14568
rect 20960 14488 20976 14552
rect 21040 14488 21056 14552
rect 20960 14472 21056 14488
rect 20960 14408 20976 14472
rect 21040 14408 21056 14472
rect 20960 14392 21056 14408
rect 20960 14328 20976 14392
rect 21040 14328 21056 14392
rect 20960 14312 21056 14328
rect 20960 14248 20976 14312
rect 21040 14248 21056 14312
rect 20960 14232 21056 14248
rect 19548 14132 19644 14168
rect 20960 14168 20976 14232
rect 21040 14168 21056 14232
rect 21379 14912 22101 14921
rect 21379 14208 21388 14912
rect 22092 14208 22101 14912
rect 21379 14199 22101 14208
rect 22372 14888 22388 14952
rect 22452 14888 22468 14952
rect 23784 14952 23880 14988
rect 22372 14872 22468 14888
rect 22372 14808 22388 14872
rect 22452 14808 22468 14872
rect 22372 14792 22468 14808
rect 22372 14728 22388 14792
rect 22452 14728 22468 14792
rect 22372 14712 22468 14728
rect 22372 14648 22388 14712
rect 22452 14648 22468 14712
rect 22372 14632 22468 14648
rect 22372 14568 22388 14632
rect 22452 14568 22468 14632
rect 22372 14552 22468 14568
rect 22372 14488 22388 14552
rect 22452 14488 22468 14552
rect 22372 14472 22468 14488
rect 22372 14408 22388 14472
rect 22452 14408 22468 14472
rect 22372 14392 22468 14408
rect 22372 14328 22388 14392
rect 22452 14328 22468 14392
rect 22372 14312 22468 14328
rect 22372 14248 22388 14312
rect 22452 14248 22468 14312
rect 22372 14232 22468 14248
rect 20960 14132 21056 14168
rect 22372 14168 22388 14232
rect 22452 14168 22468 14232
rect 22791 14912 23513 14921
rect 22791 14208 22800 14912
rect 23504 14208 23513 14912
rect 22791 14199 23513 14208
rect 23784 14888 23800 14952
rect 23864 14888 23880 14952
rect 23784 14872 23880 14888
rect 23784 14808 23800 14872
rect 23864 14808 23880 14872
rect 23784 14792 23880 14808
rect 23784 14728 23800 14792
rect 23864 14728 23880 14792
rect 23784 14712 23880 14728
rect 23784 14648 23800 14712
rect 23864 14648 23880 14712
rect 23784 14632 23880 14648
rect 23784 14568 23800 14632
rect 23864 14568 23880 14632
rect 23784 14552 23880 14568
rect 23784 14488 23800 14552
rect 23864 14488 23880 14552
rect 23784 14472 23880 14488
rect 23784 14408 23800 14472
rect 23864 14408 23880 14472
rect 23784 14392 23880 14408
rect 23784 14328 23800 14392
rect 23864 14328 23880 14392
rect 23784 14312 23880 14328
rect 23784 14248 23800 14312
rect 23864 14248 23880 14312
rect 23784 14232 23880 14248
rect 22372 14132 22468 14168
rect 23784 14168 23800 14232
rect 23864 14168 23880 14232
rect 23784 14132 23880 14168
rect -22812 13832 -22716 13868
rect -23805 13792 -23083 13801
rect -23805 13088 -23796 13792
rect -23092 13088 -23083 13792
rect -23805 13079 -23083 13088
rect -22812 13768 -22796 13832
rect -22732 13768 -22716 13832
rect -21400 13832 -21304 13868
rect -22812 13752 -22716 13768
rect -22812 13688 -22796 13752
rect -22732 13688 -22716 13752
rect -22812 13672 -22716 13688
rect -22812 13608 -22796 13672
rect -22732 13608 -22716 13672
rect -22812 13592 -22716 13608
rect -22812 13528 -22796 13592
rect -22732 13528 -22716 13592
rect -22812 13512 -22716 13528
rect -22812 13448 -22796 13512
rect -22732 13448 -22716 13512
rect -22812 13432 -22716 13448
rect -22812 13368 -22796 13432
rect -22732 13368 -22716 13432
rect -22812 13352 -22716 13368
rect -22812 13288 -22796 13352
rect -22732 13288 -22716 13352
rect -22812 13272 -22716 13288
rect -22812 13208 -22796 13272
rect -22732 13208 -22716 13272
rect -22812 13192 -22716 13208
rect -22812 13128 -22796 13192
rect -22732 13128 -22716 13192
rect -22812 13112 -22716 13128
rect -22812 13048 -22796 13112
rect -22732 13048 -22716 13112
rect -22393 13792 -21671 13801
rect -22393 13088 -22384 13792
rect -21680 13088 -21671 13792
rect -22393 13079 -21671 13088
rect -21400 13768 -21384 13832
rect -21320 13768 -21304 13832
rect -19988 13832 -19892 13868
rect -21400 13752 -21304 13768
rect -21400 13688 -21384 13752
rect -21320 13688 -21304 13752
rect -21400 13672 -21304 13688
rect -21400 13608 -21384 13672
rect -21320 13608 -21304 13672
rect -21400 13592 -21304 13608
rect -21400 13528 -21384 13592
rect -21320 13528 -21304 13592
rect -21400 13512 -21304 13528
rect -21400 13448 -21384 13512
rect -21320 13448 -21304 13512
rect -21400 13432 -21304 13448
rect -21400 13368 -21384 13432
rect -21320 13368 -21304 13432
rect -21400 13352 -21304 13368
rect -21400 13288 -21384 13352
rect -21320 13288 -21304 13352
rect -21400 13272 -21304 13288
rect -21400 13208 -21384 13272
rect -21320 13208 -21304 13272
rect -21400 13192 -21304 13208
rect -21400 13128 -21384 13192
rect -21320 13128 -21304 13192
rect -21400 13112 -21304 13128
rect -22812 13012 -22716 13048
rect -21400 13048 -21384 13112
rect -21320 13048 -21304 13112
rect -20981 13792 -20259 13801
rect -20981 13088 -20972 13792
rect -20268 13088 -20259 13792
rect -20981 13079 -20259 13088
rect -19988 13768 -19972 13832
rect -19908 13768 -19892 13832
rect -18576 13832 -18480 13868
rect -19988 13752 -19892 13768
rect -19988 13688 -19972 13752
rect -19908 13688 -19892 13752
rect -19988 13672 -19892 13688
rect -19988 13608 -19972 13672
rect -19908 13608 -19892 13672
rect -19988 13592 -19892 13608
rect -19988 13528 -19972 13592
rect -19908 13528 -19892 13592
rect -19988 13512 -19892 13528
rect -19988 13448 -19972 13512
rect -19908 13448 -19892 13512
rect -19988 13432 -19892 13448
rect -19988 13368 -19972 13432
rect -19908 13368 -19892 13432
rect -19988 13352 -19892 13368
rect -19988 13288 -19972 13352
rect -19908 13288 -19892 13352
rect -19988 13272 -19892 13288
rect -19988 13208 -19972 13272
rect -19908 13208 -19892 13272
rect -19988 13192 -19892 13208
rect -19988 13128 -19972 13192
rect -19908 13128 -19892 13192
rect -19988 13112 -19892 13128
rect -21400 13012 -21304 13048
rect -19988 13048 -19972 13112
rect -19908 13048 -19892 13112
rect -19569 13792 -18847 13801
rect -19569 13088 -19560 13792
rect -18856 13088 -18847 13792
rect -19569 13079 -18847 13088
rect -18576 13768 -18560 13832
rect -18496 13768 -18480 13832
rect -17164 13832 -17068 13868
rect -18576 13752 -18480 13768
rect -18576 13688 -18560 13752
rect -18496 13688 -18480 13752
rect -18576 13672 -18480 13688
rect -18576 13608 -18560 13672
rect -18496 13608 -18480 13672
rect -18576 13592 -18480 13608
rect -18576 13528 -18560 13592
rect -18496 13528 -18480 13592
rect -18576 13512 -18480 13528
rect -18576 13448 -18560 13512
rect -18496 13448 -18480 13512
rect -18576 13432 -18480 13448
rect -18576 13368 -18560 13432
rect -18496 13368 -18480 13432
rect -18576 13352 -18480 13368
rect -18576 13288 -18560 13352
rect -18496 13288 -18480 13352
rect -18576 13272 -18480 13288
rect -18576 13208 -18560 13272
rect -18496 13208 -18480 13272
rect -18576 13192 -18480 13208
rect -18576 13128 -18560 13192
rect -18496 13128 -18480 13192
rect -18576 13112 -18480 13128
rect -19988 13012 -19892 13048
rect -18576 13048 -18560 13112
rect -18496 13048 -18480 13112
rect -18157 13792 -17435 13801
rect -18157 13088 -18148 13792
rect -17444 13088 -17435 13792
rect -18157 13079 -17435 13088
rect -17164 13768 -17148 13832
rect -17084 13768 -17068 13832
rect -15752 13832 -15656 13868
rect -17164 13752 -17068 13768
rect -17164 13688 -17148 13752
rect -17084 13688 -17068 13752
rect -17164 13672 -17068 13688
rect -17164 13608 -17148 13672
rect -17084 13608 -17068 13672
rect -17164 13592 -17068 13608
rect -17164 13528 -17148 13592
rect -17084 13528 -17068 13592
rect -17164 13512 -17068 13528
rect -17164 13448 -17148 13512
rect -17084 13448 -17068 13512
rect -17164 13432 -17068 13448
rect -17164 13368 -17148 13432
rect -17084 13368 -17068 13432
rect -17164 13352 -17068 13368
rect -17164 13288 -17148 13352
rect -17084 13288 -17068 13352
rect -17164 13272 -17068 13288
rect -17164 13208 -17148 13272
rect -17084 13208 -17068 13272
rect -17164 13192 -17068 13208
rect -17164 13128 -17148 13192
rect -17084 13128 -17068 13192
rect -17164 13112 -17068 13128
rect -18576 13012 -18480 13048
rect -17164 13048 -17148 13112
rect -17084 13048 -17068 13112
rect -16745 13792 -16023 13801
rect -16745 13088 -16736 13792
rect -16032 13088 -16023 13792
rect -16745 13079 -16023 13088
rect -15752 13768 -15736 13832
rect -15672 13768 -15656 13832
rect -14340 13832 -14244 13868
rect -15752 13752 -15656 13768
rect -15752 13688 -15736 13752
rect -15672 13688 -15656 13752
rect -15752 13672 -15656 13688
rect -15752 13608 -15736 13672
rect -15672 13608 -15656 13672
rect -15752 13592 -15656 13608
rect -15752 13528 -15736 13592
rect -15672 13528 -15656 13592
rect -15752 13512 -15656 13528
rect -15752 13448 -15736 13512
rect -15672 13448 -15656 13512
rect -15752 13432 -15656 13448
rect -15752 13368 -15736 13432
rect -15672 13368 -15656 13432
rect -15752 13352 -15656 13368
rect -15752 13288 -15736 13352
rect -15672 13288 -15656 13352
rect -15752 13272 -15656 13288
rect -15752 13208 -15736 13272
rect -15672 13208 -15656 13272
rect -15752 13192 -15656 13208
rect -15752 13128 -15736 13192
rect -15672 13128 -15656 13192
rect -15752 13112 -15656 13128
rect -17164 13012 -17068 13048
rect -15752 13048 -15736 13112
rect -15672 13048 -15656 13112
rect -15333 13792 -14611 13801
rect -15333 13088 -15324 13792
rect -14620 13088 -14611 13792
rect -15333 13079 -14611 13088
rect -14340 13768 -14324 13832
rect -14260 13768 -14244 13832
rect -12928 13832 -12832 13868
rect -14340 13752 -14244 13768
rect -14340 13688 -14324 13752
rect -14260 13688 -14244 13752
rect -14340 13672 -14244 13688
rect -14340 13608 -14324 13672
rect -14260 13608 -14244 13672
rect -14340 13592 -14244 13608
rect -14340 13528 -14324 13592
rect -14260 13528 -14244 13592
rect -14340 13512 -14244 13528
rect -14340 13448 -14324 13512
rect -14260 13448 -14244 13512
rect -14340 13432 -14244 13448
rect -14340 13368 -14324 13432
rect -14260 13368 -14244 13432
rect -14340 13352 -14244 13368
rect -14340 13288 -14324 13352
rect -14260 13288 -14244 13352
rect -14340 13272 -14244 13288
rect -14340 13208 -14324 13272
rect -14260 13208 -14244 13272
rect -14340 13192 -14244 13208
rect -14340 13128 -14324 13192
rect -14260 13128 -14244 13192
rect -14340 13112 -14244 13128
rect -15752 13012 -15656 13048
rect -14340 13048 -14324 13112
rect -14260 13048 -14244 13112
rect -13921 13792 -13199 13801
rect -13921 13088 -13912 13792
rect -13208 13088 -13199 13792
rect -13921 13079 -13199 13088
rect -12928 13768 -12912 13832
rect -12848 13768 -12832 13832
rect -11516 13832 -11420 13868
rect -12928 13752 -12832 13768
rect -12928 13688 -12912 13752
rect -12848 13688 -12832 13752
rect -12928 13672 -12832 13688
rect -12928 13608 -12912 13672
rect -12848 13608 -12832 13672
rect -12928 13592 -12832 13608
rect -12928 13528 -12912 13592
rect -12848 13528 -12832 13592
rect -12928 13512 -12832 13528
rect -12928 13448 -12912 13512
rect -12848 13448 -12832 13512
rect -12928 13432 -12832 13448
rect -12928 13368 -12912 13432
rect -12848 13368 -12832 13432
rect -12928 13352 -12832 13368
rect -12928 13288 -12912 13352
rect -12848 13288 -12832 13352
rect -12928 13272 -12832 13288
rect -12928 13208 -12912 13272
rect -12848 13208 -12832 13272
rect -12928 13192 -12832 13208
rect -12928 13128 -12912 13192
rect -12848 13128 -12832 13192
rect -12928 13112 -12832 13128
rect -14340 13012 -14244 13048
rect -12928 13048 -12912 13112
rect -12848 13048 -12832 13112
rect -12509 13792 -11787 13801
rect -12509 13088 -12500 13792
rect -11796 13088 -11787 13792
rect -12509 13079 -11787 13088
rect -11516 13768 -11500 13832
rect -11436 13768 -11420 13832
rect -10104 13832 -10008 13868
rect -11516 13752 -11420 13768
rect -11516 13688 -11500 13752
rect -11436 13688 -11420 13752
rect -11516 13672 -11420 13688
rect -11516 13608 -11500 13672
rect -11436 13608 -11420 13672
rect -11516 13592 -11420 13608
rect -11516 13528 -11500 13592
rect -11436 13528 -11420 13592
rect -11516 13512 -11420 13528
rect -11516 13448 -11500 13512
rect -11436 13448 -11420 13512
rect -11516 13432 -11420 13448
rect -11516 13368 -11500 13432
rect -11436 13368 -11420 13432
rect -11516 13352 -11420 13368
rect -11516 13288 -11500 13352
rect -11436 13288 -11420 13352
rect -11516 13272 -11420 13288
rect -11516 13208 -11500 13272
rect -11436 13208 -11420 13272
rect -11516 13192 -11420 13208
rect -11516 13128 -11500 13192
rect -11436 13128 -11420 13192
rect -11516 13112 -11420 13128
rect -12928 13012 -12832 13048
rect -11516 13048 -11500 13112
rect -11436 13048 -11420 13112
rect -11097 13792 -10375 13801
rect -11097 13088 -11088 13792
rect -10384 13088 -10375 13792
rect -11097 13079 -10375 13088
rect -10104 13768 -10088 13832
rect -10024 13768 -10008 13832
rect -8692 13832 -8596 13868
rect -10104 13752 -10008 13768
rect -10104 13688 -10088 13752
rect -10024 13688 -10008 13752
rect -10104 13672 -10008 13688
rect -10104 13608 -10088 13672
rect -10024 13608 -10008 13672
rect -10104 13592 -10008 13608
rect -10104 13528 -10088 13592
rect -10024 13528 -10008 13592
rect -10104 13512 -10008 13528
rect -10104 13448 -10088 13512
rect -10024 13448 -10008 13512
rect -10104 13432 -10008 13448
rect -10104 13368 -10088 13432
rect -10024 13368 -10008 13432
rect -10104 13352 -10008 13368
rect -10104 13288 -10088 13352
rect -10024 13288 -10008 13352
rect -10104 13272 -10008 13288
rect -10104 13208 -10088 13272
rect -10024 13208 -10008 13272
rect -10104 13192 -10008 13208
rect -10104 13128 -10088 13192
rect -10024 13128 -10008 13192
rect -10104 13112 -10008 13128
rect -11516 13012 -11420 13048
rect -10104 13048 -10088 13112
rect -10024 13048 -10008 13112
rect -9685 13792 -8963 13801
rect -9685 13088 -9676 13792
rect -8972 13088 -8963 13792
rect -9685 13079 -8963 13088
rect -8692 13768 -8676 13832
rect -8612 13768 -8596 13832
rect -7280 13832 -7184 13868
rect -8692 13752 -8596 13768
rect -8692 13688 -8676 13752
rect -8612 13688 -8596 13752
rect -8692 13672 -8596 13688
rect -8692 13608 -8676 13672
rect -8612 13608 -8596 13672
rect -8692 13592 -8596 13608
rect -8692 13528 -8676 13592
rect -8612 13528 -8596 13592
rect -8692 13512 -8596 13528
rect -8692 13448 -8676 13512
rect -8612 13448 -8596 13512
rect -8692 13432 -8596 13448
rect -8692 13368 -8676 13432
rect -8612 13368 -8596 13432
rect -8692 13352 -8596 13368
rect -8692 13288 -8676 13352
rect -8612 13288 -8596 13352
rect -8692 13272 -8596 13288
rect -8692 13208 -8676 13272
rect -8612 13208 -8596 13272
rect -8692 13192 -8596 13208
rect -8692 13128 -8676 13192
rect -8612 13128 -8596 13192
rect -8692 13112 -8596 13128
rect -10104 13012 -10008 13048
rect -8692 13048 -8676 13112
rect -8612 13048 -8596 13112
rect -8273 13792 -7551 13801
rect -8273 13088 -8264 13792
rect -7560 13088 -7551 13792
rect -8273 13079 -7551 13088
rect -7280 13768 -7264 13832
rect -7200 13768 -7184 13832
rect -5868 13832 -5772 13868
rect -7280 13752 -7184 13768
rect -7280 13688 -7264 13752
rect -7200 13688 -7184 13752
rect -7280 13672 -7184 13688
rect -7280 13608 -7264 13672
rect -7200 13608 -7184 13672
rect -7280 13592 -7184 13608
rect -7280 13528 -7264 13592
rect -7200 13528 -7184 13592
rect -7280 13512 -7184 13528
rect -7280 13448 -7264 13512
rect -7200 13448 -7184 13512
rect -7280 13432 -7184 13448
rect -7280 13368 -7264 13432
rect -7200 13368 -7184 13432
rect -7280 13352 -7184 13368
rect -7280 13288 -7264 13352
rect -7200 13288 -7184 13352
rect -7280 13272 -7184 13288
rect -7280 13208 -7264 13272
rect -7200 13208 -7184 13272
rect -7280 13192 -7184 13208
rect -7280 13128 -7264 13192
rect -7200 13128 -7184 13192
rect -7280 13112 -7184 13128
rect -8692 13012 -8596 13048
rect -7280 13048 -7264 13112
rect -7200 13048 -7184 13112
rect -6861 13792 -6139 13801
rect -6861 13088 -6852 13792
rect -6148 13088 -6139 13792
rect -6861 13079 -6139 13088
rect -5868 13768 -5852 13832
rect -5788 13768 -5772 13832
rect -4456 13832 -4360 13868
rect -5868 13752 -5772 13768
rect -5868 13688 -5852 13752
rect -5788 13688 -5772 13752
rect -5868 13672 -5772 13688
rect -5868 13608 -5852 13672
rect -5788 13608 -5772 13672
rect -5868 13592 -5772 13608
rect -5868 13528 -5852 13592
rect -5788 13528 -5772 13592
rect -5868 13512 -5772 13528
rect -5868 13448 -5852 13512
rect -5788 13448 -5772 13512
rect -5868 13432 -5772 13448
rect -5868 13368 -5852 13432
rect -5788 13368 -5772 13432
rect -5868 13352 -5772 13368
rect -5868 13288 -5852 13352
rect -5788 13288 -5772 13352
rect -5868 13272 -5772 13288
rect -5868 13208 -5852 13272
rect -5788 13208 -5772 13272
rect -5868 13192 -5772 13208
rect -5868 13128 -5852 13192
rect -5788 13128 -5772 13192
rect -5868 13112 -5772 13128
rect -7280 13012 -7184 13048
rect -5868 13048 -5852 13112
rect -5788 13048 -5772 13112
rect -5449 13792 -4727 13801
rect -5449 13088 -5440 13792
rect -4736 13088 -4727 13792
rect -5449 13079 -4727 13088
rect -4456 13768 -4440 13832
rect -4376 13768 -4360 13832
rect -3044 13832 -2948 13868
rect -4456 13752 -4360 13768
rect -4456 13688 -4440 13752
rect -4376 13688 -4360 13752
rect -4456 13672 -4360 13688
rect -4456 13608 -4440 13672
rect -4376 13608 -4360 13672
rect -4456 13592 -4360 13608
rect -4456 13528 -4440 13592
rect -4376 13528 -4360 13592
rect -4456 13512 -4360 13528
rect -4456 13448 -4440 13512
rect -4376 13448 -4360 13512
rect -4456 13432 -4360 13448
rect -4456 13368 -4440 13432
rect -4376 13368 -4360 13432
rect -4456 13352 -4360 13368
rect -4456 13288 -4440 13352
rect -4376 13288 -4360 13352
rect -4456 13272 -4360 13288
rect -4456 13208 -4440 13272
rect -4376 13208 -4360 13272
rect -4456 13192 -4360 13208
rect -4456 13128 -4440 13192
rect -4376 13128 -4360 13192
rect -4456 13112 -4360 13128
rect -5868 13012 -5772 13048
rect -4456 13048 -4440 13112
rect -4376 13048 -4360 13112
rect -4037 13792 -3315 13801
rect -4037 13088 -4028 13792
rect -3324 13088 -3315 13792
rect -4037 13079 -3315 13088
rect -3044 13768 -3028 13832
rect -2964 13768 -2948 13832
rect -1632 13832 -1536 13868
rect -3044 13752 -2948 13768
rect -3044 13688 -3028 13752
rect -2964 13688 -2948 13752
rect -3044 13672 -2948 13688
rect -3044 13608 -3028 13672
rect -2964 13608 -2948 13672
rect -3044 13592 -2948 13608
rect -3044 13528 -3028 13592
rect -2964 13528 -2948 13592
rect -3044 13512 -2948 13528
rect -3044 13448 -3028 13512
rect -2964 13448 -2948 13512
rect -3044 13432 -2948 13448
rect -3044 13368 -3028 13432
rect -2964 13368 -2948 13432
rect -3044 13352 -2948 13368
rect -3044 13288 -3028 13352
rect -2964 13288 -2948 13352
rect -3044 13272 -2948 13288
rect -3044 13208 -3028 13272
rect -2964 13208 -2948 13272
rect -3044 13192 -2948 13208
rect -3044 13128 -3028 13192
rect -2964 13128 -2948 13192
rect -3044 13112 -2948 13128
rect -4456 13012 -4360 13048
rect -3044 13048 -3028 13112
rect -2964 13048 -2948 13112
rect -2625 13792 -1903 13801
rect -2625 13088 -2616 13792
rect -1912 13088 -1903 13792
rect -2625 13079 -1903 13088
rect -1632 13768 -1616 13832
rect -1552 13768 -1536 13832
rect -220 13832 -124 13868
rect -1632 13752 -1536 13768
rect -1632 13688 -1616 13752
rect -1552 13688 -1536 13752
rect -1632 13672 -1536 13688
rect -1632 13608 -1616 13672
rect -1552 13608 -1536 13672
rect -1632 13592 -1536 13608
rect -1632 13528 -1616 13592
rect -1552 13528 -1536 13592
rect -1632 13512 -1536 13528
rect -1632 13448 -1616 13512
rect -1552 13448 -1536 13512
rect -1632 13432 -1536 13448
rect -1632 13368 -1616 13432
rect -1552 13368 -1536 13432
rect -1632 13352 -1536 13368
rect -1632 13288 -1616 13352
rect -1552 13288 -1536 13352
rect -1632 13272 -1536 13288
rect -1632 13208 -1616 13272
rect -1552 13208 -1536 13272
rect -1632 13192 -1536 13208
rect -1632 13128 -1616 13192
rect -1552 13128 -1536 13192
rect -1632 13112 -1536 13128
rect -3044 13012 -2948 13048
rect -1632 13048 -1616 13112
rect -1552 13048 -1536 13112
rect -1213 13792 -491 13801
rect -1213 13088 -1204 13792
rect -500 13088 -491 13792
rect -1213 13079 -491 13088
rect -220 13768 -204 13832
rect -140 13768 -124 13832
rect 1192 13832 1288 13868
rect -220 13752 -124 13768
rect -220 13688 -204 13752
rect -140 13688 -124 13752
rect -220 13672 -124 13688
rect -220 13608 -204 13672
rect -140 13608 -124 13672
rect -220 13592 -124 13608
rect -220 13528 -204 13592
rect -140 13528 -124 13592
rect -220 13512 -124 13528
rect -220 13448 -204 13512
rect -140 13448 -124 13512
rect -220 13432 -124 13448
rect -220 13368 -204 13432
rect -140 13368 -124 13432
rect -220 13352 -124 13368
rect -220 13288 -204 13352
rect -140 13288 -124 13352
rect -220 13272 -124 13288
rect -220 13208 -204 13272
rect -140 13208 -124 13272
rect -220 13192 -124 13208
rect -220 13128 -204 13192
rect -140 13128 -124 13192
rect -220 13112 -124 13128
rect -1632 13012 -1536 13048
rect -220 13048 -204 13112
rect -140 13048 -124 13112
rect 199 13792 921 13801
rect 199 13088 208 13792
rect 912 13088 921 13792
rect 199 13079 921 13088
rect 1192 13768 1208 13832
rect 1272 13768 1288 13832
rect 2604 13832 2700 13868
rect 1192 13752 1288 13768
rect 1192 13688 1208 13752
rect 1272 13688 1288 13752
rect 1192 13672 1288 13688
rect 1192 13608 1208 13672
rect 1272 13608 1288 13672
rect 1192 13592 1288 13608
rect 1192 13528 1208 13592
rect 1272 13528 1288 13592
rect 1192 13512 1288 13528
rect 1192 13448 1208 13512
rect 1272 13448 1288 13512
rect 1192 13432 1288 13448
rect 1192 13368 1208 13432
rect 1272 13368 1288 13432
rect 1192 13352 1288 13368
rect 1192 13288 1208 13352
rect 1272 13288 1288 13352
rect 1192 13272 1288 13288
rect 1192 13208 1208 13272
rect 1272 13208 1288 13272
rect 1192 13192 1288 13208
rect 1192 13128 1208 13192
rect 1272 13128 1288 13192
rect 1192 13112 1288 13128
rect -220 13012 -124 13048
rect 1192 13048 1208 13112
rect 1272 13048 1288 13112
rect 1611 13792 2333 13801
rect 1611 13088 1620 13792
rect 2324 13088 2333 13792
rect 1611 13079 2333 13088
rect 2604 13768 2620 13832
rect 2684 13768 2700 13832
rect 4016 13832 4112 13868
rect 2604 13752 2700 13768
rect 2604 13688 2620 13752
rect 2684 13688 2700 13752
rect 2604 13672 2700 13688
rect 2604 13608 2620 13672
rect 2684 13608 2700 13672
rect 2604 13592 2700 13608
rect 2604 13528 2620 13592
rect 2684 13528 2700 13592
rect 2604 13512 2700 13528
rect 2604 13448 2620 13512
rect 2684 13448 2700 13512
rect 2604 13432 2700 13448
rect 2604 13368 2620 13432
rect 2684 13368 2700 13432
rect 2604 13352 2700 13368
rect 2604 13288 2620 13352
rect 2684 13288 2700 13352
rect 2604 13272 2700 13288
rect 2604 13208 2620 13272
rect 2684 13208 2700 13272
rect 2604 13192 2700 13208
rect 2604 13128 2620 13192
rect 2684 13128 2700 13192
rect 2604 13112 2700 13128
rect 1192 13012 1288 13048
rect 2604 13048 2620 13112
rect 2684 13048 2700 13112
rect 3023 13792 3745 13801
rect 3023 13088 3032 13792
rect 3736 13088 3745 13792
rect 3023 13079 3745 13088
rect 4016 13768 4032 13832
rect 4096 13768 4112 13832
rect 5428 13832 5524 13868
rect 4016 13752 4112 13768
rect 4016 13688 4032 13752
rect 4096 13688 4112 13752
rect 4016 13672 4112 13688
rect 4016 13608 4032 13672
rect 4096 13608 4112 13672
rect 4016 13592 4112 13608
rect 4016 13528 4032 13592
rect 4096 13528 4112 13592
rect 4016 13512 4112 13528
rect 4016 13448 4032 13512
rect 4096 13448 4112 13512
rect 4016 13432 4112 13448
rect 4016 13368 4032 13432
rect 4096 13368 4112 13432
rect 4016 13352 4112 13368
rect 4016 13288 4032 13352
rect 4096 13288 4112 13352
rect 4016 13272 4112 13288
rect 4016 13208 4032 13272
rect 4096 13208 4112 13272
rect 4016 13192 4112 13208
rect 4016 13128 4032 13192
rect 4096 13128 4112 13192
rect 4016 13112 4112 13128
rect 2604 13012 2700 13048
rect 4016 13048 4032 13112
rect 4096 13048 4112 13112
rect 4435 13792 5157 13801
rect 4435 13088 4444 13792
rect 5148 13088 5157 13792
rect 4435 13079 5157 13088
rect 5428 13768 5444 13832
rect 5508 13768 5524 13832
rect 6840 13832 6936 13868
rect 5428 13752 5524 13768
rect 5428 13688 5444 13752
rect 5508 13688 5524 13752
rect 5428 13672 5524 13688
rect 5428 13608 5444 13672
rect 5508 13608 5524 13672
rect 5428 13592 5524 13608
rect 5428 13528 5444 13592
rect 5508 13528 5524 13592
rect 5428 13512 5524 13528
rect 5428 13448 5444 13512
rect 5508 13448 5524 13512
rect 5428 13432 5524 13448
rect 5428 13368 5444 13432
rect 5508 13368 5524 13432
rect 5428 13352 5524 13368
rect 5428 13288 5444 13352
rect 5508 13288 5524 13352
rect 5428 13272 5524 13288
rect 5428 13208 5444 13272
rect 5508 13208 5524 13272
rect 5428 13192 5524 13208
rect 5428 13128 5444 13192
rect 5508 13128 5524 13192
rect 5428 13112 5524 13128
rect 4016 13012 4112 13048
rect 5428 13048 5444 13112
rect 5508 13048 5524 13112
rect 5847 13792 6569 13801
rect 5847 13088 5856 13792
rect 6560 13088 6569 13792
rect 5847 13079 6569 13088
rect 6840 13768 6856 13832
rect 6920 13768 6936 13832
rect 8252 13832 8348 13868
rect 6840 13752 6936 13768
rect 6840 13688 6856 13752
rect 6920 13688 6936 13752
rect 6840 13672 6936 13688
rect 6840 13608 6856 13672
rect 6920 13608 6936 13672
rect 6840 13592 6936 13608
rect 6840 13528 6856 13592
rect 6920 13528 6936 13592
rect 6840 13512 6936 13528
rect 6840 13448 6856 13512
rect 6920 13448 6936 13512
rect 6840 13432 6936 13448
rect 6840 13368 6856 13432
rect 6920 13368 6936 13432
rect 6840 13352 6936 13368
rect 6840 13288 6856 13352
rect 6920 13288 6936 13352
rect 6840 13272 6936 13288
rect 6840 13208 6856 13272
rect 6920 13208 6936 13272
rect 6840 13192 6936 13208
rect 6840 13128 6856 13192
rect 6920 13128 6936 13192
rect 6840 13112 6936 13128
rect 5428 13012 5524 13048
rect 6840 13048 6856 13112
rect 6920 13048 6936 13112
rect 7259 13792 7981 13801
rect 7259 13088 7268 13792
rect 7972 13088 7981 13792
rect 7259 13079 7981 13088
rect 8252 13768 8268 13832
rect 8332 13768 8348 13832
rect 9664 13832 9760 13868
rect 8252 13752 8348 13768
rect 8252 13688 8268 13752
rect 8332 13688 8348 13752
rect 8252 13672 8348 13688
rect 8252 13608 8268 13672
rect 8332 13608 8348 13672
rect 8252 13592 8348 13608
rect 8252 13528 8268 13592
rect 8332 13528 8348 13592
rect 8252 13512 8348 13528
rect 8252 13448 8268 13512
rect 8332 13448 8348 13512
rect 8252 13432 8348 13448
rect 8252 13368 8268 13432
rect 8332 13368 8348 13432
rect 8252 13352 8348 13368
rect 8252 13288 8268 13352
rect 8332 13288 8348 13352
rect 8252 13272 8348 13288
rect 8252 13208 8268 13272
rect 8332 13208 8348 13272
rect 8252 13192 8348 13208
rect 8252 13128 8268 13192
rect 8332 13128 8348 13192
rect 8252 13112 8348 13128
rect 6840 13012 6936 13048
rect 8252 13048 8268 13112
rect 8332 13048 8348 13112
rect 8671 13792 9393 13801
rect 8671 13088 8680 13792
rect 9384 13088 9393 13792
rect 8671 13079 9393 13088
rect 9664 13768 9680 13832
rect 9744 13768 9760 13832
rect 11076 13832 11172 13868
rect 9664 13752 9760 13768
rect 9664 13688 9680 13752
rect 9744 13688 9760 13752
rect 9664 13672 9760 13688
rect 9664 13608 9680 13672
rect 9744 13608 9760 13672
rect 9664 13592 9760 13608
rect 9664 13528 9680 13592
rect 9744 13528 9760 13592
rect 9664 13512 9760 13528
rect 9664 13448 9680 13512
rect 9744 13448 9760 13512
rect 9664 13432 9760 13448
rect 9664 13368 9680 13432
rect 9744 13368 9760 13432
rect 9664 13352 9760 13368
rect 9664 13288 9680 13352
rect 9744 13288 9760 13352
rect 9664 13272 9760 13288
rect 9664 13208 9680 13272
rect 9744 13208 9760 13272
rect 9664 13192 9760 13208
rect 9664 13128 9680 13192
rect 9744 13128 9760 13192
rect 9664 13112 9760 13128
rect 8252 13012 8348 13048
rect 9664 13048 9680 13112
rect 9744 13048 9760 13112
rect 10083 13792 10805 13801
rect 10083 13088 10092 13792
rect 10796 13088 10805 13792
rect 10083 13079 10805 13088
rect 11076 13768 11092 13832
rect 11156 13768 11172 13832
rect 12488 13832 12584 13868
rect 11076 13752 11172 13768
rect 11076 13688 11092 13752
rect 11156 13688 11172 13752
rect 11076 13672 11172 13688
rect 11076 13608 11092 13672
rect 11156 13608 11172 13672
rect 11076 13592 11172 13608
rect 11076 13528 11092 13592
rect 11156 13528 11172 13592
rect 11076 13512 11172 13528
rect 11076 13448 11092 13512
rect 11156 13448 11172 13512
rect 11076 13432 11172 13448
rect 11076 13368 11092 13432
rect 11156 13368 11172 13432
rect 11076 13352 11172 13368
rect 11076 13288 11092 13352
rect 11156 13288 11172 13352
rect 11076 13272 11172 13288
rect 11076 13208 11092 13272
rect 11156 13208 11172 13272
rect 11076 13192 11172 13208
rect 11076 13128 11092 13192
rect 11156 13128 11172 13192
rect 11076 13112 11172 13128
rect 9664 13012 9760 13048
rect 11076 13048 11092 13112
rect 11156 13048 11172 13112
rect 11495 13792 12217 13801
rect 11495 13088 11504 13792
rect 12208 13088 12217 13792
rect 11495 13079 12217 13088
rect 12488 13768 12504 13832
rect 12568 13768 12584 13832
rect 13900 13832 13996 13868
rect 12488 13752 12584 13768
rect 12488 13688 12504 13752
rect 12568 13688 12584 13752
rect 12488 13672 12584 13688
rect 12488 13608 12504 13672
rect 12568 13608 12584 13672
rect 12488 13592 12584 13608
rect 12488 13528 12504 13592
rect 12568 13528 12584 13592
rect 12488 13512 12584 13528
rect 12488 13448 12504 13512
rect 12568 13448 12584 13512
rect 12488 13432 12584 13448
rect 12488 13368 12504 13432
rect 12568 13368 12584 13432
rect 12488 13352 12584 13368
rect 12488 13288 12504 13352
rect 12568 13288 12584 13352
rect 12488 13272 12584 13288
rect 12488 13208 12504 13272
rect 12568 13208 12584 13272
rect 12488 13192 12584 13208
rect 12488 13128 12504 13192
rect 12568 13128 12584 13192
rect 12488 13112 12584 13128
rect 11076 13012 11172 13048
rect 12488 13048 12504 13112
rect 12568 13048 12584 13112
rect 12907 13792 13629 13801
rect 12907 13088 12916 13792
rect 13620 13088 13629 13792
rect 12907 13079 13629 13088
rect 13900 13768 13916 13832
rect 13980 13768 13996 13832
rect 15312 13832 15408 13868
rect 13900 13752 13996 13768
rect 13900 13688 13916 13752
rect 13980 13688 13996 13752
rect 13900 13672 13996 13688
rect 13900 13608 13916 13672
rect 13980 13608 13996 13672
rect 13900 13592 13996 13608
rect 13900 13528 13916 13592
rect 13980 13528 13996 13592
rect 13900 13512 13996 13528
rect 13900 13448 13916 13512
rect 13980 13448 13996 13512
rect 13900 13432 13996 13448
rect 13900 13368 13916 13432
rect 13980 13368 13996 13432
rect 13900 13352 13996 13368
rect 13900 13288 13916 13352
rect 13980 13288 13996 13352
rect 13900 13272 13996 13288
rect 13900 13208 13916 13272
rect 13980 13208 13996 13272
rect 13900 13192 13996 13208
rect 13900 13128 13916 13192
rect 13980 13128 13996 13192
rect 13900 13112 13996 13128
rect 12488 13012 12584 13048
rect 13900 13048 13916 13112
rect 13980 13048 13996 13112
rect 14319 13792 15041 13801
rect 14319 13088 14328 13792
rect 15032 13088 15041 13792
rect 14319 13079 15041 13088
rect 15312 13768 15328 13832
rect 15392 13768 15408 13832
rect 16724 13832 16820 13868
rect 15312 13752 15408 13768
rect 15312 13688 15328 13752
rect 15392 13688 15408 13752
rect 15312 13672 15408 13688
rect 15312 13608 15328 13672
rect 15392 13608 15408 13672
rect 15312 13592 15408 13608
rect 15312 13528 15328 13592
rect 15392 13528 15408 13592
rect 15312 13512 15408 13528
rect 15312 13448 15328 13512
rect 15392 13448 15408 13512
rect 15312 13432 15408 13448
rect 15312 13368 15328 13432
rect 15392 13368 15408 13432
rect 15312 13352 15408 13368
rect 15312 13288 15328 13352
rect 15392 13288 15408 13352
rect 15312 13272 15408 13288
rect 15312 13208 15328 13272
rect 15392 13208 15408 13272
rect 15312 13192 15408 13208
rect 15312 13128 15328 13192
rect 15392 13128 15408 13192
rect 15312 13112 15408 13128
rect 13900 13012 13996 13048
rect 15312 13048 15328 13112
rect 15392 13048 15408 13112
rect 15731 13792 16453 13801
rect 15731 13088 15740 13792
rect 16444 13088 16453 13792
rect 15731 13079 16453 13088
rect 16724 13768 16740 13832
rect 16804 13768 16820 13832
rect 18136 13832 18232 13868
rect 16724 13752 16820 13768
rect 16724 13688 16740 13752
rect 16804 13688 16820 13752
rect 16724 13672 16820 13688
rect 16724 13608 16740 13672
rect 16804 13608 16820 13672
rect 16724 13592 16820 13608
rect 16724 13528 16740 13592
rect 16804 13528 16820 13592
rect 16724 13512 16820 13528
rect 16724 13448 16740 13512
rect 16804 13448 16820 13512
rect 16724 13432 16820 13448
rect 16724 13368 16740 13432
rect 16804 13368 16820 13432
rect 16724 13352 16820 13368
rect 16724 13288 16740 13352
rect 16804 13288 16820 13352
rect 16724 13272 16820 13288
rect 16724 13208 16740 13272
rect 16804 13208 16820 13272
rect 16724 13192 16820 13208
rect 16724 13128 16740 13192
rect 16804 13128 16820 13192
rect 16724 13112 16820 13128
rect 15312 13012 15408 13048
rect 16724 13048 16740 13112
rect 16804 13048 16820 13112
rect 17143 13792 17865 13801
rect 17143 13088 17152 13792
rect 17856 13088 17865 13792
rect 17143 13079 17865 13088
rect 18136 13768 18152 13832
rect 18216 13768 18232 13832
rect 19548 13832 19644 13868
rect 18136 13752 18232 13768
rect 18136 13688 18152 13752
rect 18216 13688 18232 13752
rect 18136 13672 18232 13688
rect 18136 13608 18152 13672
rect 18216 13608 18232 13672
rect 18136 13592 18232 13608
rect 18136 13528 18152 13592
rect 18216 13528 18232 13592
rect 18136 13512 18232 13528
rect 18136 13448 18152 13512
rect 18216 13448 18232 13512
rect 18136 13432 18232 13448
rect 18136 13368 18152 13432
rect 18216 13368 18232 13432
rect 18136 13352 18232 13368
rect 18136 13288 18152 13352
rect 18216 13288 18232 13352
rect 18136 13272 18232 13288
rect 18136 13208 18152 13272
rect 18216 13208 18232 13272
rect 18136 13192 18232 13208
rect 18136 13128 18152 13192
rect 18216 13128 18232 13192
rect 18136 13112 18232 13128
rect 16724 13012 16820 13048
rect 18136 13048 18152 13112
rect 18216 13048 18232 13112
rect 18555 13792 19277 13801
rect 18555 13088 18564 13792
rect 19268 13088 19277 13792
rect 18555 13079 19277 13088
rect 19548 13768 19564 13832
rect 19628 13768 19644 13832
rect 20960 13832 21056 13868
rect 19548 13752 19644 13768
rect 19548 13688 19564 13752
rect 19628 13688 19644 13752
rect 19548 13672 19644 13688
rect 19548 13608 19564 13672
rect 19628 13608 19644 13672
rect 19548 13592 19644 13608
rect 19548 13528 19564 13592
rect 19628 13528 19644 13592
rect 19548 13512 19644 13528
rect 19548 13448 19564 13512
rect 19628 13448 19644 13512
rect 19548 13432 19644 13448
rect 19548 13368 19564 13432
rect 19628 13368 19644 13432
rect 19548 13352 19644 13368
rect 19548 13288 19564 13352
rect 19628 13288 19644 13352
rect 19548 13272 19644 13288
rect 19548 13208 19564 13272
rect 19628 13208 19644 13272
rect 19548 13192 19644 13208
rect 19548 13128 19564 13192
rect 19628 13128 19644 13192
rect 19548 13112 19644 13128
rect 18136 13012 18232 13048
rect 19548 13048 19564 13112
rect 19628 13048 19644 13112
rect 19967 13792 20689 13801
rect 19967 13088 19976 13792
rect 20680 13088 20689 13792
rect 19967 13079 20689 13088
rect 20960 13768 20976 13832
rect 21040 13768 21056 13832
rect 22372 13832 22468 13868
rect 20960 13752 21056 13768
rect 20960 13688 20976 13752
rect 21040 13688 21056 13752
rect 20960 13672 21056 13688
rect 20960 13608 20976 13672
rect 21040 13608 21056 13672
rect 20960 13592 21056 13608
rect 20960 13528 20976 13592
rect 21040 13528 21056 13592
rect 20960 13512 21056 13528
rect 20960 13448 20976 13512
rect 21040 13448 21056 13512
rect 20960 13432 21056 13448
rect 20960 13368 20976 13432
rect 21040 13368 21056 13432
rect 20960 13352 21056 13368
rect 20960 13288 20976 13352
rect 21040 13288 21056 13352
rect 20960 13272 21056 13288
rect 20960 13208 20976 13272
rect 21040 13208 21056 13272
rect 20960 13192 21056 13208
rect 20960 13128 20976 13192
rect 21040 13128 21056 13192
rect 20960 13112 21056 13128
rect 19548 13012 19644 13048
rect 20960 13048 20976 13112
rect 21040 13048 21056 13112
rect 21379 13792 22101 13801
rect 21379 13088 21388 13792
rect 22092 13088 22101 13792
rect 21379 13079 22101 13088
rect 22372 13768 22388 13832
rect 22452 13768 22468 13832
rect 23784 13832 23880 13868
rect 22372 13752 22468 13768
rect 22372 13688 22388 13752
rect 22452 13688 22468 13752
rect 22372 13672 22468 13688
rect 22372 13608 22388 13672
rect 22452 13608 22468 13672
rect 22372 13592 22468 13608
rect 22372 13528 22388 13592
rect 22452 13528 22468 13592
rect 22372 13512 22468 13528
rect 22372 13448 22388 13512
rect 22452 13448 22468 13512
rect 22372 13432 22468 13448
rect 22372 13368 22388 13432
rect 22452 13368 22468 13432
rect 22372 13352 22468 13368
rect 22372 13288 22388 13352
rect 22452 13288 22468 13352
rect 22372 13272 22468 13288
rect 22372 13208 22388 13272
rect 22452 13208 22468 13272
rect 22372 13192 22468 13208
rect 22372 13128 22388 13192
rect 22452 13128 22468 13192
rect 22372 13112 22468 13128
rect 20960 13012 21056 13048
rect 22372 13048 22388 13112
rect 22452 13048 22468 13112
rect 22791 13792 23513 13801
rect 22791 13088 22800 13792
rect 23504 13088 23513 13792
rect 22791 13079 23513 13088
rect 23784 13768 23800 13832
rect 23864 13768 23880 13832
rect 23784 13752 23880 13768
rect 23784 13688 23800 13752
rect 23864 13688 23880 13752
rect 23784 13672 23880 13688
rect 23784 13608 23800 13672
rect 23864 13608 23880 13672
rect 23784 13592 23880 13608
rect 23784 13528 23800 13592
rect 23864 13528 23880 13592
rect 23784 13512 23880 13528
rect 23784 13448 23800 13512
rect 23864 13448 23880 13512
rect 23784 13432 23880 13448
rect 23784 13368 23800 13432
rect 23864 13368 23880 13432
rect 23784 13352 23880 13368
rect 23784 13288 23800 13352
rect 23864 13288 23880 13352
rect 23784 13272 23880 13288
rect 23784 13208 23800 13272
rect 23864 13208 23880 13272
rect 23784 13192 23880 13208
rect 23784 13128 23800 13192
rect 23864 13128 23880 13192
rect 23784 13112 23880 13128
rect 22372 13012 22468 13048
rect 23784 13048 23800 13112
rect 23864 13048 23880 13112
rect 23784 13012 23880 13048
rect -22812 12712 -22716 12748
rect -23805 12672 -23083 12681
rect -23805 11968 -23796 12672
rect -23092 11968 -23083 12672
rect -23805 11959 -23083 11968
rect -22812 12648 -22796 12712
rect -22732 12648 -22716 12712
rect -21400 12712 -21304 12748
rect -22812 12632 -22716 12648
rect -22812 12568 -22796 12632
rect -22732 12568 -22716 12632
rect -22812 12552 -22716 12568
rect -22812 12488 -22796 12552
rect -22732 12488 -22716 12552
rect -22812 12472 -22716 12488
rect -22812 12408 -22796 12472
rect -22732 12408 -22716 12472
rect -22812 12392 -22716 12408
rect -22812 12328 -22796 12392
rect -22732 12328 -22716 12392
rect -22812 12312 -22716 12328
rect -22812 12248 -22796 12312
rect -22732 12248 -22716 12312
rect -22812 12232 -22716 12248
rect -22812 12168 -22796 12232
rect -22732 12168 -22716 12232
rect -22812 12152 -22716 12168
rect -22812 12088 -22796 12152
rect -22732 12088 -22716 12152
rect -22812 12072 -22716 12088
rect -22812 12008 -22796 12072
rect -22732 12008 -22716 12072
rect -22812 11992 -22716 12008
rect -22812 11928 -22796 11992
rect -22732 11928 -22716 11992
rect -22393 12672 -21671 12681
rect -22393 11968 -22384 12672
rect -21680 11968 -21671 12672
rect -22393 11959 -21671 11968
rect -21400 12648 -21384 12712
rect -21320 12648 -21304 12712
rect -19988 12712 -19892 12748
rect -21400 12632 -21304 12648
rect -21400 12568 -21384 12632
rect -21320 12568 -21304 12632
rect -21400 12552 -21304 12568
rect -21400 12488 -21384 12552
rect -21320 12488 -21304 12552
rect -21400 12472 -21304 12488
rect -21400 12408 -21384 12472
rect -21320 12408 -21304 12472
rect -21400 12392 -21304 12408
rect -21400 12328 -21384 12392
rect -21320 12328 -21304 12392
rect -21400 12312 -21304 12328
rect -21400 12248 -21384 12312
rect -21320 12248 -21304 12312
rect -21400 12232 -21304 12248
rect -21400 12168 -21384 12232
rect -21320 12168 -21304 12232
rect -21400 12152 -21304 12168
rect -21400 12088 -21384 12152
rect -21320 12088 -21304 12152
rect -21400 12072 -21304 12088
rect -21400 12008 -21384 12072
rect -21320 12008 -21304 12072
rect -21400 11992 -21304 12008
rect -22812 11892 -22716 11928
rect -21400 11928 -21384 11992
rect -21320 11928 -21304 11992
rect -20981 12672 -20259 12681
rect -20981 11968 -20972 12672
rect -20268 11968 -20259 12672
rect -20981 11959 -20259 11968
rect -19988 12648 -19972 12712
rect -19908 12648 -19892 12712
rect -18576 12712 -18480 12748
rect -19988 12632 -19892 12648
rect -19988 12568 -19972 12632
rect -19908 12568 -19892 12632
rect -19988 12552 -19892 12568
rect -19988 12488 -19972 12552
rect -19908 12488 -19892 12552
rect -19988 12472 -19892 12488
rect -19988 12408 -19972 12472
rect -19908 12408 -19892 12472
rect -19988 12392 -19892 12408
rect -19988 12328 -19972 12392
rect -19908 12328 -19892 12392
rect -19988 12312 -19892 12328
rect -19988 12248 -19972 12312
rect -19908 12248 -19892 12312
rect -19988 12232 -19892 12248
rect -19988 12168 -19972 12232
rect -19908 12168 -19892 12232
rect -19988 12152 -19892 12168
rect -19988 12088 -19972 12152
rect -19908 12088 -19892 12152
rect -19988 12072 -19892 12088
rect -19988 12008 -19972 12072
rect -19908 12008 -19892 12072
rect -19988 11992 -19892 12008
rect -21400 11892 -21304 11928
rect -19988 11928 -19972 11992
rect -19908 11928 -19892 11992
rect -19569 12672 -18847 12681
rect -19569 11968 -19560 12672
rect -18856 11968 -18847 12672
rect -19569 11959 -18847 11968
rect -18576 12648 -18560 12712
rect -18496 12648 -18480 12712
rect -17164 12712 -17068 12748
rect -18576 12632 -18480 12648
rect -18576 12568 -18560 12632
rect -18496 12568 -18480 12632
rect -18576 12552 -18480 12568
rect -18576 12488 -18560 12552
rect -18496 12488 -18480 12552
rect -18576 12472 -18480 12488
rect -18576 12408 -18560 12472
rect -18496 12408 -18480 12472
rect -18576 12392 -18480 12408
rect -18576 12328 -18560 12392
rect -18496 12328 -18480 12392
rect -18576 12312 -18480 12328
rect -18576 12248 -18560 12312
rect -18496 12248 -18480 12312
rect -18576 12232 -18480 12248
rect -18576 12168 -18560 12232
rect -18496 12168 -18480 12232
rect -18576 12152 -18480 12168
rect -18576 12088 -18560 12152
rect -18496 12088 -18480 12152
rect -18576 12072 -18480 12088
rect -18576 12008 -18560 12072
rect -18496 12008 -18480 12072
rect -18576 11992 -18480 12008
rect -19988 11892 -19892 11928
rect -18576 11928 -18560 11992
rect -18496 11928 -18480 11992
rect -18157 12672 -17435 12681
rect -18157 11968 -18148 12672
rect -17444 11968 -17435 12672
rect -18157 11959 -17435 11968
rect -17164 12648 -17148 12712
rect -17084 12648 -17068 12712
rect -15752 12712 -15656 12748
rect -17164 12632 -17068 12648
rect -17164 12568 -17148 12632
rect -17084 12568 -17068 12632
rect -17164 12552 -17068 12568
rect -17164 12488 -17148 12552
rect -17084 12488 -17068 12552
rect -17164 12472 -17068 12488
rect -17164 12408 -17148 12472
rect -17084 12408 -17068 12472
rect -17164 12392 -17068 12408
rect -17164 12328 -17148 12392
rect -17084 12328 -17068 12392
rect -17164 12312 -17068 12328
rect -17164 12248 -17148 12312
rect -17084 12248 -17068 12312
rect -17164 12232 -17068 12248
rect -17164 12168 -17148 12232
rect -17084 12168 -17068 12232
rect -17164 12152 -17068 12168
rect -17164 12088 -17148 12152
rect -17084 12088 -17068 12152
rect -17164 12072 -17068 12088
rect -17164 12008 -17148 12072
rect -17084 12008 -17068 12072
rect -17164 11992 -17068 12008
rect -18576 11892 -18480 11928
rect -17164 11928 -17148 11992
rect -17084 11928 -17068 11992
rect -16745 12672 -16023 12681
rect -16745 11968 -16736 12672
rect -16032 11968 -16023 12672
rect -16745 11959 -16023 11968
rect -15752 12648 -15736 12712
rect -15672 12648 -15656 12712
rect -14340 12712 -14244 12748
rect -15752 12632 -15656 12648
rect -15752 12568 -15736 12632
rect -15672 12568 -15656 12632
rect -15752 12552 -15656 12568
rect -15752 12488 -15736 12552
rect -15672 12488 -15656 12552
rect -15752 12472 -15656 12488
rect -15752 12408 -15736 12472
rect -15672 12408 -15656 12472
rect -15752 12392 -15656 12408
rect -15752 12328 -15736 12392
rect -15672 12328 -15656 12392
rect -15752 12312 -15656 12328
rect -15752 12248 -15736 12312
rect -15672 12248 -15656 12312
rect -15752 12232 -15656 12248
rect -15752 12168 -15736 12232
rect -15672 12168 -15656 12232
rect -15752 12152 -15656 12168
rect -15752 12088 -15736 12152
rect -15672 12088 -15656 12152
rect -15752 12072 -15656 12088
rect -15752 12008 -15736 12072
rect -15672 12008 -15656 12072
rect -15752 11992 -15656 12008
rect -17164 11892 -17068 11928
rect -15752 11928 -15736 11992
rect -15672 11928 -15656 11992
rect -15333 12672 -14611 12681
rect -15333 11968 -15324 12672
rect -14620 11968 -14611 12672
rect -15333 11959 -14611 11968
rect -14340 12648 -14324 12712
rect -14260 12648 -14244 12712
rect -12928 12712 -12832 12748
rect -14340 12632 -14244 12648
rect -14340 12568 -14324 12632
rect -14260 12568 -14244 12632
rect -14340 12552 -14244 12568
rect -14340 12488 -14324 12552
rect -14260 12488 -14244 12552
rect -14340 12472 -14244 12488
rect -14340 12408 -14324 12472
rect -14260 12408 -14244 12472
rect -14340 12392 -14244 12408
rect -14340 12328 -14324 12392
rect -14260 12328 -14244 12392
rect -14340 12312 -14244 12328
rect -14340 12248 -14324 12312
rect -14260 12248 -14244 12312
rect -14340 12232 -14244 12248
rect -14340 12168 -14324 12232
rect -14260 12168 -14244 12232
rect -14340 12152 -14244 12168
rect -14340 12088 -14324 12152
rect -14260 12088 -14244 12152
rect -14340 12072 -14244 12088
rect -14340 12008 -14324 12072
rect -14260 12008 -14244 12072
rect -14340 11992 -14244 12008
rect -15752 11892 -15656 11928
rect -14340 11928 -14324 11992
rect -14260 11928 -14244 11992
rect -13921 12672 -13199 12681
rect -13921 11968 -13912 12672
rect -13208 11968 -13199 12672
rect -13921 11959 -13199 11968
rect -12928 12648 -12912 12712
rect -12848 12648 -12832 12712
rect -11516 12712 -11420 12748
rect -12928 12632 -12832 12648
rect -12928 12568 -12912 12632
rect -12848 12568 -12832 12632
rect -12928 12552 -12832 12568
rect -12928 12488 -12912 12552
rect -12848 12488 -12832 12552
rect -12928 12472 -12832 12488
rect -12928 12408 -12912 12472
rect -12848 12408 -12832 12472
rect -12928 12392 -12832 12408
rect -12928 12328 -12912 12392
rect -12848 12328 -12832 12392
rect -12928 12312 -12832 12328
rect -12928 12248 -12912 12312
rect -12848 12248 -12832 12312
rect -12928 12232 -12832 12248
rect -12928 12168 -12912 12232
rect -12848 12168 -12832 12232
rect -12928 12152 -12832 12168
rect -12928 12088 -12912 12152
rect -12848 12088 -12832 12152
rect -12928 12072 -12832 12088
rect -12928 12008 -12912 12072
rect -12848 12008 -12832 12072
rect -12928 11992 -12832 12008
rect -14340 11892 -14244 11928
rect -12928 11928 -12912 11992
rect -12848 11928 -12832 11992
rect -12509 12672 -11787 12681
rect -12509 11968 -12500 12672
rect -11796 11968 -11787 12672
rect -12509 11959 -11787 11968
rect -11516 12648 -11500 12712
rect -11436 12648 -11420 12712
rect -10104 12712 -10008 12748
rect -11516 12632 -11420 12648
rect -11516 12568 -11500 12632
rect -11436 12568 -11420 12632
rect -11516 12552 -11420 12568
rect -11516 12488 -11500 12552
rect -11436 12488 -11420 12552
rect -11516 12472 -11420 12488
rect -11516 12408 -11500 12472
rect -11436 12408 -11420 12472
rect -11516 12392 -11420 12408
rect -11516 12328 -11500 12392
rect -11436 12328 -11420 12392
rect -11516 12312 -11420 12328
rect -11516 12248 -11500 12312
rect -11436 12248 -11420 12312
rect -11516 12232 -11420 12248
rect -11516 12168 -11500 12232
rect -11436 12168 -11420 12232
rect -11516 12152 -11420 12168
rect -11516 12088 -11500 12152
rect -11436 12088 -11420 12152
rect -11516 12072 -11420 12088
rect -11516 12008 -11500 12072
rect -11436 12008 -11420 12072
rect -11516 11992 -11420 12008
rect -12928 11892 -12832 11928
rect -11516 11928 -11500 11992
rect -11436 11928 -11420 11992
rect -11097 12672 -10375 12681
rect -11097 11968 -11088 12672
rect -10384 11968 -10375 12672
rect -11097 11959 -10375 11968
rect -10104 12648 -10088 12712
rect -10024 12648 -10008 12712
rect -8692 12712 -8596 12748
rect -10104 12632 -10008 12648
rect -10104 12568 -10088 12632
rect -10024 12568 -10008 12632
rect -10104 12552 -10008 12568
rect -10104 12488 -10088 12552
rect -10024 12488 -10008 12552
rect -10104 12472 -10008 12488
rect -10104 12408 -10088 12472
rect -10024 12408 -10008 12472
rect -10104 12392 -10008 12408
rect -10104 12328 -10088 12392
rect -10024 12328 -10008 12392
rect -10104 12312 -10008 12328
rect -10104 12248 -10088 12312
rect -10024 12248 -10008 12312
rect -10104 12232 -10008 12248
rect -10104 12168 -10088 12232
rect -10024 12168 -10008 12232
rect -10104 12152 -10008 12168
rect -10104 12088 -10088 12152
rect -10024 12088 -10008 12152
rect -10104 12072 -10008 12088
rect -10104 12008 -10088 12072
rect -10024 12008 -10008 12072
rect -10104 11992 -10008 12008
rect -11516 11892 -11420 11928
rect -10104 11928 -10088 11992
rect -10024 11928 -10008 11992
rect -9685 12672 -8963 12681
rect -9685 11968 -9676 12672
rect -8972 11968 -8963 12672
rect -9685 11959 -8963 11968
rect -8692 12648 -8676 12712
rect -8612 12648 -8596 12712
rect -7280 12712 -7184 12748
rect -8692 12632 -8596 12648
rect -8692 12568 -8676 12632
rect -8612 12568 -8596 12632
rect -8692 12552 -8596 12568
rect -8692 12488 -8676 12552
rect -8612 12488 -8596 12552
rect -8692 12472 -8596 12488
rect -8692 12408 -8676 12472
rect -8612 12408 -8596 12472
rect -8692 12392 -8596 12408
rect -8692 12328 -8676 12392
rect -8612 12328 -8596 12392
rect -8692 12312 -8596 12328
rect -8692 12248 -8676 12312
rect -8612 12248 -8596 12312
rect -8692 12232 -8596 12248
rect -8692 12168 -8676 12232
rect -8612 12168 -8596 12232
rect -8692 12152 -8596 12168
rect -8692 12088 -8676 12152
rect -8612 12088 -8596 12152
rect -8692 12072 -8596 12088
rect -8692 12008 -8676 12072
rect -8612 12008 -8596 12072
rect -8692 11992 -8596 12008
rect -10104 11892 -10008 11928
rect -8692 11928 -8676 11992
rect -8612 11928 -8596 11992
rect -8273 12672 -7551 12681
rect -8273 11968 -8264 12672
rect -7560 11968 -7551 12672
rect -8273 11959 -7551 11968
rect -7280 12648 -7264 12712
rect -7200 12648 -7184 12712
rect -5868 12712 -5772 12748
rect -7280 12632 -7184 12648
rect -7280 12568 -7264 12632
rect -7200 12568 -7184 12632
rect -7280 12552 -7184 12568
rect -7280 12488 -7264 12552
rect -7200 12488 -7184 12552
rect -7280 12472 -7184 12488
rect -7280 12408 -7264 12472
rect -7200 12408 -7184 12472
rect -7280 12392 -7184 12408
rect -7280 12328 -7264 12392
rect -7200 12328 -7184 12392
rect -7280 12312 -7184 12328
rect -7280 12248 -7264 12312
rect -7200 12248 -7184 12312
rect -7280 12232 -7184 12248
rect -7280 12168 -7264 12232
rect -7200 12168 -7184 12232
rect -7280 12152 -7184 12168
rect -7280 12088 -7264 12152
rect -7200 12088 -7184 12152
rect -7280 12072 -7184 12088
rect -7280 12008 -7264 12072
rect -7200 12008 -7184 12072
rect -7280 11992 -7184 12008
rect -8692 11892 -8596 11928
rect -7280 11928 -7264 11992
rect -7200 11928 -7184 11992
rect -6861 12672 -6139 12681
rect -6861 11968 -6852 12672
rect -6148 11968 -6139 12672
rect -6861 11959 -6139 11968
rect -5868 12648 -5852 12712
rect -5788 12648 -5772 12712
rect -4456 12712 -4360 12748
rect -5868 12632 -5772 12648
rect -5868 12568 -5852 12632
rect -5788 12568 -5772 12632
rect -5868 12552 -5772 12568
rect -5868 12488 -5852 12552
rect -5788 12488 -5772 12552
rect -5868 12472 -5772 12488
rect -5868 12408 -5852 12472
rect -5788 12408 -5772 12472
rect -5868 12392 -5772 12408
rect -5868 12328 -5852 12392
rect -5788 12328 -5772 12392
rect -5868 12312 -5772 12328
rect -5868 12248 -5852 12312
rect -5788 12248 -5772 12312
rect -5868 12232 -5772 12248
rect -5868 12168 -5852 12232
rect -5788 12168 -5772 12232
rect -5868 12152 -5772 12168
rect -5868 12088 -5852 12152
rect -5788 12088 -5772 12152
rect -5868 12072 -5772 12088
rect -5868 12008 -5852 12072
rect -5788 12008 -5772 12072
rect -5868 11992 -5772 12008
rect -7280 11892 -7184 11928
rect -5868 11928 -5852 11992
rect -5788 11928 -5772 11992
rect -5449 12672 -4727 12681
rect -5449 11968 -5440 12672
rect -4736 11968 -4727 12672
rect -5449 11959 -4727 11968
rect -4456 12648 -4440 12712
rect -4376 12648 -4360 12712
rect -3044 12712 -2948 12748
rect -4456 12632 -4360 12648
rect -4456 12568 -4440 12632
rect -4376 12568 -4360 12632
rect -4456 12552 -4360 12568
rect -4456 12488 -4440 12552
rect -4376 12488 -4360 12552
rect -4456 12472 -4360 12488
rect -4456 12408 -4440 12472
rect -4376 12408 -4360 12472
rect -4456 12392 -4360 12408
rect -4456 12328 -4440 12392
rect -4376 12328 -4360 12392
rect -4456 12312 -4360 12328
rect -4456 12248 -4440 12312
rect -4376 12248 -4360 12312
rect -4456 12232 -4360 12248
rect -4456 12168 -4440 12232
rect -4376 12168 -4360 12232
rect -4456 12152 -4360 12168
rect -4456 12088 -4440 12152
rect -4376 12088 -4360 12152
rect -4456 12072 -4360 12088
rect -4456 12008 -4440 12072
rect -4376 12008 -4360 12072
rect -4456 11992 -4360 12008
rect -5868 11892 -5772 11928
rect -4456 11928 -4440 11992
rect -4376 11928 -4360 11992
rect -4037 12672 -3315 12681
rect -4037 11968 -4028 12672
rect -3324 11968 -3315 12672
rect -4037 11959 -3315 11968
rect -3044 12648 -3028 12712
rect -2964 12648 -2948 12712
rect -1632 12712 -1536 12748
rect -3044 12632 -2948 12648
rect -3044 12568 -3028 12632
rect -2964 12568 -2948 12632
rect -3044 12552 -2948 12568
rect -3044 12488 -3028 12552
rect -2964 12488 -2948 12552
rect -3044 12472 -2948 12488
rect -3044 12408 -3028 12472
rect -2964 12408 -2948 12472
rect -3044 12392 -2948 12408
rect -3044 12328 -3028 12392
rect -2964 12328 -2948 12392
rect -3044 12312 -2948 12328
rect -3044 12248 -3028 12312
rect -2964 12248 -2948 12312
rect -3044 12232 -2948 12248
rect -3044 12168 -3028 12232
rect -2964 12168 -2948 12232
rect -3044 12152 -2948 12168
rect -3044 12088 -3028 12152
rect -2964 12088 -2948 12152
rect -3044 12072 -2948 12088
rect -3044 12008 -3028 12072
rect -2964 12008 -2948 12072
rect -3044 11992 -2948 12008
rect -4456 11892 -4360 11928
rect -3044 11928 -3028 11992
rect -2964 11928 -2948 11992
rect -2625 12672 -1903 12681
rect -2625 11968 -2616 12672
rect -1912 11968 -1903 12672
rect -2625 11959 -1903 11968
rect -1632 12648 -1616 12712
rect -1552 12648 -1536 12712
rect -220 12712 -124 12748
rect -1632 12632 -1536 12648
rect -1632 12568 -1616 12632
rect -1552 12568 -1536 12632
rect -1632 12552 -1536 12568
rect -1632 12488 -1616 12552
rect -1552 12488 -1536 12552
rect -1632 12472 -1536 12488
rect -1632 12408 -1616 12472
rect -1552 12408 -1536 12472
rect -1632 12392 -1536 12408
rect -1632 12328 -1616 12392
rect -1552 12328 -1536 12392
rect -1632 12312 -1536 12328
rect -1632 12248 -1616 12312
rect -1552 12248 -1536 12312
rect -1632 12232 -1536 12248
rect -1632 12168 -1616 12232
rect -1552 12168 -1536 12232
rect -1632 12152 -1536 12168
rect -1632 12088 -1616 12152
rect -1552 12088 -1536 12152
rect -1632 12072 -1536 12088
rect -1632 12008 -1616 12072
rect -1552 12008 -1536 12072
rect -1632 11992 -1536 12008
rect -3044 11892 -2948 11928
rect -1632 11928 -1616 11992
rect -1552 11928 -1536 11992
rect -1213 12672 -491 12681
rect -1213 11968 -1204 12672
rect -500 11968 -491 12672
rect -1213 11959 -491 11968
rect -220 12648 -204 12712
rect -140 12648 -124 12712
rect 1192 12712 1288 12748
rect -220 12632 -124 12648
rect -220 12568 -204 12632
rect -140 12568 -124 12632
rect -220 12552 -124 12568
rect -220 12488 -204 12552
rect -140 12488 -124 12552
rect -220 12472 -124 12488
rect -220 12408 -204 12472
rect -140 12408 -124 12472
rect -220 12392 -124 12408
rect -220 12328 -204 12392
rect -140 12328 -124 12392
rect -220 12312 -124 12328
rect -220 12248 -204 12312
rect -140 12248 -124 12312
rect -220 12232 -124 12248
rect -220 12168 -204 12232
rect -140 12168 -124 12232
rect -220 12152 -124 12168
rect -220 12088 -204 12152
rect -140 12088 -124 12152
rect -220 12072 -124 12088
rect -220 12008 -204 12072
rect -140 12008 -124 12072
rect -220 11992 -124 12008
rect -1632 11892 -1536 11928
rect -220 11928 -204 11992
rect -140 11928 -124 11992
rect 199 12672 921 12681
rect 199 11968 208 12672
rect 912 11968 921 12672
rect 199 11959 921 11968
rect 1192 12648 1208 12712
rect 1272 12648 1288 12712
rect 2604 12712 2700 12748
rect 1192 12632 1288 12648
rect 1192 12568 1208 12632
rect 1272 12568 1288 12632
rect 1192 12552 1288 12568
rect 1192 12488 1208 12552
rect 1272 12488 1288 12552
rect 1192 12472 1288 12488
rect 1192 12408 1208 12472
rect 1272 12408 1288 12472
rect 1192 12392 1288 12408
rect 1192 12328 1208 12392
rect 1272 12328 1288 12392
rect 1192 12312 1288 12328
rect 1192 12248 1208 12312
rect 1272 12248 1288 12312
rect 1192 12232 1288 12248
rect 1192 12168 1208 12232
rect 1272 12168 1288 12232
rect 1192 12152 1288 12168
rect 1192 12088 1208 12152
rect 1272 12088 1288 12152
rect 1192 12072 1288 12088
rect 1192 12008 1208 12072
rect 1272 12008 1288 12072
rect 1192 11992 1288 12008
rect -220 11892 -124 11928
rect 1192 11928 1208 11992
rect 1272 11928 1288 11992
rect 1611 12672 2333 12681
rect 1611 11968 1620 12672
rect 2324 11968 2333 12672
rect 1611 11959 2333 11968
rect 2604 12648 2620 12712
rect 2684 12648 2700 12712
rect 4016 12712 4112 12748
rect 2604 12632 2700 12648
rect 2604 12568 2620 12632
rect 2684 12568 2700 12632
rect 2604 12552 2700 12568
rect 2604 12488 2620 12552
rect 2684 12488 2700 12552
rect 2604 12472 2700 12488
rect 2604 12408 2620 12472
rect 2684 12408 2700 12472
rect 2604 12392 2700 12408
rect 2604 12328 2620 12392
rect 2684 12328 2700 12392
rect 2604 12312 2700 12328
rect 2604 12248 2620 12312
rect 2684 12248 2700 12312
rect 2604 12232 2700 12248
rect 2604 12168 2620 12232
rect 2684 12168 2700 12232
rect 2604 12152 2700 12168
rect 2604 12088 2620 12152
rect 2684 12088 2700 12152
rect 2604 12072 2700 12088
rect 2604 12008 2620 12072
rect 2684 12008 2700 12072
rect 2604 11992 2700 12008
rect 1192 11892 1288 11928
rect 2604 11928 2620 11992
rect 2684 11928 2700 11992
rect 3023 12672 3745 12681
rect 3023 11968 3032 12672
rect 3736 11968 3745 12672
rect 3023 11959 3745 11968
rect 4016 12648 4032 12712
rect 4096 12648 4112 12712
rect 5428 12712 5524 12748
rect 4016 12632 4112 12648
rect 4016 12568 4032 12632
rect 4096 12568 4112 12632
rect 4016 12552 4112 12568
rect 4016 12488 4032 12552
rect 4096 12488 4112 12552
rect 4016 12472 4112 12488
rect 4016 12408 4032 12472
rect 4096 12408 4112 12472
rect 4016 12392 4112 12408
rect 4016 12328 4032 12392
rect 4096 12328 4112 12392
rect 4016 12312 4112 12328
rect 4016 12248 4032 12312
rect 4096 12248 4112 12312
rect 4016 12232 4112 12248
rect 4016 12168 4032 12232
rect 4096 12168 4112 12232
rect 4016 12152 4112 12168
rect 4016 12088 4032 12152
rect 4096 12088 4112 12152
rect 4016 12072 4112 12088
rect 4016 12008 4032 12072
rect 4096 12008 4112 12072
rect 4016 11992 4112 12008
rect 2604 11892 2700 11928
rect 4016 11928 4032 11992
rect 4096 11928 4112 11992
rect 4435 12672 5157 12681
rect 4435 11968 4444 12672
rect 5148 11968 5157 12672
rect 4435 11959 5157 11968
rect 5428 12648 5444 12712
rect 5508 12648 5524 12712
rect 6840 12712 6936 12748
rect 5428 12632 5524 12648
rect 5428 12568 5444 12632
rect 5508 12568 5524 12632
rect 5428 12552 5524 12568
rect 5428 12488 5444 12552
rect 5508 12488 5524 12552
rect 5428 12472 5524 12488
rect 5428 12408 5444 12472
rect 5508 12408 5524 12472
rect 5428 12392 5524 12408
rect 5428 12328 5444 12392
rect 5508 12328 5524 12392
rect 5428 12312 5524 12328
rect 5428 12248 5444 12312
rect 5508 12248 5524 12312
rect 5428 12232 5524 12248
rect 5428 12168 5444 12232
rect 5508 12168 5524 12232
rect 5428 12152 5524 12168
rect 5428 12088 5444 12152
rect 5508 12088 5524 12152
rect 5428 12072 5524 12088
rect 5428 12008 5444 12072
rect 5508 12008 5524 12072
rect 5428 11992 5524 12008
rect 4016 11892 4112 11928
rect 5428 11928 5444 11992
rect 5508 11928 5524 11992
rect 5847 12672 6569 12681
rect 5847 11968 5856 12672
rect 6560 11968 6569 12672
rect 5847 11959 6569 11968
rect 6840 12648 6856 12712
rect 6920 12648 6936 12712
rect 8252 12712 8348 12748
rect 6840 12632 6936 12648
rect 6840 12568 6856 12632
rect 6920 12568 6936 12632
rect 6840 12552 6936 12568
rect 6840 12488 6856 12552
rect 6920 12488 6936 12552
rect 6840 12472 6936 12488
rect 6840 12408 6856 12472
rect 6920 12408 6936 12472
rect 6840 12392 6936 12408
rect 6840 12328 6856 12392
rect 6920 12328 6936 12392
rect 6840 12312 6936 12328
rect 6840 12248 6856 12312
rect 6920 12248 6936 12312
rect 6840 12232 6936 12248
rect 6840 12168 6856 12232
rect 6920 12168 6936 12232
rect 6840 12152 6936 12168
rect 6840 12088 6856 12152
rect 6920 12088 6936 12152
rect 6840 12072 6936 12088
rect 6840 12008 6856 12072
rect 6920 12008 6936 12072
rect 6840 11992 6936 12008
rect 5428 11892 5524 11928
rect 6840 11928 6856 11992
rect 6920 11928 6936 11992
rect 7259 12672 7981 12681
rect 7259 11968 7268 12672
rect 7972 11968 7981 12672
rect 7259 11959 7981 11968
rect 8252 12648 8268 12712
rect 8332 12648 8348 12712
rect 9664 12712 9760 12748
rect 8252 12632 8348 12648
rect 8252 12568 8268 12632
rect 8332 12568 8348 12632
rect 8252 12552 8348 12568
rect 8252 12488 8268 12552
rect 8332 12488 8348 12552
rect 8252 12472 8348 12488
rect 8252 12408 8268 12472
rect 8332 12408 8348 12472
rect 8252 12392 8348 12408
rect 8252 12328 8268 12392
rect 8332 12328 8348 12392
rect 8252 12312 8348 12328
rect 8252 12248 8268 12312
rect 8332 12248 8348 12312
rect 8252 12232 8348 12248
rect 8252 12168 8268 12232
rect 8332 12168 8348 12232
rect 8252 12152 8348 12168
rect 8252 12088 8268 12152
rect 8332 12088 8348 12152
rect 8252 12072 8348 12088
rect 8252 12008 8268 12072
rect 8332 12008 8348 12072
rect 8252 11992 8348 12008
rect 6840 11892 6936 11928
rect 8252 11928 8268 11992
rect 8332 11928 8348 11992
rect 8671 12672 9393 12681
rect 8671 11968 8680 12672
rect 9384 11968 9393 12672
rect 8671 11959 9393 11968
rect 9664 12648 9680 12712
rect 9744 12648 9760 12712
rect 11076 12712 11172 12748
rect 9664 12632 9760 12648
rect 9664 12568 9680 12632
rect 9744 12568 9760 12632
rect 9664 12552 9760 12568
rect 9664 12488 9680 12552
rect 9744 12488 9760 12552
rect 9664 12472 9760 12488
rect 9664 12408 9680 12472
rect 9744 12408 9760 12472
rect 9664 12392 9760 12408
rect 9664 12328 9680 12392
rect 9744 12328 9760 12392
rect 9664 12312 9760 12328
rect 9664 12248 9680 12312
rect 9744 12248 9760 12312
rect 9664 12232 9760 12248
rect 9664 12168 9680 12232
rect 9744 12168 9760 12232
rect 9664 12152 9760 12168
rect 9664 12088 9680 12152
rect 9744 12088 9760 12152
rect 9664 12072 9760 12088
rect 9664 12008 9680 12072
rect 9744 12008 9760 12072
rect 9664 11992 9760 12008
rect 8252 11892 8348 11928
rect 9664 11928 9680 11992
rect 9744 11928 9760 11992
rect 10083 12672 10805 12681
rect 10083 11968 10092 12672
rect 10796 11968 10805 12672
rect 10083 11959 10805 11968
rect 11076 12648 11092 12712
rect 11156 12648 11172 12712
rect 12488 12712 12584 12748
rect 11076 12632 11172 12648
rect 11076 12568 11092 12632
rect 11156 12568 11172 12632
rect 11076 12552 11172 12568
rect 11076 12488 11092 12552
rect 11156 12488 11172 12552
rect 11076 12472 11172 12488
rect 11076 12408 11092 12472
rect 11156 12408 11172 12472
rect 11076 12392 11172 12408
rect 11076 12328 11092 12392
rect 11156 12328 11172 12392
rect 11076 12312 11172 12328
rect 11076 12248 11092 12312
rect 11156 12248 11172 12312
rect 11076 12232 11172 12248
rect 11076 12168 11092 12232
rect 11156 12168 11172 12232
rect 11076 12152 11172 12168
rect 11076 12088 11092 12152
rect 11156 12088 11172 12152
rect 11076 12072 11172 12088
rect 11076 12008 11092 12072
rect 11156 12008 11172 12072
rect 11076 11992 11172 12008
rect 9664 11892 9760 11928
rect 11076 11928 11092 11992
rect 11156 11928 11172 11992
rect 11495 12672 12217 12681
rect 11495 11968 11504 12672
rect 12208 11968 12217 12672
rect 11495 11959 12217 11968
rect 12488 12648 12504 12712
rect 12568 12648 12584 12712
rect 13900 12712 13996 12748
rect 12488 12632 12584 12648
rect 12488 12568 12504 12632
rect 12568 12568 12584 12632
rect 12488 12552 12584 12568
rect 12488 12488 12504 12552
rect 12568 12488 12584 12552
rect 12488 12472 12584 12488
rect 12488 12408 12504 12472
rect 12568 12408 12584 12472
rect 12488 12392 12584 12408
rect 12488 12328 12504 12392
rect 12568 12328 12584 12392
rect 12488 12312 12584 12328
rect 12488 12248 12504 12312
rect 12568 12248 12584 12312
rect 12488 12232 12584 12248
rect 12488 12168 12504 12232
rect 12568 12168 12584 12232
rect 12488 12152 12584 12168
rect 12488 12088 12504 12152
rect 12568 12088 12584 12152
rect 12488 12072 12584 12088
rect 12488 12008 12504 12072
rect 12568 12008 12584 12072
rect 12488 11992 12584 12008
rect 11076 11892 11172 11928
rect 12488 11928 12504 11992
rect 12568 11928 12584 11992
rect 12907 12672 13629 12681
rect 12907 11968 12916 12672
rect 13620 11968 13629 12672
rect 12907 11959 13629 11968
rect 13900 12648 13916 12712
rect 13980 12648 13996 12712
rect 15312 12712 15408 12748
rect 13900 12632 13996 12648
rect 13900 12568 13916 12632
rect 13980 12568 13996 12632
rect 13900 12552 13996 12568
rect 13900 12488 13916 12552
rect 13980 12488 13996 12552
rect 13900 12472 13996 12488
rect 13900 12408 13916 12472
rect 13980 12408 13996 12472
rect 13900 12392 13996 12408
rect 13900 12328 13916 12392
rect 13980 12328 13996 12392
rect 13900 12312 13996 12328
rect 13900 12248 13916 12312
rect 13980 12248 13996 12312
rect 13900 12232 13996 12248
rect 13900 12168 13916 12232
rect 13980 12168 13996 12232
rect 13900 12152 13996 12168
rect 13900 12088 13916 12152
rect 13980 12088 13996 12152
rect 13900 12072 13996 12088
rect 13900 12008 13916 12072
rect 13980 12008 13996 12072
rect 13900 11992 13996 12008
rect 12488 11892 12584 11928
rect 13900 11928 13916 11992
rect 13980 11928 13996 11992
rect 14319 12672 15041 12681
rect 14319 11968 14328 12672
rect 15032 11968 15041 12672
rect 14319 11959 15041 11968
rect 15312 12648 15328 12712
rect 15392 12648 15408 12712
rect 16724 12712 16820 12748
rect 15312 12632 15408 12648
rect 15312 12568 15328 12632
rect 15392 12568 15408 12632
rect 15312 12552 15408 12568
rect 15312 12488 15328 12552
rect 15392 12488 15408 12552
rect 15312 12472 15408 12488
rect 15312 12408 15328 12472
rect 15392 12408 15408 12472
rect 15312 12392 15408 12408
rect 15312 12328 15328 12392
rect 15392 12328 15408 12392
rect 15312 12312 15408 12328
rect 15312 12248 15328 12312
rect 15392 12248 15408 12312
rect 15312 12232 15408 12248
rect 15312 12168 15328 12232
rect 15392 12168 15408 12232
rect 15312 12152 15408 12168
rect 15312 12088 15328 12152
rect 15392 12088 15408 12152
rect 15312 12072 15408 12088
rect 15312 12008 15328 12072
rect 15392 12008 15408 12072
rect 15312 11992 15408 12008
rect 13900 11892 13996 11928
rect 15312 11928 15328 11992
rect 15392 11928 15408 11992
rect 15731 12672 16453 12681
rect 15731 11968 15740 12672
rect 16444 11968 16453 12672
rect 15731 11959 16453 11968
rect 16724 12648 16740 12712
rect 16804 12648 16820 12712
rect 18136 12712 18232 12748
rect 16724 12632 16820 12648
rect 16724 12568 16740 12632
rect 16804 12568 16820 12632
rect 16724 12552 16820 12568
rect 16724 12488 16740 12552
rect 16804 12488 16820 12552
rect 16724 12472 16820 12488
rect 16724 12408 16740 12472
rect 16804 12408 16820 12472
rect 16724 12392 16820 12408
rect 16724 12328 16740 12392
rect 16804 12328 16820 12392
rect 16724 12312 16820 12328
rect 16724 12248 16740 12312
rect 16804 12248 16820 12312
rect 16724 12232 16820 12248
rect 16724 12168 16740 12232
rect 16804 12168 16820 12232
rect 16724 12152 16820 12168
rect 16724 12088 16740 12152
rect 16804 12088 16820 12152
rect 16724 12072 16820 12088
rect 16724 12008 16740 12072
rect 16804 12008 16820 12072
rect 16724 11992 16820 12008
rect 15312 11892 15408 11928
rect 16724 11928 16740 11992
rect 16804 11928 16820 11992
rect 17143 12672 17865 12681
rect 17143 11968 17152 12672
rect 17856 11968 17865 12672
rect 17143 11959 17865 11968
rect 18136 12648 18152 12712
rect 18216 12648 18232 12712
rect 19548 12712 19644 12748
rect 18136 12632 18232 12648
rect 18136 12568 18152 12632
rect 18216 12568 18232 12632
rect 18136 12552 18232 12568
rect 18136 12488 18152 12552
rect 18216 12488 18232 12552
rect 18136 12472 18232 12488
rect 18136 12408 18152 12472
rect 18216 12408 18232 12472
rect 18136 12392 18232 12408
rect 18136 12328 18152 12392
rect 18216 12328 18232 12392
rect 18136 12312 18232 12328
rect 18136 12248 18152 12312
rect 18216 12248 18232 12312
rect 18136 12232 18232 12248
rect 18136 12168 18152 12232
rect 18216 12168 18232 12232
rect 18136 12152 18232 12168
rect 18136 12088 18152 12152
rect 18216 12088 18232 12152
rect 18136 12072 18232 12088
rect 18136 12008 18152 12072
rect 18216 12008 18232 12072
rect 18136 11992 18232 12008
rect 16724 11892 16820 11928
rect 18136 11928 18152 11992
rect 18216 11928 18232 11992
rect 18555 12672 19277 12681
rect 18555 11968 18564 12672
rect 19268 11968 19277 12672
rect 18555 11959 19277 11968
rect 19548 12648 19564 12712
rect 19628 12648 19644 12712
rect 20960 12712 21056 12748
rect 19548 12632 19644 12648
rect 19548 12568 19564 12632
rect 19628 12568 19644 12632
rect 19548 12552 19644 12568
rect 19548 12488 19564 12552
rect 19628 12488 19644 12552
rect 19548 12472 19644 12488
rect 19548 12408 19564 12472
rect 19628 12408 19644 12472
rect 19548 12392 19644 12408
rect 19548 12328 19564 12392
rect 19628 12328 19644 12392
rect 19548 12312 19644 12328
rect 19548 12248 19564 12312
rect 19628 12248 19644 12312
rect 19548 12232 19644 12248
rect 19548 12168 19564 12232
rect 19628 12168 19644 12232
rect 19548 12152 19644 12168
rect 19548 12088 19564 12152
rect 19628 12088 19644 12152
rect 19548 12072 19644 12088
rect 19548 12008 19564 12072
rect 19628 12008 19644 12072
rect 19548 11992 19644 12008
rect 18136 11892 18232 11928
rect 19548 11928 19564 11992
rect 19628 11928 19644 11992
rect 19967 12672 20689 12681
rect 19967 11968 19976 12672
rect 20680 11968 20689 12672
rect 19967 11959 20689 11968
rect 20960 12648 20976 12712
rect 21040 12648 21056 12712
rect 22372 12712 22468 12748
rect 20960 12632 21056 12648
rect 20960 12568 20976 12632
rect 21040 12568 21056 12632
rect 20960 12552 21056 12568
rect 20960 12488 20976 12552
rect 21040 12488 21056 12552
rect 20960 12472 21056 12488
rect 20960 12408 20976 12472
rect 21040 12408 21056 12472
rect 20960 12392 21056 12408
rect 20960 12328 20976 12392
rect 21040 12328 21056 12392
rect 20960 12312 21056 12328
rect 20960 12248 20976 12312
rect 21040 12248 21056 12312
rect 20960 12232 21056 12248
rect 20960 12168 20976 12232
rect 21040 12168 21056 12232
rect 20960 12152 21056 12168
rect 20960 12088 20976 12152
rect 21040 12088 21056 12152
rect 20960 12072 21056 12088
rect 20960 12008 20976 12072
rect 21040 12008 21056 12072
rect 20960 11992 21056 12008
rect 19548 11892 19644 11928
rect 20960 11928 20976 11992
rect 21040 11928 21056 11992
rect 21379 12672 22101 12681
rect 21379 11968 21388 12672
rect 22092 11968 22101 12672
rect 21379 11959 22101 11968
rect 22372 12648 22388 12712
rect 22452 12648 22468 12712
rect 23784 12712 23880 12748
rect 22372 12632 22468 12648
rect 22372 12568 22388 12632
rect 22452 12568 22468 12632
rect 22372 12552 22468 12568
rect 22372 12488 22388 12552
rect 22452 12488 22468 12552
rect 22372 12472 22468 12488
rect 22372 12408 22388 12472
rect 22452 12408 22468 12472
rect 22372 12392 22468 12408
rect 22372 12328 22388 12392
rect 22452 12328 22468 12392
rect 22372 12312 22468 12328
rect 22372 12248 22388 12312
rect 22452 12248 22468 12312
rect 22372 12232 22468 12248
rect 22372 12168 22388 12232
rect 22452 12168 22468 12232
rect 22372 12152 22468 12168
rect 22372 12088 22388 12152
rect 22452 12088 22468 12152
rect 22372 12072 22468 12088
rect 22372 12008 22388 12072
rect 22452 12008 22468 12072
rect 22372 11992 22468 12008
rect 20960 11892 21056 11928
rect 22372 11928 22388 11992
rect 22452 11928 22468 11992
rect 22791 12672 23513 12681
rect 22791 11968 22800 12672
rect 23504 11968 23513 12672
rect 22791 11959 23513 11968
rect 23784 12648 23800 12712
rect 23864 12648 23880 12712
rect 23784 12632 23880 12648
rect 23784 12568 23800 12632
rect 23864 12568 23880 12632
rect 23784 12552 23880 12568
rect 23784 12488 23800 12552
rect 23864 12488 23880 12552
rect 23784 12472 23880 12488
rect 23784 12408 23800 12472
rect 23864 12408 23880 12472
rect 23784 12392 23880 12408
rect 23784 12328 23800 12392
rect 23864 12328 23880 12392
rect 23784 12312 23880 12328
rect 23784 12248 23800 12312
rect 23864 12248 23880 12312
rect 23784 12232 23880 12248
rect 23784 12168 23800 12232
rect 23864 12168 23880 12232
rect 23784 12152 23880 12168
rect 23784 12088 23800 12152
rect 23864 12088 23880 12152
rect 23784 12072 23880 12088
rect 23784 12008 23800 12072
rect 23864 12008 23880 12072
rect 23784 11992 23880 12008
rect 22372 11892 22468 11928
rect 23784 11928 23800 11992
rect 23864 11928 23880 11992
rect 23784 11892 23880 11928
rect -22812 11592 -22716 11628
rect -23805 11552 -23083 11561
rect -23805 10848 -23796 11552
rect -23092 10848 -23083 11552
rect -23805 10839 -23083 10848
rect -22812 11528 -22796 11592
rect -22732 11528 -22716 11592
rect -21400 11592 -21304 11628
rect -22812 11512 -22716 11528
rect -22812 11448 -22796 11512
rect -22732 11448 -22716 11512
rect -22812 11432 -22716 11448
rect -22812 11368 -22796 11432
rect -22732 11368 -22716 11432
rect -22812 11352 -22716 11368
rect -22812 11288 -22796 11352
rect -22732 11288 -22716 11352
rect -22812 11272 -22716 11288
rect -22812 11208 -22796 11272
rect -22732 11208 -22716 11272
rect -22812 11192 -22716 11208
rect -22812 11128 -22796 11192
rect -22732 11128 -22716 11192
rect -22812 11112 -22716 11128
rect -22812 11048 -22796 11112
rect -22732 11048 -22716 11112
rect -22812 11032 -22716 11048
rect -22812 10968 -22796 11032
rect -22732 10968 -22716 11032
rect -22812 10952 -22716 10968
rect -22812 10888 -22796 10952
rect -22732 10888 -22716 10952
rect -22812 10872 -22716 10888
rect -22812 10808 -22796 10872
rect -22732 10808 -22716 10872
rect -22393 11552 -21671 11561
rect -22393 10848 -22384 11552
rect -21680 10848 -21671 11552
rect -22393 10839 -21671 10848
rect -21400 11528 -21384 11592
rect -21320 11528 -21304 11592
rect -19988 11592 -19892 11628
rect -21400 11512 -21304 11528
rect -21400 11448 -21384 11512
rect -21320 11448 -21304 11512
rect -21400 11432 -21304 11448
rect -21400 11368 -21384 11432
rect -21320 11368 -21304 11432
rect -21400 11352 -21304 11368
rect -21400 11288 -21384 11352
rect -21320 11288 -21304 11352
rect -21400 11272 -21304 11288
rect -21400 11208 -21384 11272
rect -21320 11208 -21304 11272
rect -21400 11192 -21304 11208
rect -21400 11128 -21384 11192
rect -21320 11128 -21304 11192
rect -21400 11112 -21304 11128
rect -21400 11048 -21384 11112
rect -21320 11048 -21304 11112
rect -21400 11032 -21304 11048
rect -21400 10968 -21384 11032
rect -21320 10968 -21304 11032
rect -21400 10952 -21304 10968
rect -21400 10888 -21384 10952
rect -21320 10888 -21304 10952
rect -21400 10872 -21304 10888
rect -22812 10772 -22716 10808
rect -21400 10808 -21384 10872
rect -21320 10808 -21304 10872
rect -20981 11552 -20259 11561
rect -20981 10848 -20972 11552
rect -20268 10848 -20259 11552
rect -20981 10839 -20259 10848
rect -19988 11528 -19972 11592
rect -19908 11528 -19892 11592
rect -18576 11592 -18480 11628
rect -19988 11512 -19892 11528
rect -19988 11448 -19972 11512
rect -19908 11448 -19892 11512
rect -19988 11432 -19892 11448
rect -19988 11368 -19972 11432
rect -19908 11368 -19892 11432
rect -19988 11352 -19892 11368
rect -19988 11288 -19972 11352
rect -19908 11288 -19892 11352
rect -19988 11272 -19892 11288
rect -19988 11208 -19972 11272
rect -19908 11208 -19892 11272
rect -19988 11192 -19892 11208
rect -19988 11128 -19972 11192
rect -19908 11128 -19892 11192
rect -19988 11112 -19892 11128
rect -19988 11048 -19972 11112
rect -19908 11048 -19892 11112
rect -19988 11032 -19892 11048
rect -19988 10968 -19972 11032
rect -19908 10968 -19892 11032
rect -19988 10952 -19892 10968
rect -19988 10888 -19972 10952
rect -19908 10888 -19892 10952
rect -19988 10872 -19892 10888
rect -21400 10772 -21304 10808
rect -19988 10808 -19972 10872
rect -19908 10808 -19892 10872
rect -19569 11552 -18847 11561
rect -19569 10848 -19560 11552
rect -18856 10848 -18847 11552
rect -19569 10839 -18847 10848
rect -18576 11528 -18560 11592
rect -18496 11528 -18480 11592
rect -17164 11592 -17068 11628
rect -18576 11512 -18480 11528
rect -18576 11448 -18560 11512
rect -18496 11448 -18480 11512
rect -18576 11432 -18480 11448
rect -18576 11368 -18560 11432
rect -18496 11368 -18480 11432
rect -18576 11352 -18480 11368
rect -18576 11288 -18560 11352
rect -18496 11288 -18480 11352
rect -18576 11272 -18480 11288
rect -18576 11208 -18560 11272
rect -18496 11208 -18480 11272
rect -18576 11192 -18480 11208
rect -18576 11128 -18560 11192
rect -18496 11128 -18480 11192
rect -18576 11112 -18480 11128
rect -18576 11048 -18560 11112
rect -18496 11048 -18480 11112
rect -18576 11032 -18480 11048
rect -18576 10968 -18560 11032
rect -18496 10968 -18480 11032
rect -18576 10952 -18480 10968
rect -18576 10888 -18560 10952
rect -18496 10888 -18480 10952
rect -18576 10872 -18480 10888
rect -19988 10772 -19892 10808
rect -18576 10808 -18560 10872
rect -18496 10808 -18480 10872
rect -18157 11552 -17435 11561
rect -18157 10848 -18148 11552
rect -17444 10848 -17435 11552
rect -18157 10839 -17435 10848
rect -17164 11528 -17148 11592
rect -17084 11528 -17068 11592
rect -15752 11592 -15656 11628
rect -17164 11512 -17068 11528
rect -17164 11448 -17148 11512
rect -17084 11448 -17068 11512
rect -17164 11432 -17068 11448
rect -17164 11368 -17148 11432
rect -17084 11368 -17068 11432
rect -17164 11352 -17068 11368
rect -17164 11288 -17148 11352
rect -17084 11288 -17068 11352
rect -17164 11272 -17068 11288
rect -17164 11208 -17148 11272
rect -17084 11208 -17068 11272
rect -17164 11192 -17068 11208
rect -17164 11128 -17148 11192
rect -17084 11128 -17068 11192
rect -17164 11112 -17068 11128
rect -17164 11048 -17148 11112
rect -17084 11048 -17068 11112
rect -17164 11032 -17068 11048
rect -17164 10968 -17148 11032
rect -17084 10968 -17068 11032
rect -17164 10952 -17068 10968
rect -17164 10888 -17148 10952
rect -17084 10888 -17068 10952
rect -17164 10872 -17068 10888
rect -18576 10772 -18480 10808
rect -17164 10808 -17148 10872
rect -17084 10808 -17068 10872
rect -16745 11552 -16023 11561
rect -16745 10848 -16736 11552
rect -16032 10848 -16023 11552
rect -16745 10839 -16023 10848
rect -15752 11528 -15736 11592
rect -15672 11528 -15656 11592
rect -14340 11592 -14244 11628
rect -15752 11512 -15656 11528
rect -15752 11448 -15736 11512
rect -15672 11448 -15656 11512
rect -15752 11432 -15656 11448
rect -15752 11368 -15736 11432
rect -15672 11368 -15656 11432
rect -15752 11352 -15656 11368
rect -15752 11288 -15736 11352
rect -15672 11288 -15656 11352
rect -15752 11272 -15656 11288
rect -15752 11208 -15736 11272
rect -15672 11208 -15656 11272
rect -15752 11192 -15656 11208
rect -15752 11128 -15736 11192
rect -15672 11128 -15656 11192
rect -15752 11112 -15656 11128
rect -15752 11048 -15736 11112
rect -15672 11048 -15656 11112
rect -15752 11032 -15656 11048
rect -15752 10968 -15736 11032
rect -15672 10968 -15656 11032
rect -15752 10952 -15656 10968
rect -15752 10888 -15736 10952
rect -15672 10888 -15656 10952
rect -15752 10872 -15656 10888
rect -17164 10772 -17068 10808
rect -15752 10808 -15736 10872
rect -15672 10808 -15656 10872
rect -15333 11552 -14611 11561
rect -15333 10848 -15324 11552
rect -14620 10848 -14611 11552
rect -15333 10839 -14611 10848
rect -14340 11528 -14324 11592
rect -14260 11528 -14244 11592
rect -12928 11592 -12832 11628
rect -14340 11512 -14244 11528
rect -14340 11448 -14324 11512
rect -14260 11448 -14244 11512
rect -14340 11432 -14244 11448
rect -14340 11368 -14324 11432
rect -14260 11368 -14244 11432
rect -14340 11352 -14244 11368
rect -14340 11288 -14324 11352
rect -14260 11288 -14244 11352
rect -14340 11272 -14244 11288
rect -14340 11208 -14324 11272
rect -14260 11208 -14244 11272
rect -14340 11192 -14244 11208
rect -14340 11128 -14324 11192
rect -14260 11128 -14244 11192
rect -14340 11112 -14244 11128
rect -14340 11048 -14324 11112
rect -14260 11048 -14244 11112
rect -14340 11032 -14244 11048
rect -14340 10968 -14324 11032
rect -14260 10968 -14244 11032
rect -14340 10952 -14244 10968
rect -14340 10888 -14324 10952
rect -14260 10888 -14244 10952
rect -14340 10872 -14244 10888
rect -15752 10772 -15656 10808
rect -14340 10808 -14324 10872
rect -14260 10808 -14244 10872
rect -13921 11552 -13199 11561
rect -13921 10848 -13912 11552
rect -13208 10848 -13199 11552
rect -13921 10839 -13199 10848
rect -12928 11528 -12912 11592
rect -12848 11528 -12832 11592
rect -11516 11592 -11420 11628
rect -12928 11512 -12832 11528
rect -12928 11448 -12912 11512
rect -12848 11448 -12832 11512
rect -12928 11432 -12832 11448
rect -12928 11368 -12912 11432
rect -12848 11368 -12832 11432
rect -12928 11352 -12832 11368
rect -12928 11288 -12912 11352
rect -12848 11288 -12832 11352
rect -12928 11272 -12832 11288
rect -12928 11208 -12912 11272
rect -12848 11208 -12832 11272
rect -12928 11192 -12832 11208
rect -12928 11128 -12912 11192
rect -12848 11128 -12832 11192
rect -12928 11112 -12832 11128
rect -12928 11048 -12912 11112
rect -12848 11048 -12832 11112
rect -12928 11032 -12832 11048
rect -12928 10968 -12912 11032
rect -12848 10968 -12832 11032
rect -12928 10952 -12832 10968
rect -12928 10888 -12912 10952
rect -12848 10888 -12832 10952
rect -12928 10872 -12832 10888
rect -14340 10772 -14244 10808
rect -12928 10808 -12912 10872
rect -12848 10808 -12832 10872
rect -12509 11552 -11787 11561
rect -12509 10848 -12500 11552
rect -11796 10848 -11787 11552
rect -12509 10839 -11787 10848
rect -11516 11528 -11500 11592
rect -11436 11528 -11420 11592
rect -10104 11592 -10008 11628
rect -11516 11512 -11420 11528
rect -11516 11448 -11500 11512
rect -11436 11448 -11420 11512
rect -11516 11432 -11420 11448
rect -11516 11368 -11500 11432
rect -11436 11368 -11420 11432
rect -11516 11352 -11420 11368
rect -11516 11288 -11500 11352
rect -11436 11288 -11420 11352
rect -11516 11272 -11420 11288
rect -11516 11208 -11500 11272
rect -11436 11208 -11420 11272
rect -11516 11192 -11420 11208
rect -11516 11128 -11500 11192
rect -11436 11128 -11420 11192
rect -11516 11112 -11420 11128
rect -11516 11048 -11500 11112
rect -11436 11048 -11420 11112
rect -11516 11032 -11420 11048
rect -11516 10968 -11500 11032
rect -11436 10968 -11420 11032
rect -11516 10952 -11420 10968
rect -11516 10888 -11500 10952
rect -11436 10888 -11420 10952
rect -11516 10872 -11420 10888
rect -12928 10772 -12832 10808
rect -11516 10808 -11500 10872
rect -11436 10808 -11420 10872
rect -11097 11552 -10375 11561
rect -11097 10848 -11088 11552
rect -10384 10848 -10375 11552
rect -11097 10839 -10375 10848
rect -10104 11528 -10088 11592
rect -10024 11528 -10008 11592
rect -8692 11592 -8596 11628
rect -10104 11512 -10008 11528
rect -10104 11448 -10088 11512
rect -10024 11448 -10008 11512
rect -10104 11432 -10008 11448
rect -10104 11368 -10088 11432
rect -10024 11368 -10008 11432
rect -10104 11352 -10008 11368
rect -10104 11288 -10088 11352
rect -10024 11288 -10008 11352
rect -10104 11272 -10008 11288
rect -10104 11208 -10088 11272
rect -10024 11208 -10008 11272
rect -10104 11192 -10008 11208
rect -10104 11128 -10088 11192
rect -10024 11128 -10008 11192
rect -10104 11112 -10008 11128
rect -10104 11048 -10088 11112
rect -10024 11048 -10008 11112
rect -10104 11032 -10008 11048
rect -10104 10968 -10088 11032
rect -10024 10968 -10008 11032
rect -10104 10952 -10008 10968
rect -10104 10888 -10088 10952
rect -10024 10888 -10008 10952
rect -10104 10872 -10008 10888
rect -11516 10772 -11420 10808
rect -10104 10808 -10088 10872
rect -10024 10808 -10008 10872
rect -9685 11552 -8963 11561
rect -9685 10848 -9676 11552
rect -8972 10848 -8963 11552
rect -9685 10839 -8963 10848
rect -8692 11528 -8676 11592
rect -8612 11528 -8596 11592
rect -7280 11592 -7184 11628
rect -8692 11512 -8596 11528
rect -8692 11448 -8676 11512
rect -8612 11448 -8596 11512
rect -8692 11432 -8596 11448
rect -8692 11368 -8676 11432
rect -8612 11368 -8596 11432
rect -8692 11352 -8596 11368
rect -8692 11288 -8676 11352
rect -8612 11288 -8596 11352
rect -8692 11272 -8596 11288
rect -8692 11208 -8676 11272
rect -8612 11208 -8596 11272
rect -8692 11192 -8596 11208
rect -8692 11128 -8676 11192
rect -8612 11128 -8596 11192
rect -8692 11112 -8596 11128
rect -8692 11048 -8676 11112
rect -8612 11048 -8596 11112
rect -8692 11032 -8596 11048
rect -8692 10968 -8676 11032
rect -8612 10968 -8596 11032
rect -8692 10952 -8596 10968
rect -8692 10888 -8676 10952
rect -8612 10888 -8596 10952
rect -8692 10872 -8596 10888
rect -10104 10772 -10008 10808
rect -8692 10808 -8676 10872
rect -8612 10808 -8596 10872
rect -8273 11552 -7551 11561
rect -8273 10848 -8264 11552
rect -7560 10848 -7551 11552
rect -8273 10839 -7551 10848
rect -7280 11528 -7264 11592
rect -7200 11528 -7184 11592
rect -5868 11592 -5772 11628
rect -7280 11512 -7184 11528
rect -7280 11448 -7264 11512
rect -7200 11448 -7184 11512
rect -7280 11432 -7184 11448
rect -7280 11368 -7264 11432
rect -7200 11368 -7184 11432
rect -7280 11352 -7184 11368
rect -7280 11288 -7264 11352
rect -7200 11288 -7184 11352
rect -7280 11272 -7184 11288
rect -7280 11208 -7264 11272
rect -7200 11208 -7184 11272
rect -7280 11192 -7184 11208
rect -7280 11128 -7264 11192
rect -7200 11128 -7184 11192
rect -7280 11112 -7184 11128
rect -7280 11048 -7264 11112
rect -7200 11048 -7184 11112
rect -7280 11032 -7184 11048
rect -7280 10968 -7264 11032
rect -7200 10968 -7184 11032
rect -7280 10952 -7184 10968
rect -7280 10888 -7264 10952
rect -7200 10888 -7184 10952
rect -7280 10872 -7184 10888
rect -8692 10772 -8596 10808
rect -7280 10808 -7264 10872
rect -7200 10808 -7184 10872
rect -6861 11552 -6139 11561
rect -6861 10848 -6852 11552
rect -6148 10848 -6139 11552
rect -6861 10839 -6139 10848
rect -5868 11528 -5852 11592
rect -5788 11528 -5772 11592
rect -4456 11592 -4360 11628
rect -5868 11512 -5772 11528
rect -5868 11448 -5852 11512
rect -5788 11448 -5772 11512
rect -5868 11432 -5772 11448
rect -5868 11368 -5852 11432
rect -5788 11368 -5772 11432
rect -5868 11352 -5772 11368
rect -5868 11288 -5852 11352
rect -5788 11288 -5772 11352
rect -5868 11272 -5772 11288
rect -5868 11208 -5852 11272
rect -5788 11208 -5772 11272
rect -5868 11192 -5772 11208
rect -5868 11128 -5852 11192
rect -5788 11128 -5772 11192
rect -5868 11112 -5772 11128
rect -5868 11048 -5852 11112
rect -5788 11048 -5772 11112
rect -5868 11032 -5772 11048
rect -5868 10968 -5852 11032
rect -5788 10968 -5772 11032
rect -5868 10952 -5772 10968
rect -5868 10888 -5852 10952
rect -5788 10888 -5772 10952
rect -5868 10872 -5772 10888
rect -7280 10772 -7184 10808
rect -5868 10808 -5852 10872
rect -5788 10808 -5772 10872
rect -5449 11552 -4727 11561
rect -5449 10848 -5440 11552
rect -4736 10848 -4727 11552
rect -5449 10839 -4727 10848
rect -4456 11528 -4440 11592
rect -4376 11528 -4360 11592
rect -3044 11592 -2948 11628
rect -4456 11512 -4360 11528
rect -4456 11448 -4440 11512
rect -4376 11448 -4360 11512
rect -4456 11432 -4360 11448
rect -4456 11368 -4440 11432
rect -4376 11368 -4360 11432
rect -4456 11352 -4360 11368
rect -4456 11288 -4440 11352
rect -4376 11288 -4360 11352
rect -4456 11272 -4360 11288
rect -4456 11208 -4440 11272
rect -4376 11208 -4360 11272
rect -4456 11192 -4360 11208
rect -4456 11128 -4440 11192
rect -4376 11128 -4360 11192
rect -4456 11112 -4360 11128
rect -4456 11048 -4440 11112
rect -4376 11048 -4360 11112
rect -4456 11032 -4360 11048
rect -4456 10968 -4440 11032
rect -4376 10968 -4360 11032
rect -4456 10952 -4360 10968
rect -4456 10888 -4440 10952
rect -4376 10888 -4360 10952
rect -4456 10872 -4360 10888
rect -5868 10772 -5772 10808
rect -4456 10808 -4440 10872
rect -4376 10808 -4360 10872
rect -4037 11552 -3315 11561
rect -4037 10848 -4028 11552
rect -3324 10848 -3315 11552
rect -4037 10839 -3315 10848
rect -3044 11528 -3028 11592
rect -2964 11528 -2948 11592
rect -1632 11592 -1536 11628
rect -3044 11512 -2948 11528
rect -3044 11448 -3028 11512
rect -2964 11448 -2948 11512
rect -3044 11432 -2948 11448
rect -3044 11368 -3028 11432
rect -2964 11368 -2948 11432
rect -3044 11352 -2948 11368
rect -3044 11288 -3028 11352
rect -2964 11288 -2948 11352
rect -3044 11272 -2948 11288
rect -3044 11208 -3028 11272
rect -2964 11208 -2948 11272
rect -3044 11192 -2948 11208
rect -3044 11128 -3028 11192
rect -2964 11128 -2948 11192
rect -3044 11112 -2948 11128
rect -3044 11048 -3028 11112
rect -2964 11048 -2948 11112
rect -3044 11032 -2948 11048
rect -3044 10968 -3028 11032
rect -2964 10968 -2948 11032
rect -3044 10952 -2948 10968
rect -3044 10888 -3028 10952
rect -2964 10888 -2948 10952
rect -3044 10872 -2948 10888
rect -4456 10772 -4360 10808
rect -3044 10808 -3028 10872
rect -2964 10808 -2948 10872
rect -2625 11552 -1903 11561
rect -2625 10848 -2616 11552
rect -1912 10848 -1903 11552
rect -2625 10839 -1903 10848
rect -1632 11528 -1616 11592
rect -1552 11528 -1536 11592
rect -220 11592 -124 11628
rect -1632 11512 -1536 11528
rect -1632 11448 -1616 11512
rect -1552 11448 -1536 11512
rect -1632 11432 -1536 11448
rect -1632 11368 -1616 11432
rect -1552 11368 -1536 11432
rect -1632 11352 -1536 11368
rect -1632 11288 -1616 11352
rect -1552 11288 -1536 11352
rect -1632 11272 -1536 11288
rect -1632 11208 -1616 11272
rect -1552 11208 -1536 11272
rect -1632 11192 -1536 11208
rect -1632 11128 -1616 11192
rect -1552 11128 -1536 11192
rect -1632 11112 -1536 11128
rect -1632 11048 -1616 11112
rect -1552 11048 -1536 11112
rect -1632 11032 -1536 11048
rect -1632 10968 -1616 11032
rect -1552 10968 -1536 11032
rect -1632 10952 -1536 10968
rect -1632 10888 -1616 10952
rect -1552 10888 -1536 10952
rect -1632 10872 -1536 10888
rect -3044 10772 -2948 10808
rect -1632 10808 -1616 10872
rect -1552 10808 -1536 10872
rect -1213 11552 -491 11561
rect -1213 10848 -1204 11552
rect -500 10848 -491 11552
rect -1213 10839 -491 10848
rect -220 11528 -204 11592
rect -140 11528 -124 11592
rect 1192 11592 1288 11628
rect -220 11512 -124 11528
rect -220 11448 -204 11512
rect -140 11448 -124 11512
rect -220 11432 -124 11448
rect -220 11368 -204 11432
rect -140 11368 -124 11432
rect -220 11352 -124 11368
rect -220 11288 -204 11352
rect -140 11288 -124 11352
rect -220 11272 -124 11288
rect -220 11208 -204 11272
rect -140 11208 -124 11272
rect -220 11192 -124 11208
rect -220 11128 -204 11192
rect -140 11128 -124 11192
rect -220 11112 -124 11128
rect -220 11048 -204 11112
rect -140 11048 -124 11112
rect -220 11032 -124 11048
rect -220 10968 -204 11032
rect -140 10968 -124 11032
rect -220 10952 -124 10968
rect -220 10888 -204 10952
rect -140 10888 -124 10952
rect -220 10872 -124 10888
rect -1632 10772 -1536 10808
rect -220 10808 -204 10872
rect -140 10808 -124 10872
rect 199 11552 921 11561
rect 199 10848 208 11552
rect 912 10848 921 11552
rect 199 10839 921 10848
rect 1192 11528 1208 11592
rect 1272 11528 1288 11592
rect 2604 11592 2700 11628
rect 1192 11512 1288 11528
rect 1192 11448 1208 11512
rect 1272 11448 1288 11512
rect 1192 11432 1288 11448
rect 1192 11368 1208 11432
rect 1272 11368 1288 11432
rect 1192 11352 1288 11368
rect 1192 11288 1208 11352
rect 1272 11288 1288 11352
rect 1192 11272 1288 11288
rect 1192 11208 1208 11272
rect 1272 11208 1288 11272
rect 1192 11192 1288 11208
rect 1192 11128 1208 11192
rect 1272 11128 1288 11192
rect 1192 11112 1288 11128
rect 1192 11048 1208 11112
rect 1272 11048 1288 11112
rect 1192 11032 1288 11048
rect 1192 10968 1208 11032
rect 1272 10968 1288 11032
rect 1192 10952 1288 10968
rect 1192 10888 1208 10952
rect 1272 10888 1288 10952
rect 1192 10872 1288 10888
rect -220 10772 -124 10808
rect 1192 10808 1208 10872
rect 1272 10808 1288 10872
rect 1611 11552 2333 11561
rect 1611 10848 1620 11552
rect 2324 10848 2333 11552
rect 1611 10839 2333 10848
rect 2604 11528 2620 11592
rect 2684 11528 2700 11592
rect 4016 11592 4112 11628
rect 2604 11512 2700 11528
rect 2604 11448 2620 11512
rect 2684 11448 2700 11512
rect 2604 11432 2700 11448
rect 2604 11368 2620 11432
rect 2684 11368 2700 11432
rect 2604 11352 2700 11368
rect 2604 11288 2620 11352
rect 2684 11288 2700 11352
rect 2604 11272 2700 11288
rect 2604 11208 2620 11272
rect 2684 11208 2700 11272
rect 2604 11192 2700 11208
rect 2604 11128 2620 11192
rect 2684 11128 2700 11192
rect 2604 11112 2700 11128
rect 2604 11048 2620 11112
rect 2684 11048 2700 11112
rect 2604 11032 2700 11048
rect 2604 10968 2620 11032
rect 2684 10968 2700 11032
rect 2604 10952 2700 10968
rect 2604 10888 2620 10952
rect 2684 10888 2700 10952
rect 2604 10872 2700 10888
rect 1192 10772 1288 10808
rect 2604 10808 2620 10872
rect 2684 10808 2700 10872
rect 3023 11552 3745 11561
rect 3023 10848 3032 11552
rect 3736 10848 3745 11552
rect 3023 10839 3745 10848
rect 4016 11528 4032 11592
rect 4096 11528 4112 11592
rect 5428 11592 5524 11628
rect 4016 11512 4112 11528
rect 4016 11448 4032 11512
rect 4096 11448 4112 11512
rect 4016 11432 4112 11448
rect 4016 11368 4032 11432
rect 4096 11368 4112 11432
rect 4016 11352 4112 11368
rect 4016 11288 4032 11352
rect 4096 11288 4112 11352
rect 4016 11272 4112 11288
rect 4016 11208 4032 11272
rect 4096 11208 4112 11272
rect 4016 11192 4112 11208
rect 4016 11128 4032 11192
rect 4096 11128 4112 11192
rect 4016 11112 4112 11128
rect 4016 11048 4032 11112
rect 4096 11048 4112 11112
rect 4016 11032 4112 11048
rect 4016 10968 4032 11032
rect 4096 10968 4112 11032
rect 4016 10952 4112 10968
rect 4016 10888 4032 10952
rect 4096 10888 4112 10952
rect 4016 10872 4112 10888
rect 2604 10772 2700 10808
rect 4016 10808 4032 10872
rect 4096 10808 4112 10872
rect 4435 11552 5157 11561
rect 4435 10848 4444 11552
rect 5148 10848 5157 11552
rect 4435 10839 5157 10848
rect 5428 11528 5444 11592
rect 5508 11528 5524 11592
rect 6840 11592 6936 11628
rect 5428 11512 5524 11528
rect 5428 11448 5444 11512
rect 5508 11448 5524 11512
rect 5428 11432 5524 11448
rect 5428 11368 5444 11432
rect 5508 11368 5524 11432
rect 5428 11352 5524 11368
rect 5428 11288 5444 11352
rect 5508 11288 5524 11352
rect 5428 11272 5524 11288
rect 5428 11208 5444 11272
rect 5508 11208 5524 11272
rect 5428 11192 5524 11208
rect 5428 11128 5444 11192
rect 5508 11128 5524 11192
rect 5428 11112 5524 11128
rect 5428 11048 5444 11112
rect 5508 11048 5524 11112
rect 5428 11032 5524 11048
rect 5428 10968 5444 11032
rect 5508 10968 5524 11032
rect 5428 10952 5524 10968
rect 5428 10888 5444 10952
rect 5508 10888 5524 10952
rect 5428 10872 5524 10888
rect 4016 10772 4112 10808
rect 5428 10808 5444 10872
rect 5508 10808 5524 10872
rect 5847 11552 6569 11561
rect 5847 10848 5856 11552
rect 6560 10848 6569 11552
rect 5847 10839 6569 10848
rect 6840 11528 6856 11592
rect 6920 11528 6936 11592
rect 8252 11592 8348 11628
rect 6840 11512 6936 11528
rect 6840 11448 6856 11512
rect 6920 11448 6936 11512
rect 6840 11432 6936 11448
rect 6840 11368 6856 11432
rect 6920 11368 6936 11432
rect 6840 11352 6936 11368
rect 6840 11288 6856 11352
rect 6920 11288 6936 11352
rect 6840 11272 6936 11288
rect 6840 11208 6856 11272
rect 6920 11208 6936 11272
rect 6840 11192 6936 11208
rect 6840 11128 6856 11192
rect 6920 11128 6936 11192
rect 6840 11112 6936 11128
rect 6840 11048 6856 11112
rect 6920 11048 6936 11112
rect 6840 11032 6936 11048
rect 6840 10968 6856 11032
rect 6920 10968 6936 11032
rect 6840 10952 6936 10968
rect 6840 10888 6856 10952
rect 6920 10888 6936 10952
rect 6840 10872 6936 10888
rect 5428 10772 5524 10808
rect 6840 10808 6856 10872
rect 6920 10808 6936 10872
rect 7259 11552 7981 11561
rect 7259 10848 7268 11552
rect 7972 10848 7981 11552
rect 7259 10839 7981 10848
rect 8252 11528 8268 11592
rect 8332 11528 8348 11592
rect 9664 11592 9760 11628
rect 8252 11512 8348 11528
rect 8252 11448 8268 11512
rect 8332 11448 8348 11512
rect 8252 11432 8348 11448
rect 8252 11368 8268 11432
rect 8332 11368 8348 11432
rect 8252 11352 8348 11368
rect 8252 11288 8268 11352
rect 8332 11288 8348 11352
rect 8252 11272 8348 11288
rect 8252 11208 8268 11272
rect 8332 11208 8348 11272
rect 8252 11192 8348 11208
rect 8252 11128 8268 11192
rect 8332 11128 8348 11192
rect 8252 11112 8348 11128
rect 8252 11048 8268 11112
rect 8332 11048 8348 11112
rect 8252 11032 8348 11048
rect 8252 10968 8268 11032
rect 8332 10968 8348 11032
rect 8252 10952 8348 10968
rect 8252 10888 8268 10952
rect 8332 10888 8348 10952
rect 8252 10872 8348 10888
rect 6840 10772 6936 10808
rect 8252 10808 8268 10872
rect 8332 10808 8348 10872
rect 8671 11552 9393 11561
rect 8671 10848 8680 11552
rect 9384 10848 9393 11552
rect 8671 10839 9393 10848
rect 9664 11528 9680 11592
rect 9744 11528 9760 11592
rect 11076 11592 11172 11628
rect 9664 11512 9760 11528
rect 9664 11448 9680 11512
rect 9744 11448 9760 11512
rect 9664 11432 9760 11448
rect 9664 11368 9680 11432
rect 9744 11368 9760 11432
rect 9664 11352 9760 11368
rect 9664 11288 9680 11352
rect 9744 11288 9760 11352
rect 9664 11272 9760 11288
rect 9664 11208 9680 11272
rect 9744 11208 9760 11272
rect 9664 11192 9760 11208
rect 9664 11128 9680 11192
rect 9744 11128 9760 11192
rect 9664 11112 9760 11128
rect 9664 11048 9680 11112
rect 9744 11048 9760 11112
rect 9664 11032 9760 11048
rect 9664 10968 9680 11032
rect 9744 10968 9760 11032
rect 9664 10952 9760 10968
rect 9664 10888 9680 10952
rect 9744 10888 9760 10952
rect 9664 10872 9760 10888
rect 8252 10772 8348 10808
rect 9664 10808 9680 10872
rect 9744 10808 9760 10872
rect 10083 11552 10805 11561
rect 10083 10848 10092 11552
rect 10796 10848 10805 11552
rect 10083 10839 10805 10848
rect 11076 11528 11092 11592
rect 11156 11528 11172 11592
rect 12488 11592 12584 11628
rect 11076 11512 11172 11528
rect 11076 11448 11092 11512
rect 11156 11448 11172 11512
rect 11076 11432 11172 11448
rect 11076 11368 11092 11432
rect 11156 11368 11172 11432
rect 11076 11352 11172 11368
rect 11076 11288 11092 11352
rect 11156 11288 11172 11352
rect 11076 11272 11172 11288
rect 11076 11208 11092 11272
rect 11156 11208 11172 11272
rect 11076 11192 11172 11208
rect 11076 11128 11092 11192
rect 11156 11128 11172 11192
rect 11076 11112 11172 11128
rect 11076 11048 11092 11112
rect 11156 11048 11172 11112
rect 11076 11032 11172 11048
rect 11076 10968 11092 11032
rect 11156 10968 11172 11032
rect 11076 10952 11172 10968
rect 11076 10888 11092 10952
rect 11156 10888 11172 10952
rect 11076 10872 11172 10888
rect 9664 10772 9760 10808
rect 11076 10808 11092 10872
rect 11156 10808 11172 10872
rect 11495 11552 12217 11561
rect 11495 10848 11504 11552
rect 12208 10848 12217 11552
rect 11495 10839 12217 10848
rect 12488 11528 12504 11592
rect 12568 11528 12584 11592
rect 13900 11592 13996 11628
rect 12488 11512 12584 11528
rect 12488 11448 12504 11512
rect 12568 11448 12584 11512
rect 12488 11432 12584 11448
rect 12488 11368 12504 11432
rect 12568 11368 12584 11432
rect 12488 11352 12584 11368
rect 12488 11288 12504 11352
rect 12568 11288 12584 11352
rect 12488 11272 12584 11288
rect 12488 11208 12504 11272
rect 12568 11208 12584 11272
rect 12488 11192 12584 11208
rect 12488 11128 12504 11192
rect 12568 11128 12584 11192
rect 12488 11112 12584 11128
rect 12488 11048 12504 11112
rect 12568 11048 12584 11112
rect 12488 11032 12584 11048
rect 12488 10968 12504 11032
rect 12568 10968 12584 11032
rect 12488 10952 12584 10968
rect 12488 10888 12504 10952
rect 12568 10888 12584 10952
rect 12488 10872 12584 10888
rect 11076 10772 11172 10808
rect 12488 10808 12504 10872
rect 12568 10808 12584 10872
rect 12907 11552 13629 11561
rect 12907 10848 12916 11552
rect 13620 10848 13629 11552
rect 12907 10839 13629 10848
rect 13900 11528 13916 11592
rect 13980 11528 13996 11592
rect 15312 11592 15408 11628
rect 13900 11512 13996 11528
rect 13900 11448 13916 11512
rect 13980 11448 13996 11512
rect 13900 11432 13996 11448
rect 13900 11368 13916 11432
rect 13980 11368 13996 11432
rect 13900 11352 13996 11368
rect 13900 11288 13916 11352
rect 13980 11288 13996 11352
rect 13900 11272 13996 11288
rect 13900 11208 13916 11272
rect 13980 11208 13996 11272
rect 13900 11192 13996 11208
rect 13900 11128 13916 11192
rect 13980 11128 13996 11192
rect 13900 11112 13996 11128
rect 13900 11048 13916 11112
rect 13980 11048 13996 11112
rect 13900 11032 13996 11048
rect 13900 10968 13916 11032
rect 13980 10968 13996 11032
rect 13900 10952 13996 10968
rect 13900 10888 13916 10952
rect 13980 10888 13996 10952
rect 13900 10872 13996 10888
rect 12488 10772 12584 10808
rect 13900 10808 13916 10872
rect 13980 10808 13996 10872
rect 14319 11552 15041 11561
rect 14319 10848 14328 11552
rect 15032 10848 15041 11552
rect 14319 10839 15041 10848
rect 15312 11528 15328 11592
rect 15392 11528 15408 11592
rect 16724 11592 16820 11628
rect 15312 11512 15408 11528
rect 15312 11448 15328 11512
rect 15392 11448 15408 11512
rect 15312 11432 15408 11448
rect 15312 11368 15328 11432
rect 15392 11368 15408 11432
rect 15312 11352 15408 11368
rect 15312 11288 15328 11352
rect 15392 11288 15408 11352
rect 15312 11272 15408 11288
rect 15312 11208 15328 11272
rect 15392 11208 15408 11272
rect 15312 11192 15408 11208
rect 15312 11128 15328 11192
rect 15392 11128 15408 11192
rect 15312 11112 15408 11128
rect 15312 11048 15328 11112
rect 15392 11048 15408 11112
rect 15312 11032 15408 11048
rect 15312 10968 15328 11032
rect 15392 10968 15408 11032
rect 15312 10952 15408 10968
rect 15312 10888 15328 10952
rect 15392 10888 15408 10952
rect 15312 10872 15408 10888
rect 13900 10772 13996 10808
rect 15312 10808 15328 10872
rect 15392 10808 15408 10872
rect 15731 11552 16453 11561
rect 15731 10848 15740 11552
rect 16444 10848 16453 11552
rect 15731 10839 16453 10848
rect 16724 11528 16740 11592
rect 16804 11528 16820 11592
rect 18136 11592 18232 11628
rect 16724 11512 16820 11528
rect 16724 11448 16740 11512
rect 16804 11448 16820 11512
rect 16724 11432 16820 11448
rect 16724 11368 16740 11432
rect 16804 11368 16820 11432
rect 16724 11352 16820 11368
rect 16724 11288 16740 11352
rect 16804 11288 16820 11352
rect 16724 11272 16820 11288
rect 16724 11208 16740 11272
rect 16804 11208 16820 11272
rect 16724 11192 16820 11208
rect 16724 11128 16740 11192
rect 16804 11128 16820 11192
rect 16724 11112 16820 11128
rect 16724 11048 16740 11112
rect 16804 11048 16820 11112
rect 16724 11032 16820 11048
rect 16724 10968 16740 11032
rect 16804 10968 16820 11032
rect 16724 10952 16820 10968
rect 16724 10888 16740 10952
rect 16804 10888 16820 10952
rect 16724 10872 16820 10888
rect 15312 10772 15408 10808
rect 16724 10808 16740 10872
rect 16804 10808 16820 10872
rect 17143 11552 17865 11561
rect 17143 10848 17152 11552
rect 17856 10848 17865 11552
rect 17143 10839 17865 10848
rect 18136 11528 18152 11592
rect 18216 11528 18232 11592
rect 19548 11592 19644 11628
rect 18136 11512 18232 11528
rect 18136 11448 18152 11512
rect 18216 11448 18232 11512
rect 18136 11432 18232 11448
rect 18136 11368 18152 11432
rect 18216 11368 18232 11432
rect 18136 11352 18232 11368
rect 18136 11288 18152 11352
rect 18216 11288 18232 11352
rect 18136 11272 18232 11288
rect 18136 11208 18152 11272
rect 18216 11208 18232 11272
rect 18136 11192 18232 11208
rect 18136 11128 18152 11192
rect 18216 11128 18232 11192
rect 18136 11112 18232 11128
rect 18136 11048 18152 11112
rect 18216 11048 18232 11112
rect 18136 11032 18232 11048
rect 18136 10968 18152 11032
rect 18216 10968 18232 11032
rect 18136 10952 18232 10968
rect 18136 10888 18152 10952
rect 18216 10888 18232 10952
rect 18136 10872 18232 10888
rect 16724 10772 16820 10808
rect 18136 10808 18152 10872
rect 18216 10808 18232 10872
rect 18555 11552 19277 11561
rect 18555 10848 18564 11552
rect 19268 10848 19277 11552
rect 18555 10839 19277 10848
rect 19548 11528 19564 11592
rect 19628 11528 19644 11592
rect 20960 11592 21056 11628
rect 19548 11512 19644 11528
rect 19548 11448 19564 11512
rect 19628 11448 19644 11512
rect 19548 11432 19644 11448
rect 19548 11368 19564 11432
rect 19628 11368 19644 11432
rect 19548 11352 19644 11368
rect 19548 11288 19564 11352
rect 19628 11288 19644 11352
rect 19548 11272 19644 11288
rect 19548 11208 19564 11272
rect 19628 11208 19644 11272
rect 19548 11192 19644 11208
rect 19548 11128 19564 11192
rect 19628 11128 19644 11192
rect 19548 11112 19644 11128
rect 19548 11048 19564 11112
rect 19628 11048 19644 11112
rect 19548 11032 19644 11048
rect 19548 10968 19564 11032
rect 19628 10968 19644 11032
rect 19548 10952 19644 10968
rect 19548 10888 19564 10952
rect 19628 10888 19644 10952
rect 19548 10872 19644 10888
rect 18136 10772 18232 10808
rect 19548 10808 19564 10872
rect 19628 10808 19644 10872
rect 19967 11552 20689 11561
rect 19967 10848 19976 11552
rect 20680 10848 20689 11552
rect 19967 10839 20689 10848
rect 20960 11528 20976 11592
rect 21040 11528 21056 11592
rect 22372 11592 22468 11628
rect 20960 11512 21056 11528
rect 20960 11448 20976 11512
rect 21040 11448 21056 11512
rect 20960 11432 21056 11448
rect 20960 11368 20976 11432
rect 21040 11368 21056 11432
rect 20960 11352 21056 11368
rect 20960 11288 20976 11352
rect 21040 11288 21056 11352
rect 20960 11272 21056 11288
rect 20960 11208 20976 11272
rect 21040 11208 21056 11272
rect 20960 11192 21056 11208
rect 20960 11128 20976 11192
rect 21040 11128 21056 11192
rect 20960 11112 21056 11128
rect 20960 11048 20976 11112
rect 21040 11048 21056 11112
rect 20960 11032 21056 11048
rect 20960 10968 20976 11032
rect 21040 10968 21056 11032
rect 20960 10952 21056 10968
rect 20960 10888 20976 10952
rect 21040 10888 21056 10952
rect 20960 10872 21056 10888
rect 19548 10772 19644 10808
rect 20960 10808 20976 10872
rect 21040 10808 21056 10872
rect 21379 11552 22101 11561
rect 21379 10848 21388 11552
rect 22092 10848 22101 11552
rect 21379 10839 22101 10848
rect 22372 11528 22388 11592
rect 22452 11528 22468 11592
rect 23784 11592 23880 11628
rect 22372 11512 22468 11528
rect 22372 11448 22388 11512
rect 22452 11448 22468 11512
rect 22372 11432 22468 11448
rect 22372 11368 22388 11432
rect 22452 11368 22468 11432
rect 22372 11352 22468 11368
rect 22372 11288 22388 11352
rect 22452 11288 22468 11352
rect 22372 11272 22468 11288
rect 22372 11208 22388 11272
rect 22452 11208 22468 11272
rect 22372 11192 22468 11208
rect 22372 11128 22388 11192
rect 22452 11128 22468 11192
rect 22372 11112 22468 11128
rect 22372 11048 22388 11112
rect 22452 11048 22468 11112
rect 22372 11032 22468 11048
rect 22372 10968 22388 11032
rect 22452 10968 22468 11032
rect 22372 10952 22468 10968
rect 22372 10888 22388 10952
rect 22452 10888 22468 10952
rect 22372 10872 22468 10888
rect 20960 10772 21056 10808
rect 22372 10808 22388 10872
rect 22452 10808 22468 10872
rect 22791 11552 23513 11561
rect 22791 10848 22800 11552
rect 23504 10848 23513 11552
rect 22791 10839 23513 10848
rect 23784 11528 23800 11592
rect 23864 11528 23880 11592
rect 23784 11512 23880 11528
rect 23784 11448 23800 11512
rect 23864 11448 23880 11512
rect 23784 11432 23880 11448
rect 23784 11368 23800 11432
rect 23864 11368 23880 11432
rect 23784 11352 23880 11368
rect 23784 11288 23800 11352
rect 23864 11288 23880 11352
rect 23784 11272 23880 11288
rect 23784 11208 23800 11272
rect 23864 11208 23880 11272
rect 23784 11192 23880 11208
rect 23784 11128 23800 11192
rect 23864 11128 23880 11192
rect 23784 11112 23880 11128
rect 23784 11048 23800 11112
rect 23864 11048 23880 11112
rect 23784 11032 23880 11048
rect 23784 10968 23800 11032
rect 23864 10968 23880 11032
rect 23784 10952 23880 10968
rect 23784 10888 23800 10952
rect 23864 10888 23880 10952
rect 23784 10872 23880 10888
rect 22372 10772 22468 10808
rect 23784 10808 23800 10872
rect 23864 10808 23880 10872
rect 23784 10772 23880 10808
rect -22812 10472 -22716 10508
rect -23805 10432 -23083 10441
rect -23805 9728 -23796 10432
rect -23092 9728 -23083 10432
rect -23805 9719 -23083 9728
rect -22812 10408 -22796 10472
rect -22732 10408 -22716 10472
rect -21400 10472 -21304 10508
rect -22812 10392 -22716 10408
rect -22812 10328 -22796 10392
rect -22732 10328 -22716 10392
rect -22812 10312 -22716 10328
rect -22812 10248 -22796 10312
rect -22732 10248 -22716 10312
rect -22812 10232 -22716 10248
rect -22812 10168 -22796 10232
rect -22732 10168 -22716 10232
rect -22812 10152 -22716 10168
rect -22812 10088 -22796 10152
rect -22732 10088 -22716 10152
rect -22812 10072 -22716 10088
rect -22812 10008 -22796 10072
rect -22732 10008 -22716 10072
rect -22812 9992 -22716 10008
rect -22812 9928 -22796 9992
rect -22732 9928 -22716 9992
rect -22812 9912 -22716 9928
rect -22812 9848 -22796 9912
rect -22732 9848 -22716 9912
rect -22812 9832 -22716 9848
rect -22812 9768 -22796 9832
rect -22732 9768 -22716 9832
rect -22812 9752 -22716 9768
rect -22812 9688 -22796 9752
rect -22732 9688 -22716 9752
rect -22393 10432 -21671 10441
rect -22393 9728 -22384 10432
rect -21680 9728 -21671 10432
rect -22393 9719 -21671 9728
rect -21400 10408 -21384 10472
rect -21320 10408 -21304 10472
rect -19988 10472 -19892 10508
rect -21400 10392 -21304 10408
rect -21400 10328 -21384 10392
rect -21320 10328 -21304 10392
rect -21400 10312 -21304 10328
rect -21400 10248 -21384 10312
rect -21320 10248 -21304 10312
rect -21400 10232 -21304 10248
rect -21400 10168 -21384 10232
rect -21320 10168 -21304 10232
rect -21400 10152 -21304 10168
rect -21400 10088 -21384 10152
rect -21320 10088 -21304 10152
rect -21400 10072 -21304 10088
rect -21400 10008 -21384 10072
rect -21320 10008 -21304 10072
rect -21400 9992 -21304 10008
rect -21400 9928 -21384 9992
rect -21320 9928 -21304 9992
rect -21400 9912 -21304 9928
rect -21400 9848 -21384 9912
rect -21320 9848 -21304 9912
rect -21400 9832 -21304 9848
rect -21400 9768 -21384 9832
rect -21320 9768 -21304 9832
rect -21400 9752 -21304 9768
rect -22812 9652 -22716 9688
rect -21400 9688 -21384 9752
rect -21320 9688 -21304 9752
rect -20981 10432 -20259 10441
rect -20981 9728 -20972 10432
rect -20268 9728 -20259 10432
rect -20981 9719 -20259 9728
rect -19988 10408 -19972 10472
rect -19908 10408 -19892 10472
rect -18576 10472 -18480 10508
rect -19988 10392 -19892 10408
rect -19988 10328 -19972 10392
rect -19908 10328 -19892 10392
rect -19988 10312 -19892 10328
rect -19988 10248 -19972 10312
rect -19908 10248 -19892 10312
rect -19988 10232 -19892 10248
rect -19988 10168 -19972 10232
rect -19908 10168 -19892 10232
rect -19988 10152 -19892 10168
rect -19988 10088 -19972 10152
rect -19908 10088 -19892 10152
rect -19988 10072 -19892 10088
rect -19988 10008 -19972 10072
rect -19908 10008 -19892 10072
rect -19988 9992 -19892 10008
rect -19988 9928 -19972 9992
rect -19908 9928 -19892 9992
rect -19988 9912 -19892 9928
rect -19988 9848 -19972 9912
rect -19908 9848 -19892 9912
rect -19988 9832 -19892 9848
rect -19988 9768 -19972 9832
rect -19908 9768 -19892 9832
rect -19988 9752 -19892 9768
rect -21400 9652 -21304 9688
rect -19988 9688 -19972 9752
rect -19908 9688 -19892 9752
rect -19569 10432 -18847 10441
rect -19569 9728 -19560 10432
rect -18856 9728 -18847 10432
rect -19569 9719 -18847 9728
rect -18576 10408 -18560 10472
rect -18496 10408 -18480 10472
rect -17164 10472 -17068 10508
rect -18576 10392 -18480 10408
rect -18576 10328 -18560 10392
rect -18496 10328 -18480 10392
rect -18576 10312 -18480 10328
rect -18576 10248 -18560 10312
rect -18496 10248 -18480 10312
rect -18576 10232 -18480 10248
rect -18576 10168 -18560 10232
rect -18496 10168 -18480 10232
rect -18576 10152 -18480 10168
rect -18576 10088 -18560 10152
rect -18496 10088 -18480 10152
rect -18576 10072 -18480 10088
rect -18576 10008 -18560 10072
rect -18496 10008 -18480 10072
rect -18576 9992 -18480 10008
rect -18576 9928 -18560 9992
rect -18496 9928 -18480 9992
rect -18576 9912 -18480 9928
rect -18576 9848 -18560 9912
rect -18496 9848 -18480 9912
rect -18576 9832 -18480 9848
rect -18576 9768 -18560 9832
rect -18496 9768 -18480 9832
rect -18576 9752 -18480 9768
rect -19988 9652 -19892 9688
rect -18576 9688 -18560 9752
rect -18496 9688 -18480 9752
rect -18157 10432 -17435 10441
rect -18157 9728 -18148 10432
rect -17444 9728 -17435 10432
rect -18157 9719 -17435 9728
rect -17164 10408 -17148 10472
rect -17084 10408 -17068 10472
rect -15752 10472 -15656 10508
rect -17164 10392 -17068 10408
rect -17164 10328 -17148 10392
rect -17084 10328 -17068 10392
rect -17164 10312 -17068 10328
rect -17164 10248 -17148 10312
rect -17084 10248 -17068 10312
rect -17164 10232 -17068 10248
rect -17164 10168 -17148 10232
rect -17084 10168 -17068 10232
rect -17164 10152 -17068 10168
rect -17164 10088 -17148 10152
rect -17084 10088 -17068 10152
rect -17164 10072 -17068 10088
rect -17164 10008 -17148 10072
rect -17084 10008 -17068 10072
rect -17164 9992 -17068 10008
rect -17164 9928 -17148 9992
rect -17084 9928 -17068 9992
rect -17164 9912 -17068 9928
rect -17164 9848 -17148 9912
rect -17084 9848 -17068 9912
rect -17164 9832 -17068 9848
rect -17164 9768 -17148 9832
rect -17084 9768 -17068 9832
rect -17164 9752 -17068 9768
rect -18576 9652 -18480 9688
rect -17164 9688 -17148 9752
rect -17084 9688 -17068 9752
rect -16745 10432 -16023 10441
rect -16745 9728 -16736 10432
rect -16032 9728 -16023 10432
rect -16745 9719 -16023 9728
rect -15752 10408 -15736 10472
rect -15672 10408 -15656 10472
rect -14340 10472 -14244 10508
rect -15752 10392 -15656 10408
rect -15752 10328 -15736 10392
rect -15672 10328 -15656 10392
rect -15752 10312 -15656 10328
rect -15752 10248 -15736 10312
rect -15672 10248 -15656 10312
rect -15752 10232 -15656 10248
rect -15752 10168 -15736 10232
rect -15672 10168 -15656 10232
rect -15752 10152 -15656 10168
rect -15752 10088 -15736 10152
rect -15672 10088 -15656 10152
rect -15752 10072 -15656 10088
rect -15752 10008 -15736 10072
rect -15672 10008 -15656 10072
rect -15752 9992 -15656 10008
rect -15752 9928 -15736 9992
rect -15672 9928 -15656 9992
rect -15752 9912 -15656 9928
rect -15752 9848 -15736 9912
rect -15672 9848 -15656 9912
rect -15752 9832 -15656 9848
rect -15752 9768 -15736 9832
rect -15672 9768 -15656 9832
rect -15752 9752 -15656 9768
rect -17164 9652 -17068 9688
rect -15752 9688 -15736 9752
rect -15672 9688 -15656 9752
rect -15333 10432 -14611 10441
rect -15333 9728 -15324 10432
rect -14620 9728 -14611 10432
rect -15333 9719 -14611 9728
rect -14340 10408 -14324 10472
rect -14260 10408 -14244 10472
rect -12928 10472 -12832 10508
rect -14340 10392 -14244 10408
rect -14340 10328 -14324 10392
rect -14260 10328 -14244 10392
rect -14340 10312 -14244 10328
rect -14340 10248 -14324 10312
rect -14260 10248 -14244 10312
rect -14340 10232 -14244 10248
rect -14340 10168 -14324 10232
rect -14260 10168 -14244 10232
rect -14340 10152 -14244 10168
rect -14340 10088 -14324 10152
rect -14260 10088 -14244 10152
rect -14340 10072 -14244 10088
rect -14340 10008 -14324 10072
rect -14260 10008 -14244 10072
rect -14340 9992 -14244 10008
rect -14340 9928 -14324 9992
rect -14260 9928 -14244 9992
rect -14340 9912 -14244 9928
rect -14340 9848 -14324 9912
rect -14260 9848 -14244 9912
rect -14340 9832 -14244 9848
rect -14340 9768 -14324 9832
rect -14260 9768 -14244 9832
rect -14340 9752 -14244 9768
rect -15752 9652 -15656 9688
rect -14340 9688 -14324 9752
rect -14260 9688 -14244 9752
rect -13921 10432 -13199 10441
rect -13921 9728 -13912 10432
rect -13208 9728 -13199 10432
rect -13921 9719 -13199 9728
rect -12928 10408 -12912 10472
rect -12848 10408 -12832 10472
rect -11516 10472 -11420 10508
rect -12928 10392 -12832 10408
rect -12928 10328 -12912 10392
rect -12848 10328 -12832 10392
rect -12928 10312 -12832 10328
rect -12928 10248 -12912 10312
rect -12848 10248 -12832 10312
rect -12928 10232 -12832 10248
rect -12928 10168 -12912 10232
rect -12848 10168 -12832 10232
rect -12928 10152 -12832 10168
rect -12928 10088 -12912 10152
rect -12848 10088 -12832 10152
rect -12928 10072 -12832 10088
rect -12928 10008 -12912 10072
rect -12848 10008 -12832 10072
rect -12928 9992 -12832 10008
rect -12928 9928 -12912 9992
rect -12848 9928 -12832 9992
rect -12928 9912 -12832 9928
rect -12928 9848 -12912 9912
rect -12848 9848 -12832 9912
rect -12928 9832 -12832 9848
rect -12928 9768 -12912 9832
rect -12848 9768 -12832 9832
rect -12928 9752 -12832 9768
rect -14340 9652 -14244 9688
rect -12928 9688 -12912 9752
rect -12848 9688 -12832 9752
rect -12509 10432 -11787 10441
rect -12509 9728 -12500 10432
rect -11796 9728 -11787 10432
rect -12509 9719 -11787 9728
rect -11516 10408 -11500 10472
rect -11436 10408 -11420 10472
rect -10104 10472 -10008 10508
rect -11516 10392 -11420 10408
rect -11516 10328 -11500 10392
rect -11436 10328 -11420 10392
rect -11516 10312 -11420 10328
rect -11516 10248 -11500 10312
rect -11436 10248 -11420 10312
rect -11516 10232 -11420 10248
rect -11516 10168 -11500 10232
rect -11436 10168 -11420 10232
rect -11516 10152 -11420 10168
rect -11516 10088 -11500 10152
rect -11436 10088 -11420 10152
rect -11516 10072 -11420 10088
rect -11516 10008 -11500 10072
rect -11436 10008 -11420 10072
rect -11516 9992 -11420 10008
rect -11516 9928 -11500 9992
rect -11436 9928 -11420 9992
rect -11516 9912 -11420 9928
rect -11516 9848 -11500 9912
rect -11436 9848 -11420 9912
rect -11516 9832 -11420 9848
rect -11516 9768 -11500 9832
rect -11436 9768 -11420 9832
rect -11516 9752 -11420 9768
rect -12928 9652 -12832 9688
rect -11516 9688 -11500 9752
rect -11436 9688 -11420 9752
rect -11097 10432 -10375 10441
rect -11097 9728 -11088 10432
rect -10384 9728 -10375 10432
rect -11097 9719 -10375 9728
rect -10104 10408 -10088 10472
rect -10024 10408 -10008 10472
rect -8692 10472 -8596 10508
rect -10104 10392 -10008 10408
rect -10104 10328 -10088 10392
rect -10024 10328 -10008 10392
rect -10104 10312 -10008 10328
rect -10104 10248 -10088 10312
rect -10024 10248 -10008 10312
rect -10104 10232 -10008 10248
rect -10104 10168 -10088 10232
rect -10024 10168 -10008 10232
rect -10104 10152 -10008 10168
rect -10104 10088 -10088 10152
rect -10024 10088 -10008 10152
rect -10104 10072 -10008 10088
rect -10104 10008 -10088 10072
rect -10024 10008 -10008 10072
rect -10104 9992 -10008 10008
rect -10104 9928 -10088 9992
rect -10024 9928 -10008 9992
rect -10104 9912 -10008 9928
rect -10104 9848 -10088 9912
rect -10024 9848 -10008 9912
rect -10104 9832 -10008 9848
rect -10104 9768 -10088 9832
rect -10024 9768 -10008 9832
rect -10104 9752 -10008 9768
rect -11516 9652 -11420 9688
rect -10104 9688 -10088 9752
rect -10024 9688 -10008 9752
rect -9685 10432 -8963 10441
rect -9685 9728 -9676 10432
rect -8972 9728 -8963 10432
rect -9685 9719 -8963 9728
rect -8692 10408 -8676 10472
rect -8612 10408 -8596 10472
rect -7280 10472 -7184 10508
rect -8692 10392 -8596 10408
rect -8692 10328 -8676 10392
rect -8612 10328 -8596 10392
rect -8692 10312 -8596 10328
rect -8692 10248 -8676 10312
rect -8612 10248 -8596 10312
rect -8692 10232 -8596 10248
rect -8692 10168 -8676 10232
rect -8612 10168 -8596 10232
rect -8692 10152 -8596 10168
rect -8692 10088 -8676 10152
rect -8612 10088 -8596 10152
rect -8692 10072 -8596 10088
rect -8692 10008 -8676 10072
rect -8612 10008 -8596 10072
rect -8692 9992 -8596 10008
rect -8692 9928 -8676 9992
rect -8612 9928 -8596 9992
rect -8692 9912 -8596 9928
rect -8692 9848 -8676 9912
rect -8612 9848 -8596 9912
rect -8692 9832 -8596 9848
rect -8692 9768 -8676 9832
rect -8612 9768 -8596 9832
rect -8692 9752 -8596 9768
rect -10104 9652 -10008 9688
rect -8692 9688 -8676 9752
rect -8612 9688 -8596 9752
rect -8273 10432 -7551 10441
rect -8273 9728 -8264 10432
rect -7560 9728 -7551 10432
rect -8273 9719 -7551 9728
rect -7280 10408 -7264 10472
rect -7200 10408 -7184 10472
rect -5868 10472 -5772 10508
rect -7280 10392 -7184 10408
rect -7280 10328 -7264 10392
rect -7200 10328 -7184 10392
rect -7280 10312 -7184 10328
rect -7280 10248 -7264 10312
rect -7200 10248 -7184 10312
rect -7280 10232 -7184 10248
rect -7280 10168 -7264 10232
rect -7200 10168 -7184 10232
rect -7280 10152 -7184 10168
rect -7280 10088 -7264 10152
rect -7200 10088 -7184 10152
rect -7280 10072 -7184 10088
rect -7280 10008 -7264 10072
rect -7200 10008 -7184 10072
rect -7280 9992 -7184 10008
rect -7280 9928 -7264 9992
rect -7200 9928 -7184 9992
rect -7280 9912 -7184 9928
rect -7280 9848 -7264 9912
rect -7200 9848 -7184 9912
rect -7280 9832 -7184 9848
rect -7280 9768 -7264 9832
rect -7200 9768 -7184 9832
rect -7280 9752 -7184 9768
rect -8692 9652 -8596 9688
rect -7280 9688 -7264 9752
rect -7200 9688 -7184 9752
rect -6861 10432 -6139 10441
rect -6861 9728 -6852 10432
rect -6148 9728 -6139 10432
rect -6861 9719 -6139 9728
rect -5868 10408 -5852 10472
rect -5788 10408 -5772 10472
rect -4456 10472 -4360 10508
rect -5868 10392 -5772 10408
rect -5868 10328 -5852 10392
rect -5788 10328 -5772 10392
rect -5868 10312 -5772 10328
rect -5868 10248 -5852 10312
rect -5788 10248 -5772 10312
rect -5868 10232 -5772 10248
rect -5868 10168 -5852 10232
rect -5788 10168 -5772 10232
rect -5868 10152 -5772 10168
rect -5868 10088 -5852 10152
rect -5788 10088 -5772 10152
rect -5868 10072 -5772 10088
rect -5868 10008 -5852 10072
rect -5788 10008 -5772 10072
rect -5868 9992 -5772 10008
rect -5868 9928 -5852 9992
rect -5788 9928 -5772 9992
rect -5868 9912 -5772 9928
rect -5868 9848 -5852 9912
rect -5788 9848 -5772 9912
rect -5868 9832 -5772 9848
rect -5868 9768 -5852 9832
rect -5788 9768 -5772 9832
rect -5868 9752 -5772 9768
rect -7280 9652 -7184 9688
rect -5868 9688 -5852 9752
rect -5788 9688 -5772 9752
rect -5449 10432 -4727 10441
rect -5449 9728 -5440 10432
rect -4736 9728 -4727 10432
rect -5449 9719 -4727 9728
rect -4456 10408 -4440 10472
rect -4376 10408 -4360 10472
rect -3044 10472 -2948 10508
rect -4456 10392 -4360 10408
rect -4456 10328 -4440 10392
rect -4376 10328 -4360 10392
rect -4456 10312 -4360 10328
rect -4456 10248 -4440 10312
rect -4376 10248 -4360 10312
rect -4456 10232 -4360 10248
rect -4456 10168 -4440 10232
rect -4376 10168 -4360 10232
rect -4456 10152 -4360 10168
rect -4456 10088 -4440 10152
rect -4376 10088 -4360 10152
rect -4456 10072 -4360 10088
rect -4456 10008 -4440 10072
rect -4376 10008 -4360 10072
rect -4456 9992 -4360 10008
rect -4456 9928 -4440 9992
rect -4376 9928 -4360 9992
rect -4456 9912 -4360 9928
rect -4456 9848 -4440 9912
rect -4376 9848 -4360 9912
rect -4456 9832 -4360 9848
rect -4456 9768 -4440 9832
rect -4376 9768 -4360 9832
rect -4456 9752 -4360 9768
rect -5868 9652 -5772 9688
rect -4456 9688 -4440 9752
rect -4376 9688 -4360 9752
rect -4037 10432 -3315 10441
rect -4037 9728 -4028 10432
rect -3324 9728 -3315 10432
rect -4037 9719 -3315 9728
rect -3044 10408 -3028 10472
rect -2964 10408 -2948 10472
rect -1632 10472 -1536 10508
rect -3044 10392 -2948 10408
rect -3044 10328 -3028 10392
rect -2964 10328 -2948 10392
rect -3044 10312 -2948 10328
rect -3044 10248 -3028 10312
rect -2964 10248 -2948 10312
rect -3044 10232 -2948 10248
rect -3044 10168 -3028 10232
rect -2964 10168 -2948 10232
rect -3044 10152 -2948 10168
rect -3044 10088 -3028 10152
rect -2964 10088 -2948 10152
rect -3044 10072 -2948 10088
rect -3044 10008 -3028 10072
rect -2964 10008 -2948 10072
rect -3044 9992 -2948 10008
rect -3044 9928 -3028 9992
rect -2964 9928 -2948 9992
rect -3044 9912 -2948 9928
rect -3044 9848 -3028 9912
rect -2964 9848 -2948 9912
rect -3044 9832 -2948 9848
rect -3044 9768 -3028 9832
rect -2964 9768 -2948 9832
rect -3044 9752 -2948 9768
rect -4456 9652 -4360 9688
rect -3044 9688 -3028 9752
rect -2964 9688 -2948 9752
rect -2625 10432 -1903 10441
rect -2625 9728 -2616 10432
rect -1912 9728 -1903 10432
rect -2625 9719 -1903 9728
rect -1632 10408 -1616 10472
rect -1552 10408 -1536 10472
rect -220 10472 -124 10508
rect -1632 10392 -1536 10408
rect -1632 10328 -1616 10392
rect -1552 10328 -1536 10392
rect -1632 10312 -1536 10328
rect -1632 10248 -1616 10312
rect -1552 10248 -1536 10312
rect -1632 10232 -1536 10248
rect -1632 10168 -1616 10232
rect -1552 10168 -1536 10232
rect -1632 10152 -1536 10168
rect -1632 10088 -1616 10152
rect -1552 10088 -1536 10152
rect -1632 10072 -1536 10088
rect -1632 10008 -1616 10072
rect -1552 10008 -1536 10072
rect -1632 9992 -1536 10008
rect -1632 9928 -1616 9992
rect -1552 9928 -1536 9992
rect -1632 9912 -1536 9928
rect -1632 9848 -1616 9912
rect -1552 9848 -1536 9912
rect -1632 9832 -1536 9848
rect -1632 9768 -1616 9832
rect -1552 9768 -1536 9832
rect -1632 9752 -1536 9768
rect -3044 9652 -2948 9688
rect -1632 9688 -1616 9752
rect -1552 9688 -1536 9752
rect -1213 10432 -491 10441
rect -1213 9728 -1204 10432
rect -500 9728 -491 10432
rect -1213 9719 -491 9728
rect -220 10408 -204 10472
rect -140 10408 -124 10472
rect 1192 10472 1288 10508
rect -220 10392 -124 10408
rect -220 10328 -204 10392
rect -140 10328 -124 10392
rect -220 10312 -124 10328
rect -220 10248 -204 10312
rect -140 10248 -124 10312
rect -220 10232 -124 10248
rect -220 10168 -204 10232
rect -140 10168 -124 10232
rect -220 10152 -124 10168
rect -220 10088 -204 10152
rect -140 10088 -124 10152
rect -220 10072 -124 10088
rect -220 10008 -204 10072
rect -140 10008 -124 10072
rect -220 9992 -124 10008
rect -220 9928 -204 9992
rect -140 9928 -124 9992
rect -220 9912 -124 9928
rect -220 9848 -204 9912
rect -140 9848 -124 9912
rect -220 9832 -124 9848
rect -220 9768 -204 9832
rect -140 9768 -124 9832
rect -220 9752 -124 9768
rect -1632 9652 -1536 9688
rect -220 9688 -204 9752
rect -140 9688 -124 9752
rect 199 10432 921 10441
rect 199 9728 208 10432
rect 912 9728 921 10432
rect 199 9719 921 9728
rect 1192 10408 1208 10472
rect 1272 10408 1288 10472
rect 2604 10472 2700 10508
rect 1192 10392 1288 10408
rect 1192 10328 1208 10392
rect 1272 10328 1288 10392
rect 1192 10312 1288 10328
rect 1192 10248 1208 10312
rect 1272 10248 1288 10312
rect 1192 10232 1288 10248
rect 1192 10168 1208 10232
rect 1272 10168 1288 10232
rect 1192 10152 1288 10168
rect 1192 10088 1208 10152
rect 1272 10088 1288 10152
rect 1192 10072 1288 10088
rect 1192 10008 1208 10072
rect 1272 10008 1288 10072
rect 1192 9992 1288 10008
rect 1192 9928 1208 9992
rect 1272 9928 1288 9992
rect 1192 9912 1288 9928
rect 1192 9848 1208 9912
rect 1272 9848 1288 9912
rect 1192 9832 1288 9848
rect 1192 9768 1208 9832
rect 1272 9768 1288 9832
rect 1192 9752 1288 9768
rect -220 9652 -124 9688
rect 1192 9688 1208 9752
rect 1272 9688 1288 9752
rect 1611 10432 2333 10441
rect 1611 9728 1620 10432
rect 2324 9728 2333 10432
rect 1611 9719 2333 9728
rect 2604 10408 2620 10472
rect 2684 10408 2700 10472
rect 4016 10472 4112 10508
rect 2604 10392 2700 10408
rect 2604 10328 2620 10392
rect 2684 10328 2700 10392
rect 2604 10312 2700 10328
rect 2604 10248 2620 10312
rect 2684 10248 2700 10312
rect 2604 10232 2700 10248
rect 2604 10168 2620 10232
rect 2684 10168 2700 10232
rect 2604 10152 2700 10168
rect 2604 10088 2620 10152
rect 2684 10088 2700 10152
rect 2604 10072 2700 10088
rect 2604 10008 2620 10072
rect 2684 10008 2700 10072
rect 2604 9992 2700 10008
rect 2604 9928 2620 9992
rect 2684 9928 2700 9992
rect 2604 9912 2700 9928
rect 2604 9848 2620 9912
rect 2684 9848 2700 9912
rect 2604 9832 2700 9848
rect 2604 9768 2620 9832
rect 2684 9768 2700 9832
rect 2604 9752 2700 9768
rect 1192 9652 1288 9688
rect 2604 9688 2620 9752
rect 2684 9688 2700 9752
rect 3023 10432 3745 10441
rect 3023 9728 3032 10432
rect 3736 9728 3745 10432
rect 3023 9719 3745 9728
rect 4016 10408 4032 10472
rect 4096 10408 4112 10472
rect 5428 10472 5524 10508
rect 4016 10392 4112 10408
rect 4016 10328 4032 10392
rect 4096 10328 4112 10392
rect 4016 10312 4112 10328
rect 4016 10248 4032 10312
rect 4096 10248 4112 10312
rect 4016 10232 4112 10248
rect 4016 10168 4032 10232
rect 4096 10168 4112 10232
rect 4016 10152 4112 10168
rect 4016 10088 4032 10152
rect 4096 10088 4112 10152
rect 4016 10072 4112 10088
rect 4016 10008 4032 10072
rect 4096 10008 4112 10072
rect 4016 9992 4112 10008
rect 4016 9928 4032 9992
rect 4096 9928 4112 9992
rect 4016 9912 4112 9928
rect 4016 9848 4032 9912
rect 4096 9848 4112 9912
rect 4016 9832 4112 9848
rect 4016 9768 4032 9832
rect 4096 9768 4112 9832
rect 4016 9752 4112 9768
rect 2604 9652 2700 9688
rect 4016 9688 4032 9752
rect 4096 9688 4112 9752
rect 4435 10432 5157 10441
rect 4435 9728 4444 10432
rect 5148 9728 5157 10432
rect 4435 9719 5157 9728
rect 5428 10408 5444 10472
rect 5508 10408 5524 10472
rect 6840 10472 6936 10508
rect 5428 10392 5524 10408
rect 5428 10328 5444 10392
rect 5508 10328 5524 10392
rect 5428 10312 5524 10328
rect 5428 10248 5444 10312
rect 5508 10248 5524 10312
rect 5428 10232 5524 10248
rect 5428 10168 5444 10232
rect 5508 10168 5524 10232
rect 5428 10152 5524 10168
rect 5428 10088 5444 10152
rect 5508 10088 5524 10152
rect 5428 10072 5524 10088
rect 5428 10008 5444 10072
rect 5508 10008 5524 10072
rect 5428 9992 5524 10008
rect 5428 9928 5444 9992
rect 5508 9928 5524 9992
rect 5428 9912 5524 9928
rect 5428 9848 5444 9912
rect 5508 9848 5524 9912
rect 5428 9832 5524 9848
rect 5428 9768 5444 9832
rect 5508 9768 5524 9832
rect 5428 9752 5524 9768
rect 4016 9652 4112 9688
rect 5428 9688 5444 9752
rect 5508 9688 5524 9752
rect 5847 10432 6569 10441
rect 5847 9728 5856 10432
rect 6560 9728 6569 10432
rect 5847 9719 6569 9728
rect 6840 10408 6856 10472
rect 6920 10408 6936 10472
rect 8252 10472 8348 10508
rect 6840 10392 6936 10408
rect 6840 10328 6856 10392
rect 6920 10328 6936 10392
rect 6840 10312 6936 10328
rect 6840 10248 6856 10312
rect 6920 10248 6936 10312
rect 6840 10232 6936 10248
rect 6840 10168 6856 10232
rect 6920 10168 6936 10232
rect 6840 10152 6936 10168
rect 6840 10088 6856 10152
rect 6920 10088 6936 10152
rect 6840 10072 6936 10088
rect 6840 10008 6856 10072
rect 6920 10008 6936 10072
rect 6840 9992 6936 10008
rect 6840 9928 6856 9992
rect 6920 9928 6936 9992
rect 6840 9912 6936 9928
rect 6840 9848 6856 9912
rect 6920 9848 6936 9912
rect 6840 9832 6936 9848
rect 6840 9768 6856 9832
rect 6920 9768 6936 9832
rect 6840 9752 6936 9768
rect 5428 9652 5524 9688
rect 6840 9688 6856 9752
rect 6920 9688 6936 9752
rect 7259 10432 7981 10441
rect 7259 9728 7268 10432
rect 7972 9728 7981 10432
rect 7259 9719 7981 9728
rect 8252 10408 8268 10472
rect 8332 10408 8348 10472
rect 9664 10472 9760 10508
rect 8252 10392 8348 10408
rect 8252 10328 8268 10392
rect 8332 10328 8348 10392
rect 8252 10312 8348 10328
rect 8252 10248 8268 10312
rect 8332 10248 8348 10312
rect 8252 10232 8348 10248
rect 8252 10168 8268 10232
rect 8332 10168 8348 10232
rect 8252 10152 8348 10168
rect 8252 10088 8268 10152
rect 8332 10088 8348 10152
rect 8252 10072 8348 10088
rect 8252 10008 8268 10072
rect 8332 10008 8348 10072
rect 8252 9992 8348 10008
rect 8252 9928 8268 9992
rect 8332 9928 8348 9992
rect 8252 9912 8348 9928
rect 8252 9848 8268 9912
rect 8332 9848 8348 9912
rect 8252 9832 8348 9848
rect 8252 9768 8268 9832
rect 8332 9768 8348 9832
rect 8252 9752 8348 9768
rect 6840 9652 6936 9688
rect 8252 9688 8268 9752
rect 8332 9688 8348 9752
rect 8671 10432 9393 10441
rect 8671 9728 8680 10432
rect 9384 9728 9393 10432
rect 8671 9719 9393 9728
rect 9664 10408 9680 10472
rect 9744 10408 9760 10472
rect 11076 10472 11172 10508
rect 9664 10392 9760 10408
rect 9664 10328 9680 10392
rect 9744 10328 9760 10392
rect 9664 10312 9760 10328
rect 9664 10248 9680 10312
rect 9744 10248 9760 10312
rect 9664 10232 9760 10248
rect 9664 10168 9680 10232
rect 9744 10168 9760 10232
rect 9664 10152 9760 10168
rect 9664 10088 9680 10152
rect 9744 10088 9760 10152
rect 9664 10072 9760 10088
rect 9664 10008 9680 10072
rect 9744 10008 9760 10072
rect 9664 9992 9760 10008
rect 9664 9928 9680 9992
rect 9744 9928 9760 9992
rect 9664 9912 9760 9928
rect 9664 9848 9680 9912
rect 9744 9848 9760 9912
rect 9664 9832 9760 9848
rect 9664 9768 9680 9832
rect 9744 9768 9760 9832
rect 9664 9752 9760 9768
rect 8252 9652 8348 9688
rect 9664 9688 9680 9752
rect 9744 9688 9760 9752
rect 10083 10432 10805 10441
rect 10083 9728 10092 10432
rect 10796 9728 10805 10432
rect 10083 9719 10805 9728
rect 11076 10408 11092 10472
rect 11156 10408 11172 10472
rect 12488 10472 12584 10508
rect 11076 10392 11172 10408
rect 11076 10328 11092 10392
rect 11156 10328 11172 10392
rect 11076 10312 11172 10328
rect 11076 10248 11092 10312
rect 11156 10248 11172 10312
rect 11076 10232 11172 10248
rect 11076 10168 11092 10232
rect 11156 10168 11172 10232
rect 11076 10152 11172 10168
rect 11076 10088 11092 10152
rect 11156 10088 11172 10152
rect 11076 10072 11172 10088
rect 11076 10008 11092 10072
rect 11156 10008 11172 10072
rect 11076 9992 11172 10008
rect 11076 9928 11092 9992
rect 11156 9928 11172 9992
rect 11076 9912 11172 9928
rect 11076 9848 11092 9912
rect 11156 9848 11172 9912
rect 11076 9832 11172 9848
rect 11076 9768 11092 9832
rect 11156 9768 11172 9832
rect 11076 9752 11172 9768
rect 9664 9652 9760 9688
rect 11076 9688 11092 9752
rect 11156 9688 11172 9752
rect 11495 10432 12217 10441
rect 11495 9728 11504 10432
rect 12208 9728 12217 10432
rect 11495 9719 12217 9728
rect 12488 10408 12504 10472
rect 12568 10408 12584 10472
rect 13900 10472 13996 10508
rect 12488 10392 12584 10408
rect 12488 10328 12504 10392
rect 12568 10328 12584 10392
rect 12488 10312 12584 10328
rect 12488 10248 12504 10312
rect 12568 10248 12584 10312
rect 12488 10232 12584 10248
rect 12488 10168 12504 10232
rect 12568 10168 12584 10232
rect 12488 10152 12584 10168
rect 12488 10088 12504 10152
rect 12568 10088 12584 10152
rect 12488 10072 12584 10088
rect 12488 10008 12504 10072
rect 12568 10008 12584 10072
rect 12488 9992 12584 10008
rect 12488 9928 12504 9992
rect 12568 9928 12584 9992
rect 12488 9912 12584 9928
rect 12488 9848 12504 9912
rect 12568 9848 12584 9912
rect 12488 9832 12584 9848
rect 12488 9768 12504 9832
rect 12568 9768 12584 9832
rect 12488 9752 12584 9768
rect 11076 9652 11172 9688
rect 12488 9688 12504 9752
rect 12568 9688 12584 9752
rect 12907 10432 13629 10441
rect 12907 9728 12916 10432
rect 13620 9728 13629 10432
rect 12907 9719 13629 9728
rect 13900 10408 13916 10472
rect 13980 10408 13996 10472
rect 15312 10472 15408 10508
rect 13900 10392 13996 10408
rect 13900 10328 13916 10392
rect 13980 10328 13996 10392
rect 13900 10312 13996 10328
rect 13900 10248 13916 10312
rect 13980 10248 13996 10312
rect 13900 10232 13996 10248
rect 13900 10168 13916 10232
rect 13980 10168 13996 10232
rect 13900 10152 13996 10168
rect 13900 10088 13916 10152
rect 13980 10088 13996 10152
rect 13900 10072 13996 10088
rect 13900 10008 13916 10072
rect 13980 10008 13996 10072
rect 13900 9992 13996 10008
rect 13900 9928 13916 9992
rect 13980 9928 13996 9992
rect 13900 9912 13996 9928
rect 13900 9848 13916 9912
rect 13980 9848 13996 9912
rect 13900 9832 13996 9848
rect 13900 9768 13916 9832
rect 13980 9768 13996 9832
rect 13900 9752 13996 9768
rect 12488 9652 12584 9688
rect 13900 9688 13916 9752
rect 13980 9688 13996 9752
rect 14319 10432 15041 10441
rect 14319 9728 14328 10432
rect 15032 9728 15041 10432
rect 14319 9719 15041 9728
rect 15312 10408 15328 10472
rect 15392 10408 15408 10472
rect 16724 10472 16820 10508
rect 15312 10392 15408 10408
rect 15312 10328 15328 10392
rect 15392 10328 15408 10392
rect 15312 10312 15408 10328
rect 15312 10248 15328 10312
rect 15392 10248 15408 10312
rect 15312 10232 15408 10248
rect 15312 10168 15328 10232
rect 15392 10168 15408 10232
rect 15312 10152 15408 10168
rect 15312 10088 15328 10152
rect 15392 10088 15408 10152
rect 15312 10072 15408 10088
rect 15312 10008 15328 10072
rect 15392 10008 15408 10072
rect 15312 9992 15408 10008
rect 15312 9928 15328 9992
rect 15392 9928 15408 9992
rect 15312 9912 15408 9928
rect 15312 9848 15328 9912
rect 15392 9848 15408 9912
rect 15312 9832 15408 9848
rect 15312 9768 15328 9832
rect 15392 9768 15408 9832
rect 15312 9752 15408 9768
rect 13900 9652 13996 9688
rect 15312 9688 15328 9752
rect 15392 9688 15408 9752
rect 15731 10432 16453 10441
rect 15731 9728 15740 10432
rect 16444 9728 16453 10432
rect 15731 9719 16453 9728
rect 16724 10408 16740 10472
rect 16804 10408 16820 10472
rect 18136 10472 18232 10508
rect 16724 10392 16820 10408
rect 16724 10328 16740 10392
rect 16804 10328 16820 10392
rect 16724 10312 16820 10328
rect 16724 10248 16740 10312
rect 16804 10248 16820 10312
rect 16724 10232 16820 10248
rect 16724 10168 16740 10232
rect 16804 10168 16820 10232
rect 16724 10152 16820 10168
rect 16724 10088 16740 10152
rect 16804 10088 16820 10152
rect 16724 10072 16820 10088
rect 16724 10008 16740 10072
rect 16804 10008 16820 10072
rect 16724 9992 16820 10008
rect 16724 9928 16740 9992
rect 16804 9928 16820 9992
rect 16724 9912 16820 9928
rect 16724 9848 16740 9912
rect 16804 9848 16820 9912
rect 16724 9832 16820 9848
rect 16724 9768 16740 9832
rect 16804 9768 16820 9832
rect 16724 9752 16820 9768
rect 15312 9652 15408 9688
rect 16724 9688 16740 9752
rect 16804 9688 16820 9752
rect 17143 10432 17865 10441
rect 17143 9728 17152 10432
rect 17856 9728 17865 10432
rect 17143 9719 17865 9728
rect 18136 10408 18152 10472
rect 18216 10408 18232 10472
rect 19548 10472 19644 10508
rect 18136 10392 18232 10408
rect 18136 10328 18152 10392
rect 18216 10328 18232 10392
rect 18136 10312 18232 10328
rect 18136 10248 18152 10312
rect 18216 10248 18232 10312
rect 18136 10232 18232 10248
rect 18136 10168 18152 10232
rect 18216 10168 18232 10232
rect 18136 10152 18232 10168
rect 18136 10088 18152 10152
rect 18216 10088 18232 10152
rect 18136 10072 18232 10088
rect 18136 10008 18152 10072
rect 18216 10008 18232 10072
rect 18136 9992 18232 10008
rect 18136 9928 18152 9992
rect 18216 9928 18232 9992
rect 18136 9912 18232 9928
rect 18136 9848 18152 9912
rect 18216 9848 18232 9912
rect 18136 9832 18232 9848
rect 18136 9768 18152 9832
rect 18216 9768 18232 9832
rect 18136 9752 18232 9768
rect 16724 9652 16820 9688
rect 18136 9688 18152 9752
rect 18216 9688 18232 9752
rect 18555 10432 19277 10441
rect 18555 9728 18564 10432
rect 19268 9728 19277 10432
rect 18555 9719 19277 9728
rect 19548 10408 19564 10472
rect 19628 10408 19644 10472
rect 20960 10472 21056 10508
rect 19548 10392 19644 10408
rect 19548 10328 19564 10392
rect 19628 10328 19644 10392
rect 19548 10312 19644 10328
rect 19548 10248 19564 10312
rect 19628 10248 19644 10312
rect 19548 10232 19644 10248
rect 19548 10168 19564 10232
rect 19628 10168 19644 10232
rect 19548 10152 19644 10168
rect 19548 10088 19564 10152
rect 19628 10088 19644 10152
rect 19548 10072 19644 10088
rect 19548 10008 19564 10072
rect 19628 10008 19644 10072
rect 19548 9992 19644 10008
rect 19548 9928 19564 9992
rect 19628 9928 19644 9992
rect 19548 9912 19644 9928
rect 19548 9848 19564 9912
rect 19628 9848 19644 9912
rect 19548 9832 19644 9848
rect 19548 9768 19564 9832
rect 19628 9768 19644 9832
rect 19548 9752 19644 9768
rect 18136 9652 18232 9688
rect 19548 9688 19564 9752
rect 19628 9688 19644 9752
rect 19967 10432 20689 10441
rect 19967 9728 19976 10432
rect 20680 9728 20689 10432
rect 19967 9719 20689 9728
rect 20960 10408 20976 10472
rect 21040 10408 21056 10472
rect 22372 10472 22468 10508
rect 20960 10392 21056 10408
rect 20960 10328 20976 10392
rect 21040 10328 21056 10392
rect 20960 10312 21056 10328
rect 20960 10248 20976 10312
rect 21040 10248 21056 10312
rect 20960 10232 21056 10248
rect 20960 10168 20976 10232
rect 21040 10168 21056 10232
rect 20960 10152 21056 10168
rect 20960 10088 20976 10152
rect 21040 10088 21056 10152
rect 20960 10072 21056 10088
rect 20960 10008 20976 10072
rect 21040 10008 21056 10072
rect 20960 9992 21056 10008
rect 20960 9928 20976 9992
rect 21040 9928 21056 9992
rect 20960 9912 21056 9928
rect 20960 9848 20976 9912
rect 21040 9848 21056 9912
rect 20960 9832 21056 9848
rect 20960 9768 20976 9832
rect 21040 9768 21056 9832
rect 20960 9752 21056 9768
rect 19548 9652 19644 9688
rect 20960 9688 20976 9752
rect 21040 9688 21056 9752
rect 21379 10432 22101 10441
rect 21379 9728 21388 10432
rect 22092 9728 22101 10432
rect 21379 9719 22101 9728
rect 22372 10408 22388 10472
rect 22452 10408 22468 10472
rect 23784 10472 23880 10508
rect 22372 10392 22468 10408
rect 22372 10328 22388 10392
rect 22452 10328 22468 10392
rect 22372 10312 22468 10328
rect 22372 10248 22388 10312
rect 22452 10248 22468 10312
rect 22372 10232 22468 10248
rect 22372 10168 22388 10232
rect 22452 10168 22468 10232
rect 22372 10152 22468 10168
rect 22372 10088 22388 10152
rect 22452 10088 22468 10152
rect 22372 10072 22468 10088
rect 22372 10008 22388 10072
rect 22452 10008 22468 10072
rect 22372 9992 22468 10008
rect 22372 9928 22388 9992
rect 22452 9928 22468 9992
rect 22372 9912 22468 9928
rect 22372 9848 22388 9912
rect 22452 9848 22468 9912
rect 22372 9832 22468 9848
rect 22372 9768 22388 9832
rect 22452 9768 22468 9832
rect 22372 9752 22468 9768
rect 20960 9652 21056 9688
rect 22372 9688 22388 9752
rect 22452 9688 22468 9752
rect 22791 10432 23513 10441
rect 22791 9728 22800 10432
rect 23504 9728 23513 10432
rect 22791 9719 23513 9728
rect 23784 10408 23800 10472
rect 23864 10408 23880 10472
rect 23784 10392 23880 10408
rect 23784 10328 23800 10392
rect 23864 10328 23880 10392
rect 23784 10312 23880 10328
rect 23784 10248 23800 10312
rect 23864 10248 23880 10312
rect 23784 10232 23880 10248
rect 23784 10168 23800 10232
rect 23864 10168 23880 10232
rect 23784 10152 23880 10168
rect 23784 10088 23800 10152
rect 23864 10088 23880 10152
rect 23784 10072 23880 10088
rect 23784 10008 23800 10072
rect 23864 10008 23880 10072
rect 23784 9992 23880 10008
rect 23784 9928 23800 9992
rect 23864 9928 23880 9992
rect 23784 9912 23880 9928
rect 23784 9848 23800 9912
rect 23864 9848 23880 9912
rect 23784 9832 23880 9848
rect 23784 9768 23800 9832
rect 23864 9768 23880 9832
rect 23784 9752 23880 9768
rect 22372 9652 22468 9688
rect 23784 9688 23800 9752
rect 23864 9688 23880 9752
rect 23784 9652 23880 9688
rect -22812 9352 -22716 9388
rect -23805 9312 -23083 9321
rect -23805 8608 -23796 9312
rect -23092 8608 -23083 9312
rect -23805 8599 -23083 8608
rect -22812 9288 -22796 9352
rect -22732 9288 -22716 9352
rect -21400 9352 -21304 9388
rect -22812 9272 -22716 9288
rect -22812 9208 -22796 9272
rect -22732 9208 -22716 9272
rect -22812 9192 -22716 9208
rect -22812 9128 -22796 9192
rect -22732 9128 -22716 9192
rect -22812 9112 -22716 9128
rect -22812 9048 -22796 9112
rect -22732 9048 -22716 9112
rect -22812 9032 -22716 9048
rect -22812 8968 -22796 9032
rect -22732 8968 -22716 9032
rect -22812 8952 -22716 8968
rect -22812 8888 -22796 8952
rect -22732 8888 -22716 8952
rect -22812 8872 -22716 8888
rect -22812 8808 -22796 8872
rect -22732 8808 -22716 8872
rect -22812 8792 -22716 8808
rect -22812 8728 -22796 8792
rect -22732 8728 -22716 8792
rect -22812 8712 -22716 8728
rect -22812 8648 -22796 8712
rect -22732 8648 -22716 8712
rect -22812 8632 -22716 8648
rect -22812 8568 -22796 8632
rect -22732 8568 -22716 8632
rect -22393 9312 -21671 9321
rect -22393 8608 -22384 9312
rect -21680 8608 -21671 9312
rect -22393 8599 -21671 8608
rect -21400 9288 -21384 9352
rect -21320 9288 -21304 9352
rect -19988 9352 -19892 9388
rect -21400 9272 -21304 9288
rect -21400 9208 -21384 9272
rect -21320 9208 -21304 9272
rect -21400 9192 -21304 9208
rect -21400 9128 -21384 9192
rect -21320 9128 -21304 9192
rect -21400 9112 -21304 9128
rect -21400 9048 -21384 9112
rect -21320 9048 -21304 9112
rect -21400 9032 -21304 9048
rect -21400 8968 -21384 9032
rect -21320 8968 -21304 9032
rect -21400 8952 -21304 8968
rect -21400 8888 -21384 8952
rect -21320 8888 -21304 8952
rect -21400 8872 -21304 8888
rect -21400 8808 -21384 8872
rect -21320 8808 -21304 8872
rect -21400 8792 -21304 8808
rect -21400 8728 -21384 8792
rect -21320 8728 -21304 8792
rect -21400 8712 -21304 8728
rect -21400 8648 -21384 8712
rect -21320 8648 -21304 8712
rect -21400 8632 -21304 8648
rect -22812 8532 -22716 8568
rect -21400 8568 -21384 8632
rect -21320 8568 -21304 8632
rect -20981 9312 -20259 9321
rect -20981 8608 -20972 9312
rect -20268 8608 -20259 9312
rect -20981 8599 -20259 8608
rect -19988 9288 -19972 9352
rect -19908 9288 -19892 9352
rect -18576 9352 -18480 9388
rect -19988 9272 -19892 9288
rect -19988 9208 -19972 9272
rect -19908 9208 -19892 9272
rect -19988 9192 -19892 9208
rect -19988 9128 -19972 9192
rect -19908 9128 -19892 9192
rect -19988 9112 -19892 9128
rect -19988 9048 -19972 9112
rect -19908 9048 -19892 9112
rect -19988 9032 -19892 9048
rect -19988 8968 -19972 9032
rect -19908 8968 -19892 9032
rect -19988 8952 -19892 8968
rect -19988 8888 -19972 8952
rect -19908 8888 -19892 8952
rect -19988 8872 -19892 8888
rect -19988 8808 -19972 8872
rect -19908 8808 -19892 8872
rect -19988 8792 -19892 8808
rect -19988 8728 -19972 8792
rect -19908 8728 -19892 8792
rect -19988 8712 -19892 8728
rect -19988 8648 -19972 8712
rect -19908 8648 -19892 8712
rect -19988 8632 -19892 8648
rect -21400 8532 -21304 8568
rect -19988 8568 -19972 8632
rect -19908 8568 -19892 8632
rect -19569 9312 -18847 9321
rect -19569 8608 -19560 9312
rect -18856 8608 -18847 9312
rect -19569 8599 -18847 8608
rect -18576 9288 -18560 9352
rect -18496 9288 -18480 9352
rect -17164 9352 -17068 9388
rect -18576 9272 -18480 9288
rect -18576 9208 -18560 9272
rect -18496 9208 -18480 9272
rect -18576 9192 -18480 9208
rect -18576 9128 -18560 9192
rect -18496 9128 -18480 9192
rect -18576 9112 -18480 9128
rect -18576 9048 -18560 9112
rect -18496 9048 -18480 9112
rect -18576 9032 -18480 9048
rect -18576 8968 -18560 9032
rect -18496 8968 -18480 9032
rect -18576 8952 -18480 8968
rect -18576 8888 -18560 8952
rect -18496 8888 -18480 8952
rect -18576 8872 -18480 8888
rect -18576 8808 -18560 8872
rect -18496 8808 -18480 8872
rect -18576 8792 -18480 8808
rect -18576 8728 -18560 8792
rect -18496 8728 -18480 8792
rect -18576 8712 -18480 8728
rect -18576 8648 -18560 8712
rect -18496 8648 -18480 8712
rect -18576 8632 -18480 8648
rect -19988 8532 -19892 8568
rect -18576 8568 -18560 8632
rect -18496 8568 -18480 8632
rect -18157 9312 -17435 9321
rect -18157 8608 -18148 9312
rect -17444 8608 -17435 9312
rect -18157 8599 -17435 8608
rect -17164 9288 -17148 9352
rect -17084 9288 -17068 9352
rect -15752 9352 -15656 9388
rect -17164 9272 -17068 9288
rect -17164 9208 -17148 9272
rect -17084 9208 -17068 9272
rect -17164 9192 -17068 9208
rect -17164 9128 -17148 9192
rect -17084 9128 -17068 9192
rect -17164 9112 -17068 9128
rect -17164 9048 -17148 9112
rect -17084 9048 -17068 9112
rect -17164 9032 -17068 9048
rect -17164 8968 -17148 9032
rect -17084 8968 -17068 9032
rect -17164 8952 -17068 8968
rect -17164 8888 -17148 8952
rect -17084 8888 -17068 8952
rect -17164 8872 -17068 8888
rect -17164 8808 -17148 8872
rect -17084 8808 -17068 8872
rect -17164 8792 -17068 8808
rect -17164 8728 -17148 8792
rect -17084 8728 -17068 8792
rect -17164 8712 -17068 8728
rect -17164 8648 -17148 8712
rect -17084 8648 -17068 8712
rect -17164 8632 -17068 8648
rect -18576 8532 -18480 8568
rect -17164 8568 -17148 8632
rect -17084 8568 -17068 8632
rect -16745 9312 -16023 9321
rect -16745 8608 -16736 9312
rect -16032 8608 -16023 9312
rect -16745 8599 -16023 8608
rect -15752 9288 -15736 9352
rect -15672 9288 -15656 9352
rect -14340 9352 -14244 9388
rect -15752 9272 -15656 9288
rect -15752 9208 -15736 9272
rect -15672 9208 -15656 9272
rect -15752 9192 -15656 9208
rect -15752 9128 -15736 9192
rect -15672 9128 -15656 9192
rect -15752 9112 -15656 9128
rect -15752 9048 -15736 9112
rect -15672 9048 -15656 9112
rect -15752 9032 -15656 9048
rect -15752 8968 -15736 9032
rect -15672 8968 -15656 9032
rect -15752 8952 -15656 8968
rect -15752 8888 -15736 8952
rect -15672 8888 -15656 8952
rect -15752 8872 -15656 8888
rect -15752 8808 -15736 8872
rect -15672 8808 -15656 8872
rect -15752 8792 -15656 8808
rect -15752 8728 -15736 8792
rect -15672 8728 -15656 8792
rect -15752 8712 -15656 8728
rect -15752 8648 -15736 8712
rect -15672 8648 -15656 8712
rect -15752 8632 -15656 8648
rect -17164 8532 -17068 8568
rect -15752 8568 -15736 8632
rect -15672 8568 -15656 8632
rect -15333 9312 -14611 9321
rect -15333 8608 -15324 9312
rect -14620 8608 -14611 9312
rect -15333 8599 -14611 8608
rect -14340 9288 -14324 9352
rect -14260 9288 -14244 9352
rect -12928 9352 -12832 9388
rect -14340 9272 -14244 9288
rect -14340 9208 -14324 9272
rect -14260 9208 -14244 9272
rect -14340 9192 -14244 9208
rect -14340 9128 -14324 9192
rect -14260 9128 -14244 9192
rect -14340 9112 -14244 9128
rect -14340 9048 -14324 9112
rect -14260 9048 -14244 9112
rect -14340 9032 -14244 9048
rect -14340 8968 -14324 9032
rect -14260 8968 -14244 9032
rect -14340 8952 -14244 8968
rect -14340 8888 -14324 8952
rect -14260 8888 -14244 8952
rect -14340 8872 -14244 8888
rect -14340 8808 -14324 8872
rect -14260 8808 -14244 8872
rect -14340 8792 -14244 8808
rect -14340 8728 -14324 8792
rect -14260 8728 -14244 8792
rect -14340 8712 -14244 8728
rect -14340 8648 -14324 8712
rect -14260 8648 -14244 8712
rect -14340 8632 -14244 8648
rect -15752 8532 -15656 8568
rect -14340 8568 -14324 8632
rect -14260 8568 -14244 8632
rect -13921 9312 -13199 9321
rect -13921 8608 -13912 9312
rect -13208 8608 -13199 9312
rect -13921 8599 -13199 8608
rect -12928 9288 -12912 9352
rect -12848 9288 -12832 9352
rect -11516 9352 -11420 9388
rect -12928 9272 -12832 9288
rect -12928 9208 -12912 9272
rect -12848 9208 -12832 9272
rect -12928 9192 -12832 9208
rect -12928 9128 -12912 9192
rect -12848 9128 -12832 9192
rect -12928 9112 -12832 9128
rect -12928 9048 -12912 9112
rect -12848 9048 -12832 9112
rect -12928 9032 -12832 9048
rect -12928 8968 -12912 9032
rect -12848 8968 -12832 9032
rect -12928 8952 -12832 8968
rect -12928 8888 -12912 8952
rect -12848 8888 -12832 8952
rect -12928 8872 -12832 8888
rect -12928 8808 -12912 8872
rect -12848 8808 -12832 8872
rect -12928 8792 -12832 8808
rect -12928 8728 -12912 8792
rect -12848 8728 -12832 8792
rect -12928 8712 -12832 8728
rect -12928 8648 -12912 8712
rect -12848 8648 -12832 8712
rect -12928 8632 -12832 8648
rect -14340 8532 -14244 8568
rect -12928 8568 -12912 8632
rect -12848 8568 -12832 8632
rect -12509 9312 -11787 9321
rect -12509 8608 -12500 9312
rect -11796 8608 -11787 9312
rect -12509 8599 -11787 8608
rect -11516 9288 -11500 9352
rect -11436 9288 -11420 9352
rect -10104 9352 -10008 9388
rect -11516 9272 -11420 9288
rect -11516 9208 -11500 9272
rect -11436 9208 -11420 9272
rect -11516 9192 -11420 9208
rect -11516 9128 -11500 9192
rect -11436 9128 -11420 9192
rect -11516 9112 -11420 9128
rect -11516 9048 -11500 9112
rect -11436 9048 -11420 9112
rect -11516 9032 -11420 9048
rect -11516 8968 -11500 9032
rect -11436 8968 -11420 9032
rect -11516 8952 -11420 8968
rect -11516 8888 -11500 8952
rect -11436 8888 -11420 8952
rect -11516 8872 -11420 8888
rect -11516 8808 -11500 8872
rect -11436 8808 -11420 8872
rect -11516 8792 -11420 8808
rect -11516 8728 -11500 8792
rect -11436 8728 -11420 8792
rect -11516 8712 -11420 8728
rect -11516 8648 -11500 8712
rect -11436 8648 -11420 8712
rect -11516 8632 -11420 8648
rect -12928 8532 -12832 8568
rect -11516 8568 -11500 8632
rect -11436 8568 -11420 8632
rect -11097 9312 -10375 9321
rect -11097 8608 -11088 9312
rect -10384 8608 -10375 9312
rect -11097 8599 -10375 8608
rect -10104 9288 -10088 9352
rect -10024 9288 -10008 9352
rect -8692 9352 -8596 9388
rect -10104 9272 -10008 9288
rect -10104 9208 -10088 9272
rect -10024 9208 -10008 9272
rect -10104 9192 -10008 9208
rect -10104 9128 -10088 9192
rect -10024 9128 -10008 9192
rect -10104 9112 -10008 9128
rect -10104 9048 -10088 9112
rect -10024 9048 -10008 9112
rect -10104 9032 -10008 9048
rect -10104 8968 -10088 9032
rect -10024 8968 -10008 9032
rect -10104 8952 -10008 8968
rect -10104 8888 -10088 8952
rect -10024 8888 -10008 8952
rect -10104 8872 -10008 8888
rect -10104 8808 -10088 8872
rect -10024 8808 -10008 8872
rect -10104 8792 -10008 8808
rect -10104 8728 -10088 8792
rect -10024 8728 -10008 8792
rect -10104 8712 -10008 8728
rect -10104 8648 -10088 8712
rect -10024 8648 -10008 8712
rect -10104 8632 -10008 8648
rect -11516 8532 -11420 8568
rect -10104 8568 -10088 8632
rect -10024 8568 -10008 8632
rect -9685 9312 -8963 9321
rect -9685 8608 -9676 9312
rect -8972 8608 -8963 9312
rect -9685 8599 -8963 8608
rect -8692 9288 -8676 9352
rect -8612 9288 -8596 9352
rect -7280 9352 -7184 9388
rect -8692 9272 -8596 9288
rect -8692 9208 -8676 9272
rect -8612 9208 -8596 9272
rect -8692 9192 -8596 9208
rect -8692 9128 -8676 9192
rect -8612 9128 -8596 9192
rect -8692 9112 -8596 9128
rect -8692 9048 -8676 9112
rect -8612 9048 -8596 9112
rect -8692 9032 -8596 9048
rect -8692 8968 -8676 9032
rect -8612 8968 -8596 9032
rect -8692 8952 -8596 8968
rect -8692 8888 -8676 8952
rect -8612 8888 -8596 8952
rect -8692 8872 -8596 8888
rect -8692 8808 -8676 8872
rect -8612 8808 -8596 8872
rect -8692 8792 -8596 8808
rect -8692 8728 -8676 8792
rect -8612 8728 -8596 8792
rect -8692 8712 -8596 8728
rect -8692 8648 -8676 8712
rect -8612 8648 -8596 8712
rect -8692 8632 -8596 8648
rect -10104 8532 -10008 8568
rect -8692 8568 -8676 8632
rect -8612 8568 -8596 8632
rect -8273 9312 -7551 9321
rect -8273 8608 -8264 9312
rect -7560 8608 -7551 9312
rect -8273 8599 -7551 8608
rect -7280 9288 -7264 9352
rect -7200 9288 -7184 9352
rect -5868 9352 -5772 9388
rect -7280 9272 -7184 9288
rect -7280 9208 -7264 9272
rect -7200 9208 -7184 9272
rect -7280 9192 -7184 9208
rect -7280 9128 -7264 9192
rect -7200 9128 -7184 9192
rect -7280 9112 -7184 9128
rect -7280 9048 -7264 9112
rect -7200 9048 -7184 9112
rect -7280 9032 -7184 9048
rect -7280 8968 -7264 9032
rect -7200 8968 -7184 9032
rect -7280 8952 -7184 8968
rect -7280 8888 -7264 8952
rect -7200 8888 -7184 8952
rect -7280 8872 -7184 8888
rect -7280 8808 -7264 8872
rect -7200 8808 -7184 8872
rect -7280 8792 -7184 8808
rect -7280 8728 -7264 8792
rect -7200 8728 -7184 8792
rect -7280 8712 -7184 8728
rect -7280 8648 -7264 8712
rect -7200 8648 -7184 8712
rect -7280 8632 -7184 8648
rect -8692 8532 -8596 8568
rect -7280 8568 -7264 8632
rect -7200 8568 -7184 8632
rect -6861 9312 -6139 9321
rect -6861 8608 -6852 9312
rect -6148 8608 -6139 9312
rect -6861 8599 -6139 8608
rect -5868 9288 -5852 9352
rect -5788 9288 -5772 9352
rect -4456 9352 -4360 9388
rect -5868 9272 -5772 9288
rect -5868 9208 -5852 9272
rect -5788 9208 -5772 9272
rect -5868 9192 -5772 9208
rect -5868 9128 -5852 9192
rect -5788 9128 -5772 9192
rect -5868 9112 -5772 9128
rect -5868 9048 -5852 9112
rect -5788 9048 -5772 9112
rect -5868 9032 -5772 9048
rect -5868 8968 -5852 9032
rect -5788 8968 -5772 9032
rect -5868 8952 -5772 8968
rect -5868 8888 -5852 8952
rect -5788 8888 -5772 8952
rect -5868 8872 -5772 8888
rect -5868 8808 -5852 8872
rect -5788 8808 -5772 8872
rect -5868 8792 -5772 8808
rect -5868 8728 -5852 8792
rect -5788 8728 -5772 8792
rect -5868 8712 -5772 8728
rect -5868 8648 -5852 8712
rect -5788 8648 -5772 8712
rect -5868 8632 -5772 8648
rect -7280 8532 -7184 8568
rect -5868 8568 -5852 8632
rect -5788 8568 -5772 8632
rect -5449 9312 -4727 9321
rect -5449 8608 -5440 9312
rect -4736 8608 -4727 9312
rect -5449 8599 -4727 8608
rect -4456 9288 -4440 9352
rect -4376 9288 -4360 9352
rect -3044 9352 -2948 9388
rect -4456 9272 -4360 9288
rect -4456 9208 -4440 9272
rect -4376 9208 -4360 9272
rect -4456 9192 -4360 9208
rect -4456 9128 -4440 9192
rect -4376 9128 -4360 9192
rect -4456 9112 -4360 9128
rect -4456 9048 -4440 9112
rect -4376 9048 -4360 9112
rect -4456 9032 -4360 9048
rect -4456 8968 -4440 9032
rect -4376 8968 -4360 9032
rect -4456 8952 -4360 8968
rect -4456 8888 -4440 8952
rect -4376 8888 -4360 8952
rect -4456 8872 -4360 8888
rect -4456 8808 -4440 8872
rect -4376 8808 -4360 8872
rect -4456 8792 -4360 8808
rect -4456 8728 -4440 8792
rect -4376 8728 -4360 8792
rect -4456 8712 -4360 8728
rect -4456 8648 -4440 8712
rect -4376 8648 -4360 8712
rect -4456 8632 -4360 8648
rect -5868 8532 -5772 8568
rect -4456 8568 -4440 8632
rect -4376 8568 -4360 8632
rect -4037 9312 -3315 9321
rect -4037 8608 -4028 9312
rect -3324 8608 -3315 9312
rect -4037 8599 -3315 8608
rect -3044 9288 -3028 9352
rect -2964 9288 -2948 9352
rect -1632 9352 -1536 9388
rect -3044 9272 -2948 9288
rect -3044 9208 -3028 9272
rect -2964 9208 -2948 9272
rect -3044 9192 -2948 9208
rect -3044 9128 -3028 9192
rect -2964 9128 -2948 9192
rect -3044 9112 -2948 9128
rect -3044 9048 -3028 9112
rect -2964 9048 -2948 9112
rect -3044 9032 -2948 9048
rect -3044 8968 -3028 9032
rect -2964 8968 -2948 9032
rect -3044 8952 -2948 8968
rect -3044 8888 -3028 8952
rect -2964 8888 -2948 8952
rect -3044 8872 -2948 8888
rect -3044 8808 -3028 8872
rect -2964 8808 -2948 8872
rect -3044 8792 -2948 8808
rect -3044 8728 -3028 8792
rect -2964 8728 -2948 8792
rect -3044 8712 -2948 8728
rect -3044 8648 -3028 8712
rect -2964 8648 -2948 8712
rect -3044 8632 -2948 8648
rect -4456 8532 -4360 8568
rect -3044 8568 -3028 8632
rect -2964 8568 -2948 8632
rect -2625 9312 -1903 9321
rect -2625 8608 -2616 9312
rect -1912 8608 -1903 9312
rect -2625 8599 -1903 8608
rect -1632 9288 -1616 9352
rect -1552 9288 -1536 9352
rect -220 9352 -124 9388
rect -1632 9272 -1536 9288
rect -1632 9208 -1616 9272
rect -1552 9208 -1536 9272
rect -1632 9192 -1536 9208
rect -1632 9128 -1616 9192
rect -1552 9128 -1536 9192
rect -1632 9112 -1536 9128
rect -1632 9048 -1616 9112
rect -1552 9048 -1536 9112
rect -1632 9032 -1536 9048
rect -1632 8968 -1616 9032
rect -1552 8968 -1536 9032
rect -1632 8952 -1536 8968
rect -1632 8888 -1616 8952
rect -1552 8888 -1536 8952
rect -1632 8872 -1536 8888
rect -1632 8808 -1616 8872
rect -1552 8808 -1536 8872
rect -1632 8792 -1536 8808
rect -1632 8728 -1616 8792
rect -1552 8728 -1536 8792
rect -1632 8712 -1536 8728
rect -1632 8648 -1616 8712
rect -1552 8648 -1536 8712
rect -1632 8632 -1536 8648
rect -3044 8532 -2948 8568
rect -1632 8568 -1616 8632
rect -1552 8568 -1536 8632
rect -1213 9312 -491 9321
rect -1213 8608 -1204 9312
rect -500 8608 -491 9312
rect -1213 8599 -491 8608
rect -220 9288 -204 9352
rect -140 9288 -124 9352
rect 1192 9352 1288 9388
rect -220 9272 -124 9288
rect -220 9208 -204 9272
rect -140 9208 -124 9272
rect -220 9192 -124 9208
rect -220 9128 -204 9192
rect -140 9128 -124 9192
rect -220 9112 -124 9128
rect -220 9048 -204 9112
rect -140 9048 -124 9112
rect -220 9032 -124 9048
rect -220 8968 -204 9032
rect -140 8968 -124 9032
rect -220 8952 -124 8968
rect -220 8888 -204 8952
rect -140 8888 -124 8952
rect -220 8872 -124 8888
rect -220 8808 -204 8872
rect -140 8808 -124 8872
rect -220 8792 -124 8808
rect -220 8728 -204 8792
rect -140 8728 -124 8792
rect -220 8712 -124 8728
rect -220 8648 -204 8712
rect -140 8648 -124 8712
rect -220 8632 -124 8648
rect -1632 8532 -1536 8568
rect -220 8568 -204 8632
rect -140 8568 -124 8632
rect 199 9312 921 9321
rect 199 8608 208 9312
rect 912 8608 921 9312
rect 199 8599 921 8608
rect 1192 9288 1208 9352
rect 1272 9288 1288 9352
rect 2604 9352 2700 9388
rect 1192 9272 1288 9288
rect 1192 9208 1208 9272
rect 1272 9208 1288 9272
rect 1192 9192 1288 9208
rect 1192 9128 1208 9192
rect 1272 9128 1288 9192
rect 1192 9112 1288 9128
rect 1192 9048 1208 9112
rect 1272 9048 1288 9112
rect 1192 9032 1288 9048
rect 1192 8968 1208 9032
rect 1272 8968 1288 9032
rect 1192 8952 1288 8968
rect 1192 8888 1208 8952
rect 1272 8888 1288 8952
rect 1192 8872 1288 8888
rect 1192 8808 1208 8872
rect 1272 8808 1288 8872
rect 1192 8792 1288 8808
rect 1192 8728 1208 8792
rect 1272 8728 1288 8792
rect 1192 8712 1288 8728
rect 1192 8648 1208 8712
rect 1272 8648 1288 8712
rect 1192 8632 1288 8648
rect -220 8532 -124 8568
rect 1192 8568 1208 8632
rect 1272 8568 1288 8632
rect 1611 9312 2333 9321
rect 1611 8608 1620 9312
rect 2324 8608 2333 9312
rect 1611 8599 2333 8608
rect 2604 9288 2620 9352
rect 2684 9288 2700 9352
rect 4016 9352 4112 9388
rect 2604 9272 2700 9288
rect 2604 9208 2620 9272
rect 2684 9208 2700 9272
rect 2604 9192 2700 9208
rect 2604 9128 2620 9192
rect 2684 9128 2700 9192
rect 2604 9112 2700 9128
rect 2604 9048 2620 9112
rect 2684 9048 2700 9112
rect 2604 9032 2700 9048
rect 2604 8968 2620 9032
rect 2684 8968 2700 9032
rect 2604 8952 2700 8968
rect 2604 8888 2620 8952
rect 2684 8888 2700 8952
rect 2604 8872 2700 8888
rect 2604 8808 2620 8872
rect 2684 8808 2700 8872
rect 2604 8792 2700 8808
rect 2604 8728 2620 8792
rect 2684 8728 2700 8792
rect 2604 8712 2700 8728
rect 2604 8648 2620 8712
rect 2684 8648 2700 8712
rect 2604 8632 2700 8648
rect 1192 8532 1288 8568
rect 2604 8568 2620 8632
rect 2684 8568 2700 8632
rect 3023 9312 3745 9321
rect 3023 8608 3032 9312
rect 3736 8608 3745 9312
rect 3023 8599 3745 8608
rect 4016 9288 4032 9352
rect 4096 9288 4112 9352
rect 5428 9352 5524 9388
rect 4016 9272 4112 9288
rect 4016 9208 4032 9272
rect 4096 9208 4112 9272
rect 4016 9192 4112 9208
rect 4016 9128 4032 9192
rect 4096 9128 4112 9192
rect 4016 9112 4112 9128
rect 4016 9048 4032 9112
rect 4096 9048 4112 9112
rect 4016 9032 4112 9048
rect 4016 8968 4032 9032
rect 4096 8968 4112 9032
rect 4016 8952 4112 8968
rect 4016 8888 4032 8952
rect 4096 8888 4112 8952
rect 4016 8872 4112 8888
rect 4016 8808 4032 8872
rect 4096 8808 4112 8872
rect 4016 8792 4112 8808
rect 4016 8728 4032 8792
rect 4096 8728 4112 8792
rect 4016 8712 4112 8728
rect 4016 8648 4032 8712
rect 4096 8648 4112 8712
rect 4016 8632 4112 8648
rect 2604 8532 2700 8568
rect 4016 8568 4032 8632
rect 4096 8568 4112 8632
rect 4435 9312 5157 9321
rect 4435 8608 4444 9312
rect 5148 8608 5157 9312
rect 4435 8599 5157 8608
rect 5428 9288 5444 9352
rect 5508 9288 5524 9352
rect 6840 9352 6936 9388
rect 5428 9272 5524 9288
rect 5428 9208 5444 9272
rect 5508 9208 5524 9272
rect 5428 9192 5524 9208
rect 5428 9128 5444 9192
rect 5508 9128 5524 9192
rect 5428 9112 5524 9128
rect 5428 9048 5444 9112
rect 5508 9048 5524 9112
rect 5428 9032 5524 9048
rect 5428 8968 5444 9032
rect 5508 8968 5524 9032
rect 5428 8952 5524 8968
rect 5428 8888 5444 8952
rect 5508 8888 5524 8952
rect 5428 8872 5524 8888
rect 5428 8808 5444 8872
rect 5508 8808 5524 8872
rect 5428 8792 5524 8808
rect 5428 8728 5444 8792
rect 5508 8728 5524 8792
rect 5428 8712 5524 8728
rect 5428 8648 5444 8712
rect 5508 8648 5524 8712
rect 5428 8632 5524 8648
rect 4016 8532 4112 8568
rect 5428 8568 5444 8632
rect 5508 8568 5524 8632
rect 5847 9312 6569 9321
rect 5847 8608 5856 9312
rect 6560 8608 6569 9312
rect 5847 8599 6569 8608
rect 6840 9288 6856 9352
rect 6920 9288 6936 9352
rect 8252 9352 8348 9388
rect 6840 9272 6936 9288
rect 6840 9208 6856 9272
rect 6920 9208 6936 9272
rect 6840 9192 6936 9208
rect 6840 9128 6856 9192
rect 6920 9128 6936 9192
rect 6840 9112 6936 9128
rect 6840 9048 6856 9112
rect 6920 9048 6936 9112
rect 6840 9032 6936 9048
rect 6840 8968 6856 9032
rect 6920 8968 6936 9032
rect 6840 8952 6936 8968
rect 6840 8888 6856 8952
rect 6920 8888 6936 8952
rect 6840 8872 6936 8888
rect 6840 8808 6856 8872
rect 6920 8808 6936 8872
rect 6840 8792 6936 8808
rect 6840 8728 6856 8792
rect 6920 8728 6936 8792
rect 6840 8712 6936 8728
rect 6840 8648 6856 8712
rect 6920 8648 6936 8712
rect 6840 8632 6936 8648
rect 5428 8532 5524 8568
rect 6840 8568 6856 8632
rect 6920 8568 6936 8632
rect 7259 9312 7981 9321
rect 7259 8608 7268 9312
rect 7972 8608 7981 9312
rect 7259 8599 7981 8608
rect 8252 9288 8268 9352
rect 8332 9288 8348 9352
rect 9664 9352 9760 9388
rect 8252 9272 8348 9288
rect 8252 9208 8268 9272
rect 8332 9208 8348 9272
rect 8252 9192 8348 9208
rect 8252 9128 8268 9192
rect 8332 9128 8348 9192
rect 8252 9112 8348 9128
rect 8252 9048 8268 9112
rect 8332 9048 8348 9112
rect 8252 9032 8348 9048
rect 8252 8968 8268 9032
rect 8332 8968 8348 9032
rect 8252 8952 8348 8968
rect 8252 8888 8268 8952
rect 8332 8888 8348 8952
rect 8252 8872 8348 8888
rect 8252 8808 8268 8872
rect 8332 8808 8348 8872
rect 8252 8792 8348 8808
rect 8252 8728 8268 8792
rect 8332 8728 8348 8792
rect 8252 8712 8348 8728
rect 8252 8648 8268 8712
rect 8332 8648 8348 8712
rect 8252 8632 8348 8648
rect 6840 8532 6936 8568
rect 8252 8568 8268 8632
rect 8332 8568 8348 8632
rect 8671 9312 9393 9321
rect 8671 8608 8680 9312
rect 9384 8608 9393 9312
rect 8671 8599 9393 8608
rect 9664 9288 9680 9352
rect 9744 9288 9760 9352
rect 11076 9352 11172 9388
rect 9664 9272 9760 9288
rect 9664 9208 9680 9272
rect 9744 9208 9760 9272
rect 9664 9192 9760 9208
rect 9664 9128 9680 9192
rect 9744 9128 9760 9192
rect 9664 9112 9760 9128
rect 9664 9048 9680 9112
rect 9744 9048 9760 9112
rect 9664 9032 9760 9048
rect 9664 8968 9680 9032
rect 9744 8968 9760 9032
rect 9664 8952 9760 8968
rect 9664 8888 9680 8952
rect 9744 8888 9760 8952
rect 9664 8872 9760 8888
rect 9664 8808 9680 8872
rect 9744 8808 9760 8872
rect 9664 8792 9760 8808
rect 9664 8728 9680 8792
rect 9744 8728 9760 8792
rect 9664 8712 9760 8728
rect 9664 8648 9680 8712
rect 9744 8648 9760 8712
rect 9664 8632 9760 8648
rect 8252 8532 8348 8568
rect 9664 8568 9680 8632
rect 9744 8568 9760 8632
rect 10083 9312 10805 9321
rect 10083 8608 10092 9312
rect 10796 8608 10805 9312
rect 10083 8599 10805 8608
rect 11076 9288 11092 9352
rect 11156 9288 11172 9352
rect 12488 9352 12584 9388
rect 11076 9272 11172 9288
rect 11076 9208 11092 9272
rect 11156 9208 11172 9272
rect 11076 9192 11172 9208
rect 11076 9128 11092 9192
rect 11156 9128 11172 9192
rect 11076 9112 11172 9128
rect 11076 9048 11092 9112
rect 11156 9048 11172 9112
rect 11076 9032 11172 9048
rect 11076 8968 11092 9032
rect 11156 8968 11172 9032
rect 11076 8952 11172 8968
rect 11076 8888 11092 8952
rect 11156 8888 11172 8952
rect 11076 8872 11172 8888
rect 11076 8808 11092 8872
rect 11156 8808 11172 8872
rect 11076 8792 11172 8808
rect 11076 8728 11092 8792
rect 11156 8728 11172 8792
rect 11076 8712 11172 8728
rect 11076 8648 11092 8712
rect 11156 8648 11172 8712
rect 11076 8632 11172 8648
rect 9664 8532 9760 8568
rect 11076 8568 11092 8632
rect 11156 8568 11172 8632
rect 11495 9312 12217 9321
rect 11495 8608 11504 9312
rect 12208 8608 12217 9312
rect 11495 8599 12217 8608
rect 12488 9288 12504 9352
rect 12568 9288 12584 9352
rect 13900 9352 13996 9388
rect 12488 9272 12584 9288
rect 12488 9208 12504 9272
rect 12568 9208 12584 9272
rect 12488 9192 12584 9208
rect 12488 9128 12504 9192
rect 12568 9128 12584 9192
rect 12488 9112 12584 9128
rect 12488 9048 12504 9112
rect 12568 9048 12584 9112
rect 12488 9032 12584 9048
rect 12488 8968 12504 9032
rect 12568 8968 12584 9032
rect 12488 8952 12584 8968
rect 12488 8888 12504 8952
rect 12568 8888 12584 8952
rect 12488 8872 12584 8888
rect 12488 8808 12504 8872
rect 12568 8808 12584 8872
rect 12488 8792 12584 8808
rect 12488 8728 12504 8792
rect 12568 8728 12584 8792
rect 12488 8712 12584 8728
rect 12488 8648 12504 8712
rect 12568 8648 12584 8712
rect 12488 8632 12584 8648
rect 11076 8532 11172 8568
rect 12488 8568 12504 8632
rect 12568 8568 12584 8632
rect 12907 9312 13629 9321
rect 12907 8608 12916 9312
rect 13620 8608 13629 9312
rect 12907 8599 13629 8608
rect 13900 9288 13916 9352
rect 13980 9288 13996 9352
rect 15312 9352 15408 9388
rect 13900 9272 13996 9288
rect 13900 9208 13916 9272
rect 13980 9208 13996 9272
rect 13900 9192 13996 9208
rect 13900 9128 13916 9192
rect 13980 9128 13996 9192
rect 13900 9112 13996 9128
rect 13900 9048 13916 9112
rect 13980 9048 13996 9112
rect 13900 9032 13996 9048
rect 13900 8968 13916 9032
rect 13980 8968 13996 9032
rect 13900 8952 13996 8968
rect 13900 8888 13916 8952
rect 13980 8888 13996 8952
rect 13900 8872 13996 8888
rect 13900 8808 13916 8872
rect 13980 8808 13996 8872
rect 13900 8792 13996 8808
rect 13900 8728 13916 8792
rect 13980 8728 13996 8792
rect 13900 8712 13996 8728
rect 13900 8648 13916 8712
rect 13980 8648 13996 8712
rect 13900 8632 13996 8648
rect 12488 8532 12584 8568
rect 13900 8568 13916 8632
rect 13980 8568 13996 8632
rect 14319 9312 15041 9321
rect 14319 8608 14328 9312
rect 15032 8608 15041 9312
rect 14319 8599 15041 8608
rect 15312 9288 15328 9352
rect 15392 9288 15408 9352
rect 16724 9352 16820 9388
rect 15312 9272 15408 9288
rect 15312 9208 15328 9272
rect 15392 9208 15408 9272
rect 15312 9192 15408 9208
rect 15312 9128 15328 9192
rect 15392 9128 15408 9192
rect 15312 9112 15408 9128
rect 15312 9048 15328 9112
rect 15392 9048 15408 9112
rect 15312 9032 15408 9048
rect 15312 8968 15328 9032
rect 15392 8968 15408 9032
rect 15312 8952 15408 8968
rect 15312 8888 15328 8952
rect 15392 8888 15408 8952
rect 15312 8872 15408 8888
rect 15312 8808 15328 8872
rect 15392 8808 15408 8872
rect 15312 8792 15408 8808
rect 15312 8728 15328 8792
rect 15392 8728 15408 8792
rect 15312 8712 15408 8728
rect 15312 8648 15328 8712
rect 15392 8648 15408 8712
rect 15312 8632 15408 8648
rect 13900 8532 13996 8568
rect 15312 8568 15328 8632
rect 15392 8568 15408 8632
rect 15731 9312 16453 9321
rect 15731 8608 15740 9312
rect 16444 8608 16453 9312
rect 15731 8599 16453 8608
rect 16724 9288 16740 9352
rect 16804 9288 16820 9352
rect 18136 9352 18232 9388
rect 16724 9272 16820 9288
rect 16724 9208 16740 9272
rect 16804 9208 16820 9272
rect 16724 9192 16820 9208
rect 16724 9128 16740 9192
rect 16804 9128 16820 9192
rect 16724 9112 16820 9128
rect 16724 9048 16740 9112
rect 16804 9048 16820 9112
rect 16724 9032 16820 9048
rect 16724 8968 16740 9032
rect 16804 8968 16820 9032
rect 16724 8952 16820 8968
rect 16724 8888 16740 8952
rect 16804 8888 16820 8952
rect 16724 8872 16820 8888
rect 16724 8808 16740 8872
rect 16804 8808 16820 8872
rect 16724 8792 16820 8808
rect 16724 8728 16740 8792
rect 16804 8728 16820 8792
rect 16724 8712 16820 8728
rect 16724 8648 16740 8712
rect 16804 8648 16820 8712
rect 16724 8632 16820 8648
rect 15312 8532 15408 8568
rect 16724 8568 16740 8632
rect 16804 8568 16820 8632
rect 17143 9312 17865 9321
rect 17143 8608 17152 9312
rect 17856 8608 17865 9312
rect 17143 8599 17865 8608
rect 18136 9288 18152 9352
rect 18216 9288 18232 9352
rect 19548 9352 19644 9388
rect 18136 9272 18232 9288
rect 18136 9208 18152 9272
rect 18216 9208 18232 9272
rect 18136 9192 18232 9208
rect 18136 9128 18152 9192
rect 18216 9128 18232 9192
rect 18136 9112 18232 9128
rect 18136 9048 18152 9112
rect 18216 9048 18232 9112
rect 18136 9032 18232 9048
rect 18136 8968 18152 9032
rect 18216 8968 18232 9032
rect 18136 8952 18232 8968
rect 18136 8888 18152 8952
rect 18216 8888 18232 8952
rect 18136 8872 18232 8888
rect 18136 8808 18152 8872
rect 18216 8808 18232 8872
rect 18136 8792 18232 8808
rect 18136 8728 18152 8792
rect 18216 8728 18232 8792
rect 18136 8712 18232 8728
rect 18136 8648 18152 8712
rect 18216 8648 18232 8712
rect 18136 8632 18232 8648
rect 16724 8532 16820 8568
rect 18136 8568 18152 8632
rect 18216 8568 18232 8632
rect 18555 9312 19277 9321
rect 18555 8608 18564 9312
rect 19268 8608 19277 9312
rect 18555 8599 19277 8608
rect 19548 9288 19564 9352
rect 19628 9288 19644 9352
rect 20960 9352 21056 9388
rect 19548 9272 19644 9288
rect 19548 9208 19564 9272
rect 19628 9208 19644 9272
rect 19548 9192 19644 9208
rect 19548 9128 19564 9192
rect 19628 9128 19644 9192
rect 19548 9112 19644 9128
rect 19548 9048 19564 9112
rect 19628 9048 19644 9112
rect 19548 9032 19644 9048
rect 19548 8968 19564 9032
rect 19628 8968 19644 9032
rect 19548 8952 19644 8968
rect 19548 8888 19564 8952
rect 19628 8888 19644 8952
rect 19548 8872 19644 8888
rect 19548 8808 19564 8872
rect 19628 8808 19644 8872
rect 19548 8792 19644 8808
rect 19548 8728 19564 8792
rect 19628 8728 19644 8792
rect 19548 8712 19644 8728
rect 19548 8648 19564 8712
rect 19628 8648 19644 8712
rect 19548 8632 19644 8648
rect 18136 8532 18232 8568
rect 19548 8568 19564 8632
rect 19628 8568 19644 8632
rect 19967 9312 20689 9321
rect 19967 8608 19976 9312
rect 20680 8608 20689 9312
rect 19967 8599 20689 8608
rect 20960 9288 20976 9352
rect 21040 9288 21056 9352
rect 22372 9352 22468 9388
rect 20960 9272 21056 9288
rect 20960 9208 20976 9272
rect 21040 9208 21056 9272
rect 20960 9192 21056 9208
rect 20960 9128 20976 9192
rect 21040 9128 21056 9192
rect 20960 9112 21056 9128
rect 20960 9048 20976 9112
rect 21040 9048 21056 9112
rect 20960 9032 21056 9048
rect 20960 8968 20976 9032
rect 21040 8968 21056 9032
rect 20960 8952 21056 8968
rect 20960 8888 20976 8952
rect 21040 8888 21056 8952
rect 20960 8872 21056 8888
rect 20960 8808 20976 8872
rect 21040 8808 21056 8872
rect 20960 8792 21056 8808
rect 20960 8728 20976 8792
rect 21040 8728 21056 8792
rect 20960 8712 21056 8728
rect 20960 8648 20976 8712
rect 21040 8648 21056 8712
rect 20960 8632 21056 8648
rect 19548 8532 19644 8568
rect 20960 8568 20976 8632
rect 21040 8568 21056 8632
rect 21379 9312 22101 9321
rect 21379 8608 21388 9312
rect 22092 8608 22101 9312
rect 21379 8599 22101 8608
rect 22372 9288 22388 9352
rect 22452 9288 22468 9352
rect 23784 9352 23880 9388
rect 22372 9272 22468 9288
rect 22372 9208 22388 9272
rect 22452 9208 22468 9272
rect 22372 9192 22468 9208
rect 22372 9128 22388 9192
rect 22452 9128 22468 9192
rect 22372 9112 22468 9128
rect 22372 9048 22388 9112
rect 22452 9048 22468 9112
rect 22372 9032 22468 9048
rect 22372 8968 22388 9032
rect 22452 8968 22468 9032
rect 22372 8952 22468 8968
rect 22372 8888 22388 8952
rect 22452 8888 22468 8952
rect 22372 8872 22468 8888
rect 22372 8808 22388 8872
rect 22452 8808 22468 8872
rect 22372 8792 22468 8808
rect 22372 8728 22388 8792
rect 22452 8728 22468 8792
rect 22372 8712 22468 8728
rect 22372 8648 22388 8712
rect 22452 8648 22468 8712
rect 22372 8632 22468 8648
rect 20960 8532 21056 8568
rect 22372 8568 22388 8632
rect 22452 8568 22468 8632
rect 22791 9312 23513 9321
rect 22791 8608 22800 9312
rect 23504 8608 23513 9312
rect 22791 8599 23513 8608
rect 23784 9288 23800 9352
rect 23864 9288 23880 9352
rect 23784 9272 23880 9288
rect 23784 9208 23800 9272
rect 23864 9208 23880 9272
rect 23784 9192 23880 9208
rect 23784 9128 23800 9192
rect 23864 9128 23880 9192
rect 23784 9112 23880 9128
rect 23784 9048 23800 9112
rect 23864 9048 23880 9112
rect 23784 9032 23880 9048
rect 23784 8968 23800 9032
rect 23864 8968 23880 9032
rect 23784 8952 23880 8968
rect 23784 8888 23800 8952
rect 23864 8888 23880 8952
rect 23784 8872 23880 8888
rect 23784 8808 23800 8872
rect 23864 8808 23880 8872
rect 23784 8792 23880 8808
rect 23784 8728 23800 8792
rect 23864 8728 23880 8792
rect 23784 8712 23880 8728
rect 23784 8648 23800 8712
rect 23864 8648 23880 8712
rect 23784 8632 23880 8648
rect 22372 8532 22468 8568
rect 23784 8568 23800 8632
rect 23864 8568 23880 8632
rect 23784 8532 23880 8568
rect -22812 8232 -22716 8268
rect -23805 8192 -23083 8201
rect -23805 7488 -23796 8192
rect -23092 7488 -23083 8192
rect -23805 7479 -23083 7488
rect -22812 8168 -22796 8232
rect -22732 8168 -22716 8232
rect -21400 8232 -21304 8268
rect -22812 8152 -22716 8168
rect -22812 8088 -22796 8152
rect -22732 8088 -22716 8152
rect -22812 8072 -22716 8088
rect -22812 8008 -22796 8072
rect -22732 8008 -22716 8072
rect -22812 7992 -22716 8008
rect -22812 7928 -22796 7992
rect -22732 7928 -22716 7992
rect -22812 7912 -22716 7928
rect -22812 7848 -22796 7912
rect -22732 7848 -22716 7912
rect -22812 7832 -22716 7848
rect -22812 7768 -22796 7832
rect -22732 7768 -22716 7832
rect -22812 7752 -22716 7768
rect -22812 7688 -22796 7752
rect -22732 7688 -22716 7752
rect -22812 7672 -22716 7688
rect -22812 7608 -22796 7672
rect -22732 7608 -22716 7672
rect -22812 7592 -22716 7608
rect -22812 7528 -22796 7592
rect -22732 7528 -22716 7592
rect -22812 7512 -22716 7528
rect -22812 7448 -22796 7512
rect -22732 7448 -22716 7512
rect -22393 8192 -21671 8201
rect -22393 7488 -22384 8192
rect -21680 7488 -21671 8192
rect -22393 7479 -21671 7488
rect -21400 8168 -21384 8232
rect -21320 8168 -21304 8232
rect -19988 8232 -19892 8268
rect -21400 8152 -21304 8168
rect -21400 8088 -21384 8152
rect -21320 8088 -21304 8152
rect -21400 8072 -21304 8088
rect -21400 8008 -21384 8072
rect -21320 8008 -21304 8072
rect -21400 7992 -21304 8008
rect -21400 7928 -21384 7992
rect -21320 7928 -21304 7992
rect -21400 7912 -21304 7928
rect -21400 7848 -21384 7912
rect -21320 7848 -21304 7912
rect -21400 7832 -21304 7848
rect -21400 7768 -21384 7832
rect -21320 7768 -21304 7832
rect -21400 7752 -21304 7768
rect -21400 7688 -21384 7752
rect -21320 7688 -21304 7752
rect -21400 7672 -21304 7688
rect -21400 7608 -21384 7672
rect -21320 7608 -21304 7672
rect -21400 7592 -21304 7608
rect -21400 7528 -21384 7592
rect -21320 7528 -21304 7592
rect -21400 7512 -21304 7528
rect -22812 7412 -22716 7448
rect -21400 7448 -21384 7512
rect -21320 7448 -21304 7512
rect -20981 8192 -20259 8201
rect -20981 7488 -20972 8192
rect -20268 7488 -20259 8192
rect -20981 7479 -20259 7488
rect -19988 8168 -19972 8232
rect -19908 8168 -19892 8232
rect -18576 8232 -18480 8268
rect -19988 8152 -19892 8168
rect -19988 8088 -19972 8152
rect -19908 8088 -19892 8152
rect -19988 8072 -19892 8088
rect -19988 8008 -19972 8072
rect -19908 8008 -19892 8072
rect -19988 7992 -19892 8008
rect -19988 7928 -19972 7992
rect -19908 7928 -19892 7992
rect -19988 7912 -19892 7928
rect -19988 7848 -19972 7912
rect -19908 7848 -19892 7912
rect -19988 7832 -19892 7848
rect -19988 7768 -19972 7832
rect -19908 7768 -19892 7832
rect -19988 7752 -19892 7768
rect -19988 7688 -19972 7752
rect -19908 7688 -19892 7752
rect -19988 7672 -19892 7688
rect -19988 7608 -19972 7672
rect -19908 7608 -19892 7672
rect -19988 7592 -19892 7608
rect -19988 7528 -19972 7592
rect -19908 7528 -19892 7592
rect -19988 7512 -19892 7528
rect -21400 7412 -21304 7448
rect -19988 7448 -19972 7512
rect -19908 7448 -19892 7512
rect -19569 8192 -18847 8201
rect -19569 7488 -19560 8192
rect -18856 7488 -18847 8192
rect -19569 7479 -18847 7488
rect -18576 8168 -18560 8232
rect -18496 8168 -18480 8232
rect -17164 8232 -17068 8268
rect -18576 8152 -18480 8168
rect -18576 8088 -18560 8152
rect -18496 8088 -18480 8152
rect -18576 8072 -18480 8088
rect -18576 8008 -18560 8072
rect -18496 8008 -18480 8072
rect -18576 7992 -18480 8008
rect -18576 7928 -18560 7992
rect -18496 7928 -18480 7992
rect -18576 7912 -18480 7928
rect -18576 7848 -18560 7912
rect -18496 7848 -18480 7912
rect -18576 7832 -18480 7848
rect -18576 7768 -18560 7832
rect -18496 7768 -18480 7832
rect -18576 7752 -18480 7768
rect -18576 7688 -18560 7752
rect -18496 7688 -18480 7752
rect -18576 7672 -18480 7688
rect -18576 7608 -18560 7672
rect -18496 7608 -18480 7672
rect -18576 7592 -18480 7608
rect -18576 7528 -18560 7592
rect -18496 7528 -18480 7592
rect -18576 7512 -18480 7528
rect -19988 7412 -19892 7448
rect -18576 7448 -18560 7512
rect -18496 7448 -18480 7512
rect -18157 8192 -17435 8201
rect -18157 7488 -18148 8192
rect -17444 7488 -17435 8192
rect -18157 7479 -17435 7488
rect -17164 8168 -17148 8232
rect -17084 8168 -17068 8232
rect -15752 8232 -15656 8268
rect -17164 8152 -17068 8168
rect -17164 8088 -17148 8152
rect -17084 8088 -17068 8152
rect -17164 8072 -17068 8088
rect -17164 8008 -17148 8072
rect -17084 8008 -17068 8072
rect -17164 7992 -17068 8008
rect -17164 7928 -17148 7992
rect -17084 7928 -17068 7992
rect -17164 7912 -17068 7928
rect -17164 7848 -17148 7912
rect -17084 7848 -17068 7912
rect -17164 7832 -17068 7848
rect -17164 7768 -17148 7832
rect -17084 7768 -17068 7832
rect -17164 7752 -17068 7768
rect -17164 7688 -17148 7752
rect -17084 7688 -17068 7752
rect -17164 7672 -17068 7688
rect -17164 7608 -17148 7672
rect -17084 7608 -17068 7672
rect -17164 7592 -17068 7608
rect -17164 7528 -17148 7592
rect -17084 7528 -17068 7592
rect -17164 7512 -17068 7528
rect -18576 7412 -18480 7448
rect -17164 7448 -17148 7512
rect -17084 7448 -17068 7512
rect -16745 8192 -16023 8201
rect -16745 7488 -16736 8192
rect -16032 7488 -16023 8192
rect -16745 7479 -16023 7488
rect -15752 8168 -15736 8232
rect -15672 8168 -15656 8232
rect -14340 8232 -14244 8268
rect -15752 8152 -15656 8168
rect -15752 8088 -15736 8152
rect -15672 8088 -15656 8152
rect -15752 8072 -15656 8088
rect -15752 8008 -15736 8072
rect -15672 8008 -15656 8072
rect -15752 7992 -15656 8008
rect -15752 7928 -15736 7992
rect -15672 7928 -15656 7992
rect -15752 7912 -15656 7928
rect -15752 7848 -15736 7912
rect -15672 7848 -15656 7912
rect -15752 7832 -15656 7848
rect -15752 7768 -15736 7832
rect -15672 7768 -15656 7832
rect -15752 7752 -15656 7768
rect -15752 7688 -15736 7752
rect -15672 7688 -15656 7752
rect -15752 7672 -15656 7688
rect -15752 7608 -15736 7672
rect -15672 7608 -15656 7672
rect -15752 7592 -15656 7608
rect -15752 7528 -15736 7592
rect -15672 7528 -15656 7592
rect -15752 7512 -15656 7528
rect -17164 7412 -17068 7448
rect -15752 7448 -15736 7512
rect -15672 7448 -15656 7512
rect -15333 8192 -14611 8201
rect -15333 7488 -15324 8192
rect -14620 7488 -14611 8192
rect -15333 7479 -14611 7488
rect -14340 8168 -14324 8232
rect -14260 8168 -14244 8232
rect -12928 8232 -12832 8268
rect -14340 8152 -14244 8168
rect -14340 8088 -14324 8152
rect -14260 8088 -14244 8152
rect -14340 8072 -14244 8088
rect -14340 8008 -14324 8072
rect -14260 8008 -14244 8072
rect -14340 7992 -14244 8008
rect -14340 7928 -14324 7992
rect -14260 7928 -14244 7992
rect -14340 7912 -14244 7928
rect -14340 7848 -14324 7912
rect -14260 7848 -14244 7912
rect -14340 7832 -14244 7848
rect -14340 7768 -14324 7832
rect -14260 7768 -14244 7832
rect -14340 7752 -14244 7768
rect -14340 7688 -14324 7752
rect -14260 7688 -14244 7752
rect -14340 7672 -14244 7688
rect -14340 7608 -14324 7672
rect -14260 7608 -14244 7672
rect -14340 7592 -14244 7608
rect -14340 7528 -14324 7592
rect -14260 7528 -14244 7592
rect -14340 7512 -14244 7528
rect -15752 7412 -15656 7448
rect -14340 7448 -14324 7512
rect -14260 7448 -14244 7512
rect -13921 8192 -13199 8201
rect -13921 7488 -13912 8192
rect -13208 7488 -13199 8192
rect -13921 7479 -13199 7488
rect -12928 8168 -12912 8232
rect -12848 8168 -12832 8232
rect -11516 8232 -11420 8268
rect -12928 8152 -12832 8168
rect -12928 8088 -12912 8152
rect -12848 8088 -12832 8152
rect -12928 8072 -12832 8088
rect -12928 8008 -12912 8072
rect -12848 8008 -12832 8072
rect -12928 7992 -12832 8008
rect -12928 7928 -12912 7992
rect -12848 7928 -12832 7992
rect -12928 7912 -12832 7928
rect -12928 7848 -12912 7912
rect -12848 7848 -12832 7912
rect -12928 7832 -12832 7848
rect -12928 7768 -12912 7832
rect -12848 7768 -12832 7832
rect -12928 7752 -12832 7768
rect -12928 7688 -12912 7752
rect -12848 7688 -12832 7752
rect -12928 7672 -12832 7688
rect -12928 7608 -12912 7672
rect -12848 7608 -12832 7672
rect -12928 7592 -12832 7608
rect -12928 7528 -12912 7592
rect -12848 7528 -12832 7592
rect -12928 7512 -12832 7528
rect -14340 7412 -14244 7448
rect -12928 7448 -12912 7512
rect -12848 7448 -12832 7512
rect -12509 8192 -11787 8201
rect -12509 7488 -12500 8192
rect -11796 7488 -11787 8192
rect -12509 7479 -11787 7488
rect -11516 8168 -11500 8232
rect -11436 8168 -11420 8232
rect -10104 8232 -10008 8268
rect -11516 8152 -11420 8168
rect -11516 8088 -11500 8152
rect -11436 8088 -11420 8152
rect -11516 8072 -11420 8088
rect -11516 8008 -11500 8072
rect -11436 8008 -11420 8072
rect -11516 7992 -11420 8008
rect -11516 7928 -11500 7992
rect -11436 7928 -11420 7992
rect -11516 7912 -11420 7928
rect -11516 7848 -11500 7912
rect -11436 7848 -11420 7912
rect -11516 7832 -11420 7848
rect -11516 7768 -11500 7832
rect -11436 7768 -11420 7832
rect -11516 7752 -11420 7768
rect -11516 7688 -11500 7752
rect -11436 7688 -11420 7752
rect -11516 7672 -11420 7688
rect -11516 7608 -11500 7672
rect -11436 7608 -11420 7672
rect -11516 7592 -11420 7608
rect -11516 7528 -11500 7592
rect -11436 7528 -11420 7592
rect -11516 7512 -11420 7528
rect -12928 7412 -12832 7448
rect -11516 7448 -11500 7512
rect -11436 7448 -11420 7512
rect -11097 8192 -10375 8201
rect -11097 7488 -11088 8192
rect -10384 7488 -10375 8192
rect -11097 7479 -10375 7488
rect -10104 8168 -10088 8232
rect -10024 8168 -10008 8232
rect -8692 8232 -8596 8268
rect -10104 8152 -10008 8168
rect -10104 8088 -10088 8152
rect -10024 8088 -10008 8152
rect -10104 8072 -10008 8088
rect -10104 8008 -10088 8072
rect -10024 8008 -10008 8072
rect -10104 7992 -10008 8008
rect -10104 7928 -10088 7992
rect -10024 7928 -10008 7992
rect -10104 7912 -10008 7928
rect -10104 7848 -10088 7912
rect -10024 7848 -10008 7912
rect -10104 7832 -10008 7848
rect -10104 7768 -10088 7832
rect -10024 7768 -10008 7832
rect -10104 7752 -10008 7768
rect -10104 7688 -10088 7752
rect -10024 7688 -10008 7752
rect -10104 7672 -10008 7688
rect -10104 7608 -10088 7672
rect -10024 7608 -10008 7672
rect -10104 7592 -10008 7608
rect -10104 7528 -10088 7592
rect -10024 7528 -10008 7592
rect -10104 7512 -10008 7528
rect -11516 7412 -11420 7448
rect -10104 7448 -10088 7512
rect -10024 7448 -10008 7512
rect -9685 8192 -8963 8201
rect -9685 7488 -9676 8192
rect -8972 7488 -8963 8192
rect -9685 7479 -8963 7488
rect -8692 8168 -8676 8232
rect -8612 8168 -8596 8232
rect -7280 8232 -7184 8268
rect -8692 8152 -8596 8168
rect -8692 8088 -8676 8152
rect -8612 8088 -8596 8152
rect -8692 8072 -8596 8088
rect -8692 8008 -8676 8072
rect -8612 8008 -8596 8072
rect -8692 7992 -8596 8008
rect -8692 7928 -8676 7992
rect -8612 7928 -8596 7992
rect -8692 7912 -8596 7928
rect -8692 7848 -8676 7912
rect -8612 7848 -8596 7912
rect -8692 7832 -8596 7848
rect -8692 7768 -8676 7832
rect -8612 7768 -8596 7832
rect -8692 7752 -8596 7768
rect -8692 7688 -8676 7752
rect -8612 7688 -8596 7752
rect -8692 7672 -8596 7688
rect -8692 7608 -8676 7672
rect -8612 7608 -8596 7672
rect -8692 7592 -8596 7608
rect -8692 7528 -8676 7592
rect -8612 7528 -8596 7592
rect -8692 7512 -8596 7528
rect -10104 7412 -10008 7448
rect -8692 7448 -8676 7512
rect -8612 7448 -8596 7512
rect -8273 8192 -7551 8201
rect -8273 7488 -8264 8192
rect -7560 7488 -7551 8192
rect -8273 7479 -7551 7488
rect -7280 8168 -7264 8232
rect -7200 8168 -7184 8232
rect -5868 8232 -5772 8268
rect -7280 8152 -7184 8168
rect -7280 8088 -7264 8152
rect -7200 8088 -7184 8152
rect -7280 8072 -7184 8088
rect -7280 8008 -7264 8072
rect -7200 8008 -7184 8072
rect -7280 7992 -7184 8008
rect -7280 7928 -7264 7992
rect -7200 7928 -7184 7992
rect -7280 7912 -7184 7928
rect -7280 7848 -7264 7912
rect -7200 7848 -7184 7912
rect -7280 7832 -7184 7848
rect -7280 7768 -7264 7832
rect -7200 7768 -7184 7832
rect -7280 7752 -7184 7768
rect -7280 7688 -7264 7752
rect -7200 7688 -7184 7752
rect -7280 7672 -7184 7688
rect -7280 7608 -7264 7672
rect -7200 7608 -7184 7672
rect -7280 7592 -7184 7608
rect -7280 7528 -7264 7592
rect -7200 7528 -7184 7592
rect -7280 7512 -7184 7528
rect -8692 7412 -8596 7448
rect -7280 7448 -7264 7512
rect -7200 7448 -7184 7512
rect -6861 8192 -6139 8201
rect -6861 7488 -6852 8192
rect -6148 7488 -6139 8192
rect -6861 7479 -6139 7488
rect -5868 8168 -5852 8232
rect -5788 8168 -5772 8232
rect -4456 8232 -4360 8268
rect -5868 8152 -5772 8168
rect -5868 8088 -5852 8152
rect -5788 8088 -5772 8152
rect -5868 8072 -5772 8088
rect -5868 8008 -5852 8072
rect -5788 8008 -5772 8072
rect -5868 7992 -5772 8008
rect -5868 7928 -5852 7992
rect -5788 7928 -5772 7992
rect -5868 7912 -5772 7928
rect -5868 7848 -5852 7912
rect -5788 7848 -5772 7912
rect -5868 7832 -5772 7848
rect -5868 7768 -5852 7832
rect -5788 7768 -5772 7832
rect -5868 7752 -5772 7768
rect -5868 7688 -5852 7752
rect -5788 7688 -5772 7752
rect -5868 7672 -5772 7688
rect -5868 7608 -5852 7672
rect -5788 7608 -5772 7672
rect -5868 7592 -5772 7608
rect -5868 7528 -5852 7592
rect -5788 7528 -5772 7592
rect -5868 7512 -5772 7528
rect -7280 7412 -7184 7448
rect -5868 7448 -5852 7512
rect -5788 7448 -5772 7512
rect -5449 8192 -4727 8201
rect -5449 7488 -5440 8192
rect -4736 7488 -4727 8192
rect -5449 7479 -4727 7488
rect -4456 8168 -4440 8232
rect -4376 8168 -4360 8232
rect -3044 8232 -2948 8268
rect -4456 8152 -4360 8168
rect -4456 8088 -4440 8152
rect -4376 8088 -4360 8152
rect -4456 8072 -4360 8088
rect -4456 8008 -4440 8072
rect -4376 8008 -4360 8072
rect -4456 7992 -4360 8008
rect -4456 7928 -4440 7992
rect -4376 7928 -4360 7992
rect -4456 7912 -4360 7928
rect -4456 7848 -4440 7912
rect -4376 7848 -4360 7912
rect -4456 7832 -4360 7848
rect -4456 7768 -4440 7832
rect -4376 7768 -4360 7832
rect -4456 7752 -4360 7768
rect -4456 7688 -4440 7752
rect -4376 7688 -4360 7752
rect -4456 7672 -4360 7688
rect -4456 7608 -4440 7672
rect -4376 7608 -4360 7672
rect -4456 7592 -4360 7608
rect -4456 7528 -4440 7592
rect -4376 7528 -4360 7592
rect -4456 7512 -4360 7528
rect -5868 7412 -5772 7448
rect -4456 7448 -4440 7512
rect -4376 7448 -4360 7512
rect -4037 8192 -3315 8201
rect -4037 7488 -4028 8192
rect -3324 7488 -3315 8192
rect -4037 7479 -3315 7488
rect -3044 8168 -3028 8232
rect -2964 8168 -2948 8232
rect -1632 8232 -1536 8268
rect -3044 8152 -2948 8168
rect -3044 8088 -3028 8152
rect -2964 8088 -2948 8152
rect -3044 8072 -2948 8088
rect -3044 8008 -3028 8072
rect -2964 8008 -2948 8072
rect -3044 7992 -2948 8008
rect -3044 7928 -3028 7992
rect -2964 7928 -2948 7992
rect -3044 7912 -2948 7928
rect -3044 7848 -3028 7912
rect -2964 7848 -2948 7912
rect -3044 7832 -2948 7848
rect -3044 7768 -3028 7832
rect -2964 7768 -2948 7832
rect -3044 7752 -2948 7768
rect -3044 7688 -3028 7752
rect -2964 7688 -2948 7752
rect -3044 7672 -2948 7688
rect -3044 7608 -3028 7672
rect -2964 7608 -2948 7672
rect -3044 7592 -2948 7608
rect -3044 7528 -3028 7592
rect -2964 7528 -2948 7592
rect -3044 7512 -2948 7528
rect -4456 7412 -4360 7448
rect -3044 7448 -3028 7512
rect -2964 7448 -2948 7512
rect -2625 8192 -1903 8201
rect -2625 7488 -2616 8192
rect -1912 7488 -1903 8192
rect -2625 7479 -1903 7488
rect -1632 8168 -1616 8232
rect -1552 8168 -1536 8232
rect -220 8232 -124 8268
rect -1632 8152 -1536 8168
rect -1632 8088 -1616 8152
rect -1552 8088 -1536 8152
rect -1632 8072 -1536 8088
rect -1632 8008 -1616 8072
rect -1552 8008 -1536 8072
rect -1632 7992 -1536 8008
rect -1632 7928 -1616 7992
rect -1552 7928 -1536 7992
rect -1632 7912 -1536 7928
rect -1632 7848 -1616 7912
rect -1552 7848 -1536 7912
rect -1632 7832 -1536 7848
rect -1632 7768 -1616 7832
rect -1552 7768 -1536 7832
rect -1632 7752 -1536 7768
rect -1632 7688 -1616 7752
rect -1552 7688 -1536 7752
rect -1632 7672 -1536 7688
rect -1632 7608 -1616 7672
rect -1552 7608 -1536 7672
rect -1632 7592 -1536 7608
rect -1632 7528 -1616 7592
rect -1552 7528 -1536 7592
rect -1632 7512 -1536 7528
rect -3044 7412 -2948 7448
rect -1632 7448 -1616 7512
rect -1552 7448 -1536 7512
rect -1213 8192 -491 8201
rect -1213 7488 -1204 8192
rect -500 7488 -491 8192
rect -1213 7479 -491 7488
rect -220 8168 -204 8232
rect -140 8168 -124 8232
rect 1192 8232 1288 8268
rect -220 8152 -124 8168
rect -220 8088 -204 8152
rect -140 8088 -124 8152
rect -220 8072 -124 8088
rect -220 8008 -204 8072
rect -140 8008 -124 8072
rect -220 7992 -124 8008
rect -220 7928 -204 7992
rect -140 7928 -124 7992
rect -220 7912 -124 7928
rect -220 7848 -204 7912
rect -140 7848 -124 7912
rect -220 7832 -124 7848
rect -220 7768 -204 7832
rect -140 7768 -124 7832
rect -220 7752 -124 7768
rect -220 7688 -204 7752
rect -140 7688 -124 7752
rect -220 7672 -124 7688
rect -220 7608 -204 7672
rect -140 7608 -124 7672
rect -220 7592 -124 7608
rect -220 7528 -204 7592
rect -140 7528 -124 7592
rect -220 7512 -124 7528
rect -1632 7412 -1536 7448
rect -220 7448 -204 7512
rect -140 7448 -124 7512
rect 199 8192 921 8201
rect 199 7488 208 8192
rect 912 7488 921 8192
rect 199 7479 921 7488
rect 1192 8168 1208 8232
rect 1272 8168 1288 8232
rect 2604 8232 2700 8268
rect 1192 8152 1288 8168
rect 1192 8088 1208 8152
rect 1272 8088 1288 8152
rect 1192 8072 1288 8088
rect 1192 8008 1208 8072
rect 1272 8008 1288 8072
rect 1192 7992 1288 8008
rect 1192 7928 1208 7992
rect 1272 7928 1288 7992
rect 1192 7912 1288 7928
rect 1192 7848 1208 7912
rect 1272 7848 1288 7912
rect 1192 7832 1288 7848
rect 1192 7768 1208 7832
rect 1272 7768 1288 7832
rect 1192 7752 1288 7768
rect 1192 7688 1208 7752
rect 1272 7688 1288 7752
rect 1192 7672 1288 7688
rect 1192 7608 1208 7672
rect 1272 7608 1288 7672
rect 1192 7592 1288 7608
rect 1192 7528 1208 7592
rect 1272 7528 1288 7592
rect 1192 7512 1288 7528
rect -220 7412 -124 7448
rect 1192 7448 1208 7512
rect 1272 7448 1288 7512
rect 1611 8192 2333 8201
rect 1611 7488 1620 8192
rect 2324 7488 2333 8192
rect 1611 7479 2333 7488
rect 2604 8168 2620 8232
rect 2684 8168 2700 8232
rect 4016 8232 4112 8268
rect 2604 8152 2700 8168
rect 2604 8088 2620 8152
rect 2684 8088 2700 8152
rect 2604 8072 2700 8088
rect 2604 8008 2620 8072
rect 2684 8008 2700 8072
rect 2604 7992 2700 8008
rect 2604 7928 2620 7992
rect 2684 7928 2700 7992
rect 2604 7912 2700 7928
rect 2604 7848 2620 7912
rect 2684 7848 2700 7912
rect 2604 7832 2700 7848
rect 2604 7768 2620 7832
rect 2684 7768 2700 7832
rect 2604 7752 2700 7768
rect 2604 7688 2620 7752
rect 2684 7688 2700 7752
rect 2604 7672 2700 7688
rect 2604 7608 2620 7672
rect 2684 7608 2700 7672
rect 2604 7592 2700 7608
rect 2604 7528 2620 7592
rect 2684 7528 2700 7592
rect 2604 7512 2700 7528
rect 1192 7412 1288 7448
rect 2604 7448 2620 7512
rect 2684 7448 2700 7512
rect 3023 8192 3745 8201
rect 3023 7488 3032 8192
rect 3736 7488 3745 8192
rect 3023 7479 3745 7488
rect 4016 8168 4032 8232
rect 4096 8168 4112 8232
rect 5428 8232 5524 8268
rect 4016 8152 4112 8168
rect 4016 8088 4032 8152
rect 4096 8088 4112 8152
rect 4016 8072 4112 8088
rect 4016 8008 4032 8072
rect 4096 8008 4112 8072
rect 4016 7992 4112 8008
rect 4016 7928 4032 7992
rect 4096 7928 4112 7992
rect 4016 7912 4112 7928
rect 4016 7848 4032 7912
rect 4096 7848 4112 7912
rect 4016 7832 4112 7848
rect 4016 7768 4032 7832
rect 4096 7768 4112 7832
rect 4016 7752 4112 7768
rect 4016 7688 4032 7752
rect 4096 7688 4112 7752
rect 4016 7672 4112 7688
rect 4016 7608 4032 7672
rect 4096 7608 4112 7672
rect 4016 7592 4112 7608
rect 4016 7528 4032 7592
rect 4096 7528 4112 7592
rect 4016 7512 4112 7528
rect 2604 7412 2700 7448
rect 4016 7448 4032 7512
rect 4096 7448 4112 7512
rect 4435 8192 5157 8201
rect 4435 7488 4444 8192
rect 5148 7488 5157 8192
rect 4435 7479 5157 7488
rect 5428 8168 5444 8232
rect 5508 8168 5524 8232
rect 6840 8232 6936 8268
rect 5428 8152 5524 8168
rect 5428 8088 5444 8152
rect 5508 8088 5524 8152
rect 5428 8072 5524 8088
rect 5428 8008 5444 8072
rect 5508 8008 5524 8072
rect 5428 7992 5524 8008
rect 5428 7928 5444 7992
rect 5508 7928 5524 7992
rect 5428 7912 5524 7928
rect 5428 7848 5444 7912
rect 5508 7848 5524 7912
rect 5428 7832 5524 7848
rect 5428 7768 5444 7832
rect 5508 7768 5524 7832
rect 5428 7752 5524 7768
rect 5428 7688 5444 7752
rect 5508 7688 5524 7752
rect 5428 7672 5524 7688
rect 5428 7608 5444 7672
rect 5508 7608 5524 7672
rect 5428 7592 5524 7608
rect 5428 7528 5444 7592
rect 5508 7528 5524 7592
rect 5428 7512 5524 7528
rect 4016 7412 4112 7448
rect 5428 7448 5444 7512
rect 5508 7448 5524 7512
rect 5847 8192 6569 8201
rect 5847 7488 5856 8192
rect 6560 7488 6569 8192
rect 5847 7479 6569 7488
rect 6840 8168 6856 8232
rect 6920 8168 6936 8232
rect 8252 8232 8348 8268
rect 6840 8152 6936 8168
rect 6840 8088 6856 8152
rect 6920 8088 6936 8152
rect 6840 8072 6936 8088
rect 6840 8008 6856 8072
rect 6920 8008 6936 8072
rect 6840 7992 6936 8008
rect 6840 7928 6856 7992
rect 6920 7928 6936 7992
rect 6840 7912 6936 7928
rect 6840 7848 6856 7912
rect 6920 7848 6936 7912
rect 6840 7832 6936 7848
rect 6840 7768 6856 7832
rect 6920 7768 6936 7832
rect 6840 7752 6936 7768
rect 6840 7688 6856 7752
rect 6920 7688 6936 7752
rect 6840 7672 6936 7688
rect 6840 7608 6856 7672
rect 6920 7608 6936 7672
rect 6840 7592 6936 7608
rect 6840 7528 6856 7592
rect 6920 7528 6936 7592
rect 6840 7512 6936 7528
rect 5428 7412 5524 7448
rect 6840 7448 6856 7512
rect 6920 7448 6936 7512
rect 7259 8192 7981 8201
rect 7259 7488 7268 8192
rect 7972 7488 7981 8192
rect 7259 7479 7981 7488
rect 8252 8168 8268 8232
rect 8332 8168 8348 8232
rect 9664 8232 9760 8268
rect 8252 8152 8348 8168
rect 8252 8088 8268 8152
rect 8332 8088 8348 8152
rect 8252 8072 8348 8088
rect 8252 8008 8268 8072
rect 8332 8008 8348 8072
rect 8252 7992 8348 8008
rect 8252 7928 8268 7992
rect 8332 7928 8348 7992
rect 8252 7912 8348 7928
rect 8252 7848 8268 7912
rect 8332 7848 8348 7912
rect 8252 7832 8348 7848
rect 8252 7768 8268 7832
rect 8332 7768 8348 7832
rect 8252 7752 8348 7768
rect 8252 7688 8268 7752
rect 8332 7688 8348 7752
rect 8252 7672 8348 7688
rect 8252 7608 8268 7672
rect 8332 7608 8348 7672
rect 8252 7592 8348 7608
rect 8252 7528 8268 7592
rect 8332 7528 8348 7592
rect 8252 7512 8348 7528
rect 6840 7412 6936 7448
rect 8252 7448 8268 7512
rect 8332 7448 8348 7512
rect 8671 8192 9393 8201
rect 8671 7488 8680 8192
rect 9384 7488 9393 8192
rect 8671 7479 9393 7488
rect 9664 8168 9680 8232
rect 9744 8168 9760 8232
rect 11076 8232 11172 8268
rect 9664 8152 9760 8168
rect 9664 8088 9680 8152
rect 9744 8088 9760 8152
rect 9664 8072 9760 8088
rect 9664 8008 9680 8072
rect 9744 8008 9760 8072
rect 9664 7992 9760 8008
rect 9664 7928 9680 7992
rect 9744 7928 9760 7992
rect 9664 7912 9760 7928
rect 9664 7848 9680 7912
rect 9744 7848 9760 7912
rect 9664 7832 9760 7848
rect 9664 7768 9680 7832
rect 9744 7768 9760 7832
rect 9664 7752 9760 7768
rect 9664 7688 9680 7752
rect 9744 7688 9760 7752
rect 9664 7672 9760 7688
rect 9664 7608 9680 7672
rect 9744 7608 9760 7672
rect 9664 7592 9760 7608
rect 9664 7528 9680 7592
rect 9744 7528 9760 7592
rect 9664 7512 9760 7528
rect 8252 7412 8348 7448
rect 9664 7448 9680 7512
rect 9744 7448 9760 7512
rect 10083 8192 10805 8201
rect 10083 7488 10092 8192
rect 10796 7488 10805 8192
rect 10083 7479 10805 7488
rect 11076 8168 11092 8232
rect 11156 8168 11172 8232
rect 12488 8232 12584 8268
rect 11076 8152 11172 8168
rect 11076 8088 11092 8152
rect 11156 8088 11172 8152
rect 11076 8072 11172 8088
rect 11076 8008 11092 8072
rect 11156 8008 11172 8072
rect 11076 7992 11172 8008
rect 11076 7928 11092 7992
rect 11156 7928 11172 7992
rect 11076 7912 11172 7928
rect 11076 7848 11092 7912
rect 11156 7848 11172 7912
rect 11076 7832 11172 7848
rect 11076 7768 11092 7832
rect 11156 7768 11172 7832
rect 11076 7752 11172 7768
rect 11076 7688 11092 7752
rect 11156 7688 11172 7752
rect 11076 7672 11172 7688
rect 11076 7608 11092 7672
rect 11156 7608 11172 7672
rect 11076 7592 11172 7608
rect 11076 7528 11092 7592
rect 11156 7528 11172 7592
rect 11076 7512 11172 7528
rect 9664 7412 9760 7448
rect 11076 7448 11092 7512
rect 11156 7448 11172 7512
rect 11495 8192 12217 8201
rect 11495 7488 11504 8192
rect 12208 7488 12217 8192
rect 11495 7479 12217 7488
rect 12488 8168 12504 8232
rect 12568 8168 12584 8232
rect 13900 8232 13996 8268
rect 12488 8152 12584 8168
rect 12488 8088 12504 8152
rect 12568 8088 12584 8152
rect 12488 8072 12584 8088
rect 12488 8008 12504 8072
rect 12568 8008 12584 8072
rect 12488 7992 12584 8008
rect 12488 7928 12504 7992
rect 12568 7928 12584 7992
rect 12488 7912 12584 7928
rect 12488 7848 12504 7912
rect 12568 7848 12584 7912
rect 12488 7832 12584 7848
rect 12488 7768 12504 7832
rect 12568 7768 12584 7832
rect 12488 7752 12584 7768
rect 12488 7688 12504 7752
rect 12568 7688 12584 7752
rect 12488 7672 12584 7688
rect 12488 7608 12504 7672
rect 12568 7608 12584 7672
rect 12488 7592 12584 7608
rect 12488 7528 12504 7592
rect 12568 7528 12584 7592
rect 12488 7512 12584 7528
rect 11076 7412 11172 7448
rect 12488 7448 12504 7512
rect 12568 7448 12584 7512
rect 12907 8192 13629 8201
rect 12907 7488 12916 8192
rect 13620 7488 13629 8192
rect 12907 7479 13629 7488
rect 13900 8168 13916 8232
rect 13980 8168 13996 8232
rect 15312 8232 15408 8268
rect 13900 8152 13996 8168
rect 13900 8088 13916 8152
rect 13980 8088 13996 8152
rect 13900 8072 13996 8088
rect 13900 8008 13916 8072
rect 13980 8008 13996 8072
rect 13900 7992 13996 8008
rect 13900 7928 13916 7992
rect 13980 7928 13996 7992
rect 13900 7912 13996 7928
rect 13900 7848 13916 7912
rect 13980 7848 13996 7912
rect 13900 7832 13996 7848
rect 13900 7768 13916 7832
rect 13980 7768 13996 7832
rect 13900 7752 13996 7768
rect 13900 7688 13916 7752
rect 13980 7688 13996 7752
rect 13900 7672 13996 7688
rect 13900 7608 13916 7672
rect 13980 7608 13996 7672
rect 13900 7592 13996 7608
rect 13900 7528 13916 7592
rect 13980 7528 13996 7592
rect 13900 7512 13996 7528
rect 12488 7412 12584 7448
rect 13900 7448 13916 7512
rect 13980 7448 13996 7512
rect 14319 8192 15041 8201
rect 14319 7488 14328 8192
rect 15032 7488 15041 8192
rect 14319 7479 15041 7488
rect 15312 8168 15328 8232
rect 15392 8168 15408 8232
rect 16724 8232 16820 8268
rect 15312 8152 15408 8168
rect 15312 8088 15328 8152
rect 15392 8088 15408 8152
rect 15312 8072 15408 8088
rect 15312 8008 15328 8072
rect 15392 8008 15408 8072
rect 15312 7992 15408 8008
rect 15312 7928 15328 7992
rect 15392 7928 15408 7992
rect 15312 7912 15408 7928
rect 15312 7848 15328 7912
rect 15392 7848 15408 7912
rect 15312 7832 15408 7848
rect 15312 7768 15328 7832
rect 15392 7768 15408 7832
rect 15312 7752 15408 7768
rect 15312 7688 15328 7752
rect 15392 7688 15408 7752
rect 15312 7672 15408 7688
rect 15312 7608 15328 7672
rect 15392 7608 15408 7672
rect 15312 7592 15408 7608
rect 15312 7528 15328 7592
rect 15392 7528 15408 7592
rect 15312 7512 15408 7528
rect 13900 7412 13996 7448
rect 15312 7448 15328 7512
rect 15392 7448 15408 7512
rect 15731 8192 16453 8201
rect 15731 7488 15740 8192
rect 16444 7488 16453 8192
rect 15731 7479 16453 7488
rect 16724 8168 16740 8232
rect 16804 8168 16820 8232
rect 18136 8232 18232 8268
rect 16724 8152 16820 8168
rect 16724 8088 16740 8152
rect 16804 8088 16820 8152
rect 16724 8072 16820 8088
rect 16724 8008 16740 8072
rect 16804 8008 16820 8072
rect 16724 7992 16820 8008
rect 16724 7928 16740 7992
rect 16804 7928 16820 7992
rect 16724 7912 16820 7928
rect 16724 7848 16740 7912
rect 16804 7848 16820 7912
rect 16724 7832 16820 7848
rect 16724 7768 16740 7832
rect 16804 7768 16820 7832
rect 16724 7752 16820 7768
rect 16724 7688 16740 7752
rect 16804 7688 16820 7752
rect 16724 7672 16820 7688
rect 16724 7608 16740 7672
rect 16804 7608 16820 7672
rect 16724 7592 16820 7608
rect 16724 7528 16740 7592
rect 16804 7528 16820 7592
rect 16724 7512 16820 7528
rect 15312 7412 15408 7448
rect 16724 7448 16740 7512
rect 16804 7448 16820 7512
rect 17143 8192 17865 8201
rect 17143 7488 17152 8192
rect 17856 7488 17865 8192
rect 17143 7479 17865 7488
rect 18136 8168 18152 8232
rect 18216 8168 18232 8232
rect 19548 8232 19644 8268
rect 18136 8152 18232 8168
rect 18136 8088 18152 8152
rect 18216 8088 18232 8152
rect 18136 8072 18232 8088
rect 18136 8008 18152 8072
rect 18216 8008 18232 8072
rect 18136 7992 18232 8008
rect 18136 7928 18152 7992
rect 18216 7928 18232 7992
rect 18136 7912 18232 7928
rect 18136 7848 18152 7912
rect 18216 7848 18232 7912
rect 18136 7832 18232 7848
rect 18136 7768 18152 7832
rect 18216 7768 18232 7832
rect 18136 7752 18232 7768
rect 18136 7688 18152 7752
rect 18216 7688 18232 7752
rect 18136 7672 18232 7688
rect 18136 7608 18152 7672
rect 18216 7608 18232 7672
rect 18136 7592 18232 7608
rect 18136 7528 18152 7592
rect 18216 7528 18232 7592
rect 18136 7512 18232 7528
rect 16724 7412 16820 7448
rect 18136 7448 18152 7512
rect 18216 7448 18232 7512
rect 18555 8192 19277 8201
rect 18555 7488 18564 8192
rect 19268 7488 19277 8192
rect 18555 7479 19277 7488
rect 19548 8168 19564 8232
rect 19628 8168 19644 8232
rect 20960 8232 21056 8268
rect 19548 8152 19644 8168
rect 19548 8088 19564 8152
rect 19628 8088 19644 8152
rect 19548 8072 19644 8088
rect 19548 8008 19564 8072
rect 19628 8008 19644 8072
rect 19548 7992 19644 8008
rect 19548 7928 19564 7992
rect 19628 7928 19644 7992
rect 19548 7912 19644 7928
rect 19548 7848 19564 7912
rect 19628 7848 19644 7912
rect 19548 7832 19644 7848
rect 19548 7768 19564 7832
rect 19628 7768 19644 7832
rect 19548 7752 19644 7768
rect 19548 7688 19564 7752
rect 19628 7688 19644 7752
rect 19548 7672 19644 7688
rect 19548 7608 19564 7672
rect 19628 7608 19644 7672
rect 19548 7592 19644 7608
rect 19548 7528 19564 7592
rect 19628 7528 19644 7592
rect 19548 7512 19644 7528
rect 18136 7412 18232 7448
rect 19548 7448 19564 7512
rect 19628 7448 19644 7512
rect 19967 8192 20689 8201
rect 19967 7488 19976 8192
rect 20680 7488 20689 8192
rect 19967 7479 20689 7488
rect 20960 8168 20976 8232
rect 21040 8168 21056 8232
rect 22372 8232 22468 8268
rect 20960 8152 21056 8168
rect 20960 8088 20976 8152
rect 21040 8088 21056 8152
rect 20960 8072 21056 8088
rect 20960 8008 20976 8072
rect 21040 8008 21056 8072
rect 20960 7992 21056 8008
rect 20960 7928 20976 7992
rect 21040 7928 21056 7992
rect 20960 7912 21056 7928
rect 20960 7848 20976 7912
rect 21040 7848 21056 7912
rect 20960 7832 21056 7848
rect 20960 7768 20976 7832
rect 21040 7768 21056 7832
rect 20960 7752 21056 7768
rect 20960 7688 20976 7752
rect 21040 7688 21056 7752
rect 20960 7672 21056 7688
rect 20960 7608 20976 7672
rect 21040 7608 21056 7672
rect 20960 7592 21056 7608
rect 20960 7528 20976 7592
rect 21040 7528 21056 7592
rect 20960 7512 21056 7528
rect 19548 7412 19644 7448
rect 20960 7448 20976 7512
rect 21040 7448 21056 7512
rect 21379 8192 22101 8201
rect 21379 7488 21388 8192
rect 22092 7488 22101 8192
rect 21379 7479 22101 7488
rect 22372 8168 22388 8232
rect 22452 8168 22468 8232
rect 23784 8232 23880 8268
rect 22372 8152 22468 8168
rect 22372 8088 22388 8152
rect 22452 8088 22468 8152
rect 22372 8072 22468 8088
rect 22372 8008 22388 8072
rect 22452 8008 22468 8072
rect 22372 7992 22468 8008
rect 22372 7928 22388 7992
rect 22452 7928 22468 7992
rect 22372 7912 22468 7928
rect 22372 7848 22388 7912
rect 22452 7848 22468 7912
rect 22372 7832 22468 7848
rect 22372 7768 22388 7832
rect 22452 7768 22468 7832
rect 22372 7752 22468 7768
rect 22372 7688 22388 7752
rect 22452 7688 22468 7752
rect 22372 7672 22468 7688
rect 22372 7608 22388 7672
rect 22452 7608 22468 7672
rect 22372 7592 22468 7608
rect 22372 7528 22388 7592
rect 22452 7528 22468 7592
rect 22372 7512 22468 7528
rect 20960 7412 21056 7448
rect 22372 7448 22388 7512
rect 22452 7448 22468 7512
rect 22791 8192 23513 8201
rect 22791 7488 22800 8192
rect 23504 7488 23513 8192
rect 22791 7479 23513 7488
rect 23784 8168 23800 8232
rect 23864 8168 23880 8232
rect 23784 8152 23880 8168
rect 23784 8088 23800 8152
rect 23864 8088 23880 8152
rect 23784 8072 23880 8088
rect 23784 8008 23800 8072
rect 23864 8008 23880 8072
rect 23784 7992 23880 8008
rect 23784 7928 23800 7992
rect 23864 7928 23880 7992
rect 23784 7912 23880 7928
rect 23784 7848 23800 7912
rect 23864 7848 23880 7912
rect 23784 7832 23880 7848
rect 23784 7768 23800 7832
rect 23864 7768 23880 7832
rect 23784 7752 23880 7768
rect 23784 7688 23800 7752
rect 23864 7688 23880 7752
rect 23784 7672 23880 7688
rect 23784 7608 23800 7672
rect 23864 7608 23880 7672
rect 23784 7592 23880 7608
rect 23784 7528 23800 7592
rect 23864 7528 23880 7592
rect 23784 7512 23880 7528
rect 22372 7412 22468 7448
rect 23784 7448 23800 7512
rect 23864 7448 23880 7512
rect 23784 7412 23880 7448
rect -22812 7112 -22716 7148
rect -23805 7072 -23083 7081
rect -23805 6368 -23796 7072
rect -23092 6368 -23083 7072
rect -23805 6359 -23083 6368
rect -22812 7048 -22796 7112
rect -22732 7048 -22716 7112
rect -21400 7112 -21304 7148
rect -22812 7032 -22716 7048
rect -22812 6968 -22796 7032
rect -22732 6968 -22716 7032
rect -22812 6952 -22716 6968
rect -22812 6888 -22796 6952
rect -22732 6888 -22716 6952
rect -22812 6872 -22716 6888
rect -22812 6808 -22796 6872
rect -22732 6808 -22716 6872
rect -22812 6792 -22716 6808
rect -22812 6728 -22796 6792
rect -22732 6728 -22716 6792
rect -22812 6712 -22716 6728
rect -22812 6648 -22796 6712
rect -22732 6648 -22716 6712
rect -22812 6632 -22716 6648
rect -22812 6568 -22796 6632
rect -22732 6568 -22716 6632
rect -22812 6552 -22716 6568
rect -22812 6488 -22796 6552
rect -22732 6488 -22716 6552
rect -22812 6472 -22716 6488
rect -22812 6408 -22796 6472
rect -22732 6408 -22716 6472
rect -22812 6392 -22716 6408
rect -22812 6328 -22796 6392
rect -22732 6328 -22716 6392
rect -22393 7072 -21671 7081
rect -22393 6368 -22384 7072
rect -21680 6368 -21671 7072
rect -22393 6359 -21671 6368
rect -21400 7048 -21384 7112
rect -21320 7048 -21304 7112
rect -19988 7112 -19892 7148
rect -21400 7032 -21304 7048
rect -21400 6968 -21384 7032
rect -21320 6968 -21304 7032
rect -21400 6952 -21304 6968
rect -21400 6888 -21384 6952
rect -21320 6888 -21304 6952
rect -21400 6872 -21304 6888
rect -21400 6808 -21384 6872
rect -21320 6808 -21304 6872
rect -21400 6792 -21304 6808
rect -21400 6728 -21384 6792
rect -21320 6728 -21304 6792
rect -21400 6712 -21304 6728
rect -21400 6648 -21384 6712
rect -21320 6648 -21304 6712
rect -21400 6632 -21304 6648
rect -21400 6568 -21384 6632
rect -21320 6568 -21304 6632
rect -21400 6552 -21304 6568
rect -21400 6488 -21384 6552
rect -21320 6488 -21304 6552
rect -21400 6472 -21304 6488
rect -21400 6408 -21384 6472
rect -21320 6408 -21304 6472
rect -21400 6392 -21304 6408
rect -22812 6292 -22716 6328
rect -21400 6328 -21384 6392
rect -21320 6328 -21304 6392
rect -20981 7072 -20259 7081
rect -20981 6368 -20972 7072
rect -20268 6368 -20259 7072
rect -20981 6359 -20259 6368
rect -19988 7048 -19972 7112
rect -19908 7048 -19892 7112
rect -18576 7112 -18480 7148
rect -19988 7032 -19892 7048
rect -19988 6968 -19972 7032
rect -19908 6968 -19892 7032
rect -19988 6952 -19892 6968
rect -19988 6888 -19972 6952
rect -19908 6888 -19892 6952
rect -19988 6872 -19892 6888
rect -19988 6808 -19972 6872
rect -19908 6808 -19892 6872
rect -19988 6792 -19892 6808
rect -19988 6728 -19972 6792
rect -19908 6728 -19892 6792
rect -19988 6712 -19892 6728
rect -19988 6648 -19972 6712
rect -19908 6648 -19892 6712
rect -19988 6632 -19892 6648
rect -19988 6568 -19972 6632
rect -19908 6568 -19892 6632
rect -19988 6552 -19892 6568
rect -19988 6488 -19972 6552
rect -19908 6488 -19892 6552
rect -19988 6472 -19892 6488
rect -19988 6408 -19972 6472
rect -19908 6408 -19892 6472
rect -19988 6392 -19892 6408
rect -21400 6292 -21304 6328
rect -19988 6328 -19972 6392
rect -19908 6328 -19892 6392
rect -19569 7072 -18847 7081
rect -19569 6368 -19560 7072
rect -18856 6368 -18847 7072
rect -19569 6359 -18847 6368
rect -18576 7048 -18560 7112
rect -18496 7048 -18480 7112
rect -17164 7112 -17068 7148
rect -18576 7032 -18480 7048
rect -18576 6968 -18560 7032
rect -18496 6968 -18480 7032
rect -18576 6952 -18480 6968
rect -18576 6888 -18560 6952
rect -18496 6888 -18480 6952
rect -18576 6872 -18480 6888
rect -18576 6808 -18560 6872
rect -18496 6808 -18480 6872
rect -18576 6792 -18480 6808
rect -18576 6728 -18560 6792
rect -18496 6728 -18480 6792
rect -18576 6712 -18480 6728
rect -18576 6648 -18560 6712
rect -18496 6648 -18480 6712
rect -18576 6632 -18480 6648
rect -18576 6568 -18560 6632
rect -18496 6568 -18480 6632
rect -18576 6552 -18480 6568
rect -18576 6488 -18560 6552
rect -18496 6488 -18480 6552
rect -18576 6472 -18480 6488
rect -18576 6408 -18560 6472
rect -18496 6408 -18480 6472
rect -18576 6392 -18480 6408
rect -19988 6292 -19892 6328
rect -18576 6328 -18560 6392
rect -18496 6328 -18480 6392
rect -18157 7072 -17435 7081
rect -18157 6368 -18148 7072
rect -17444 6368 -17435 7072
rect -18157 6359 -17435 6368
rect -17164 7048 -17148 7112
rect -17084 7048 -17068 7112
rect -15752 7112 -15656 7148
rect -17164 7032 -17068 7048
rect -17164 6968 -17148 7032
rect -17084 6968 -17068 7032
rect -17164 6952 -17068 6968
rect -17164 6888 -17148 6952
rect -17084 6888 -17068 6952
rect -17164 6872 -17068 6888
rect -17164 6808 -17148 6872
rect -17084 6808 -17068 6872
rect -17164 6792 -17068 6808
rect -17164 6728 -17148 6792
rect -17084 6728 -17068 6792
rect -17164 6712 -17068 6728
rect -17164 6648 -17148 6712
rect -17084 6648 -17068 6712
rect -17164 6632 -17068 6648
rect -17164 6568 -17148 6632
rect -17084 6568 -17068 6632
rect -17164 6552 -17068 6568
rect -17164 6488 -17148 6552
rect -17084 6488 -17068 6552
rect -17164 6472 -17068 6488
rect -17164 6408 -17148 6472
rect -17084 6408 -17068 6472
rect -17164 6392 -17068 6408
rect -18576 6292 -18480 6328
rect -17164 6328 -17148 6392
rect -17084 6328 -17068 6392
rect -16745 7072 -16023 7081
rect -16745 6368 -16736 7072
rect -16032 6368 -16023 7072
rect -16745 6359 -16023 6368
rect -15752 7048 -15736 7112
rect -15672 7048 -15656 7112
rect -14340 7112 -14244 7148
rect -15752 7032 -15656 7048
rect -15752 6968 -15736 7032
rect -15672 6968 -15656 7032
rect -15752 6952 -15656 6968
rect -15752 6888 -15736 6952
rect -15672 6888 -15656 6952
rect -15752 6872 -15656 6888
rect -15752 6808 -15736 6872
rect -15672 6808 -15656 6872
rect -15752 6792 -15656 6808
rect -15752 6728 -15736 6792
rect -15672 6728 -15656 6792
rect -15752 6712 -15656 6728
rect -15752 6648 -15736 6712
rect -15672 6648 -15656 6712
rect -15752 6632 -15656 6648
rect -15752 6568 -15736 6632
rect -15672 6568 -15656 6632
rect -15752 6552 -15656 6568
rect -15752 6488 -15736 6552
rect -15672 6488 -15656 6552
rect -15752 6472 -15656 6488
rect -15752 6408 -15736 6472
rect -15672 6408 -15656 6472
rect -15752 6392 -15656 6408
rect -17164 6292 -17068 6328
rect -15752 6328 -15736 6392
rect -15672 6328 -15656 6392
rect -15333 7072 -14611 7081
rect -15333 6368 -15324 7072
rect -14620 6368 -14611 7072
rect -15333 6359 -14611 6368
rect -14340 7048 -14324 7112
rect -14260 7048 -14244 7112
rect -12928 7112 -12832 7148
rect -14340 7032 -14244 7048
rect -14340 6968 -14324 7032
rect -14260 6968 -14244 7032
rect -14340 6952 -14244 6968
rect -14340 6888 -14324 6952
rect -14260 6888 -14244 6952
rect -14340 6872 -14244 6888
rect -14340 6808 -14324 6872
rect -14260 6808 -14244 6872
rect -14340 6792 -14244 6808
rect -14340 6728 -14324 6792
rect -14260 6728 -14244 6792
rect -14340 6712 -14244 6728
rect -14340 6648 -14324 6712
rect -14260 6648 -14244 6712
rect -14340 6632 -14244 6648
rect -14340 6568 -14324 6632
rect -14260 6568 -14244 6632
rect -14340 6552 -14244 6568
rect -14340 6488 -14324 6552
rect -14260 6488 -14244 6552
rect -14340 6472 -14244 6488
rect -14340 6408 -14324 6472
rect -14260 6408 -14244 6472
rect -14340 6392 -14244 6408
rect -15752 6292 -15656 6328
rect -14340 6328 -14324 6392
rect -14260 6328 -14244 6392
rect -13921 7072 -13199 7081
rect -13921 6368 -13912 7072
rect -13208 6368 -13199 7072
rect -13921 6359 -13199 6368
rect -12928 7048 -12912 7112
rect -12848 7048 -12832 7112
rect -11516 7112 -11420 7148
rect -12928 7032 -12832 7048
rect -12928 6968 -12912 7032
rect -12848 6968 -12832 7032
rect -12928 6952 -12832 6968
rect -12928 6888 -12912 6952
rect -12848 6888 -12832 6952
rect -12928 6872 -12832 6888
rect -12928 6808 -12912 6872
rect -12848 6808 -12832 6872
rect -12928 6792 -12832 6808
rect -12928 6728 -12912 6792
rect -12848 6728 -12832 6792
rect -12928 6712 -12832 6728
rect -12928 6648 -12912 6712
rect -12848 6648 -12832 6712
rect -12928 6632 -12832 6648
rect -12928 6568 -12912 6632
rect -12848 6568 -12832 6632
rect -12928 6552 -12832 6568
rect -12928 6488 -12912 6552
rect -12848 6488 -12832 6552
rect -12928 6472 -12832 6488
rect -12928 6408 -12912 6472
rect -12848 6408 -12832 6472
rect -12928 6392 -12832 6408
rect -14340 6292 -14244 6328
rect -12928 6328 -12912 6392
rect -12848 6328 -12832 6392
rect -12509 7072 -11787 7081
rect -12509 6368 -12500 7072
rect -11796 6368 -11787 7072
rect -12509 6359 -11787 6368
rect -11516 7048 -11500 7112
rect -11436 7048 -11420 7112
rect -10104 7112 -10008 7148
rect -11516 7032 -11420 7048
rect -11516 6968 -11500 7032
rect -11436 6968 -11420 7032
rect -11516 6952 -11420 6968
rect -11516 6888 -11500 6952
rect -11436 6888 -11420 6952
rect -11516 6872 -11420 6888
rect -11516 6808 -11500 6872
rect -11436 6808 -11420 6872
rect -11516 6792 -11420 6808
rect -11516 6728 -11500 6792
rect -11436 6728 -11420 6792
rect -11516 6712 -11420 6728
rect -11516 6648 -11500 6712
rect -11436 6648 -11420 6712
rect -11516 6632 -11420 6648
rect -11516 6568 -11500 6632
rect -11436 6568 -11420 6632
rect -11516 6552 -11420 6568
rect -11516 6488 -11500 6552
rect -11436 6488 -11420 6552
rect -11516 6472 -11420 6488
rect -11516 6408 -11500 6472
rect -11436 6408 -11420 6472
rect -11516 6392 -11420 6408
rect -12928 6292 -12832 6328
rect -11516 6328 -11500 6392
rect -11436 6328 -11420 6392
rect -11097 7072 -10375 7081
rect -11097 6368 -11088 7072
rect -10384 6368 -10375 7072
rect -11097 6359 -10375 6368
rect -10104 7048 -10088 7112
rect -10024 7048 -10008 7112
rect -8692 7112 -8596 7148
rect -10104 7032 -10008 7048
rect -10104 6968 -10088 7032
rect -10024 6968 -10008 7032
rect -10104 6952 -10008 6968
rect -10104 6888 -10088 6952
rect -10024 6888 -10008 6952
rect -10104 6872 -10008 6888
rect -10104 6808 -10088 6872
rect -10024 6808 -10008 6872
rect -10104 6792 -10008 6808
rect -10104 6728 -10088 6792
rect -10024 6728 -10008 6792
rect -10104 6712 -10008 6728
rect -10104 6648 -10088 6712
rect -10024 6648 -10008 6712
rect -10104 6632 -10008 6648
rect -10104 6568 -10088 6632
rect -10024 6568 -10008 6632
rect -10104 6552 -10008 6568
rect -10104 6488 -10088 6552
rect -10024 6488 -10008 6552
rect -10104 6472 -10008 6488
rect -10104 6408 -10088 6472
rect -10024 6408 -10008 6472
rect -10104 6392 -10008 6408
rect -11516 6292 -11420 6328
rect -10104 6328 -10088 6392
rect -10024 6328 -10008 6392
rect -9685 7072 -8963 7081
rect -9685 6368 -9676 7072
rect -8972 6368 -8963 7072
rect -9685 6359 -8963 6368
rect -8692 7048 -8676 7112
rect -8612 7048 -8596 7112
rect -7280 7112 -7184 7148
rect -8692 7032 -8596 7048
rect -8692 6968 -8676 7032
rect -8612 6968 -8596 7032
rect -8692 6952 -8596 6968
rect -8692 6888 -8676 6952
rect -8612 6888 -8596 6952
rect -8692 6872 -8596 6888
rect -8692 6808 -8676 6872
rect -8612 6808 -8596 6872
rect -8692 6792 -8596 6808
rect -8692 6728 -8676 6792
rect -8612 6728 -8596 6792
rect -8692 6712 -8596 6728
rect -8692 6648 -8676 6712
rect -8612 6648 -8596 6712
rect -8692 6632 -8596 6648
rect -8692 6568 -8676 6632
rect -8612 6568 -8596 6632
rect -8692 6552 -8596 6568
rect -8692 6488 -8676 6552
rect -8612 6488 -8596 6552
rect -8692 6472 -8596 6488
rect -8692 6408 -8676 6472
rect -8612 6408 -8596 6472
rect -8692 6392 -8596 6408
rect -10104 6292 -10008 6328
rect -8692 6328 -8676 6392
rect -8612 6328 -8596 6392
rect -8273 7072 -7551 7081
rect -8273 6368 -8264 7072
rect -7560 6368 -7551 7072
rect -8273 6359 -7551 6368
rect -7280 7048 -7264 7112
rect -7200 7048 -7184 7112
rect -5868 7112 -5772 7148
rect -7280 7032 -7184 7048
rect -7280 6968 -7264 7032
rect -7200 6968 -7184 7032
rect -7280 6952 -7184 6968
rect -7280 6888 -7264 6952
rect -7200 6888 -7184 6952
rect -7280 6872 -7184 6888
rect -7280 6808 -7264 6872
rect -7200 6808 -7184 6872
rect -7280 6792 -7184 6808
rect -7280 6728 -7264 6792
rect -7200 6728 -7184 6792
rect -7280 6712 -7184 6728
rect -7280 6648 -7264 6712
rect -7200 6648 -7184 6712
rect -7280 6632 -7184 6648
rect -7280 6568 -7264 6632
rect -7200 6568 -7184 6632
rect -7280 6552 -7184 6568
rect -7280 6488 -7264 6552
rect -7200 6488 -7184 6552
rect -7280 6472 -7184 6488
rect -7280 6408 -7264 6472
rect -7200 6408 -7184 6472
rect -7280 6392 -7184 6408
rect -8692 6292 -8596 6328
rect -7280 6328 -7264 6392
rect -7200 6328 -7184 6392
rect -6861 7072 -6139 7081
rect -6861 6368 -6852 7072
rect -6148 6368 -6139 7072
rect -6861 6359 -6139 6368
rect -5868 7048 -5852 7112
rect -5788 7048 -5772 7112
rect -4456 7112 -4360 7148
rect -5868 7032 -5772 7048
rect -5868 6968 -5852 7032
rect -5788 6968 -5772 7032
rect -5868 6952 -5772 6968
rect -5868 6888 -5852 6952
rect -5788 6888 -5772 6952
rect -5868 6872 -5772 6888
rect -5868 6808 -5852 6872
rect -5788 6808 -5772 6872
rect -5868 6792 -5772 6808
rect -5868 6728 -5852 6792
rect -5788 6728 -5772 6792
rect -5868 6712 -5772 6728
rect -5868 6648 -5852 6712
rect -5788 6648 -5772 6712
rect -5868 6632 -5772 6648
rect -5868 6568 -5852 6632
rect -5788 6568 -5772 6632
rect -5868 6552 -5772 6568
rect -5868 6488 -5852 6552
rect -5788 6488 -5772 6552
rect -5868 6472 -5772 6488
rect -5868 6408 -5852 6472
rect -5788 6408 -5772 6472
rect -5868 6392 -5772 6408
rect -7280 6292 -7184 6328
rect -5868 6328 -5852 6392
rect -5788 6328 -5772 6392
rect -5449 7072 -4727 7081
rect -5449 6368 -5440 7072
rect -4736 6368 -4727 7072
rect -5449 6359 -4727 6368
rect -4456 7048 -4440 7112
rect -4376 7048 -4360 7112
rect -3044 7112 -2948 7148
rect -4456 7032 -4360 7048
rect -4456 6968 -4440 7032
rect -4376 6968 -4360 7032
rect -4456 6952 -4360 6968
rect -4456 6888 -4440 6952
rect -4376 6888 -4360 6952
rect -4456 6872 -4360 6888
rect -4456 6808 -4440 6872
rect -4376 6808 -4360 6872
rect -4456 6792 -4360 6808
rect -4456 6728 -4440 6792
rect -4376 6728 -4360 6792
rect -4456 6712 -4360 6728
rect -4456 6648 -4440 6712
rect -4376 6648 -4360 6712
rect -4456 6632 -4360 6648
rect -4456 6568 -4440 6632
rect -4376 6568 -4360 6632
rect -4456 6552 -4360 6568
rect -4456 6488 -4440 6552
rect -4376 6488 -4360 6552
rect -4456 6472 -4360 6488
rect -4456 6408 -4440 6472
rect -4376 6408 -4360 6472
rect -4456 6392 -4360 6408
rect -5868 6292 -5772 6328
rect -4456 6328 -4440 6392
rect -4376 6328 -4360 6392
rect -4037 7072 -3315 7081
rect -4037 6368 -4028 7072
rect -3324 6368 -3315 7072
rect -4037 6359 -3315 6368
rect -3044 7048 -3028 7112
rect -2964 7048 -2948 7112
rect -1632 7112 -1536 7148
rect -3044 7032 -2948 7048
rect -3044 6968 -3028 7032
rect -2964 6968 -2948 7032
rect -3044 6952 -2948 6968
rect -3044 6888 -3028 6952
rect -2964 6888 -2948 6952
rect -3044 6872 -2948 6888
rect -3044 6808 -3028 6872
rect -2964 6808 -2948 6872
rect -3044 6792 -2948 6808
rect -3044 6728 -3028 6792
rect -2964 6728 -2948 6792
rect -3044 6712 -2948 6728
rect -3044 6648 -3028 6712
rect -2964 6648 -2948 6712
rect -3044 6632 -2948 6648
rect -3044 6568 -3028 6632
rect -2964 6568 -2948 6632
rect -3044 6552 -2948 6568
rect -3044 6488 -3028 6552
rect -2964 6488 -2948 6552
rect -3044 6472 -2948 6488
rect -3044 6408 -3028 6472
rect -2964 6408 -2948 6472
rect -3044 6392 -2948 6408
rect -4456 6292 -4360 6328
rect -3044 6328 -3028 6392
rect -2964 6328 -2948 6392
rect -2625 7072 -1903 7081
rect -2625 6368 -2616 7072
rect -1912 6368 -1903 7072
rect -2625 6359 -1903 6368
rect -1632 7048 -1616 7112
rect -1552 7048 -1536 7112
rect -220 7112 -124 7148
rect -1632 7032 -1536 7048
rect -1632 6968 -1616 7032
rect -1552 6968 -1536 7032
rect -1632 6952 -1536 6968
rect -1632 6888 -1616 6952
rect -1552 6888 -1536 6952
rect -1632 6872 -1536 6888
rect -1632 6808 -1616 6872
rect -1552 6808 -1536 6872
rect -1632 6792 -1536 6808
rect -1632 6728 -1616 6792
rect -1552 6728 -1536 6792
rect -1632 6712 -1536 6728
rect -1632 6648 -1616 6712
rect -1552 6648 -1536 6712
rect -1632 6632 -1536 6648
rect -1632 6568 -1616 6632
rect -1552 6568 -1536 6632
rect -1632 6552 -1536 6568
rect -1632 6488 -1616 6552
rect -1552 6488 -1536 6552
rect -1632 6472 -1536 6488
rect -1632 6408 -1616 6472
rect -1552 6408 -1536 6472
rect -1632 6392 -1536 6408
rect -3044 6292 -2948 6328
rect -1632 6328 -1616 6392
rect -1552 6328 -1536 6392
rect -1213 7072 -491 7081
rect -1213 6368 -1204 7072
rect -500 6368 -491 7072
rect -1213 6359 -491 6368
rect -220 7048 -204 7112
rect -140 7048 -124 7112
rect 1192 7112 1288 7148
rect -220 7032 -124 7048
rect -220 6968 -204 7032
rect -140 6968 -124 7032
rect -220 6952 -124 6968
rect -220 6888 -204 6952
rect -140 6888 -124 6952
rect -220 6872 -124 6888
rect -220 6808 -204 6872
rect -140 6808 -124 6872
rect -220 6792 -124 6808
rect -220 6728 -204 6792
rect -140 6728 -124 6792
rect -220 6712 -124 6728
rect -220 6648 -204 6712
rect -140 6648 -124 6712
rect -220 6632 -124 6648
rect -220 6568 -204 6632
rect -140 6568 -124 6632
rect -220 6552 -124 6568
rect -220 6488 -204 6552
rect -140 6488 -124 6552
rect -220 6472 -124 6488
rect -220 6408 -204 6472
rect -140 6408 -124 6472
rect -220 6392 -124 6408
rect -1632 6292 -1536 6328
rect -220 6328 -204 6392
rect -140 6328 -124 6392
rect 199 7072 921 7081
rect 199 6368 208 7072
rect 912 6368 921 7072
rect 199 6359 921 6368
rect 1192 7048 1208 7112
rect 1272 7048 1288 7112
rect 2604 7112 2700 7148
rect 1192 7032 1288 7048
rect 1192 6968 1208 7032
rect 1272 6968 1288 7032
rect 1192 6952 1288 6968
rect 1192 6888 1208 6952
rect 1272 6888 1288 6952
rect 1192 6872 1288 6888
rect 1192 6808 1208 6872
rect 1272 6808 1288 6872
rect 1192 6792 1288 6808
rect 1192 6728 1208 6792
rect 1272 6728 1288 6792
rect 1192 6712 1288 6728
rect 1192 6648 1208 6712
rect 1272 6648 1288 6712
rect 1192 6632 1288 6648
rect 1192 6568 1208 6632
rect 1272 6568 1288 6632
rect 1192 6552 1288 6568
rect 1192 6488 1208 6552
rect 1272 6488 1288 6552
rect 1192 6472 1288 6488
rect 1192 6408 1208 6472
rect 1272 6408 1288 6472
rect 1192 6392 1288 6408
rect -220 6292 -124 6328
rect 1192 6328 1208 6392
rect 1272 6328 1288 6392
rect 1611 7072 2333 7081
rect 1611 6368 1620 7072
rect 2324 6368 2333 7072
rect 1611 6359 2333 6368
rect 2604 7048 2620 7112
rect 2684 7048 2700 7112
rect 4016 7112 4112 7148
rect 2604 7032 2700 7048
rect 2604 6968 2620 7032
rect 2684 6968 2700 7032
rect 2604 6952 2700 6968
rect 2604 6888 2620 6952
rect 2684 6888 2700 6952
rect 2604 6872 2700 6888
rect 2604 6808 2620 6872
rect 2684 6808 2700 6872
rect 2604 6792 2700 6808
rect 2604 6728 2620 6792
rect 2684 6728 2700 6792
rect 2604 6712 2700 6728
rect 2604 6648 2620 6712
rect 2684 6648 2700 6712
rect 2604 6632 2700 6648
rect 2604 6568 2620 6632
rect 2684 6568 2700 6632
rect 2604 6552 2700 6568
rect 2604 6488 2620 6552
rect 2684 6488 2700 6552
rect 2604 6472 2700 6488
rect 2604 6408 2620 6472
rect 2684 6408 2700 6472
rect 2604 6392 2700 6408
rect 1192 6292 1288 6328
rect 2604 6328 2620 6392
rect 2684 6328 2700 6392
rect 3023 7072 3745 7081
rect 3023 6368 3032 7072
rect 3736 6368 3745 7072
rect 3023 6359 3745 6368
rect 4016 7048 4032 7112
rect 4096 7048 4112 7112
rect 5428 7112 5524 7148
rect 4016 7032 4112 7048
rect 4016 6968 4032 7032
rect 4096 6968 4112 7032
rect 4016 6952 4112 6968
rect 4016 6888 4032 6952
rect 4096 6888 4112 6952
rect 4016 6872 4112 6888
rect 4016 6808 4032 6872
rect 4096 6808 4112 6872
rect 4016 6792 4112 6808
rect 4016 6728 4032 6792
rect 4096 6728 4112 6792
rect 4016 6712 4112 6728
rect 4016 6648 4032 6712
rect 4096 6648 4112 6712
rect 4016 6632 4112 6648
rect 4016 6568 4032 6632
rect 4096 6568 4112 6632
rect 4016 6552 4112 6568
rect 4016 6488 4032 6552
rect 4096 6488 4112 6552
rect 4016 6472 4112 6488
rect 4016 6408 4032 6472
rect 4096 6408 4112 6472
rect 4016 6392 4112 6408
rect 2604 6292 2700 6328
rect 4016 6328 4032 6392
rect 4096 6328 4112 6392
rect 4435 7072 5157 7081
rect 4435 6368 4444 7072
rect 5148 6368 5157 7072
rect 4435 6359 5157 6368
rect 5428 7048 5444 7112
rect 5508 7048 5524 7112
rect 6840 7112 6936 7148
rect 5428 7032 5524 7048
rect 5428 6968 5444 7032
rect 5508 6968 5524 7032
rect 5428 6952 5524 6968
rect 5428 6888 5444 6952
rect 5508 6888 5524 6952
rect 5428 6872 5524 6888
rect 5428 6808 5444 6872
rect 5508 6808 5524 6872
rect 5428 6792 5524 6808
rect 5428 6728 5444 6792
rect 5508 6728 5524 6792
rect 5428 6712 5524 6728
rect 5428 6648 5444 6712
rect 5508 6648 5524 6712
rect 5428 6632 5524 6648
rect 5428 6568 5444 6632
rect 5508 6568 5524 6632
rect 5428 6552 5524 6568
rect 5428 6488 5444 6552
rect 5508 6488 5524 6552
rect 5428 6472 5524 6488
rect 5428 6408 5444 6472
rect 5508 6408 5524 6472
rect 5428 6392 5524 6408
rect 4016 6292 4112 6328
rect 5428 6328 5444 6392
rect 5508 6328 5524 6392
rect 5847 7072 6569 7081
rect 5847 6368 5856 7072
rect 6560 6368 6569 7072
rect 5847 6359 6569 6368
rect 6840 7048 6856 7112
rect 6920 7048 6936 7112
rect 8252 7112 8348 7148
rect 6840 7032 6936 7048
rect 6840 6968 6856 7032
rect 6920 6968 6936 7032
rect 6840 6952 6936 6968
rect 6840 6888 6856 6952
rect 6920 6888 6936 6952
rect 6840 6872 6936 6888
rect 6840 6808 6856 6872
rect 6920 6808 6936 6872
rect 6840 6792 6936 6808
rect 6840 6728 6856 6792
rect 6920 6728 6936 6792
rect 6840 6712 6936 6728
rect 6840 6648 6856 6712
rect 6920 6648 6936 6712
rect 6840 6632 6936 6648
rect 6840 6568 6856 6632
rect 6920 6568 6936 6632
rect 6840 6552 6936 6568
rect 6840 6488 6856 6552
rect 6920 6488 6936 6552
rect 6840 6472 6936 6488
rect 6840 6408 6856 6472
rect 6920 6408 6936 6472
rect 6840 6392 6936 6408
rect 5428 6292 5524 6328
rect 6840 6328 6856 6392
rect 6920 6328 6936 6392
rect 7259 7072 7981 7081
rect 7259 6368 7268 7072
rect 7972 6368 7981 7072
rect 7259 6359 7981 6368
rect 8252 7048 8268 7112
rect 8332 7048 8348 7112
rect 9664 7112 9760 7148
rect 8252 7032 8348 7048
rect 8252 6968 8268 7032
rect 8332 6968 8348 7032
rect 8252 6952 8348 6968
rect 8252 6888 8268 6952
rect 8332 6888 8348 6952
rect 8252 6872 8348 6888
rect 8252 6808 8268 6872
rect 8332 6808 8348 6872
rect 8252 6792 8348 6808
rect 8252 6728 8268 6792
rect 8332 6728 8348 6792
rect 8252 6712 8348 6728
rect 8252 6648 8268 6712
rect 8332 6648 8348 6712
rect 8252 6632 8348 6648
rect 8252 6568 8268 6632
rect 8332 6568 8348 6632
rect 8252 6552 8348 6568
rect 8252 6488 8268 6552
rect 8332 6488 8348 6552
rect 8252 6472 8348 6488
rect 8252 6408 8268 6472
rect 8332 6408 8348 6472
rect 8252 6392 8348 6408
rect 6840 6292 6936 6328
rect 8252 6328 8268 6392
rect 8332 6328 8348 6392
rect 8671 7072 9393 7081
rect 8671 6368 8680 7072
rect 9384 6368 9393 7072
rect 8671 6359 9393 6368
rect 9664 7048 9680 7112
rect 9744 7048 9760 7112
rect 11076 7112 11172 7148
rect 9664 7032 9760 7048
rect 9664 6968 9680 7032
rect 9744 6968 9760 7032
rect 9664 6952 9760 6968
rect 9664 6888 9680 6952
rect 9744 6888 9760 6952
rect 9664 6872 9760 6888
rect 9664 6808 9680 6872
rect 9744 6808 9760 6872
rect 9664 6792 9760 6808
rect 9664 6728 9680 6792
rect 9744 6728 9760 6792
rect 9664 6712 9760 6728
rect 9664 6648 9680 6712
rect 9744 6648 9760 6712
rect 9664 6632 9760 6648
rect 9664 6568 9680 6632
rect 9744 6568 9760 6632
rect 9664 6552 9760 6568
rect 9664 6488 9680 6552
rect 9744 6488 9760 6552
rect 9664 6472 9760 6488
rect 9664 6408 9680 6472
rect 9744 6408 9760 6472
rect 9664 6392 9760 6408
rect 8252 6292 8348 6328
rect 9664 6328 9680 6392
rect 9744 6328 9760 6392
rect 10083 7072 10805 7081
rect 10083 6368 10092 7072
rect 10796 6368 10805 7072
rect 10083 6359 10805 6368
rect 11076 7048 11092 7112
rect 11156 7048 11172 7112
rect 12488 7112 12584 7148
rect 11076 7032 11172 7048
rect 11076 6968 11092 7032
rect 11156 6968 11172 7032
rect 11076 6952 11172 6968
rect 11076 6888 11092 6952
rect 11156 6888 11172 6952
rect 11076 6872 11172 6888
rect 11076 6808 11092 6872
rect 11156 6808 11172 6872
rect 11076 6792 11172 6808
rect 11076 6728 11092 6792
rect 11156 6728 11172 6792
rect 11076 6712 11172 6728
rect 11076 6648 11092 6712
rect 11156 6648 11172 6712
rect 11076 6632 11172 6648
rect 11076 6568 11092 6632
rect 11156 6568 11172 6632
rect 11076 6552 11172 6568
rect 11076 6488 11092 6552
rect 11156 6488 11172 6552
rect 11076 6472 11172 6488
rect 11076 6408 11092 6472
rect 11156 6408 11172 6472
rect 11076 6392 11172 6408
rect 9664 6292 9760 6328
rect 11076 6328 11092 6392
rect 11156 6328 11172 6392
rect 11495 7072 12217 7081
rect 11495 6368 11504 7072
rect 12208 6368 12217 7072
rect 11495 6359 12217 6368
rect 12488 7048 12504 7112
rect 12568 7048 12584 7112
rect 13900 7112 13996 7148
rect 12488 7032 12584 7048
rect 12488 6968 12504 7032
rect 12568 6968 12584 7032
rect 12488 6952 12584 6968
rect 12488 6888 12504 6952
rect 12568 6888 12584 6952
rect 12488 6872 12584 6888
rect 12488 6808 12504 6872
rect 12568 6808 12584 6872
rect 12488 6792 12584 6808
rect 12488 6728 12504 6792
rect 12568 6728 12584 6792
rect 12488 6712 12584 6728
rect 12488 6648 12504 6712
rect 12568 6648 12584 6712
rect 12488 6632 12584 6648
rect 12488 6568 12504 6632
rect 12568 6568 12584 6632
rect 12488 6552 12584 6568
rect 12488 6488 12504 6552
rect 12568 6488 12584 6552
rect 12488 6472 12584 6488
rect 12488 6408 12504 6472
rect 12568 6408 12584 6472
rect 12488 6392 12584 6408
rect 11076 6292 11172 6328
rect 12488 6328 12504 6392
rect 12568 6328 12584 6392
rect 12907 7072 13629 7081
rect 12907 6368 12916 7072
rect 13620 6368 13629 7072
rect 12907 6359 13629 6368
rect 13900 7048 13916 7112
rect 13980 7048 13996 7112
rect 15312 7112 15408 7148
rect 13900 7032 13996 7048
rect 13900 6968 13916 7032
rect 13980 6968 13996 7032
rect 13900 6952 13996 6968
rect 13900 6888 13916 6952
rect 13980 6888 13996 6952
rect 13900 6872 13996 6888
rect 13900 6808 13916 6872
rect 13980 6808 13996 6872
rect 13900 6792 13996 6808
rect 13900 6728 13916 6792
rect 13980 6728 13996 6792
rect 13900 6712 13996 6728
rect 13900 6648 13916 6712
rect 13980 6648 13996 6712
rect 13900 6632 13996 6648
rect 13900 6568 13916 6632
rect 13980 6568 13996 6632
rect 13900 6552 13996 6568
rect 13900 6488 13916 6552
rect 13980 6488 13996 6552
rect 13900 6472 13996 6488
rect 13900 6408 13916 6472
rect 13980 6408 13996 6472
rect 13900 6392 13996 6408
rect 12488 6292 12584 6328
rect 13900 6328 13916 6392
rect 13980 6328 13996 6392
rect 14319 7072 15041 7081
rect 14319 6368 14328 7072
rect 15032 6368 15041 7072
rect 14319 6359 15041 6368
rect 15312 7048 15328 7112
rect 15392 7048 15408 7112
rect 16724 7112 16820 7148
rect 15312 7032 15408 7048
rect 15312 6968 15328 7032
rect 15392 6968 15408 7032
rect 15312 6952 15408 6968
rect 15312 6888 15328 6952
rect 15392 6888 15408 6952
rect 15312 6872 15408 6888
rect 15312 6808 15328 6872
rect 15392 6808 15408 6872
rect 15312 6792 15408 6808
rect 15312 6728 15328 6792
rect 15392 6728 15408 6792
rect 15312 6712 15408 6728
rect 15312 6648 15328 6712
rect 15392 6648 15408 6712
rect 15312 6632 15408 6648
rect 15312 6568 15328 6632
rect 15392 6568 15408 6632
rect 15312 6552 15408 6568
rect 15312 6488 15328 6552
rect 15392 6488 15408 6552
rect 15312 6472 15408 6488
rect 15312 6408 15328 6472
rect 15392 6408 15408 6472
rect 15312 6392 15408 6408
rect 13900 6292 13996 6328
rect 15312 6328 15328 6392
rect 15392 6328 15408 6392
rect 15731 7072 16453 7081
rect 15731 6368 15740 7072
rect 16444 6368 16453 7072
rect 15731 6359 16453 6368
rect 16724 7048 16740 7112
rect 16804 7048 16820 7112
rect 18136 7112 18232 7148
rect 16724 7032 16820 7048
rect 16724 6968 16740 7032
rect 16804 6968 16820 7032
rect 16724 6952 16820 6968
rect 16724 6888 16740 6952
rect 16804 6888 16820 6952
rect 16724 6872 16820 6888
rect 16724 6808 16740 6872
rect 16804 6808 16820 6872
rect 16724 6792 16820 6808
rect 16724 6728 16740 6792
rect 16804 6728 16820 6792
rect 16724 6712 16820 6728
rect 16724 6648 16740 6712
rect 16804 6648 16820 6712
rect 16724 6632 16820 6648
rect 16724 6568 16740 6632
rect 16804 6568 16820 6632
rect 16724 6552 16820 6568
rect 16724 6488 16740 6552
rect 16804 6488 16820 6552
rect 16724 6472 16820 6488
rect 16724 6408 16740 6472
rect 16804 6408 16820 6472
rect 16724 6392 16820 6408
rect 15312 6292 15408 6328
rect 16724 6328 16740 6392
rect 16804 6328 16820 6392
rect 17143 7072 17865 7081
rect 17143 6368 17152 7072
rect 17856 6368 17865 7072
rect 17143 6359 17865 6368
rect 18136 7048 18152 7112
rect 18216 7048 18232 7112
rect 19548 7112 19644 7148
rect 18136 7032 18232 7048
rect 18136 6968 18152 7032
rect 18216 6968 18232 7032
rect 18136 6952 18232 6968
rect 18136 6888 18152 6952
rect 18216 6888 18232 6952
rect 18136 6872 18232 6888
rect 18136 6808 18152 6872
rect 18216 6808 18232 6872
rect 18136 6792 18232 6808
rect 18136 6728 18152 6792
rect 18216 6728 18232 6792
rect 18136 6712 18232 6728
rect 18136 6648 18152 6712
rect 18216 6648 18232 6712
rect 18136 6632 18232 6648
rect 18136 6568 18152 6632
rect 18216 6568 18232 6632
rect 18136 6552 18232 6568
rect 18136 6488 18152 6552
rect 18216 6488 18232 6552
rect 18136 6472 18232 6488
rect 18136 6408 18152 6472
rect 18216 6408 18232 6472
rect 18136 6392 18232 6408
rect 16724 6292 16820 6328
rect 18136 6328 18152 6392
rect 18216 6328 18232 6392
rect 18555 7072 19277 7081
rect 18555 6368 18564 7072
rect 19268 6368 19277 7072
rect 18555 6359 19277 6368
rect 19548 7048 19564 7112
rect 19628 7048 19644 7112
rect 20960 7112 21056 7148
rect 19548 7032 19644 7048
rect 19548 6968 19564 7032
rect 19628 6968 19644 7032
rect 19548 6952 19644 6968
rect 19548 6888 19564 6952
rect 19628 6888 19644 6952
rect 19548 6872 19644 6888
rect 19548 6808 19564 6872
rect 19628 6808 19644 6872
rect 19548 6792 19644 6808
rect 19548 6728 19564 6792
rect 19628 6728 19644 6792
rect 19548 6712 19644 6728
rect 19548 6648 19564 6712
rect 19628 6648 19644 6712
rect 19548 6632 19644 6648
rect 19548 6568 19564 6632
rect 19628 6568 19644 6632
rect 19548 6552 19644 6568
rect 19548 6488 19564 6552
rect 19628 6488 19644 6552
rect 19548 6472 19644 6488
rect 19548 6408 19564 6472
rect 19628 6408 19644 6472
rect 19548 6392 19644 6408
rect 18136 6292 18232 6328
rect 19548 6328 19564 6392
rect 19628 6328 19644 6392
rect 19967 7072 20689 7081
rect 19967 6368 19976 7072
rect 20680 6368 20689 7072
rect 19967 6359 20689 6368
rect 20960 7048 20976 7112
rect 21040 7048 21056 7112
rect 22372 7112 22468 7148
rect 20960 7032 21056 7048
rect 20960 6968 20976 7032
rect 21040 6968 21056 7032
rect 20960 6952 21056 6968
rect 20960 6888 20976 6952
rect 21040 6888 21056 6952
rect 20960 6872 21056 6888
rect 20960 6808 20976 6872
rect 21040 6808 21056 6872
rect 20960 6792 21056 6808
rect 20960 6728 20976 6792
rect 21040 6728 21056 6792
rect 20960 6712 21056 6728
rect 20960 6648 20976 6712
rect 21040 6648 21056 6712
rect 20960 6632 21056 6648
rect 20960 6568 20976 6632
rect 21040 6568 21056 6632
rect 20960 6552 21056 6568
rect 20960 6488 20976 6552
rect 21040 6488 21056 6552
rect 20960 6472 21056 6488
rect 20960 6408 20976 6472
rect 21040 6408 21056 6472
rect 20960 6392 21056 6408
rect 19548 6292 19644 6328
rect 20960 6328 20976 6392
rect 21040 6328 21056 6392
rect 21379 7072 22101 7081
rect 21379 6368 21388 7072
rect 22092 6368 22101 7072
rect 21379 6359 22101 6368
rect 22372 7048 22388 7112
rect 22452 7048 22468 7112
rect 23784 7112 23880 7148
rect 22372 7032 22468 7048
rect 22372 6968 22388 7032
rect 22452 6968 22468 7032
rect 22372 6952 22468 6968
rect 22372 6888 22388 6952
rect 22452 6888 22468 6952
rect 22372 6872 22468 6888
rect 22372 6808 22388 6872
rect 22452 6808 22468 6872
rect 22372 6792 22468 6808
rect 22372 6728 22388 6792
rect 22452 6728 22468 6792
rect 22372 6712 22468 6728
rect 22372 6648 22388 6712
rect 22452 6648 22468 6712
rect 22372 6632 22468 6648
rect 22372 6568 22388 6632
rect 22452 6568 22468 6632
rect 22372 6552 22468 6568
rect 22372 6488 22388 6552
rect 22452 6488 22468 6552
rect 22372 6472 22468 6488
rect 22372 6408 22388 6472
rect 22452 6408 22468 6472
rect 22372 6392 22468 6408
rect 20960 6292 21056 6328
rect 22372 6328 22388 6392
rect 22452 6328 22468 6392
rect 22791 7072 23513 7081
rect 22791 6368 22800 7072
rect 23504 6368 23513 7072
rect 22791 6359 23513 6368
rect 23784 7048 23800 7112
rect 23864 7048 23880 7112
rect 23784 7032 23880 7048
rect 23784 6968 23800 7032
rect 23864 6968 23880 7032
rect 23784 6952 23880 6968
rect 23784 6888 23800 6952
rect 23864 6888 23880 6952
rect 23784 6872 23880 6888
rect 23784 6808 23800 6872
rect 23864 6808 23880 6872
rect 23784 6792 23880 6808
rect 23784 6728 23800 6792
rect 23864 6728 23880 6792
rect 23784 6712 23880 6728
rect 23784 6648 23800 6712
rect 23864 6648 23880 6712
rect 23784 6632 23880 6648
rect 23784 6568 23800 6632
rect 23864 6568 23880 6632
rect 23784 6552 23880 6568
rect 23784 6488 23800 6552
rect 23864 6488 23880 6552
rect 23784 6472 23880 6488
rect 23784 6408 23800 6472
rect 23864 6408 23880 6472
rect 23784 6392 23880 6408
rect 22372 6292 22468 6328
rect 23784 6328 23800 6392
rect 23864 6328 23880 6392
rect 23784 6292 23880 6328
rect -22812 5992 -22716 6028
rect -23805 5952 -23083 5961
rect -23805 5248 -23796 5952
rect -23092 5248 -23083 5952
rect -23805 5239 -23083 5248
rect -22812 5928 -22796 5992
rect -22732 5928 -22716 5992
rect -21400 5992 -21304 6028
rect -22812 5912 -22716 5928
rect -22812 5848 -22796 5912
rect -22732 5848 -22716 5912
rect -22812 5832 -22716 5848
rect -22812 5768 -22796 5832
rect -22732 5768 -22716 5832
rect -22812 5752 -22716 5768
rect -22812 5688 -22796 5752
rect -22732 5688 -22716 5752
rect -22812 5672 -22716 5688
rect -22812 5608 -22796 5672
rect -22732 5608 -22716 5672
rect -22812 5592 -22716 5608
rect -22812 5528 -22796 5592
rect -22732 5528 -22716 5592
rect -22812 5512 -22716 5528
rect -22812 5448 -22796 5512
rect -22732 5448 -22716 5512
rect -22812 5432 -22716 5448
rect -22812 5368 -22796 5432
rect -22732 5368 -22716 5432
rect -22812 5352 -22716 5368
rect -22812 5288 -22796 5352
rect -22732 5288 -22716 5352
rect -22812 5272 -22716 5288
rect -22812 5208 -22796 5272
rect -22732 5208 -22716 5272
rect -22393 5952 -21671 5961
rect -22393 5248 -22384 5952
rect -21680 5248 -21671 5952
rect -22393 5239 -21671 5248
rect -21400 5928 -21384 5992
rect -21320 5928 -21304 5992
rect -19988 5992 -19892 6028
rect -21400 5912 -21304 5928
rect -21400 5848 -21384 5912
rect -21320 5848 -21304 5912
rect -21400 5832 -21304 5848
rect -21400 5768 -21384 5832
rect -21320 5768 -21304 5832
rect -21400 5752 -21304 5768
rect -21400 5688 -21384 5752
rect -21320 5688 -21304 5752
rect -21400 5672 -21304 5688
rect -21400 5608 -21384 5672
rect -21320 5608 -21304 5672
rect -21400 5592 -21304 5608
rect -21400 5528 -21384 5592
rect -21320 5528 -21304 5592
rect -21400 5512 -21304 5528
rect -21400 5448 -21384 5512
rect -21320 5448 -21304 5512
rect -21400 5432 -21304 5448
rect -21400 5368 -21384 5432
rect -21320 5368 -21304 5432
rect -21400 5352 -21304 5368
rect -21400 5288 -21384 5352
rect -21320 5288 -21304 5352
rect -21400 5272 -21304 5288
rect -22812 5172 -22716 5208
rect -21400 5208 -21384 5272
rect -21320 5208 -21304 5272
rect -20981 5952 -20259 5961
rect -20981 5248 -20972 5952
rect -20268 5248 -20259 5952
rect -20981 5239 -20259 5248
rect -19988 5928 -19972 5992
rect -19908 5928 -19892 5992
rect -18576 5992 -18480 6028
rect -19988 5912 -19892 5928
rect -19988 5848 -19972 5912
rect -19908 5848 -19892 5912
rect -19988 5832 -19892 5848
rect -19988 5768 -19972 5832
rect -19908 5768 -19892 5832
rect -19988 5752 -19892 5768
rect -19988 5688 -19972 5752
rect -19908 5688 -19892 5752
rect -19988 5672 -19892 5688
rect -19988 5608 -19972 5672
rect -19908 5608 -19892 5672
rect -19988 5592 -19892 5608
rect -19988 5528 -19972 5592
rect -19908 5528 -19892 5592
rect -19988 5512 -19892 5528
rect -19988 5448 -19972 5512
rect -19908 5448 -19892 5512
rect -19988 5432 -19892 5448
rect -19988 5368 -19972 5432
rect -19908 5368 -19892 5432
rect -19988 5352 -19892 5368
rect -19988 5288 -19972 5352
rect -19908 5288 -19892 5352
rect -19988 5272 -19892 5288
rect -21400 5172 -21304 5208
rect -19988 5208 -19972 5272
rect -19908 5208 -19892 5272
rect -19569 5952 -18847 5961
rect -19569 5248 -19560 5952
rect -18856 5248 -18847 5952
rect -19569 5239 -18847 5248
rect -18576 5928 -18560 5992
rect -18496 5928 -18480 5992
rect -17164 5992 -17068 6028
rect -18576 5912 -18480 5928
rect -18576 5848 -18560 5912
rect -18496 5848 -18480 5912
rect -18576 5832 -18480 5848
rect -18576 5768 -18560 5832
rect -18496 5768 -18480 5832
rect -18576 5752 -18480 5768
rect -18576 5688 -18560 5752
rect -18496 5688 -18480 5752
rect -18576 5672 -18480 5688
rect -18576 5608 -18560 5672
rect -18496 5608 -18480 5672
rect -18576 5592 -18480 5608
rect -18576 5528 -18560 5592
rect -18496 5528 -18480 5592
rect -18576 5512 -18480 5528
rect -18576 5448 -18560 5512
rect -18496 5448 -18480 5512
rect -18576 5432 -18480 5448
rect -18576 5368 -18560 5432
rect -18496 5368 -18480 5432
rect -18576 5352 -18480 5368
rect -18576 5288 -18560 5352
rect -18496 5288 -18480 5352
rect -18576 5272 -18480 5288
rect -19988 5172 -19892 5208
rect -18576 5208 -18560 5272
rect -18496 5208 -18480 5272
rect -18157 5952 -17435 5961
rect -18157 5248 -18148 5952
rect -17444 5248 -17435 5952
rect -18157 5239 -17435 5248
rect -17164 5928 -17148 5992
rect -17084 5928 -17068 5992
rect -15752 5992 -15656 6028
rect -17164 5912 -17068 5928
rect -17164 5848 -17148 5912
rect -17084 5848 -17068 5912
rect -17164 5832 -17068 5848
rect -17164 5768 -17148 5832
rect -17084 5768 -17068 5832
rect -17164 5752 -17068 5768
rect -17164 5688 -17148 5752
rect -17084 5688 -17068 5752
rect -17164 5672 -17068 5688
rect -17164 5608 -17148 5672
rect -17084 5608 -17068 5672
rect -17164 5592 -17068 5608
rect -17164 5528 -17148 5592
rect -17084 5528 -17068 5592
rect -17164 5512 -17068 5528
rect -17164 5448 -17148 5512
rect -17084 5448 -17068 5512
rect -17164 5432 -17068 5448
rect -17164 5368 -17148 5432
rect -17084 5368 -17068 5432
rect -17164 5352 -17068 5368
rect -17164 5288 -17148 5352
rect -17084 5288 -17068 5352
rect -17164 5272 -17068 5288
rect -18576 5172 -18480 5208
rect -17164 5208 -17148 5272
rect -17084 5208 -17068 5272
rect -16745 5952 -16023 5961
rect -16745 5248 -16736 5952
rect -16032 5248 -16023 5952
rect -16745 5239 -16023 5248
rect -15752 5928 -15736 5992
rect -15672 5928 -15656 5992
rect -14340 5992 -14244 6028
rect -15752 5912 -15656 5928
rect -15752 5848 -15736 5912
rect -15672 5848 -15656 5912
rect -15752 5832 -15656 5848
rect -15752 5768 -15736 5832
rect -15672 5768 -15656 5832
rect -15752 5752 -15656 5768
rect -15752 5688 -15736 5752
rect -15672 5688 -15656 5752
rect -15752 5672 -15656 5688
rect -15752 5608 -15736 5672
rect -15672 5608 -15656 5672
rect -15752 5592 -15656 5608
rect -15752 5528 -15736 5592
rect -15672 5528 -15656 5592
rect -15752 5512 -15656 5528
rect -15752 5448 -15736 5512
rect -15672 5448 -15656 5512
rect -15752 5432 -15656 5448
rect -15752 5368 -15736 5432
rect -15672 5368 -15656 5432
rect -15752 5352 -15656 5368
rect -15752 5288 -15736 5352
rect -15672 5288 -15656 5352
rect -15752 5272 -15656 5288
rect -17164 5172 -17068 5208
rect -15752 5208 -15736 5272
rect -15672 5208 -15656 5272
rect -15333 5952 -14611 5961
rect -15333 5248 -15324 5952
rect -14620 5248 -14611 5952
rect -15333 5239 -14611 5248
rect -14340 5928 -14324 5992
rect -14260 5928 -14244 5992
rect -12928 5992 -12832 6028
rect -14340 5912 -14244 5928
rect -14340 5848 -14324 5912
rect -14260 5848 -14244 5912
rect -14340 5832 -14244 5848
rect -14340 5768 -14324 5832
rect -14260 5768 -14244 5832
rect -14340 5752 -14244 5768
rect -14340 5688 -14324 5752
rect -14260 5688 -14244 5752
rect -14340 5672 -14244 5688
rect -14340 5608 -14324 5672
rect -14260 5608 -14244 5672
rect -14340 5592 -14244 5608
rect -14340 5528 -14324 5592
rect -14260 5528 -14244 5592
rect -14340 5512 -14244 5528
rect -14340 5448 -14324 5512
rect -14260 5448 -14244 5512
rect -14340 5432 -14244 5448
rect -14340 5368 -14324 5432
rect -14260 5368 -14244 5432
rect -14340 5352 -14244 5368
rect -14340 5288 -14324 5352
rect -14260 5288 -14244 5352
rect -14340 5272 -14244 5288
rect -15752 5172 -15656 5208
rect -14340 5208 -14324 5272
rect -14260 5208 -14244 5272
rect -13921 5952 -13199 5961
rect -13921 5248 -13912 5952
rect -13208 5248 -13199 5952
rect -13921 5239 -13199 5248
rect -12928 5928 -12912 5992
rect -12848 5928 -12832 5992
rect -11516 5992 -11420 6028
rect -12928 5912 -12832 5928
rect -12928 5848 -12912 5912
rect -12848 5848 -12832 5912
rect -12928 5832 -12832 5848
rect -12928 5768 -12912 5832
rect -12848 5768 -12832 5832
rect -12928 5752 -12832 5768
rect -12928 5688 -12912 5752
rect -12848 5688 -12832 5752
rect -12928 5672 -12832 5688
rect -12928 5608 -12912 5672
rect -12848 5608 -12832 5672
rect -12928 5592 -12832 5608
rect -12928 5528 -12912 5592
rect -12848 5528 -12832 5592
rect -12928 5512 -12832 5528
rect -12928 5448 -12912 5512
rect -12848 5448 -12832 5512
rect -12928 5432 -12832 5448
rect -12928 5368 -12912 5432
rect -12848 5368 -12832 5432
rect -12928 5352 -12832 5368
rect -12928 5288 -12912 5352
rect -12848 5288 -12832 5352
rect -12928 5272 -12832 5288
rect -14340 5172 -14244 5208
rect -12928 5208 -12912 5272
rect -12848 5208 -12832 5272
rect -12509 5952 -11787 5961
rect -12509 5248 -12500 5952
rect -11796 5248 -11787 5952
rect -12509 5239 -11787 5248
rect -11516 5928 -11500 5992
rect -11436 5928 -11420 5992
rect -10104 5992 -10008 6028
rect -11516 5912 -11420 5928
rect -11516 5848 -11500 5912
rect -11436 5848 -11420 5912
rect -11516 5832 -11420 5848
rect -11516 5768 -11500 5832
rect -11436 5768 -11420 5832
rect -11516 5752 -11420 5768
rect -11516 5688 -11500 5752
rect -11436 5688 -11420 5752
rect -11516 5672 -11420 5688
rect -11516 5608 -11500 5672
rect -11436 5608 -11420 5672
rect -11516 5592 -11420 5608
rect -11516 5528 -11500 5592
rect -11436 5528 -11420 5592
rect -11516 5512 -11420 5528
rect -11516 5448 -11500 5512
rect -11436 5448 -11420 5512
rect -11516 5432 -11420 5448
rect -11516 5368 -11500 5432
rect -11436 5368 -11420 5432
rect -11516 5352 -11420 5368
rect -11516 5288 -11500 5352
rect -11436 5288 -11420 5352
rect -11516 5272 -11420 5288
rect -12928 5172 -12832 5208
rect -11516 5208 -11500 5272
rect -11436 5208 -11420 5272
rect -11097 5952 -10375 5961
rect -11097 5248 -11088 5952
rect -10384 5248 -10375 5952
rect -11097 5239 -10375 5248
rect -10104 5928 -10088 5992
rect -10024 5928 -10008 5992
rect -8692 5992 -8596 6028
rect -10104 5912 -10008 5928
rect -10104 5848 -10088 5912
rect -10024 5848 -10008 5912
rect -10104 5832 -10008 5848
rect -10104 5768 -10088 5832
rect -10024 5768 -10008 5832
rect -10104 5752 -10008 5768
rect -10104 5688 -10088 5752
rect -10024 5688 -10008 5752
rect -10104 5672 -10008 5688
rect -10104 5608 -10088 5672
rect -10024 5608 -10008 5672
rect -10104 5592 -10008 5608
rect -10104 5528 -10088 5592
rect -10024 5528 -10008 5592
rect -10104 5512 -10008 5528
rect -10104 5448 -10088 5512
rect -10024 5448 -10008 5512
rect -10104 5432 -10008 5448
rect -10104 5368 -10088 5432
rect -10024 5368 -10008 5432
rect -10104 5352 -10008 5368
rect -10104 5288 -10088 5352
rect -10024 5288 -10008 5352
rect -10104 5272 -10008 5288
rect -11516 5172 -11420 5208
rect -10104 5208 -10088 5272
rect -10024 5208 -10008 5272
rect -9685 5952 -8963 5961
rect -9685 5248 -9676 5952
rect -8972 5248 -8963 5952
rect -9685 5239 -8963 5248
rect -8692 5928 -8676 5992
rect -8612 5928 -8596 5992
rect -7280 5992 -7184 6028
rect -8692 5912 -8596 5928
rect -8692 5848 -8676 5912
rect -8612 5848 -8596 5912
rect -8692 5832 -8596 5848
rect -8692 5768 -8676 5832
rect -8612 5768 -8596 5832
rect -8692 5752 -8596 5768
rect -8692 5688 -8676 5752
rect -8612 5688 -8596 5752
rect -8692 5672 -8596 5688
rect -8692 5608 -8676 5672
rect -8612 5608 -8596 5672
rect -8692 5592 -8596 5608
rect -8692 5528 -8676 5592
rect -8612 5528 -8596 5592
rect -8692 5512 -8596 5528
rect -8692 5448 -8676 5512
rect -8612 5448 -8596 5512
rect -8692 5432 -8596 5448
rect -8692 5368 -8676 5432
rect -8612 5368 -8596 5432
rect -8692 5352 -8596 5368
rect -8692 5288 -8676 5352
rect -8612 5288 -8596 5352
rect -8692 5272 -8596 5288
rect -10104 5172 -10008 5208
rect -8692 5208 -8676 5272
rect -8612 5208 -8596 5272
rect -8273 5952 -7551 5961
rect -8273 5248 -8264 5952
rect -7560 5248 -7551 5952
rect -8273 5239 -7551 5248
rect -7280 5928 -7264 5992
rect -7200 5928 -7184 5992
rect -5868 5992 -5772 6028
rect -7280 5912 -7184 5928
rect -7280 5848 -7264 5912
rect -7200 5848 -7184 5912
rect -7280 5832 -7184 5848
rect -7280 5768 -7264 5832
rect -7200 5768 -7184 5832
rect -7280 5752 -7184 5768
rect -7280 5688 -7264 5752
rect -7200 5688 -7184 5752
rect -7280 5672 -7184 5688
rect -7280 5608 -7264 5672
rect -7200 5608 -7184 5672
rect -7280 5592 -7184 5608
rect -7280 5528 -7264 5592
rect -7200 5528 -7184 5592
rect -7280 5512 -7184 5528
rect -7280 5448 -7264 5512
rect -7200 5448 -7184 5512
rect -7280 5432 -7184 5448
rect -7280 5368 -7264 5432
rect -7200 5368 -7184 5432
rect -7280 5352 -7184 5368
rect -7280 5288 -7264 5352
rect -7200 5288 -7184 5352
rect -7280 5272 -7184 5288
rect -8692 5172 -8596 5208
rect -7280 5208 -7264 5272
rect -7200 5208 -7184 5272
rect -6861 5952 -6139 5961
rect -6861 5248 -6852 5952
rect -6148 5248 -6139 5952
rect -6861 5239 -6139 5248
rect -5868 5928 -5852 5992
rect -5788 5928 -5772 5992
rect -4456 5992 -4360 6028
rect -5868 5912 -5772 5928
rect -5868 5848 -5852 5912
rect -5788 5848 -5772 5912
rect -5868 5832 -5772 5848
rect -5868 5768 -5852 5832
rect -5788 5768 -5772 5832
rect -5868 5752 -5772 5768
rect -5868 5688 -5852 5752
rect -5788 5688 -5772 5752
rect -5868 5672 -5772 5688
rect -5868 5608 -5852 5672
rect -5788 5608 -5772 5672
rect -5868 5592 -5772 5608
rect -5868 5528 -5852 5592
rect -5788 5528 -5772 5592
rect -5868 5512 -5772 5528
rect -5868 5448 -5852 5512
rect -5788 5448 -5772 5512
rect -5868 5432 -5772 5448
rect -5868 5368 -5852 5432
rect -5788 5368 -5772 5432
rect -5868 5352 -5772 5368
rect -5868 5288 -5852 5352
rect -5788 5288 -5772 5352
rect -5868 5272 -5772 5288
rect -7280 5172 -7184 5208
rect -5868 5208 -5852 5272
rect -5788 5208 -5772 5272
rect -5449 5952 -4727 5961
rect -5449 5248 -5440 5952
rect -4736 5248 -4727 5952
rect -5449 5239 -4727 5248
rect -4456 5928 -4440 5992
rect -4376 5928 -4360 5992
rect -3044 5992 -2948 6028
rect -4456 5912 -4360 5928
rect -4456 5848 -4440 5912
rect -4376 5848 -4360 5912
rect -4456 5832 -4360 5848
rect -4456 5768 -4440 5832
rect -4376 5768 -4360 5832
rect -4456 5752 -4360 5768
rect -4456 5688 -4440 5752
rect -4376 5688 -4360 5752
rect -4456 5672 -4360 5688
rect -4456 5608 -4440 5672
rect -4376 5608 -4360 5672
rect -4456 5592 -4360 5608
rect -4456 5528 -4440 5592
rect -4376 5528 -4360 5592
rect -4456 5512 -4360 5528
rect -4456 5448 -4440 5512
rect -4376 5448 -4360 5512
rect -4456 5432 -4360 5448
rect -4456 5368 -4440 5432
rect -4376 5368 -4360 5432
rect -4456 5352 -4360 5368
rect -4456 5288 -4440 5352
rect -4376 5288 -4360 5352
rect -4456 5272 -4360 5288
rect -5868 5172 -5772 5208
rect -4456 5208 -4440 5272
rect -4376 5208 -4360 5272
rect -4037 5952 -3315 5961
rect -4037 5248 -4028 5952
rect -3324 5248 -3315 5952
rect -4037 5239 -3315 5248
rect -3044 5928 -3028 5992
rect -2964 5928 -2948 5992
rect -1632 5992 -1536 6028
rect -3044 5912 -2948 5928
rect -3044 5848 -3028 5912
rect -2964 5848 -2948 5912
rect -3044 5832 -2948 5848
rect -3044 5768 -3028 5832
rect -2964 5768 -2948 5832
rect -3044 5752 -2948 5768
rect -3044 5688 -3028 5752
rect -2964 5688 -2948 5752
rect -3044 5672 -2948 5688
rect -3044 5608 -3028 5672
rect -2964 5608 -2948 5672
rect -3044 5592 -2948 5608
rect -3044 5528 -3028 5592
rect -2964 5528 -2948 5592
rect -3044 5512 -2948 5528
rect -3044 5448 -3028 5512
rect -2964 5448 -2948 5512
rect -3044 5432 -2948 5448
rect -3044 5368 -3028 5432
rect -2964 5368 -2948 5432
rect -3044 5352 -2948 5368
rect -3044 5288 -3028 5352
rect -2964 5288 -2948 5352
rect -3044 5272 -2948 5288
rect -4456 5172 -4360 5208
rect -3044 5208 -3028 5272
rect -2964 5208 -2948 5272
rect -2625 5952 -1903 5961
rect -2625 5248 -2616 5952
rect -1912 5248 -1903 5952
rect -2625 5239 -1903 5248
rect -1632 5928 -1616 5992
rect -1552 5928 -1536 5992
rect -220 5992 -124 6028
rect -1632 5912 -1536 5928
rect -1632 5848 -1616 5912
rect -1552 5848 -1536 5912
rect -1632 5832 -1536 5848
rect -1632 5768 -1616 5832
rect -1552 5768 -1536 5832
rect -1632 5752 -1536 5768
rect -1632 5688 -1616 5752
rect -1552 5688 -1536 5752
rect -1632 5672 -1536 5688
rect -1632 5608 -1616 5672
rect -1552 5608 -1536 5672
rect -1632 5592 -1536 5608
rect -1632 5528 -1616 5592
rect -1552 5528 -1536 5592
rect -1632 5512 -1536 5528
rect -1632 5448 -1616 5512
rect -1552 5448 -1536 5512
rect -1632 5432 -1536 5448
rect -1632 5368 -1616 5432
rect -1552 5368 -1536 5432
rect -1632 5352 -1536 5368
rect -1632 5288 -1616 5352
rect -1552 5288 -1536 5352
rect -1632 5272 -1536 5288
rect -3044 5172 -2948 5208
rect -1632 5208 -1616 5272
rect -1552 5208 -1536 5272
rect -1213 5952 -491 5961
rect -1213 5248 -1204 5952
rect -500 5248 -491 5952
rect -1213 5239 -491 5248
rect -220 5928 -204 5992
rect -140 5928 -124 5992
rect 1192 5992 1288 6028
rect -220 5912 -124 5928
rect -220 5848 -204 5912
rect -140 5848 -124 5912
rect -220 5832 -124 5848
rect -220 5768 -204 5832
rect -140 5768 -124 5832
rect -220 5752 -124 5768
rect -220 5688 -204 5752
rect -140 5688 -124 5752
rect -220 5672 -124 5688
rect -220 5608 -204 5672
rect -140 5608 -124 5672
rect -220 5592 -124 5608
rect -220 5528 -204 5592
rect -140 5528 -124 5592
rect -220 5512 -124 5528
rect -220 5448 -204 5512
rect -140 5448 -124 5512
rect -220 5432 -124 5448
rect -220 5368 -204 5432
rect -140 5368 -124 5432
rect -220 5352 -124 5368
rect -220 5288 -204 5352
rect -140 5288 -124 5352
rect -220 5272 -124 5288
rect -1632 5172 -1536 5208
rect -220 5208 -204 5272
rect -140 5208 -124 5272
rect 199 5952 921 5961
rect 199 5248 208 5952
rect 912 5248 921 5952
rect 199 5239 921 5248
rect 1192 5928 1208 5992
rect 1272 5928 1288 5992
rect 2604 5992 2700 6028
rect 1192 5912 1288 5928
rect 1192 5848 1208 5912
rect 1272 5848 1288 5912
rect 1192 5832 1288 5848
rect 1192 5768 1208 5832
rect 1272 5768 1288 5832
rect 1192 5752 1288 5768
rect 1192 5688 1208 5752
rect 1272 5688 1288 5752
rect 1192 5672 1288 5688
rect 1192 5608 1208 5672
rect 1272 5608 1288 5672
rect 1192 5592 1288 5608
rect 1192 5528 1208 5592
rect 1272 5528 1288 5592
rect 1192 5512 1288 5528
rect 1192 5448 1208 5512
rect 1272 5448 1288 5512
rect 1192 5432 1288 5448
rect 1192 5368 1208 5432
rect 1272 5368 1288 5432
rect 1192 5352 1288 5368
rect 1192 5288 1208 5352
rect 1272 5288 1288 5352
rect 1192 5272 1288 5288
rect -220 5172 -124 5208
rect 1192 5208 1208 5272
rect 1272 5208 1288 5272
rect 1611 5952 2333 5961
rect 1611 5248 1620 5952
rect 2324 5248 2333 5952
rect 1611 5239 2333 5248
rect 2604 5928 2620 5992
rect 2684 5928 2700 5992
rect 4016 5992 4112 6028
rect 2604 5912 2700 5928
rect 2604 5848 2620 5912
rect 2684 5848 2700 5912
rect 2604 5832 2700 5848
rect 2604 5768 2620 5832
rect 2684 5768 2700 5832
rect 2604 5752 2700 5768
rect 2604 5688 2620 5752
rect 2684 5688 2700 5752
rect 2604 5672 2700 5688
rect 2604 5608 2620 5672
rect 2684 5608 2700 5672
rect 2604 5592 2700 5608
rect 2604 5528 2620 5592
rect 2684 5528 2700 5592
rect 2604 5512 2700 5528
rect 2604 5448 2620 5512
rect 2684 5448 2700 5512
rect 2604 5432 2700 5448
rect 2604 5368 2620 5432
rect 2684 5368 2700 5432
rect 2604 5352 2700 5368
rect 2604 5288 2620 5352
rect 2684 5288 2700 5352
rect 2604 5272 2700 5288
rect 1192 5172 1288 5208
rect 2604 5208 2620 5272
rect 2684 5208 2700 5272
rect 3023 5952 3745 5961
rect 3023 5248 3032 5952
rect 3736 5248 3745 5952
rect 3023 5239 3745 5248
rect 4016 5928 4032 5992
rect 4096 5928 4112 5992
rect 5428 5992 5524 6028
rect 4016 5912 4112 5928
rect 4016 5848 4032 5912
rect 4096 5848 4112 5912
rect 4016 5832 4112 5848
rect 4016 5768 4032 5832
rect 4096 5768 4112 5832
rect 4016 5752 4112 5768
rect 4016 5688 4032 5752
rect 4096 5688 4112 5752
rect 4016 5672 4112 5688
rect 4016 5608 4032 5672
rect 4096 5608 4112 5672
rect 4016 5592 4112 5608
rect 4016 5528 4032 5592
rect 4096 5528 4112 5592
rect 4016 5512 4112 5528
rect 4016 5448 4032 5512
rect 4096 5448 4112 5512
rect 4016 5432 4112 5448
rect 4016 5368 4032 5432
rect 4096 5368 4112 5432
rect 4016 5352 4112 5368
rect 4016 5288 4032 5352
rect 4096 5288 4112 5352
rect 4016 5272 4112 5288
rect 2604 5172 2700 5208
rect 4016 5208 4032 5272
rect 4096 5208 4112 5272
rect 4435 5952 5157 5961
rect 4435 5248 4444 5952
rect 5148 5248 5157 5952
rect 4435 5239 5157 5248
rect 5428 5928 5444 5992
rect 5508 5928 5524 5992
rect 6840 5992 6936 6028
rect 5428 5912 5524 5928
rect 5428 5848 5444 5912
rect 5508 5848 5524 5912
rect 5428 5832 5524 5848
rect 5428 5768 5444 5832
rect 5508 5768 5524 5832
rect 5428 5752 5524 5768
rect 5428 5688 5444 5752
rect 5508 5688 5524 5752
rect 5428 5672 5524 5688
rect 5428 5608 5444 5672
rect 5508 5608 5524 5672
rect 5428 5592 5524 5608
rect 5428 5528 5444 5592
rect 5508 5528 5524 5592
rect 5428 5512 5524 5528
rect 5428 5448 5444 5512
rect 5508 5448 5524 5512
rect 5428 5432 5524 5448
rect 5428 5368 5444 5432
rect 5508 5368 5524 5432
rect 5428 5352 5524 5368
rect 5428 5288 5444 5352
rect 5508 5288 5524 5352
rect 5428 5272 5524 5288
rect 4016 5172 4112 5208
rect 5428 5208 5444 5272
rect 5508 5208 5524 5272
rect 5847 5952 6569 5961
rect 5847 5248 5856 5952
rect 6560 5248 6569 5952
rect 5847 5239 6569 5248
rect 6840 5928 6856 5992
rect 6920 5928 6936 5992
rect 8252 5992 8348 6028
rect 6840 5912 6936 5928
rect 6840 5848 6856 5912
rect 6920 5848 6936 5912
rect 6840 5832 6936 5848
rect 6840 5768 6856 5832
rect 6920 5768 6936 5832
rect 6840 5752 6936 5768
rect 6840 5688 6856 5752
rect 6920 5688 6936 5752
rect 6840 5672 6936 5688
rect 6840 5608 6856 5672
rect 6920 5608 6936 5672
rect 6840 5592 6936 5608
rect 6840 5528 6856 5592
rect 6920 5528 6936 5592
rect 6840 5512 6936 5528
rect 6840 5448 6856 5512
rect 6920 5448 6936 5512
rect 6840 5432 6936 5448
rect 6840 5368 6856 5432
rect 6920 5368 6936 5432
rect 6840 5352 6936 5368
rect 6840 5288 6856 5352
rect 6920 5288 6936 5352
rect 6840 5272 6936 5288
rect 5428 5172 5524 5208
rect 6840 5208 6856 5272
rect 6920 5208 6936 5272
rect 7259 5952 7981 5961
rect 7259 5248 7268 5952
rect 7972 5248 7981 5952
rect 7259 5239 7981 5248
rect 8252 5928 8268 5992
rect 8332 5928 8348 5992
rect 9664 5992 9760 6028
rect 8252 5912 8348 5928
rect 8252 5848 8268 5912
rect 8332 5848 8348 5912
rect 8252 5832 8348 5848
rect 8252 5768 8268 5832
rect 8332 5768 8348 5832
rect 8252 5752 8348 5768
rect 8252 5688 8268 5752
rect 8332 5688 8348 5752
rect 8252 5672 8348 5688
rect 8252 5608 8268 5672
rect 8332 5608 8348 5672
rect 8252 5592 8348 5608
rect 8252 5528 8268 5592
rect 8332 5528 8348 5592
rect 8252 5512 8348 5528
rect 8252 5448 8268 5512
rect 8332 5448 8348 5512
rect 8252 5432 8348 5448
rect 8252 5368 8268 5432
rect 8332 5368 8348 5432
rect 8252 5352 8348 5368
rect 8252 5288 8268 5352
rect 8332 5288 8348 5352
rect 8252 5272 8348 5288
rect 6840 5172 6936 5208
rect 8252 5208 8268 5272
rect 8332 5208 8348 5272
rect 8671 5952 9393 5961
rect 8671 5248 8680 5952
rect 9384 5248 9393 5952
rect 8671 5239 9393 5248
rect 9664 5928 9680 5992
rect 9744 5928 9760 5992
rect 11076 5992 11172 6028
rect 9664 5912 9760 5928
rect 9664 5848 9680 5912
rect 9744 5848 9760 5912
rect 9664 5832 9760 5848
rect 9664 5768 9680 5832
rect 9744 5768 9760 5832
rect 9664 5752 9760 5768
rect 9664 5688 9680 5752
rect 9744 5688 9760 5752
rect 9664 5672 9760 5688
rect 9664 5608 9680 5672
rect 9744 5608 9760 5672
rect 9664 5592 9760 5608
rect 9664 5528 9680 5592
rect 9744 5528 9760 5592
rect 9664 5512 9760 5528
rect 9664 5448 9680 5512
rect 9744 5448 9760 5512
rect 9664 5432 9760 5448
rect 9664 5368 9680 5432
rect 9744 5368 9760 5432
rect 9664 5352 9760 5368
rect 9664 5288 9680 5352
rect 9744 5288 9760 5352
rect 9664 5272 9760 5288
rect 8252 5172 8348 5208
rect 9664 5208 9680 5272
rect 9744 5208 9760 5272
rect 10083 5952 10805 5961
rect 10083 5248 10092 5952
rect 10796 5248 10805 5952
rect 10083 5239 10805 5248
rect 11076 5928 11092 5992
rect 11156 5928 11172 5992
rect 12488 5992 12584 6028
rect 11076 5912 11172 5928
rect 11076 5848 11092 5912
rect 11156 5848 11172 5912
rect 11076 5832 11172 5848
rect 11076 5768 11092 5832
rect 11156 5768 11172 5832
rect 11076 5752 11172 5768
rect 11076 5688 11092 5752
rect 11156 5688 11172 5752
rect 11076 5672 11172 5688
rect 11076 5608 11092 5672
rect 11156 5608 11172 5672
rect 11076 5592 11172 5608
rect 11076 5528 11092 5592
rect 11156 5528 11172 5592
rect 11076 5512 11172 5528
rect 11076 5448 11092 5512
rect 11156 5448 11172 5512
rect 11076 5432 11172 5448
rect 11076 5368 11092 5432
rect 11156 5368 11172 5432
rect 11076 5352 11172 5368
rect 11076 5288 11092 5352
rect 11156 5288 11172 5352
rect 11076 5272 11172 5288
rect 9664 5172 9760 5208
rect 11076 5208 11092 5272
rect 11156 5208 11172 5272
rect 11495 5952 12217 5961
rect 11495 5248 11504 5952
rect 12208 5248 12217 5952
rect 11495 5239 12217 5248
rect 12488 5928 12504 5992
rect 12568 5928 12584 5992
rect 13900 5992 13996 6028
rect 12488 5912 12584 5928
rect 12488 5848 12504 5912
rect 12568 5848 12584 5912
rect 12488 5832 12584 5848
rect 12488 5768 12504 5832
rect 12568 5768 12584 5832
rect 12488 5752 12584 5768
rect 12488 5688 12504 5752
rect 12568 5688 12584 5752
rect 12488 5672 12584 5688
rect 12488 5608 12504 5672
rect 12568 5608 12584 5672
rect 12488 5592 12584 5608
rect 12488 5528 12504 5592
rect 12568 5528 12584 5592
rect 12488 5512 12584 5528
rect 12488 5448 12504 5512
rect 12568 5448 12584 5512
rect 12488 5432 12584 5448
rect 12488 5368 12504 5432
rect 12568 5368 12584 5432
rect 12488 5352 12584 5368
rect 12488 5288 12504 5352
rect 12568 5288 12584 5352
rect 12488 5272 12584 5288
rect 11076 5172 11172 5208
rect 12488 5208 12504 5272
rect 12568 5208 12584 5272
rect 12907 5952 13629 5961
rect 12907 5248 12916 5952
rect 13620 5248 13629 5952
rect 12907 5239 13629 5248
rect 13900 5928 13916 5992
rect 13980 5928 13996 5992
rect 15312 5992 15408 6028
rect 13900 5912 13996 5928
rect 13900 5848 13916 5912
rect 13980 5848 13996 5912
rect 13900 5832 13996 5848
rect 13900 5768 13916 5832
rect 13980 5768 13996 5832
rect 13900 5752 13996 5768
rect 13900 5688 13916 5752
rect 13980 5688 13996 5752
rect 13900 5672 13996 5688
rect 13900 5608 13916 5672
rect 13980 5608 13996 5672
rect 13900 5592 13996 5608
rect 13900 5528 13916 5592
rect 13980 5528 13996 5592
rect 13900 5512 13996 5528
rect 13900 5448 13916 5512
rect 13980 5448 13996 5512
rect 13900 5432 13996 5448
rect 13900 5368 13916 5432
rect 13980 5368 13996 5432
rect 13900 5352 13996 5368
rect 13900 5288 13916 5352
rect 13980 5288 13996 5352
rect 13900 5272 13996 5288
rect 12488 5172 12584 5208
rect 13900 5208 13916 5272
rect 13980 5208 13996 5272
rect 14319 5952 15041 5961
rect 14319 5248 14328 5952
rect 15032 5248 15041 5952
rect 14319 5239 15041 5248
rect 15312 5928 15328 5992
rect 15392 5928 15408 5992
rect 16724 5992 16820 6028
rect 15312 5912 15408 5928
rect 15312 5848 15328 5912
rect 15392 5848 15408 5912
rect 15312 5832 15408 5848
rect 15312 5768 15328 5832
rect 15392 5768 15408 5832
rect 15312 5752 15408 5768
rect 15312 5688 15328 5752
rect 15392 5688 15408 5752
rect 15312 5672 15408 5688
rect 15312 5608 15328 5672
rect 15392 5608 15408 5672
rect 15312 5592 15408 5608
rect 15312 5528 15328 5592
rect 15392 5528 15408 5592
rect 15312 5512 15408 5528
rect 15312 5448 15328 5512
rect 15392 5448 15408 5512
rect 15312 5432 15408 5448
rect 15312 5368 15328 5432
rect 15392 5368 15408 5432
rect 15312 5352 15408 5368
rect 15312 5288 15328 5352
rect 15392 5288 15408 5352
rect 15312 5272 15408 5288
rect 13900 5172 13996 5208
rect 15312 5208 15328 5272
rect 15392 5208 15408 5272
rect 15731 5952 16453 5961
rect 15731 5248 15740 5952
rect 16444 5248 16453 5952
rect 15731 5239 16453 5248
rect 16724 5928 16740 5992
rect 16804 5928 16820 5992
rect 18136 5992 18232 6028
rect 16724 5912 16820 5928
rect 16724 5848 16740 5912
rect 16804 5848 16820 5912
rect 16724 5832 16820 5848
rect 16724 5768 16740 5832
rect 16804 5768 16820 5832
rect 16724 5752 16820 5768
rect 16724 5688 16740 5752
rect 16804 5688 16820 5752
rect 16724 5672 16820 5688
rect 16724 5608 16740 5672
rect 16804 5608 16820 5672
rect 16724 5592 16820 5608
rect 16724 5528 16740 5592
rect 16804 5528 16820 5592
rect 16724 5512 16820 5528
rect 16724 5448 16740 5512
rect 16804 5448 16820 5512
rect 16724 5432 16820 5448
rect 16724 5368 16740 5432
rect 16804 5368 16820 5432
rect 16724 5352 16820 5368
rect 16724 5288 16740 5352
rect 16804 5288 16820 5352
rect 16724 5272 16820 5288
rect 15312 5172 15408 5208
rect 16724 5208 16740 5272
rect 16804 5208 16820 5272
rect 17143 5952 17865 5961
rect 17143 5248 17152 5952
rect 17856 5248 17865 5952
rect 17143 5239 17865 5248
rect 18136 5928 18152 5992
rect 18216 5928 18232 5992
rect 19548 5992 19644 6028
rect 18136 5912 18232 5928
rect 18136 5848 18152 5912
rect 18216 5848 18232 5912
rect 18136 5832 18232 5848
rect 18136 5768 18152 5832
rect 18216 5768 18232 5832
rect 18136 5752 18232 5768
rect 18136 5688 18152 5752
rect 18216 5688 18232 5752
rect 18136 5672 18232 5688
rect 18136 5608 18152 5672
rect 18216 5608 18232 5672
rect 18136 5592 18232 5608
rect 18136 5528 18152 5592
rect 18216 5528 18232 5592
rect 18136 5512 18232 5528
rect 18136 5448 18152 5512
rect 18216 5448 18232 5512
rect 18136 5432 18232 5448
rect 18136 5368 18152 5432
rect 18216 5368 18232 5432
rect 18136 5352 18232 5368
rect 18136 5288 18152 5352
rect 18216 5288 18232 5352
rect 18136 5272 18232 5288
rect 16724 5172 16820 5208
rect 18136 5208 18152 5272
rect 18216 5208 18232 5272
rect 18555 5952 19277 5961
rect 18555 5248 18564 5952
rect 19268 5248 19277 5952
rect 18555 5239 19277 5248
rect 19548 5928 19564 5992
rect 19628 5928 19644 5992
rect 20960 5992 21056 6028
rect 19548 5912 19644 5928
rect 19548 5848 19564 5912
rect 19628 5848 19644 5912
rect 19548 5832 19644 5848
rect 19548 5768 19564 5832
rect 19628 5768 19644 5832
rect 19548 5752 19644 5768
rect 19548 5688 19564 5752
rect 19628 5688 19644 5752
rect 19548 5672 19644 5688
rect 19548 5608 19564 5672
rect 19628 5608 19644 5672
rect 19548 5592 19644 5608
rect 19548 5528 19564 5592
rect 19628 5528 19644 5592
rect 19548 5512 19644 5528
rect 19548 5448 19564 5512
rect 19628 5448 19644 5512
rect 19548 5432 19644 5448
rect 19548 5368 19564 5432
rect 19628 5368 19644 5432
rect 19548 5352 19644 5368
rect 19548 5288 19564 5352
rect 19628 5288 19644 5352
rect 19548 5272 19644 5288
rect 18136 5172 18232 5208
rect 19548 5208 19564 5272
rect 19628 5208 19644 5272
rect 19967 5952 20689 5961
rect 19967 5248 19976 5952
rect 20680 5248 20689 5952
rect 19967 5239 20689 5248
rect 20960 5928 20976 5992
rect 21040 5928 21056 5992
rect 22372 5992 22468 6028
rect 20960 5912 21056 5928
rect 20960 5848 20976 5912
rect 21040 5848 21056 5912
rect 20960 5832 21056 5848
rect 20960 5768 20976 5832
rect 21040 5768 21056 5832
rect 20960 5752 21056 5768
rect 20960 5688 20976 5752
rect 21040 5688 21056 5752
rect 20960 5672 21056 5688
rect 20960 5608 20976 5672
rect 21040 5608 21056 5672
rect 20960 5592 21056 5608
rect 20960 5528 20976 5592
rect 21040 5528 21056 5592
rect 20960 5512 21056 5528
rect 20960 5448 20976 5512
rect 21040 5448 21056 5512
rect 20960 5432 21056 5448
rect 20960 5368 20976 5432
rect 21040 5368 21056 5432
rect 20960 5352 21056 5368
rect 20960 5288 20976 5352
rect 21040 5288 21056 5352
rect 20960 5272 21056 5288
rect 19548 5172 19644 5208
rect 20960 5208 20976 5272
rect 21040 5208 21056 5272
rect 21379 5952 22101 5961
rect 21379 5248 21388 5952
rect 22092 5248 22101 5952
rect 21379 5239 22101 5248
rect 22372 5928 22388 5992
rect 22452 5928 22468 5992
rect 23784 5992 23880 6028
rect 22372 5912 22468 5928
rect 22372 5848 22388 5912
rect 22452 5848 22468 5912
rect 22372 5832 22468 5848
rect 22372 5768 22388 5832
rect 22452 5768 22468 5832
rect 22372 5752 22468 5768
rect 22372 5688 22388 5752
rect 22452 5688 22468 5752
rect 22372 5672 22468 5688
rect 22372 5608 22388 5672
rect 22452 5608 22468 5672
rect 22372 5592 22468 5608
rect 22372 5528 22388 5592
rect 22452 5528 22468 5592
rect 22372 5512 22468 5528
rect 22372 5448 22388 5512
rect 22452 5448 22468 5512
rect 22372 5432 22468 5448
rect 22372 5368 22388 5432
rect 22452 5368 22468 5432
rect 22372 5352 22468 5368
rect 22372 5288 22388 5352
rect 22452 5288 22468 5352
rect 22372 5272 22468 5288
rect 20960 5172 21056 5208
rect 22372 5208 22388 5272
rect 22452 5208 22468 5272
rect 22791 5952 23513 5961
rect 22791 5248 22800 5952
rect 23504 5248 23513 5952
rect 22791 5239 23513 5248
rect 23784 5928 23800 5992
rect 23864 5928 23880 5992
rect 23784 5912 23880 5928
rect 23784 5848 23800 5912
rect 23864 5848 23880 5912
rect 23784 5832 23880 5848
rect 23784 5768 23800 5832
rect 23864 5768 23880 5832
rect 23784 5752 23880 5768
rect 23784 5688 23800 5752
rect 23864 5688 23880 5752
rect 23784 5672 23880 5688
rect 23784 5608 23800 5672
rect 23864 5608 23880 5672
rect 23784 5592 23880 5608
rect 23784 5528 23800 5592
rect 23864 5528 23880 5592
rect 23784 5512 23880 5528
rect 23784 5448 23800 5512
rect 23864 5448 23880 5512
rect 23784 5432 23880 5448
rect 23784 5368 23800 5432
rect 23864 5368 23880 5432
rect 23784 5352 23880 5368
rect 23784 5288 23800 5352
rect 23864 5288 23880 5352
rect 23784 5272 23880 5288
rect 22372 5172 22468 5208
rect 23784 5208 23800 5272
rect 23864 5208 23880 5272
rect 23784 5172 23880 5208
rect -22812 4872 -22716 4908
rect -23805 4832 -23083 4841
rect -23805 4128 -23796 4832
rect -23092 4128 -23083 4832
rect -23805 4119 -23083 4128
rect -22812 4808 -22796 4872
rect -22732 4808 -22716 4872
rect -21400 4872 -21304 4908
rect -22812 4792 -22716 4808
rect -22812 4728 -22796 4792
rect -22732 4728 -22716 4792
rect -22812 4712 -22716 4728
rect -22812 4648 -22796 4712
rect -22732 4648 -22716 4712
rect -22812 4632 -22716 4648
rect -22812 4568 -22796 4632
rect -22732 4568 -22716 4632
rect -22812 4552 -22716 4568
rect -22812 4488 -22796 4552
rect -22732 4488 -22716 4552
rect -22812 4472 -22716 4488
rect -22812 4408 -22796 4472
rect -22732 4408 -22716 4472
rect -22812 4392 -22716 4408
rect -22812 4328 -22796 4392
rect -22732 4328 -22716 4392
rect -22812 4312 -22716 4328
rect -22812 4248 -22796 4312
rect -22732 4248 -22716 4312
rect -22812 4232 -22716 4248
rect -22812 4168 -22796 4232
rect -22732 4168 -22716 4232
rect -22812 4152 -22716 4168
rect -22812 4088 -22796 4152
rect -22732 4088 -22716 4152
rect -22393 4832 -21671 4841
rect -22393 4128 -22384 4832
rect -21680 4128 -21671 4832
rect -22393 4119 -21671 4128
rect -21400 4808 -21384 4872
rect -21320 4808 -21304 4872
rect -19988 4872 -19892 4908
rect -21400 4792 -21304 4808
rect -21400 4728 -21384 4792
rect -21320 4728 -21304 4792
rect -21400 4712 -21304 4728
rect -21400 4648 -21384 4712
rect -21320 4648 -21304 4712
rect -21400 4632 -21304 4648
rect -21400 4568 -21384 4632
rect -21320 4568 -21304 4632
rect -21400 4552 -21304 4568
rect -21400 4488 -21384 4552
rect -21320 4488 -21304 4552
rect -21400 4472 -21304 4488
rect -21400 4408 -21384 4472
rect -21320 4408 -21304 4472
rect -21400 4392 -21304 4408
rect -21400 4328 -21384 4392
rect -21320 4328 -21304 4392
rect -21400 4312 -21304 4328
rect -21400 4248 -21384 4312
rect -21320 4248 -21304 4312
rect -21400 4232 -21304 4248
rect -21400 4168 -21384 4232
rect -21320 4168 -21304 4232
rect -21400 4152 -21304 4168
rect -22812 4052 -22716 4088
rect -21400 4088 -21384 4152
rect -21320 4088 -21304 4152
rect -20981 4832 -20259 4841
rect -20981 4128 -20972 4832
rect -20268 4128 -20259 4832
rect -20981 4119 -20259 4128
rect -19988 4808 -19972 4872
rect -19908 4808 -19892 4872
rect -18576 4872 -18480 4908
rect -19988 4792 -19892 4808
rect -19988 4728 -19972 4792
rect -19908 4728 -19892 4792
rect -19988 4712 -19892 4728
rect -19988 4648 -19972 4712
rect -19908 4648 -19892 4712
rect -19988 4632 -19892 4648
rect -19988 4568 -19972 4632
rect -19908 4568 -19892 4632
rect -19988 4552 -19892 4568
rect -19988 4488 -19972 4552
rect -19908 4488 -19892 4552
rect -19988 4472 -19892 4488
rect -19988 4408 -19972 4472
rect -19908 4408 -19892 4472
rect -19988 4392 -19892 4408
rect -19988 4328 -19972 4392
rect -19908 4328 -19892 4392
rect -19988 4312 -19892 4328
rect -19988 4248 -19972 4312
rect -19908 4248 -19892 4312
rect -19988 4232 -19892 4248
rect -19988 4168 -19972 4232
rect -19908 4168 -19892 4232
rect -19988 4152 -19892 4168
rect -21400 4052 -21304 4088
rect -19988 4088 -19972 4152
rect -19908 4088 -19892 4152
rect -19569 4832 -18847 4841
rect -19569 4128 -19560 4832
rect -18856 4128 -18847 4832
rect -19569 4119 -18847 4128
rect -18576 4808 -18560 4872
rect -18496 4808 -18480 4872
rect -17164 4872 -17068 4908
rect -18576 4792 -18480 4808
rect -18576 4728 -18560 4792
rect -18496 4728 -18480 4792
rect -18576 4712 -18480 4728
rect -18576 4648 -18560 4712
rect -18496 4648 -18480 4712
rect -18576 4632 -18480 4648
rect -18576 4568 -18560 4632
rect -18496 4568 -18480 4632
rect -18576 4552 -18480 4568
rect -18576 4488 -18560 4552
rect -18496 4488 -18480 4552
rect -18576 4472 -18480 4488
rect -18576 4408 -18560 4472
rect -18496 4408 -18480 4472
rect -18576 4392 -18480 4408
rect -18576 4328 -18560 4392
rect -18496 4328 -18480 4392
rect -18576 4312 -18480 4328
rect -18576 4248 -18560 4312
rect -18496 4248 -18480 4312
rect -18576 4232 -18480 4248
rect -18576 4168 -18560 4232
rect -18496 4168 -18480 4232
rect -18576 4152 -18480 4168
rect -19988 4052 -19892 4088
rect -18576 4088 -18560 4152
rect -18496 4088 -18480 4152
rect -18157 4832 -17435 4841
rect -18157 4128 -18148 4832
rect -17444 4128 -17435 4832
rect -18157 4119 -17435 4128
rect -17164 4808 -17148 4872
rect -17084 4808 -17068 4872
rect -15752 4872 -15656 4908
rect -17164 4792 -17068 4808
rect -17164 4728 -17148 4792
rect -17084 4728 -17068 4792
rect -17164 4712 -17068 4728
rect -17164 4648 -17148 4712
rect -17084 4648 -17068 4712
rect -17164 4632 -17068 4648
rect -17164 4568 -17148 4632
rect -17084 4568 -17068 4632
rect -17164 4552 -17068 4568
rect -17164 4488 -17148 4552
rect -17084 4488 -17068 4552
rect -17164 4472 -17068 4488
rect -17164 4408 -17148 4472
rect -17084 4408 -17068 4472
rect -17164 4392 -17068 4408
rect -17164 4328 -17148 4392
rect -17084 4328 -17068 4392
rect -17164 4312 -17068 4328
rect -17164 4248 -17148 4312
rect -17084 4248 -17068 4312
rect -17164 4232 -17068 4248
rect -17164 4168 -17148 4232
rect -17084 4168 -17068 4232
rect -17164 4152 -17068 4168
rect -18576 4052 -18480 4088
rect -17164 4088 -17148 4152
rect -17084 4088 -17068 4152
rect -16745 4832 -16023 4841
rect -16745 4128 -16736 4832
rect -16032 4128 -16023 4832
rect -16745 4119 -16023 4128
rect -15752 4808 -15736 4872
rect -15672 4808 -15656 4872
rect -14340 4872 -14244 4908
rect -15752 4792 -15656 4808
rect -15752 4728 -15736 4792
rect -15672 4728 -15656 4792
rect -15752 4712 -15656 4728
rect -15752 4648 -15736 4712
rect -15672 4648 -15656 4712
rect -15752 4632 -15656 4648
rect -15752 4568 -15736 4632
rect -15672 4568 -15656 4632
rect -15752 4552 -15656 4568
rect -15752 4488 -15736 4552
rect -15672 4488 -15656 4552
rect -15752 4472 -15656 4488
rect -15752 4408 -15736 4472
rect -15672 4408 -15656 4472
rect -15752 4392 -15656 4408
rect -15752 4328 -15736 4392
rect -15672 4328 -15656 4392
rect -15752 4312 -15656 4328
rect -15752 4248 -15736 4312
rect -15672 4248 -15656 4312
rect -15752 4232 -15656 4248
rect -15752 4168 -15736 4232
rect -15672 4168 -15656 4232
rect -15752 4152 -15656 4168
rect -17164 4052 -17068 4088
rect -15752 4088 -15736 4152
rect -15672 4088 -15656 4152
rect -15333 4832 -14611 4841
rect -15333 4128 -15324 4832
rect -14620 4128 -14611 4832
rect -15333 4119 -14611 4128
rect -14340 4808 -14324 4872
rect -14260 4808 -14244 4872
rect -12928 4872 -12832 4908
rect -14340 4792 -14244 4808
rect -14340 4728 -14324 4792
rect -14260 4728 -14244 4792
rect -14340 4712 -14244 4728
rect -14340 4648 -14324 4712
rect -14260 4648 -14244 4712
rect -14340 4632 -14244 4648
rect -14340 4568 -14324 4632
rect -14260 4568 -14244 4632
rect -14340 4552 -14244 4568
rect -14340 4488 -14324 4552
rect -14260 4488 -14244 4552
rect -14340 4472 -14244 4488
rect -14340 4408 -14324 4472
rect -14260 4408 -14244 4472
rect -14340 4392 -14244 4408
rect -14340 4328 -14324 4392
rect -14260 4328 -14244 4392
rect -14340 4312 -14244 4328
rect -14340 4248 -14324 4312
rect -14260 4248 -14244 4312
rect -14340 4232 -14244 4248
rect -14340 4168 -14324 4232
rect -14260 4168 -14244 4232
rect -14340 4152 -14244 4168
rect -15752 4052 -15656 4088
rect -14340 4088 -14324 4152
rect -14260 4088 -14244 4152
rect -13921 4832 -13199 4841
rect -13921 4128 -13912 4832
rect -13208 4128 -13199 4832
rect -13921 4119 -13199 4128
rect -12928 4808 -12912 4872
rect -12848 4808 -12832 4872
rect -11516 4872 -11420 4908
rect -12928 4792 -12832 4808
rect -12928 4728 -12912 4792
rect -12848 4728 -12832 4792
rect -12928 4712 -12832 4728
rect -12928 4648 -12912 4712
rect -12848 4648 -12832 4712
rect -12928 4632 -12832 4648
rect -12928 4568 -12912 4632
rect -12848 4568 -12832 4632
rect -12928 4552 -12832 4568
rect -12928 4488 -12912 4552
rect -12848 4488 -12832 4552
rect -12928 4472 -12832 4488
rect -12928 4408 -12912 4472
rect -12848 4408 -12832 4472
rect -12928 4392 -12832 4408
rect -12928 4328 -12912 4392
rect -12848 4328 -12832 4392
rect -12928 4312 -12832 4328
rect -12928 4248 -12912 4312
rect -12848 4248 -12832 4312
rect -12928 4232 -12832 4248
rect -12928 4168 -12912 4232
rect -12848 4168 -12832 4232
rect -12928 4152 -12832 4168
rect -14340 4052 -14244 4088
rect -12928 4088 -12912 4152
rect -12848 4088 -12832 4152
rect -12509 4832 -11787 4841
rect -12509 4128 -12500 4832
rect -11796 4128 -11787 4832
rect -12509 4119 -11787 4128
rect -11516 4808 -11500 4872
rect -11436 4808 -11420 4872
rect -10104 4872 -10008 4908
rect -11516 4792 -11420 4808
rect -11516 4728 -11500 4792
rect -11436 4728 -11420 4792
rect -11516 4712 -11420 4728
rect -11516 4648 -11500 4712
rect -11436 4648 -11420 4712
rect -11516 4632 -11420 4648
rect -11516 4568 -11500 4632
rect -11436 4568 -11420 4632
rect -11516 4552 -11420 4568
rect -11516 4488 -11500 4552
rect -11436 4488 -11420 4552
rect -11516 4472 -11420 4488
rect -11516 4408 -11500 4472
rect -11436 4408 -11420 4472
rect -11516 4392 -11420 4408
rect -11516 4328 -11500 4392
rect -11436 4328 -11420 4392
rect -11516 4312 -11420 4328
rect -11516 4248 -11500 4312
rect -11436 4248 -11420 4312
rect -11516 4232 -11420 4248
rect -11516 4168 -11500 4232
rect -11436 4168 -11420 4232
rect -11516 4152 -11420 4168
rect -12928 4052 -12832 4088
rect -11516 4088 -11500 4152
rect -11436 4088 -11420 4152
rect -11097 4832 -10375 4841
rect -11097 4128 -11088 4832
rect -10384 4128 -10375 4832
rect -11097 4119 -10375 4128
rect -10104 4808 -10088 4872
rect -10024 4808 -10008 4872
rect -8692 4872 -8596 4908
rect -10104 4792 -10008 4808
rect -10104 4728 -10088 4792
rect -10024 4728 -10008 4792
rect -10104 4712 -10008 4728
rect -10104 4648 -10088 4712
rect -10024 4648 -10008 4712
rect -10104 4632 -10008 4648
rect -10104 4568 -10088 4632
rect -10024 4568 -10008 4632
rect -10104 4552 -10008 4568
rect -10104 4488 -10088 4552
rect -10024 4488 -10008 4552
rect -10104 4472 -10008 4488
rect -10104 4408 -10088 4472
rect -10024 4408 -10008 4472
rect -10104 4392 -10008 4408
rect -10104 4328 -10088 4392
rect -10024 4328 -10008 4392
rect -10104 4312 -10008 4328
rect -10104 4248 -10088 4312
rect -10024 4248 -10008 4312
rect -10104 4232 -10008 4248
rect -10104 4168 -10088 4232
rect -10024 4168 -10008 4232
rect -10104 4152 -10008 4168
rect -11516 4052 -11420 4088
rect -10104 4088 -10088 4152
rect -10024 4088 -10008 4152
rect -9685 4832 -8963 4841
rect -9685 4128 -9676 4832
rect -8972 4128 -8963 4832
rect -9685 4119 -8963 4128
rect -8692 4808 -8676 4872
rect -8612 4808 -8596 4872
rect -7280 4872 -7184 4908
rect -8692 4792 -8596 4808
rect -8692 4728 -8676 4792
rect -8612 4728 -8596 4792
rect -8692 4712 -8596 4728
rect -8692 4648 -8676 4712
rect -8612 4648 -8596 4712
rect -8692 4632 -8596 4648
rect -8692 4568 -8676 4632
rect -8612 4568 -8596 4632
rect -8692 4552 -8596 4568
rect -8692 4488 -8676 4552
rect -8612 4488 -8596 4552
rect -8692 4472 -8596 4488
rect -8692 4408 -8676 4472
rect -8612 4408 -8596 4472
rect -8692 4392 -8596 4408
rect -8692 4328 -8676 4392
rect -8612 4328 -8596 4392
rect -8692 4312 -8596 4328
rect -8692 4248 -8676 4312
rect -8612 4248 -8596 4312
rect -8692 4232 -8596 4248
rect -8692 4168 -8676 4232
rect -8612 4168 -8596 4232
rect -8692 4152 -8596 4168
rect -10104 4052 -10008 4088
rect -8692 4088 -8676 4152
rect -8612 4088 -8596 4152
rect -8273 4832 -7551 4841
rect -8273 4128 -8264 4832
rect -7560 4128 -7551 4832
rect -8273 4119 -7551 4128
rect -7280 4808 -7264 4872
rect -7200 4808 -7184 4872
rect -5868 4872 -5772 4908
rect -7280 4792 -7184 4808
rect -7280 4728 -7264 4792
rect -7200 4728 -7184 4792
rect -7280 4712 -7184 4728
rect -7280 4648 -7264 4712
rect -7200 4648 -7184 4712
rect -7280 4632 -7184 4648
rect -7280 4568 -7264 4632
rect -7200 4568 -7184 4632
rect -7280 4552 -7184 4568
rect -7280 4488 -7264 4552
rect -7200 4488 -7184 4552
rect -7280 4472 -7184 4488
rect -7280 4408 -7264 4472
rect -7200 4408 -7184 4472
rect -7280 4392 -7184 4408
rect -7280 4328 -7264 4392
rect -7200 4328 -7184 4392
rect -7280 4312 -7184 4328
rect -7280 4248 -7264 4312
rect -7200 4248 -7184 4312
rect -7280 4232 -7184 4248
rect -7280 4168 -7264 4232
rect -7200 4168 -7184 4232
rect -7280 4152 -7184 4168
rect -8692 4052 -8596 4088
rect -7280 4088 -7264 4152
rect -7200 4088 -7184 4152
rect -6861 4832 -6139 4841
rect -6861 4128 -6852 4832
rect -6148 4128 -6139 4832
rect -6861 4119 -6139 4128
rect -5868 4808 -5852 4872
rect -5788 4808 -5772 4872
rect -4456 4872 -4360 4908
rect -5868 4792 -5772 4808
rect -5868 4728 -5852 4792
rect -5788 4728 -5772 4792
rect -5868 4712 -5772 4728
rect -5868 4648 -5852 4712
rect -5788 4648 -5772 4712
rect -5868 4632 -5772 4648
rect -5868 4568 -5852 4632
rect -5788 4568 -5772 4632
rect -5868 4552 -5772 4568
rect -5868 4488 -5852 4552
rect -5788 4488 -5772 4552
rect -5868 4472 -5772 4488
rect -5868 4408 -5852 4472
rect -5788 4408 -5772 4472
rect -5868 4392 -5772 4408
rect -5868 4328 -5852 4392
rect -5788 4328 -5772 4392
rect -5868 4312 -5772 4328
rect -5868 4248 -5852 4312
rect -5788 4248 -5772 4312
rect -5868 4232 -5772 4248
rect -5868 4168 -5852 4232
rect -5788 4168 -5772 4232
rect -5868 4152 -5772 4168
rect -7280 4052 -7184 4088
rect -5868 4088 -5852 4152
rect -5788 4088 -5772 4152
rect -5449 4832 -4727 4841
rect -5449 4128 -5440 4832
rect -4736 4128 -4727 4832
rect -5449 4119 -4727 4128
rect -4456 4808 -4440 4872
rect -4376 4808 -4360 4872
rect -3044 4872 -2948 4908
rect -4456 4792 -4360 4808
rect -4456 4728 -4440 4792
rect -4376 4728 -4360 4792
rect -4456 4712 -4360 4728
rect -4456 4648 -4440 4712
rect -4376 4648 -4360 4712
rect -4456 4632 -4360 4648
rect -4456 4568 -4440 4632
rect -4376 4568 -4360 4632
rect -4456 4552 -4360 4568
rect -4456 4488 -4440 4552
rect -4376 4488 -4360 4552
rect -4456 4472 -4360 4488
rect -4456 4408 -4440 4472
rect -4376 4408 -4360 4472
rect -4456 4392 -4360 4408
rect -4456 4328 -4440 4392
rect -4376 4328 -4360 4392
rect -4456 4312 -4360 4328
rect -4456 4248 -4440 4312
rect -4376 4248 -4360 4312
rect -4456 4232 -4360 4248
rect -4456 4168 -4440 4232
rect -4376 4168 -4360 4232
rect -4456 4152 -4360 4168
rect -5868 4052 -5772 4088
rect -4456 4088 -4440 4152
rect -4376 4088 -4360 4152
rect -4037 4832 -3315 4841
rect -4037 4128 -4028 4832
rect -3324 4128 -3315 4832
rect -4037 4119 -3315 4128
rect -3044 4808 -3028 4872
rect -2964 4808 -2948 4872
rect -1632 4872 -1536 4908
rect -3044 4792 -2948 4808
rect -3044 4728 -3028 4792
rect -2964 4728 -2948 4792
rect -3044 4712 -2948 4728
rect -3044 4648 -3028 4712
rect -2964 4648 -2948 4712
rect -3044 4632 -2948 4648
rect -3044 4568 -3028 4632
rect -2964 4568 -2948 4632
rect -3044 4552 -2948 4568
rect -3044 4488 -3028 4552
rect -2964 4488 -2948 4552
rect -3044 4472 -2948 4488
rect -3044 4408 -3028 4472
rect -2964 4408 -2948 4472
rect -3044 4392 -2948 4408
rect -3044 4328 -3028 4392
rect -2964 4328 -2948 4392
rect -3044 4312 -2948 4328
rect -3044 4248 -3028 4312
rect -2964 4248 -2948 4312
rect -3044 4232 -2948 4248
rect -3044 4168 -3028 4232
rect -2964 4168 -2948 4232
rect -3044 4152 -2948 4168
rect -4456 4052 -4360 4088
rect -3044 4088 -3028 4152
rect -2964 4088 -2948 4152
rect -2625 4832 -1903 4841
rect -2625 4128 -2616 4832
rect -1912 4128 -1903 4832
rect -2625 4119 -1903 4128
rect -1632 4808 -1616 4872
rect -1552 4808 -1536 4872
rect -220 4872 -124 4908
rect -1632 4792 -1536 4808
rect -1632 4728 -1616 4792
rect -1552 4728 -1536 4792
rect -1632 4712 -1536 4728
rect -1632 4648 -1616 4712
rect -1552 4648 -1536 4712
rect -1632 4632 -1536 4648
rect -1632 4568 -1616 4632
rect -1552 4568 -1536 4632
rect -1632 4552 -1536 4568
rect -1632 4488 -1616 4552
rect -1552 4488 -1536 4552
rect -1632 4472 -1536 4488
rect -1632 4408 -1616 4472
rect -1552 4408 -1536 4472
rect -1632 4392 -1536 4408
rect -1632 4328 -1616 4392
rect -1552 4328 -1536 4392
rect -1632 4312 -1536 4328
rect -1632 4248 -1616 4312
rect -1552 4248 -1536 4312
rect -1632 4232 -1536 4248
rect -1632 4168 -1616 4232
rect -1552 4168 -1536 4232
rect -1632 4152 -1536 4168
rect -3044 4052 -2948 4088
rect -1632 4088 -1616 4152
rect -1552 4088 -1536 4152
rect -1213 4832 -491 4841
rect -1213 4128 -1204 4832
rect -500 4128 -491 4832
rect -1213 4119 -491 4128
rect -220 4808 -204 4872
rect -140 4808 -124 4872
rect 1192 4872 1288 4908
rect -220 4792 -124 4808
rect -220 4728 -204 4792
rect -140 4728 -124 4792
rect -220 4712 -124 4728
rect -220 4648 -204 4712
rect -140 4648 -124 4712
rect -220 4632 -124 4648
rect -220 4568 -204 4632
rect -140 4568 -124 4632
rect -220 4552 -124 4568
rect -220 4488 -204 4552
rect -140 4488 -124 4552
rect -220 4472 -124 4488
rect -220 4408 -204 4472
rect -140 4408 -124 4472
rect -220 4392 -124 4408
rect -220 4328 -204 4392
rect -140 4328 -124 4392
rect -220 4312 -124 4328
rect -220 4248 -204 4312
rect -140 4248 -124 4312
rect -220 4232 -124 4248
rect -220 4168 -204 4232
rect -140 4168 -124 4232
rect -220 4152 -124 4168
rect -1632 4052 -1536 4088
rect -220 4088 -204 4152
rect -140 4088 -124 4152
rect 199 4832 921 4841
rect 199 4128 208 4832
rect 912 4128 921 4832
rect 199 4119 921 4128
rect 1192 4808 1208 4872
rect 1272 4808 1288 4872
rect 2604 4872 2700 4908
rect 1192 4792 1288 4808
rect 1192 4728 1208 4792
rect 1272 4728 1288 4792
rect 1192 4712 1288 4728
rect 1192 4648 1208 4712
rect 1272 4648 1288 4712
rect 1192 4632 1288 4648
rect 1192 4568 1208 4632
rect 1272 4568 1288 4632
rect 1192 4552 1288 4568
rect 1192 4488 1208 4552
rect 1272 4488 1288 4552
rect 1192 4472 1288 4488
rect 1192 4408 1208 4472
rect 1272 4408 1288 4472
rect 1192 4392 1288 4408
rect 1192 4328 1208 4392
rect 1272 4328 1288 4392
rect 1192 4312 1288 4328
rect 1192 4248 1208 4312
rect 1272 4248 1288 4312
rect 1192 4232 1288 4248
rect 1192 4168 1208 4232
rect 1272 4168 1288 4232
rect 1192 4152 1288 4168
rect -220 4052 -124 4088
rect 1192 4088 1208 4152
rect 1272 4088 1288 4152
rect 1611 4832 2333 4841
rect 1611 4128 1620 4832
rect 2324 4128 2333 4832
rect 1611 4119 2333 4128
rect 2604 4808 2620 4872
rect 2684 4808 2700 4872
rect 4016 4872 4112 4908
rect 2604 4792 2700 4808
rect 2604 4728 2620 4792
rect 2684 4728 2700 4792
rect 2604 4712 2700 4728
rect 2604 4648 2620 4712
rect 2684 4648 2700 4712
rect 2604 4632 2700 4648
rect 2604 4568 2620 4632
rect 2684 4568 2700 4632
rect 2604 4552 2700 4568
rect 2604 4488 2620 4552
rect 2684 4488 2700 4552
rect 2604 4472 2700 4488
rect 2604 4408 2620 4472
rect 2684 4408 2700 4472
rect 2604 4392 2700 4408
rect 2604 4328 2620 4392
rect 2684 4328 2700 4392
rect 2604 4312 2700 4328
rect 2604 4248 2620 4312
rect 2684 4248 2700 4312
rect 2604 4232 2700 4248
rect 2604 4168 2620 4232
rect 2684 4168 2700 4232
rect 2604 4152 2700 4168
rect 1192 4052 1288 4088
rect 2604 4088 2620 4152
rect 2684 4088 2700 4152
rect 3023 4832 3745 4841
rect 3023 4128 3032 4832
rect 3736 4128 3745 4832
rect 3023 4119 3745 4128
rect 4016 4808 4032 4872
rect 4096 4808 4112 4872
rect 5428 4872 5524 4908
rect 4016 4792 4112 4808
rect 4016 4728 4032 4792
rect 4096 4728 4112 4792
rect 4016 4712 4112 4728
rect 4016 4648 4032 4712
rect 4096 4648 4112 4712
rect 4016 4632 4112 4648
rect 4016 4568 4032 4632
rect 4096 4568 4112 4632
rect 4016 4552 4112 4568
rect 4016 4488 4032 4552
rect 4096 4488 4112 4552
rect 4016 4472 4112 4488
rect 4016 4408 4032 4472
rect 4096 4408 4112 4472
rect 4016 4392 4112 4408
rect 4016 4328 4032 4392
rect 4096 4328 4112 4392
rect 4016 4312 4112 4328
rect 4016 4248 4032 4312
rect 4096 4248 4112 4312
rect 4016 4232 4112 4248
rect 4016 4168 4032 4232
rect 4096 4168 4112 4232
rect 4016 4152 4112 4168
rect 2604 4052 2700 4088
rect 4016 4088 4032 4152
rect 4096 4088 4112 4152
rect 4435 4832 5157 4841
rect 4435 4128 4444 4832
rect 5148 4128 5157 4832
rect 4435 4119 5157 4128
rect 5428 4808 5444 4872
rect 5508 4808 5524 4872
rect 6840 4872 6936 4908
rect 5428 4792 5524 4808
rect 5428 4728 5444 4792
rect 5508 4728 5524 4792
rect 5428 4712 5524 4728
rect 5428 4648 5444 4712
rect 5508 4648 5524 4712
rect 5428 4632 5524 4648
rect 5428 4568 5444 4632
rect 5508 4568 5524 4632
rect 5428 4552 5524 4568
rect 5428 4488 5444 4552
rect 5508 4488 5524 4552
rect 5428 4472 5524 4488
rect 5428 4408 5444 4472
rect 5508 4408 5524 4472
rect 5428 4392 5524 4408
rect 5428 4328 5444 4392
rect 5508 4328 5524 4392
rect 5428 4312 5524 4328
rect 5428 4248 5444 4312
rect 5508 4248 5524 4312
rect 5428 4232 5524 4248
rect 5428 4168 5444 4232
rect 5508 4168 5524 4232
rect 5428 4152 5524 4168
rect 4016 4052 4112 4088
rect 5428 4088 5444 4152
rect 5508 4088 5524 4152
rect 5847 4832 6569 4841
rect 5847 4128 5856 4832
rect 6560 4128 6569 4832
rect 5847 4119 6569 4128
rect 6840 4808 6856 4872
rect 6920 4808 6936 4872
rect 8252 4872 8348 4908
rect 6840 4792 6936 4808
rect 6840 4728 6856 4792
rect 6920 4728 6936 4792
rect 6840 4712 6936 4728
rect 6840 4648 6856 4712
rect 6920 4648 6936 4712
rect 6840 4632 6936 4648
rect 6840 4568 6856 4632
rect 6920 4568 6936 4632
rect 6840 4552 6936 4568
rect 6840 4488 6856 4552
rect 6920 4488 6936 4552
rect 6840 4472 6936 4488
rect 6840 4408 6856 4472
rect 6920 4408 6936 4472
rect 6840 4392 6936 4408
rect 6840 4328 6856 4392
rect 6920 4328 6936 4392
rect 6840 4312 6936 4328
rect 6840 4248 6856 4312
rect 6920 4248 6936 4312
rect 6840 4232 6936 4248
rect 6840 4168 6856 4232
rect 6920 4168 6936 4232
rect 6840 4152 6936 4168
rect 5428 4052 5524 4088
rect 6840 4088 6856 4152
rect 6920 4088 6936 4152
rect 7259 4832 7981 4841
rect 7259 4128 7268 4832
rect 7972 4128 7981 4832
rect 7259 4119 7981 4128
rect 8252 4808 8268 4872
rect 8332 4808 8348 4872
rect 9664 4872 9760 4908
rect 8252 4792 8348 4808
rect 8252 4728 8268 4792
rect 8332 4728 8348 4792
rect 8252 4712 8348 4728
rect 8252 4648 8268 4712
rect 8332 4648 8348 4712
rect 8252 4632 8348 4648
rect 8252 4568 8268 4632
rect 8332 4568 8348 4632
rect 8252 4552 8348 4568
rect 8252 4488 8268 4552
rect 8332 4488 8348 4552
rect 8252 4472 8348 4488
rect 8252 4408 8268 4472
rect 8332 4408 8348 4472
rect 8252 4392 8348 4408
rect 8252 4328 8268 4392
rect 8332 4328 8348 4392
rect 8252 4312 8348 4328
rect 8252 4248 8268 4312
rect 8332 4248 8348 4312
rect 8252 4232 8348 4248
rect 8252 4168 8268 4232
rect 8332 4168 8348 4232
rect 8252 4152 8348 4168
rect 6840 4052 6936 4088
rect 8252 4088 8268 4152
rect 8332 4088 8348 4152
rect 8671 4832 9393 4841
rect 8671 4128 8680 4832
rect 9384 4128 9393 4832
rect 8671 4119 9393 4128
rect 9664 4808 9680 4872
rect 9744 4808 9760 4872
rect 11076 4872 11172 4908
rect 9664 4792 9760 4808
rect 9664 4728 9680 4792
rect 9744 4728 9760 4792
rect 9664 4712 9760 4728
rect 9664 4648 9680 4712
rect 9744 4648 9760 4712
rect 9664 4632 9760 4648
rect 9664 4568 9680 4632
rect 9744 4568 9760 4632
rect 9664 4552 9760 4568
rect 9664 4488 9680 4552
rect 9744 4488 9760 4552
rect 9664 4472 9760 4488
rect 9664 4408 9680 4472
rect 9744 4408 9760 4472
rect 9664 4392 9760 4408
rect 9664 4328 9680 4392
rect 9744 4328 9760 4392
rect 9664 4312 9760 4328
rect 9664 4248 9680 4312
rect 9744 4248 9760 4312
rect 9664 4232 9760 4248
rect 9664 4168 9680 4232
rect 9744 4168 9760 4232
rect 9664 4152 9760 4168
rect 8252 4052 8348 4088
rect 9664 4088 9680 4152
rect 9744 4088 9760 4152
rect 10083 4832 10805 4841
rect 10083 4128 10092 4832
rect 10796 4128 10805 4832
rect 10083 4119 10805 4128
rect 11076 4808 11092 4872
rect 11156 4808 11172 4872
rect 12488 4872 12584 4908
rect 11076 4792 11172 4808
rect 11076 4728 11092 4792
rect 11156 4728 11172 4792
rect 11076 4712 11172 4728
rect 11076 4648 11092 4712
rect 11156 4648 11172 4712
rect 11076 4632 11172 4648
rect 11076 4568 11092 4632
rect 11156 4568 11172 4632
rect 11076 4552 11172 4568
rect 11076 4488 11092 4552
rect 11156 4488 11172 4552
rect 11076 4472 11172 4488
rect 11076 4408 11092 4472
rect 11156 4408 11172 4472
rect 11076 4392 11172 4408
rect 11076 4328 11092 4392
rect 11156 4328 11172 4392
rect 11076 4312 11172 4328
rect 11076 4248 11092 4312
rect 11156 4248 11172 4312
rect 11076 4232 11172 4248
rect 11076 4168 11092 4232
rect 11156 4168 11172 4232
rect 11076 4152 11172 4168
rect 9664 4052 9760 4088
rect 11076 4088 11092 4152
rect 11156 4088 11172 4152
rect 11495 4832 12217 4841
rect 11495 4128 11504 4832
rect 12208 4128 12217 4832
rect 11495 4119 12217 4128
rect 12488 4808 12504 4872
rect 12568 4808 12584 4872
rect 13900 4872 13996 4908
rect 12488 4792 12584 4808
rect 12488 4728 12504 4792
rect 12568 4728 12584 4792
rect 12488 4712 12584 4728
rect 12488 4648 12504 4712
rect 12568 4648 12584 4712
rect 12488 4632 12584 4648
rect 12488 4568 12504 4632
rect 12568 4568 12584 4632
rect 12488 4552 12584 4568
rect 12488 4488 12504 4552
rect 12568 4488 12584 4552
rect 12488 4472 12584 4488
rect 12488 4408 12504 4472
rect 12568 4408 12584 4472
rect 12488 4392 12584 4408
rect 12488 4328 12504 4392
rect 12568 4328 12584 4392
rect 12488 4312 12584 4328
rect 12488 4248 12504 4312
rect 12568 4248 12584 4312
rect 12488 4232 12584 4248
rect 12488 4168 12504 4232
rect 12568 4168 12584 4232
rect 12488 4152 12584 4168
rect 11076 4052 11172 4088
rect 12488 4088 12504 4152
rect 12568 4088 12584 4152
rect 12907 4832 13629 4841
rect 12907 4128 12916 4832
rect 13620 4128 13629 4832
rect 12907 4119 13629 4128
rect 13900 4808 13916 4872
rect 13980 4808 13996 4872
rect 15312 4872 15408 4908
rect 13900 4792 13996 4808
rect 13900 4728 13916 4792
rect 13980 4728 13996 4792
rect 13900 4712 13996 4728
rect 13900 4648 13916 4712
rect 13980 4648 13996 4712
rect 13900 4632 13996 4648
rect 13900 4568 13916 4632
rect 13980 4568 13996 4632
rect 13900 4552 13996 4568
rect 13900 4488 13916 4552
rect 13980 4488 13996 4552
rect 13900 4472 13996 4488
rect 13900 4408 13916 4472
rect 13980 4408 13996 4472
rect 13900 4392 13996 4408
rect 13900 4328 13916 4392
rect 13980 4328 13996 4392
rect 13900 4312 13996 4328
rect 13900 4248 13916 4312
rect 13980 4248 13996 4312
rect 13900 4232 13996 4248
rect 13900 4168 13916 4232
rect 13980 4168 13996 4232
rect 13900 4152 13996 4168
rect 12488 4052 12584 4088
rect 13900 4088 13916 4152
rect 13980 4088 13996 4152
rect 14319 4832 15041 4841
rect 14319 4128 14328 4832
rect 15032 4128 15041 4832
rect 14319 4119 15041 4128
rect 15312 4808 15328 4872
rect 15392 4808 15408 4872
rect 16724 4872 16820 4908
rect 15312 4792 15408 4808
rect 15312 4728 15328 4792
rect 15392 4728 15408 4792
rect 15312 4712 15408 4728
rect 15312 4648 15328 4712
rect 15392 4648 15408 4712
rect 15312 4632 15408 4648
rect 15312 4568 15328 4632
rect 15392 4568 15408 4632
rect 15312 4552 15408 4568
rect 15312 4488 15328 4552
rect 15392 4488 15408 4552
rect 15312 4472 15408 4488
rect 15312 4408 15328 4472
rect 15392 4408 15408 4472
rect 15312 4392 15408 4408
rect 15312 4328 15328 4392
rect 15392 4328 15408 4392
rect 15312 4312 15408 4328
rect 15312 4248 15328 4312
rect 15392 4248 15408 4312
rect 15312 4232 15408 4248
rect 15312 4168 15328 4232
rect 15392 4168 15408 4232
rect 15312 4152 15408 4168
rect 13900 4052 13996 4088
rect 15312 4088 15328 4152
rect 15392 4088 15408 4152
rect 15731 4832 16453 4841
rect 15731 4128 15740 4832
rect 16444 4128 16453 4832
rect 15731 4119 16453 4128
rect 16724 4808 16740 4872
rect 16804 4808 16820 4872
rect 18136 4872 18232 4908
rect 16724 4792 16820 4808
rect 16724 4728 16740 4792
rect 16804 4728 16820 4792
rect 16724 4712 16820 4728
rect 16724 4648 16740 4712
rect 16804 4648 16820 4712
rect 16724 4632 16820 4648
rect 16724 4568 16740 4632
rect 16804 4568 16820 4632
rect 16724 4552 16820 4568
rect 16724 4488 16740 4552
rect 16804 4488 16820 4552
rect 16724 4472 16820 4488
rect 16724 4408 16740 4472
rect 16804 4408 16820 4472
rect 16724 4392 16820 4408
rect 16724 4328 16740 4392
rect 16804 4328 16820 4392
rect 16724 4312 16820 4328
rect 16724 4248 16740 4312
rect 16804 4248 16820 4312
rect 16724 4232 16820 4248
rect 16724 4168 16740 4232
rect 16804 4168 16820 4232
rect 16724 4152 16820 4168
rect 15312 4052 15408 4088
rect 16724 4088 16740 4152
rect 16804 4088 16820 4152
rect 17143 4832 17865 4841
rect 17143 4128 17152 4832
rect 17856 4128 17865 4832
rect 17143 4119 17865 4128
rect 18136 4808 18152 4872
rect 18216 4808 18232 4872
rect 19548 4872 19644 4908
rect 18136 4792 18232 4808
rect 18136 4728 18152 4792
rect 18216 4728 18232 4792
rect 18136 4712 18232 4728
rect 18136 4648 18152 4712
rect 18216 4648 18232 4712
rect 18136 4632 18232 4648
rect 18136 4568 18152 4632
rect 18216 4568 18232 4632
rect 18136 4552 18232 4568
rect 18136 4488 18152 4552
rect 18216 4488 18232 4552
rect 18136 4472 18232 4488
rect 18136 4408 18152 4472
rect 18216 4408 18232 4472
rect 18136 4392 18232 4408
rect 18136 4328 18152 4392
rect 18216 4328 18232 4392
rect 18136 4312 18232 4328
rect 18136 4248 18152 4312
rect 18216 4248 18232 4312
rect 18136 4232 18232 4248
rect 18136 4168 18152 4232
rect 18216 4168 18232 4232
rect 18136 4152 18232 4168
rect 16724 4052 16820 4088
rect 18136 4088 18152 4152
rect 18216 4088 18232 4152
rect 18555 4832 19277 4841
rect 18555 4128 18564 4832
rect 19268 4128 19277 4832
rect 18555 4119 19277 4128
rect 19548 4808 19564 4872
rect 19628 4808 19644 4872
rect 20960 4872 21056 4908
rect 19548 4792 19644 4808
rect 19548 4728 19564 4792
rect 19628 4728 19644 4792
rect 19548 4712 19644 4728
rect 19548 4648 19564 4712
rect 19628 4648 19644 4712
rect 19548 4632 19644 4648
rect 19548 4568 19564 4632
rect 19628 4568 19644 4632
rect 19548 4552 19644 4568
rect 19548 4488 19564 4552
rect 19628 4488 19644 4552
rect 19548 4472 19644 4488
rect 19548 4408 19564 4472
rect 19628 4408 19644 4472
rect 19548 4392 19644 4408
rect 19548 4328 19564 4392
rect 19628 4328 19644 4392
rect 19548 4312 19644 4328
rect 19548 4248 19564 4312
rect 19628 4248 19644 4312
rect 19548 4232 19644 4248
rect 19548 4168 19564 4232
rect 19628 4168 19644 4232
rect 19548 4152 19644 4168
rect 18136 4052 18232 4088
rect 19548 4088 19564 4152
rect 19628 4088 19644 4152
rect 19967 4832 20689 4841
rect 19967 4128 19976 4832
rect 20680 4128 20689 4832
rect 19967 4119 20689 4128
rect 20960 4808 20976 4872
rect 21040 4808 21056 4872
rect 22372 4872 22468 4908
rect 20960 4792 21056 4808
rect 20960 4728 20976 4792
rect 21040 4728 21056 4792
rect 20960 4712 21056 4728
rect 20960 4648 20976 4712
rect 21040 4648 21056 4712
rect 20960 4632 21056 4648
rect 20960 4568 20976 4632
rect 21040 4568 21056 4632
rect 20960 4552 21056 4568
rect 20960 4488 20976 4552
rect 21040 4488 21056 4552
rect 20960 4472 21056 4488
rect 20960 4408 20976 4472
rect 21040 4408 21056 4472
rect 20960 4392 21056 4408
rect 20960 4328 20976 4392
rect 21040 4328 21056 4392
rect 20960 4312 21056 4328
rect 20960 4248 20976 4312
rect 21040 4248 21056 4312
rect 20960 4232 21056 4248
rect 20960 4168 20976 4232
rect 21040 4168 21056 4232
rect 20960 4152 21056 4168
rect 19548 4052 19644 4088
rect 20960 4088 20976 4152
rect 21040 4088 21056 4152
rect 21379 4832 22101 4841
rect 21379 4128 21388 4832
rect 22092 4128 22101 4832
rect 21379 4119 22101 4128
rect 22372 4808 22388 4872
rect 22452 4808 22468 4872
rect 23784 4872 23880 4908
rect 22372 4792 22468 4808
rect 22372 4728 22388 4792
rect 22452 4728 22468 4792
rect 22372 4712 22468 4728
rect 22372 4648 22388 4712
rect 22452 4648 22468 4712
rect 22372 4632 22468 4648
rect 22372 4568 22388 4632
rect 22452 4568 22468 4632
rect 22372 4552 22468 4568
rect 22372 4488 22388 4552
rect 22452 4488 22468 4552
rect 22372 4472 22468 4488
rect 22372 4408 22388 4472
rect 22452 4408 22468 4472
rect 22372 4392 22468 4408
rect 22372 4328 22388 4392
rect 22452 4328 22468 4392
rect 22372 4312 22468 4328
rect 22372 4248 22388 4312
rect 22452 4248 22468 4312
rect 22372 4232 22468 4248
rect 22372 4168 22388 4232
rect 22452 4168 22468 4232
rect 22372 4152 22468 4168
rect 20960 4052 21056 4088
rect 22372 4088 22388 4152
rect 22452 4088 22468 4152
rect 22791 4832 23513 4841
rect 22791 4128 22800 4832
rect 23504 4128 23513 4832
rect 22791 4119 23513 4128
rect 23784 4808 23800 4872
rect 23864 4808 23880 4872
rect 23784 4792 23880 4808
rect 23784 4728 23800 4792
rect 23864 4728 23880 4792
rect 23784 4712 23880 4728
rect 23784 4648 23800 4712
rect 23864 4648 23880 4712
rect 23784 4632 23880 4648
rect 23784 4568 23800 4632
rect 23864 4568 23880 4632
rect 23784 4552 23880 4568
rect 23784 4488 23800 4552
rect 23864 4488 23880 4552
rect 23784 4472 23880 4488
rect 23784 4408 23800 4472
rect 23864 4408 23880 4472
rect 23784 4392 23880 4408
rect 23784 4328 23800 4392
rect 23864 4328 23880 4392
rect 23784 4312 23880 4328
rect 23784 4248 23800 4312
rect 23864 4248 23880 4312
rect 23784 4232 23880 4248
rect 23784 4168 23800 4232
rect 23864 4168 23880 4232
rect 23784 4152 23880 4168
rect 22372 4052 22468 4088
rect 23784 4088 23800 4152
rect 23864 4088 23880 4152
rect 23784 4052 23880 4088
rect -22812 3752 -22716 3788
rect -23805 3712 -23083 3721
rect -23805 3008 -23796 3712
rect -23092 3008 -23083 3712
rect -23805 2999 -23083 3008
rect -22812 3688 -22796 3752
rect -22732 3688 -22716 3752
rect -21400 3752 -21304 3788
rect -22812 3672 -22716 3688
rect -22812 3608 -22796 3672
rect -22732 3608 -22716 3672
rect -22812 3592 -22716 3608
rect -22812 3528 -22796 3592
rect -22732 3528 -22716 3592
rect -22812 3512 -22716 3528
rect -22812 3448 -22796 3512
rect -22732 3448 -22716 3512
rect -22812 3432 -22716 3448
rect -22812 3368 -22796 3432
rect -22732 3368 -22716 3432
rect -22812 3352 -22716 3368
rect -22812 3288 -22796 3352
rect -22732 3288 -22716 3352
rect -22812 3272 -22716 3288
rect -22812 3208 -22796 3272
rect -22732 3208 -22716 3272
rect -22812 3192 -22716 3208
rect -22812 3128 -22796 3192
rect -22732 3128 -22716 3192
rect -22812 3112 -22716 3128
rect -22812 3048 -22796 3112
rect -22732 3048 -22716 3112
rect -22812 3032 -22716 3048
rect -22812 2968 -22796 3032
rect -22732 2968 -22716 3032
rect -22393 3712 -21671 3721
rect -22393 3008 -22384 3712
rect -21680 3008 -21671 3712
rect -22393 2999 -21671 3008
rect -21400 3688 -21384 3752
rect -21320 3688 -21304 3752
rect -19988 3752 -19892 3788
rect -21400 3672 -21304 3688
rect -21400 3608 -21384 3672
rect -21320 3608 -21304 3672
rect -21400 3592 -21304 3608
rect -21400 3528 -21384 3592
rect -21320 3528 -21304 3592
rect -21400 3512 -21304 3528
rect -21400 3448 -21384 3512
rect -21320 3448 -21304 3512
rect -21400 3432 -21304 3448
rect -21400 3368 -21384 3432
rect -21320 3368 -21304 3432
rect -21400 3352 -21304 3368
rect -21400 3288 -21384 3352
rect -21320 3288 -21304 3352
rect -21400 3272 -21304 3288
rect -21400 3208 -21384 3272
rect -21320 3208 -21304 3272
rect -21400 3192 -21304 3208
rect -21400 3128 -21384 3192
rect -21320 3128 -21304 3192
rect -21400 3112 -21304 3128
rect -21400 3048 -21384 3112
rect -21320 3048 -21304 3112
rect -21400 3032 -21304 3048
rect -22812 2932 -22716 2968
rect -21400 2968 -21384 3032
rect -21320 2968 -21304 3032
rect -20981 3712 -20259 3721
rect -20981 3008 -20972 3712
rect -20268 3008 -20259 3712
rect -20981 2999 -20259 3008
rect -19988 3688 -19972 3752
rect -19908 3688 -19892 3752
rect -18576 3752 -18480 3788
rect -19988 3672 -19892 3688
rect -19988 3608 -19972 3672
rect -19908 3608 -19892 3672
rect -19988 3592 -19892 3608
rect -19988 3528 -19972 3592
rect -19908 3528 -19892 3592
rect -19988 3512 -19892 3528
rect -19988 3448 -19972 3512
rect -19908 3448 -19892 3512
rect -19988 3432 -19892 3448
rect -19988 3368 -19972 3432
rect -19908 3368 -19892 3432
rect -19988 3352 -19892 3368
rect -19988 3288 -19972 3352
rect -19908 3288 -19892 3352
rect -19988 3272 -19892 3288
rect -19988 3208 -19972 3272
rect -19908 3208 -19892 3272
rect -19988 3192 -19892 3208
rect -19988 3128 -19972 3192
rect -19908 3128 -19892 3192
rect -19988 3112 -19892 3128
rect -19988 3048 -19972 3112
rect -19908 3048 -19892 3112
rect -19988 3032 -19892 3048
rect -21400 2932 -21304 2968
rect -19988 2968 -19972 3032
rect -19908 2968 -19892 3032
rect -19569 3712 -18847 3721
rect -19569 3008 -19560 3712
rect -18856 3008 -18847 3712
rect -19569 2999 -18847 3008
rect -18576 3688 -18560 3752
rect -18496 3688 -18480 3752
rect -17164 3752 -17068 3788
rect -18576 3672 -18480 3688
rect -18576 3608 -18560 3672
rect -18496 3608 -18480 3672
rect -18576 3592 -18480 3608
rect -18576 3528 -18560 3592
rect -18496 3528 -18480 3592
rect -18576 3512 -18480 3528
rect -18576 3448 -18560 3512
rect -18496 3448 -18480 3512
rect -18576 3432 -18480 3448
rect -18576 3368 -18560 3432
rect -18496 3368 -18480 3432
rect -18576 3352 -18480 3368
rect -18576 3288 -18560 3352
rect -18496 3288 -18480 3352
rect -18576 3272 -18480 3288
rect -18576 3208 -18560 3272
rect -18496 3208 -18480 3272
rect -18576 3192 -18480 3208
rect -18576 3128 -18560 3192
rect -18496 3128 -18480 3192
rect -18576 3112 -18480 3128
rect -18576 3048 -18560 3112
rect -18496 3048 -18480 3112
rect -18576 3032 -18480 3048
rect -19988 2932 -19892 2968
rect -18576 2968 -18560 3032
rect -18496 2968 -18480 3032
rect -18157 3712 -17435 3721
rect -18157 3008 -18148 3712
rect -17444 3008 -17435 3712
rect -18157 2999 -17435 3008
rect -17164 3688 -17148 3752
rect -17084 3688 -17068 3752
rect -15752 3752 -15656 3788
rect -17164 3672 -17068 3688
rect -17164 3608 -17148 3672
rect -17084 3608 -17068 3672
rect -17164 3592 -17068 3608
rect -17164 3528 -17148 3592
rect -17084 3528 -17068 3592
rect -17164 3512 -17068 3528
rect -17164 3448 -17148 3512
rect -17084 3448 -17068 3512
rect -17164 3432 -17068 3448
rect -17164 3368 -17148 3432
rect -17084 3368 -17068 3432
rect -17164 3352 -17068 3368
rect -17164 3288 -17148 3352
rect -17084 3288 -17068 3352
rect -17164 3272 -17068 3288
rect -17164 3208 -17148 3272
rect -17084 3208 -17068 3272
rect -17164 3192 -17068 3208
rect -17164 3128 -17148 3192
rect -17084 3128 -17068 3192
rect -17164 3112 -17068 3128
rect -17164 3048 -17148 3112
rect -17084 3048 -17068 3112
rect -17164 3032 -17068 3048
rect -18576 2932 -18480 2968
rect -17164 2968 -17148 3032
rect -17084 2968 -17068 3032
rect -16745 3712 -16023 3721
rect -16745 3008 -16736 3712
rect -16032 3008 -16023 3712
rect -16745 2999 -16023 3008
rect -15752 3688 -15736 3752
rect -15672 3688 -15656 3752
rect -14340 3752 -14244 3788
rect -15752 3672 -15656 3688
rect -15752 3608 -15736 3672
rect -15672 3608 -15656 3672
rect -15752 3592 -15656 3608
rect -15752 3528 -15736 3592
rect -15672 3528 -15656 3592
rect -15752 3512 -15656 3528
rect -15752 3448 -15736 3512
rect -15672 3448 -15656 3512
rect -15752 3432 -15656 3448
rect -15752 3368 -15736 3432
rect -15672 3368 -15656 3432
rect -15752 3352 -15656 3368
rect -15752 3288 -15736 3352
rect -15672 3288 -15656 3352
rect -15752 3272 -15656 3288
rect -15752 3208 -15736 3272
rect -15672 3208 -15656 3272
rect -15752 3192 -15656 3208
rect -15752 3128 -15736 3192
rect -15672 3128 -15656 3192
rect -15752 3112 -15656 3128
rect -15752 3048 -15736 3112
rect -15672 3048 -15656 3112
rect -15752 3032 -15656 3048
rect -17164 2932 -17068 2968
rect -15752 2968 -15736 3032
rect -15672 2968 -15656 3032
rect -15333 3712 -14611 3721
rect -15333 3008 -15324 3712
rect -14620 3008 -14611 3712
rect -15333 2999 -14611 3008
rect -14340 3688 -14324 3752
rect -14260 3688 -14244 3752
rect -12928 3752 -12832 3788
rect -14340 3672 -14244 3688
rect -14340 3608 -14324 3672
rect -14260 3608 -14244 3672
rect -14340 3592 -14244 3608
rect -14340 3528 -14324 3592
rect -14260 3528 -14244 3592
rect -14340 3512 -14244 3528
rect -14340 3448 -14324 3512
rect -14260 3448 -14244 3512
rect -14340 3432 -14244 3448
rect -14340 3368 -14324 3432
rect -14260 3368 -14244 3432
rect -14340 3352 -14244 3368
rect -14340 3288 -14324 3352
rect -14260 3288 -14244 3352
rect -14340 3272 -14244 3288
rect -14340 3208 -14324 3272
rect -14260 3208 -14244 3272
rect -14340 3192 -14244 3208
rect -14340 3128 -14324 3192
rect -14260 3128 -14244 3192
rect -14340 3112 -14244 3128
rect -14340 3048 -14324 3112
rect -14260 3048 -14244 3112
rect -14340 3032 -14244 3048
rect -15752 2932 -15656 2968
rect -14340 2968 -14324 3032
rect -14260 2968 -14244 3032
rect -13921 3712 -13199 3721
rect -13921 3008 -13912 3712
rect -13208 3008 -13199 3712
rect -13921 2999 -13199 3008
rect -12928 3688 -12912 3752
rect -12848 3688 -12832 3752
rect -11516 3752 -11420 3788
rect -12928 3672 -12832 3688
rect -12928 3608 -12912 3672
rect -12848 3608 -12832 3672
rect -12928 3592 -12832 3608
rect -12928 3528 -12912 3592
rect -12848 3528 -12832 3592
rect -12928 3512 -12832 3528
rect -12928 3448 -12912 3512
rect -12848 3448 -12832 3512
rect -12928 3432 -12832 3448
rect -12928 3368 -12912 3432
rect -12848 3368 -12832 3432
rect -12928 3352 -12832 3368
rect -12928 3288 -12912 3352
rect -12848 3288 -12832 3352
rect -12928 3272 -12832 3288
rect -12928 3208 -12912 3272
rect -12848 3208 -12832 3272
rect -12928 3192 -12832 3208
rect -12928 3128 -12912 3192
rect -12848 3128 -12832 3192
rect -12928 3112 -12832 3128
rect -12928 3048 -12912 3112
rect -12848 3048 -12832 3112
rect -12928 3032 -12832 3048
rect -14340 2932 -14244 2968
rect -12928 2968 -12912 3032
rect -12848 2968 -12832 3032
rect -12509 3712 -11787 3721
rect -12509 3008 -12500 3712
rect -11796 3008 -11787 3712
rect -12509 2999 -11787 3008
rect -11516 3688 -11500 3752
rect -11436 3688 -11420 3752
rect -10104 3752 -10008 3788
rect -11516 3672 -11420 3688
rect -11516 3608 -11500 3672
rect -11436 3608 -11420 3672
rect -11516 3592 -11420 3608
rect -11516 3528 -11500 3592
rect -11436 3528 -11420 3592
rect -11516 3512 -11420 3528
rect -11516 3448 -11500 3512
rect -11436 3448 -11420 3512
rect -11516 3432 -11420 3448
rect -11516 3368 -11500 3432
rect -11436 3368 -11420 3432
rect -11516 3352 -11420 3368
rect -11516 3288 -11500 3352
rect -11436 3288 -11420 3352
rect -11516 3272 -11420 3288
rect -11516 3208 -11500 3272
rect -11436 3208 -11420 3272
rect -11516 3192 -11420 3208
rect -11516 3128 -11500 3192
rect -11436 3128 -11420 3192
rect -11516 3112 -11420 3128
rect -11516 3048 -11500 3112
rect -11436 3048 -11420 3112
rect -11516 3032 -11420 3048
rect -12928 2932 -12832 2968
rect -11516 2968 -11500 3032
rect -11436 2968 -11420 3032
rect -11097 3712 -10375 3721
rect -11097 3008 -11088 3712
rect -10384 3008 -10375 3712
rect -11097 2999 -10375 3008
rect -10104 3688 -10088 3752
rect -10024 3688 -10008 3752
rect -8692 3752 -8596 3788
rect -10104 3672 -10008 3688
rect -10104 3608 -10088 3672
rect -10024 3608 -10008 3672
rect -10104 3592 -10008 3608
rect -10104 3528 -10088 3592
rect -10024 3528 -10008 3592
rect -10104 3512 -10008 3528
rect -10104 3448 -10088 3512
rect -10024 3448 -10008 3512
rect -10104 3432 -10008 3448
rect -10104 3368 -10088 3432
rect -10024 3368 -10008 3432
rect -10104 3352 -10008 3368
rect -10104 3288 -10088 3352
rect -10024 3288 -10008 3352
rect -10104 3272 -10008 3288
rect -10104 3208 -10088 3272
rect -10024 3208 -10008 3272
rect -10104 3192 -10008 3208
rect -10104 3128 -10088 3192
rect -10024 3128 -10008 3192
rect -10104 3112 -10008 3128
rect -10104 3048 -10088 3112
rect -10024 3048 -10008 3112
rect -10104 3032 -10008 3048
rect -11516 2932 -11420 2968
rect -10104 2968 -10088 3032
rect -10024 2968 -10008 3032
rect -9685 3712 -8963 3721
rect -9685 3008 -9676 3712
rect -8972 3008 -8963 3712
rect -9685 2999 -8963 3008
rect -8692 3688 -8676 3752
rect -8612 3688 -8596 3752
rect -7280 3752 -7184 3788
rect -8692 3672 -8596 3688
rect -8692 3608 -8676 3672
rect -8612 3608 -8596 3672
rect -8692 3592 -8596 3608
rect -8692 3528 -8676 3592
rect -8612 3528 -8596 3592
rect -8692 3512 -8596 3528
rect -8692 3448 -8676 3512
rect -8612 3448 -8596 3512
rect -8692 3432 -8596 3448
rect -8692 3368 -8676 3432
rect -8612 3368 -8596 3432
rect -8692 3352 -8596 3368
rect -8692 3288 -8676 3352
rect -8612 3288 -8596 3352
rect -8692 3272 -8596 3288
rect -8692 3208 -8676 3272
rect -8612 3208 -8596 3272
rect -8692 3192 -8596 3208
rect -8692 3128 -8676 3192
rect -8612 3128 -8596 3192
rect -8692 3112 -8596 3128
rect -8692 3048 -8676 3112
rect -8612 3048 -8596 3112
rect -8692 3032 -8596 3048
rect -10104 2932 -10008 2968
rect -8692 2968 -8676 3032
rect -8612 2968 -8596 3032
rect -8273 3712 -7551 3721
rect -8273 3008 -8264 3712
rect -7560 3008 -7551 3712
rect -8273 2999 -7551 3008
rect -7280 3688 -7264 3752
rect -7200 3688 -7184 3752
rect -5868 3752 -5772 3788
rect -7280 3672 -7184 3688
rect -7280 3608 -7264 3672
rect -7200 3608 -7184 3672
rect -7280 3592 -7184 3608
rect -7280 3528 -7264 3592
rect -7200 3528 -7184 3592
rect -7280 3512 -7184 3528
rect -7280 3448 -7264 3512
rect -7200 3448 -7184 3512
rect -7280 3432 -7184 3448
rect -7280 3368 -7264 3432
rect -7200 3368 -7184 3432
rect -7280 3352 -7184 3368
rect -7280 3288 -7264 3352
rect -7200 3288 -7184 3352
rect -7280 3272 -7184 3288
rect -7280 3208 -7264 3272
rect -7200 3208 -7184 3272
rect -7280 3192 -7184 3208
rect -7280 3128 -7264 3192
rect -7200 3128 -7184 3192
rect -7280 3112 -7184 3128
rect -7280 3048 -7264 3112
rect -7200 3048 -7184 3112
rect -7280 3032 -7184 3048
rect -8692 2932 -8596 2968
rect -7280 2968 -7264 3032
rect -7200 2968 -7184 3032
rect -6861 3712 -6139 3721
rect -6861 3008 -6852 3712
rect -6148 3008 -6139 3712
rect -6861 2999 -6139 3008
rect -5868 3688 -5852 3752
rect -5788 3688 -5772 3752
rect -4456 3752 -4360 3788
rect -5868 3672 -5772 3688
rect -5868 3608 -5852 3672
rect -5788 3608 -5772 3672
rect -5868 3592 -5772 3608
rect -5868 3528 -5852 3592
rect -5788 3528 -5772 3592
rect -5868 3512 -5772 3528
rect -5868 3448 -5852 3512
rect -5788 3448 -5772 3512
rect -5868 3432 -5772 3448
rect -5868 3368 -5852 3432
rect -5788 3368 -5772 3432
rect -5868 3352 -5772 3368
rect -5868 3288 -5852 3352
rect -5788 3288 -5772 3352
rect -5868 3272 -5772 3288
rect -5868 3208 -5852 3272
rect -5788 3208 -5772 3272
rect -5868 3192 -5772 3208
rect -5868 3128 -5852 3192
rect -5788 3128 -5772 3192
rect -5868 3112 -5772 3128
rect -5868 3048 -5852 3112
rect -5788 3048 -5772 3112
rect -5868 3032 -5772 3048
rect -7280 2932 -7184 2968
rect -5868 2968 -5852 3032
rect -5788 2968 -5772 3032
rect -5449 3712 -4727 3721
rect -5449 3008 -5440 3712
rect -4736 3008 -4727 3712
rect -5449 2999 -4727 3008
rect -4456 3688 -4440 3752
rect -4376 3688 -4360 3752
rect -3044 3752 -2948 3788
rect -4456 3672 -4360 3688
rect -4456 3608 -4440 3672
rect -4376 3608 -4360 3672
rect -4456 3592 -4360 3608
rect -4456 3528 -4440 3592
rect -4376 3528 -4360 3592
rect -4456 3512 -4360 3528
rect -4456 3448 -4440 3512
rect -4376 3448 -4360 3512
rect -4456 3432 -4360 3448
rect -4456 3368 -4440 3432
rect -4376 3368 -4360 3432
rect -4456 3352 -4360 3368
rect -4456 3288 -4440 3352
rect -4376 3288 -4360 3352
rect -4456 3272 -4360 3288
rect -4456 3208 -4440 3272
rect -4376 3208 -4360 3272
rect -4456 3192 -4360 3208
rect -4456 3128 -4440 3192
rect -4376 3128 -4360 3192
rect -4456 3112 -4360 3128
rect -4456 3048 -4440 3112
rect -4376 3048 -4360 3112
rect -4456 3032 -4360 3048
rect -5868 2932 -5772 2968
rect -4456 2968 -4440 3032
rect -4376 2968 -4360 3032
rect -4037 3712 -3315 3721
rect -4037 3008 -4028 3712
rect -3324 3008 -3315 3712
rect -4037 2999 -3315 3008
rect -3044 3688 -3028 3752
rect -2964 3688 -2948 3752
rect -1632 3752 -1536 3788
rect -3044 3672 -2948 3688
rect -3044 3608 -3028 3672
rect -2964 3608 -2948 3672
rect -3044 3592 -2948 3608
rect -3044 3528 -3028 3592
rect -2964 3528 -2948 3592
rect -3044 3512 -2948 3528
rect -3044 3448 -3028 3512
rect -2964 3448 -2948 3512
rect -3044 3432 -2948 3448
rect -3044 3368 -3028 3432
rect -2964 3368 -2948 3432
rect -3044 3352 -2948 3368
rect -3044 3288 -3028 3352
rect -2964 3288 -2948 3352
rect -3044 3272 -2948 3288
rect -3044 3208 -3028 3272
rect -2964 3208 -2948 3272
rect -3044 3192 -2948 3208
rect -3044 3128 -3028 3192
rect -2964 3128 -2948 3192
rect -3044 3112 -2948 3128
rect -3044 3048 -3028 3112
rect -2964 3048 -2948 3112
rect -3044 3032 -2948 3048
rect -4456 2932 -4360 2968
rect -3044 2968 -3028 3032
rect -2964 2968 -2948 3032
rect -2625 3712 -1903 3721
rect -2625 3008 -2616 3712
rect -1912 3008 -1903 3712
rect -2625 2999 -1903 3008
rect -1632 3688 -1616 3752
rect -1552 3688 -1536 3752
rect -220 3752 -124 3788
rect -1632 3672 -1536 3688
rect -1632 3608 -1616 3672
rect -1552 3608 -1536 3672
rect -1632 3592 -1536 3608
rect -1632 3528 -1616 3592
rect -1552 3528 -1536 3592
rect -1632 3512 -1536 3528
rect -1632 3448 -1616 3512
rect -1552 3448 -1536 3512
rect -1632 3432 -1536 3448
rect -1632 3368 -1616 3432
rect -1552 3368 -1536 3432
rect -1632 3352 -1536 3368
rect -1632 3288 -1616 3352
rect -1552 3288 -1536 3352
rect -1632 3272 -1536 3288
rect -1632 3208 -1616 3272
rect -1552 3208 -1536 3272
rect -1632 3192 -1536 3208
rect -1632 3128 -1616 3192
rect -1552 3128 -1536 3192
rect -1632 3112 -1536 3128
rect -1632 3048 -1616 3112
rect -1552 3048 -1536 3112
rect -1632 3032 -1536 3048
rect -3044 2932 -2948 2968
rect -1632 2968 -1616 3032
rect -1552 2968 -1536 3032
rect -1213 3712 -491 3721
rect -1213 3008 -1204 3712
rect -500 3008 -491 3712
rect -1213 2999 -491 3008
rect -220 3688 -204 3752
rect -140 3688 -124 3752
rect 1192 3752 1288 3788
rect -220 3672 -124 3688
rect -220 3608 -204 3672
rect -140 3608 -124 3672
rect -220 3592 -124 3608
rect -220 3528 -204 3592
rect -140 3528 -124 3592
rect -220 3512 -124 3528
rect -220 3448 -204 3512
rect -140 3448 -124 3512
rect -220 3432 -124 3448
rect -220 3368 -204 3432
rect -140 3368 -124 3432
rect -220 3352 -124 3368
rect -220 3288 -204 3352
rect -140 3288 -124 3352
rect -220 3272 -124 3288
rect -220 3208 -204 3272
rect -140 3208 -124 3272
rect -220 3192 -124 3208
rect -220 3128 -204 3192
rect -140 3128 -124 3192
rect -220 3112 -124 3128
rect -220 3048 -204 3112
rect -140 3048 -124 3112
rect -220 3032 -124 3048
rect -1632 2932 -1536 2968
rect -220 2968 -204 3032
rect -140 2968 -124 3032
rect 199 3712 921 3721
rect 199 3008 208 3712
rect 912 3008 921 3712
rect 199 2999 921 3008
rect 1192 3688 1208 3752
rect 1272 3688 1288 3752
rect 2604 3752 2700 3788
rect 1192 3672 1288 3688
rect 1192 3608 1208 3672
rect 1272 3608 1288 3672
rect 1192 3592 1288 3608
rect 1192 3528 1208 3592
rect 1272 3528 1288 3592
rect 1192 3512 1288 3528
rect 1192 3448 1208 3512
rect 1272 3448 1288 3512
rect 1192 3432 1288 3448
rect 1192 3368 1208 3432
rect 1272 3368 1288 3432
rect 1192 3352 1288 3368
rect 1192 3288 1208 3352
rect 1272 3288 1288 3352
rect 1192 3272 1288 3288
rect 1192 3208 1208 3272
rect 1272 3208 1288 3272
rect 1192 3192 1288 3208
rect 1192 3128 1208 3192
rect 1272 3128 1288 3192
rect 1192 3112 1288 3128
rect 1192 3048 1208 3112
rect 1272 3048 1288 3112
rect 1192 3032 1288 3048
rect -220 2932 -124 2968
rect 1192 2968 1208 3032
rect 1272 2968 1288 3032
rect 1611 3712 2333 3721
rect 1611 3008 1620 3712
rect 2324 3008 2333 3712
rect 1611 2999 2333 3008
rect 2604 3688 2620 3752
rect 2684 3688 2700 3752
rect 4016 3752 4112 3788
rect 2604 3672 2700 3688
rect 2604 3608 2620 3672
rect 2684 3608 2700 3672
rect 2604 3592 2700 3608
rect 2604 3528 2620 3592
rect 2684 3528 2700 3592
rect 2604 3512 2700 3528
rect 2604 3448 2620 3512
rect 2684 3448 2700 3512
rect 2604 3432 2700 3448
rect 2604 3368 2620 3432
rect 2684 3368 2700 3432
rect 2604 3352 2700 3368
rect 2604 3288 2620 3352
rect 2684 3288 2700 3352
rect 2604 3272 2700 3288
rect 2604 3208 2620 3272
rect 2684 3208 2700 3272
rect 2604 3192 2700 3208
rect 2604 3128 2620 3192
rect 2684 3128 2700 3192
rect 2604 3112 2700 3128
rect 2604 3048 2620 3112
rect 2684 3048 2700 3112
rect 2604 3032 2700 3048
rect 1192 2932 1288 2968
rect 2604 2968 2620 3032
rect 2684 2968 2700 3032
rect 3023 3712 3745 3721
rect 3023 3008 3032 3712
rect 3736 3008 3745 3712
rect 3023 2999 3745 3008
rect 4016 3688 4032 3752
rect 4096 3688 4112 3752
rect 5428 3752 5524 3788
rect 4016 3672 4112 3688
rect 4016 3608 4032 3672
rect 4096 3608 4112 3672
rect 4016 3592 4112 3608
rect 4016 3528 4032 3592
rect 4096 3528 4112 3592
rect 4016 3512 4112 3528
rect 4016 3448 4032 3512
rect 4096 3448 4112 3512
rect 4016 3432 4112 3448
rect 4016 3368 4032 3432
rect 4096 3368 4112 3432
rect 4016 3352 4112 3368
rect 4016 3288 4032 3352
rect 4096 3288 4112 3352
rect 4016 3272 4112 3288
rect 4016 3208 4032 3272
rect 4096 3208 4112 3272
rect 4016 3192 4112 3208
rect 4016 3128 4032 3192
rect 4096 3128 4112 3192
rect 4016 3112 4112 3128
rect 4016 3048 4032 3112
rect 4096 3048 4112 3112
rect 4016 3032 4112 3048
rect 2604 2932 2700 2968
rect 4016 2968 4032 3032
rect 4096 2968 4112 3032
rect 4435 3712 5157 3721
rect 4435 3008 4444 3712
rect 5148 3008 5157 3712
rect 4435 2999 5157 3008
rect 5428 3688 5444 3752
rect 5508 3688 5524 3752
rect 6840 3752 6936 3788
rect 5428 3672 5524 3688
rect 5428 3608 5444 3672
rect 5508 3608 5524 3672
rect 5428 3592 5524 3608
rect 5428 3528 5444 3592
rect 5508 3528 5524 3592
rect 5428 3512 5524 3528
rect 5428 3448 5444 3512
rect 5508 3448 5524 3512
rect 5428 3432 5524 3448
rect 5428 3368 5444 3432
rect 5508 3368 5524 3432
rect 5428 3352 5524 3368
rect 5428 3288 5444 3352
rect 5508 3288 5524 3352
rect 5428 3272 5524 3288
rect 5428 3208 5444 3272
rect 5508 3208 5524 3272
rect 5428 3192 5524 3208
rect 5428 3128 5444 3192
rect 5508 3128 5524 3192
rect 5428 3112 5524 3128
rect 5428 3048 5444 3112
rect 5508 3048 5524 3112
rect 5428 3032 5524 3048
rect 4016 2932 4112 2968
rect 5428 2968 5444 3032
rect 5508 2968 5524 3032
rect 5847 3712 6569 3721
rect 5847 3008 5856 3712
rect 6560 3008 6569 3712
rect 5847 2999 6569 3008
rect 6840 3688 6856 3752
rect 6920 3688 6936 3752
rect 8252 3752 8348 3788
rect 6840 3672 6936 3688
rect 6840 3608 6856 3672
rect 6920 3608 6936 3672
rect 6840 3592 6936 3608
rect 6840 3528 6856 3592
rect 6920 3528 6936 3592
rect 6840 3512 6936 3528
rect 6840 3448 6856 3512
rect 6920 3448 6936 3512
rect 6840 3432 6936 3448
rect 6840 3368 6856 3432
rect 6920 3368 6936 3432
rect 6840 3352 6936 3368
rect 6840 3288 6856 3352
rect 6920 3288 6936 3352
rect 6840 3272 6936 3288
rect 6840 3208 6856 3272
rect 6920 3208 6936 3272
rect 6840 3192 6936 3208
rect 6840 3128 6856 3192
rect 6920 3128 6936 3192
rect 6840 3112 6936 3128
rect 6840 3048 6856 3112
rect 6920 3048 6936 3112
rect 6840 3032 6936 3048
rect 5428 2932 5524 2968
rect 6840 2968 6856 3032
rect 6920 2968 6936 3032
rect 7259 3712 7981 3721
rect 7259 3008 7268 3712
rect 7972 3008 7981 3712
rect 7259 2999 7981 3008
rect 8252 3688 8268 3752
rect 8332 3688 8348 3752
rect 9664 3752 9760 3788
rect 8252 3672 8348 3688
rect 8252 3608 8268 3672
rect 8332 3608 8348 3672
rect 8252 3592 8348 3608
rect 8252 3528 8268 3592
rect 8332 3528 8348 3592
rect 8252 3512 8348 3528
rect 8252 3448 8268 3512
rect 8332 3448 8348 3512
rect 8252 3432 8348 3448
rect 8252 3368 8268 3432
rect 8332 3368 8348 3432
rect 8252 3352 8348 3368
rect 8252 3288 8268 3352
rect 8332 3288 8348 3352
rect 8252 3272 8348 3288
rect 8252 3208 8268 3272
rect 8332 3208 8348 3272
rect 8252 3192 8348 3208
rect 8252 3128 8268 3192
rect 8332 3128 8348 3192
rect 8252 3112 8348 3128
rect 8252 3048 8268 3112
rect 8332 3048 8348 3112
rect 8252 3032 8348 3048
rect 6840 2932 6936 2968
rect 8252 2968 8268 3032
rect 8332 2968 8348 3032
rect 8671 3712 9393 3721
rect 8671 3008 8680 3712
rect 9384 3008 9393 3712
rect 8671 2999 9393 3008
rect 9664 3688 9680 3752
rect 9744 3688 9760 3752
rect 11076 3752 11172 3788
rect 9664 3672 9760 3688
rect 9664 3608 9680 3672
rect 9744 3608 9760 3672
rect 9664 3592 9760 3608
rect 9664 3528 9680 3592
rect 9744 3528 9760 3592
rect 9664 3512 9760 3528
rect 9664 3448 9680 3512
rect 9744 3448 9760 3512
rect 9664 3432 9760 3448
rect 9664 3368 9680 3432
rect 9744 3368 9760 3432
rect 9664 3352 9760 3368
rect 9664 3288 9680 3352
rect 9744 3288 9760 3352
rect 9664 3272 9760 3288
rect 9664 3208 9680 3272
rect 9744 3208 9760 3272
rect 9664 3192 9760 3208
rect 9664 3128 9680 3192
rect 9744 3128 9760 3192
rect 9664 3112 9760 3128
rect 9664 3048 9680 3112
rect 9744 3048 9760 3112
rect 9664 3032 9760 3048
rect 8252 2932 8348 2968
rect 9664 2968 9680 3032
rect 9744 2968 9760 3032
rect 10083 3712 10805 3721
rect 10083 3008 10092 3712
rect 10796 3008 10805 3712
rect 10083 2999 10805 3008
rect 11076 3688 11092 3752
rect 11156 3688 11172 3752
rect 12488 3752 12584 3788
rect 11076 3672 11172 3688
rect 11076 3608 11092 3672
rect 11156 3608 11172 3672
rect 11076 3592 11172 3608
rect 11076 3528 11092 3592
rect 11156 3528 11172 3592
rect 11076 3512 11172 3528
rect 11076 3448 11092 3512
rect 11156 3448 11172 3512
rect 11076 3432 11172 3448
rect 11076 3368 11092 3432
rect 11156 3368 11172 3432
rect 11076 3352 11172 3368
rect 11076 3288 11092 3352
rect 11156 3288 11172 3352
rect 11076 3272 11172 3288
rect 11076 3208 11092 3272
rect 11156 3208 11172 3272
rect 11076 3192 11172 3208
rect 11076 3128 11092 3192
rect 11156 3128 11172 3192
rect 11076 3112 11172 3128
rect 11076 3048 11092 3112
rect 11156 3048 11172 3112
rect 11076 3032 11172 3048
rect 9664 2932 9760 2968
rect 11076 2968 11092 3032
rect 11156 2968 11172 3032
rect 11495 3712 12217 3721
rect 11495 3008 11504 3712
rect 12208 3008 12217 3712
rect 11495 2999 12217 3008
rect 12488 3688 12504 3752
rect 12568 3688 12584 3752
rect 13900 3752 13996 3788
rect 12488 3672 12584 3688
rect 12488 3608 12504 3672
rect 12568 3608 12584 3672
rect 12488 3592 12584 3608
rect 12488 3528 12504 3592
rect 12568 3528 12584 3592
rect 12488 3512 12584 3528
rect 12488 3448 12504 3512
rect 12568 3448 12584 3512
rect 12488 3432 12584 3448
rect 12488 3368 12504 3432
rect 12568 3368 12584 3432
rect 12488 3352 12584 3368
rect 12488 3288 12504 3352
rect 12568 3288 12584 3352
rect 12488 3272 12584 3288
rect 12488 3208 12504 3272
rect 12568 3208 12584 3272
rect 12488 3192 12584 3208
rect 12488 3128 12504 3192
rect 12568 3128 12584 3192
rect 12488 3112 12584 3128
rect 12488 3048 12504 3112
rect 12568 3048 12584 3112
rect 12488 3032 12584 3048
rect 11076 2932 11172 2968
rect 12488 2968 12504 3032
rect 12568 2968 12584 3032
rect 12907 3712 13629 3721
rect 12907 3008 12916 3712
rect 13620 3008 13629 3712
rect 12907 2999 13629 3008
rect 13900 3688 13916 3752
rect 13980 3688 13996 3752
rect 15312 3752 15408 3788
rect 13900 3672 13996 3688
rect 13900 3608 13916 3672
rect 13980 3608 13996 3672
rect 13900 3592 13996 3608
rect 13900 3528 13916 3592
rect 13980 3528 13996 3592
rect 13900 3512 13996 3528
rect 13900 3448 13916 3512
rect 13980 3448 13996 3512
rect 13900 3432 13996 3448
rect 13900 3368 13916 3432
rect 13980 3368 13996 3432
rect 13900 3352 13996 3368
rect 13900 3288 13916 3352
rect 13980 3288 13996 3352
rect 13900 3272 13996 3288
rect 13900 3208 13916 3272
rect 13980 3208 13996 3272
rect 13900 3192 13996 3208
rect 13900 3128 13916 3192
rect 13980 3128 13996 3192
rect 13900 3112 13996 3128
rect 13900 3048 13916 3112
rect 13980 3048 13996 3112
rect 13900 3032 13996 3048
rect 12488 2932 12584 2968
rect 13900 2968 13916 3032
rect 13980 2968 13996 3032
rect 14319 3712 15041 3721
rect 14319 3008 14328 3712
rect 15032 3008 15041 3712
rect 14319 2999 15041 3008
rect 15312 3688 15328 3752
rect 15392 3688 15408 3752
rect 16724 3752 16820 3788
rect 15312 3672 15408 3688
rect 15312 3608 15328 3672
rect 15392 3608 15408 3672
rect 15312 3592 15408 3608
rect 15312 3528 15328 3592
rect 15392 3528 15408 3592
rect 15312 3512 15408 3528
rect 15312 3448 15328 3512
rect 15392 3448 15408 3512
rect 15312 3432 15408 3448
rect 15312 3368 15328 3432
rect 15392 3368 15408 3432
rect 15312 3352 15408 3368
rect 15312 3288 15328 3352
rect 15392 3288 15408 3352
rect 15312 3272 15408 3288
rect 15312 3208 15328 3272
rect 15392 3208 15408 3272
rect 15312 3192 15408 3208
rect 15312 3128 15328 3192
rect 15392 3128 15408 3192
rect 15312 3112 15408 3128
rect 15312 3048 15328 3112
rect 15392 3048 15408 3112
rect 15312 3032 15408 3048
rect 13900 2932 13996 2968
rect 15312 2968 15328 3032
rect 15392 2968 15408 3032
rect 15731 3712 16453 3721
rect 15731 3008 15740 3712
rect 16444 3008 16453 3712
rect 15731 2999 16453 3008
rect 16724 3688 16740 3752
rect 16804 3688 16820 3752
rect 18136 3752 18232 3788
rect 16724 3672 16820 3688
rect 16724 3608 16740 3672
rect 16804 3608 16820 3672
rect 16724 3592 16820 3608
rect 16724 3528 16740 3592
rect 16804 3528 16820 3592
rect 16724 3512 16820 3528
rect 16724 3448 16740 3512
rect 16804 3448 16820 3512
rect 16724 3432 16820 3448
rect 16724 3368 16740 3432
rect 16804 3368 16820 3432
rect 16724 3352 16820 3368
rect 16724 3288 16740 3352
rect 16804 3288 16820 3352
rect 16724 3272 16820 3288
rect 16724 3208 16740 3272
rect 16804 3208 16820 3272
rect 16724 3192 16820 3208
rect 16724 3128 16740 3192
rect 16804 3128 16820 3192
rect 16724 3112 16820 3128
rect 16724 3048 16740 3112
rect 16804 3048 16820 3112
rect 16724 3032 16820 3048
rect 15312 2932 15408 2968
rect 16724 2968 16740 3032
rect 16804 2968 16820 3032
rect 17143 3712 17865 3721
rect 17143 3008 17152 3712
rect 17856 3008 17865 3712
rect 17143 2999 17865 3008
rect 18136 3688 18152 3752
rect 18216 3688 18232 3752
rect 19548 3752 19644 3788
rect 18136 3672 18232 3688
rect 18136 3608 18152 3672
rect 18216 3608 18232 3672
rect 18136 3592 18232 3608
rect 18136 3528 18152 3592
rect 18216 3528 18232 3592
rect 18136 3512 18232 3528
rect 18136 3448 18152 3512
rect 18216 3448 18232 3512
rect 18136 3432 18232 3448
rect 18136 3368 18152 3432
rect 18216 3368 18232 3432
rect 18136 3352 18232 3368
rect 18136 3288 18152 3352
rect 18216 3288 18232 3352
rect 18136 3272 18232 3288
rect 18136 3208 18152 3272
rect 18216 3208 18232 3272
rect 18136 3192 18232 3208
rect 18136 3128 18152 3192
rect 18216 3128 18232 3192
rect 18136 3112 18232 3128
rect 18136 3048 18152 3112
rect 18216 3048 18232 3112
rect 18136 3032 18232 3048
rect 16724 2932 16820 2968
rect 18136 2968 18152 3032
rect 18216 2968 18232 3032
rect 18555 3712 19277 3721
rect 18555 3008 18564 3712
rect 19268 3008 19277 3712
rect 18555 2999 19277 3008
rect 19548 3688 19564 3752
rect 19628 3688 19644 3752
rect 20960 3752 21056 3788
rect 19548 3672 19644 3688
rect 19548 3608 19564 3672
rect 19628 3608 19644 3672
rect 19548 3592 19644 3608
rect 19548 3528 19564 3592
rect 19628 3528 19644 3592
rect 19548 3512 19644 3528
rect 19548 3448 19564 3512
rect 19628 3448 19644 3512
rect 19548 3432 19644 3448
rect 19548 3368 19564 3432
rect 19628 3368 19644 3432
rect 19548 3352 19644 3368
rect 19548 3288 19564 3352
rect 19628 3288 19644 3352
rect 19548 3272 19644 3288
rect 19548 3208 19564 3272
rect 19628 3208 19644 3272
rect 19548 3192 19644 3208
rect 19548 3128 19564 3192
rect 19628 3128 19644 3192
rect 19548 3112 19644 3128
rect 19548 3048 19564 3112
rect 19628 3048 19644 3112
rect 19548 3032 19644 3048
rect 18136 2932 18232 2968
rect 19548 2968 19564 3032
rect 19628 2968 19644 3032
rect 19967 3712 20689 3721
rect 19967 3008 19976 3712
rect 20680 3008 20689 3712
rect 19967 2999 20689 3008
rect 20960 3688 20976 3752
rect 21040 3688 21056 3752
rect 22372 3752 22468 3788
rect 20960 3672 21056 3688
rect 20960 3608 20976 3672
rect 21040 3608 21056 3672
rect 20960 3592 21056 3608
rect 20960 3528 20976 3592
rect 21040 3528 21056 3592
rect 20960 3512 21056 3528
rect 20960 3448 20976 3512
rect 21040 3448 21056 3512
rect 20960 3432 21056 3448
rect 20960 3368 20976 3432
rect 21040 3368 21056 3432
rect 20960 3352 21056 3368
rect 20960 3288 20976 3352
rect 21040 3288 21056 3352
rect 20960 3272 21056 3288
rect 20960 3208 20976 3272
rect 21040 3208 21056 3272
rect 20960 3192 21056 3208
rect 20960 3128 20976 3192
rect 21040 3128 21056 3192
rect 20960 3112 21056 3128
rect 20960 3048 20976 3112
rect 21040 3048 21056 3112
rect 20960 3032 21056 3048
rect 19548 2932 19644 2968
rect 20960 2968 20976 3032
rect 21040 2968 21056 3032
rect 21379 3712 22101 3721
rect 21379 3008 21388 3712
rect 22092 3008 22101 3712
rect 21379 2999 22101 3008
rect 22372 3688 22388 3752
rect 22452 3688 22468 3752
rect 23784 3752 23880 3788
rect 22372 3672 22468 3688
rect 22372 3608 22388 3672
rect 22452 3608 22468 3672
rect 22372 3592 22468 3608
rect 22372 3528 22388 3592
rect 22452 3528 22468 3592
rect 22372 3512 22468 3528
rect 22372 3448 22388 3512
rect 22452 3448 22468 3512
rect 22372 3432 22468 3448
rect 22372 3368 22388 3432
rect 22452 3368 22468 3432
rect 22372 3352 22468 3368
rect 22372 3288 22388 3352
rect 22452 3288 22468 3352
rect 22372 3272 22468 3288
rect 22372 3208 22388 3272
rect 22452 3208 22468 3272
rect 22372 3192 22468 3208
rect 22372 3128 22388 3192
rect 22452 3128 22468 3192
rect 22372 3112 22468 3128
rect 22372 3048 22388 3112
rect 22452 3048 22468 3112
rect 22372 3032 22468 3048
rect 20960 2932 21056 2968
rect 22372 2968 22388 3032
rect 22452 2968 22468 3032
rect 22791 3712 23513 3721
rect 22791 3008 22800 3712
rect 23504 3008 23513 3712
rect 22791 2999 23513 3008
rect 23784 3688 23800 3752
rect 23864 3688 23880 3752
rect 23784 3672 23880 3688
rect 23784 3608 23800 3672
rect 23864 3608 23880 3672
rect 23784 3592 23880 3608
rect 23784 3528 23800 3592
rect 23864 3528 23880 3592
rect 23784 3512 23880 3528
rect 23784 3448 23800 3512
rect 23864 3448 23880 3512
rect 23784 3432 23880 3448
rect 23784 3368 23800 3432
rect 23864 3368 23880 3432
rect 23784 3352 23880 3368
rect 23784 3288 23800 3352
rect 23864 3288 23880 3352
rect 23784 3272 23880 3288
rect 23784 3208 23800 3272
rect 23864 3208 23880 3272
rect 23784 3192 23880 3208
rect 23784 3128 23800 3192
rect 23864 3128 23880 3192
rect 23784 3112 23880 3128
rect 23784 3048 23800 3112
rect 23864 3048 23880 3112
rect 23784 3032 23880 3048
rect 22372 2932 22468 2968
rect 23784 2968 23800 3032
rect 23864 2968 23880 3032
rect 23784 2932 23880 2968
rect -22812 2632 -22716 2668
rect -23805 2592 -23083 2601
rect -23805 1888 -23796 2592
rect -23092 1888 -23083 2592
rect -23805 1879 -23083 1888
rect -22812 2568 -22796 2632
rect -22732 2568 -22716 2632
rect -21400 2632 -21304 2668
rect -22812 2552 -22716 2568
rect -22812 2488 -22796 2552
rect -22732 2488 -22716 2552
rect -22812 2472 -22716 2488
rect -22812 2408 -22796 2472
rect -22732 2408 -22716 2472
rect -22812 2392 -22716 2408
rect -22812 2328 -22796 2392
rect -22732 2328 -22716 2392
rect -22812 2312 -22716 2328
rect -22812 2248 -22796 2312
rect -22732 2248 -22716 2312
rect -22812 2232 -22716 2248
rect -22812 2168 -22796 2232
rect -22732 2168 -22716 2232
rect -22812 2152 -22716 2168
rect -22812 2088 -22796 2152
rect -22732 2088 -22716 2152
rect -22812 2072 -22716 2088
rect -22812 2008 -22796 2072
rect -22732 2008 -22716 2072
rect -22812 1992 -22716 2008
rect -22812 1928 -22796 1992
rect -22732 1928 -22716 1992
rect -22812 1912 -22716 1928
rect -22812 1848 -22796 1912
rect -22732 1848 -22716 1912
rect -22393 2592 -21671 2601
rect -22393 1888 -22384 2592
rect -21680 1888 -21671 2592
rect -22393 1879 -21671 1888
rect -21400 2568 -21384 2632
rect -21320 2568 -21304 2632
rect -19988 2632 -19892 2668
rect -21400 2552 -21304 2568
rect -21400 2488 -21384 2552
rect -21320 2488 -21304 2552
rect -21400 2472 -21304 2488
rect -21400 2408 -21384 2472
rect -21320 2408 -21304 2472
rect -21400 2392 -21304 2408
rect -21400 2328 -21384 2392
rect -21320 2328 -21304 2392
rect -21400 2312 -21304 2328
rect -21400 2248 -21384 2312
rect -21320 2248 -21304 2312
rect -21400 2232 -21304 2248
rect -21400 2168 -21384 2232
rect -21320 2168 -21304 2232
rect -21400 2152 -21304 2168
rect -21400 2088 -21384 2152
rect -21320 2088 -21304 2152
rect -21400 2072 -21304 2088
rect -21400 2008 -21384 2072
rect -21320 2008 -21304 2072
rect -21400 1992 -21304 2008
rect -21400 1928 -21384 1992
rect -21320 1928 -21304 1992
rect -21400 1912 -21304 1928
rect -22812 1812 -22716 1848
rect -21400 1848 -21384 1912
rect -21320 1848 -21304 1912
rect -20981 2592 -20259 2601
rect -20981 1888 -20972 2592
rect -20268 1888 -20259 2592
rect -20981 1879 -20259 1888
rect -19988 2568 -19972 2632
rect -19908 2568 -19892 2632
rect -18576 2632 -18480 2668
rect -19988 2552 -19892 2568
rect -19988 2488 -19972 2552
rect -19908 2488 -19892 2552
rect -19988 2472 -19892 2488
rect -19988 2408 -19972 2472
rect -19908 2408 -19892 2472
rect -19988 2392 -19892 2408
rect -19988 2328 -19972 2392
rect -19908 2328 -19892 2392
rect -19988 2312 -19892 2328
rect -19988 2248 -19972 2312
rect -19908 2248 -19892 2312
rect -19988 2232 -19892 2248
rect -19988 2168 -19972 2232
rect -19908 2168 -19892 2232
rect -19988 2152 -19892 2168
rect -19988 2088 -19972 2152
rect -19908 2088 -19892 2152
rect -19988 2072 -19892 2088
rect -19988 2008 -19972 2072
rect -19908 2008 -19892 2072
rect -19988 1992 -19892 2008
rect -19988 1928 -19972 1992
rect -19908 1928 -19892 1992
rect -19988 1912 -19892 1928
rect -21400 1812 -21304 1848
rect -19988 1848 -19972 1912
rect -19908 1848 -19892 1912
rect -19569 2592 -18847 2601
rect -19569 1888 -19560 2592
rect -18856 1888 -18847 2592
rect -19569 1879 -18847 1888
rect -18576 2568 -18560 2632
rect -18496 2568 -18480 2632
rect -17164 2632 -17068 2668
rect -18576 2552 -18480 2568
rect -18576 2488 -18560 2552
rect -18496 2488 -18480 2552
rect -18576 2472 -18480 2488
rect -18576 2408 -18560 2472
rect -18496 2408 -18480 2472
rect -18576 2392 -18480 2408
rect -18576 2328 -18560 2392
rect -18496 2328 -18480 2392
rect -18576 2312 -18480 2328
rect -18576 2248 -18560 2312
rect -18496 2248 -18480 2312
rect -18576 2232 -18480 2248
rect -18576 2168 -18560 2232
rect -18496 2168 -18480 2232
rect -18576 2152 -18480 2168
rect -18576 2088 -18560 2152
rect -18496 2088 -18480 2152
rect -18576 2072 -18480 2088
rect -18576 2008 -18560 2072
rect -18496 2008 -18480 2072
rect -18576 1992 -18480 2008
rect -18576 1928 -18560 1992
rect -18496 1928 -18480 1992
rect -18576 1912 -18480 1928
rect -19988 1812 -19892 1848
rect -18576 1848 -18560 1912
rect -18496 1848 -18480 1912
rect -18157 2592 -17435 2601
rect -18157 1888 -18148 2592
rect -17444 1888 -17435 2592
rect -18157 1879 -17435 1888
rect -17164 2568 -17148 2632
rect -17084 2568 -17068 2632
rect -15752 2632 -15656 2668
rect -17164 2552 -17068 2568
rect -17164 2488 -17148 2552
rect -17084 2488 -17068 2552
rect -17164 2472 -17068 2488
rect -17164 2408 -17148 2472
rect -17084 2408 -17068 2472
rect -17164 2392 -17068 2408
rect -17164 2328 -17148 2392
rect -17084 2328 -17068 2392
rect -17164 2312 -17068 2328
rect -17164 2248 -17148 2312
rect -17084 2248 -17068 2312
rect -17164 2232 -17068 2248
rect -17164 2168 -17148 2232
rect -17084 2168 -17068 2232
rect -17164 2152 -17068 2168
rect -17164 2088 -17148 2152
rect -17084 2088 -17068 2152
rect -17164 2072 -17068 2088
rect -17164 2008 -17148 2072
rect -17084 2008 -17068 2072
rect -17164 1992 -17068 2008
rect -17164 1928 -17148 1992
rect -17084 1928 -17068 1992
rect -17164 1912 -17068 1928
rect -18576 1812 -18480 1848
rect -17164 1848 -17148 1912
rect -17084 1848 -17068 1912
rect -16745 2592 -16023 2601
rect -16745 1888 -16736 2592
rect -16032 1888 -16023 2592
rect -16745 1879 -16023 1888
rect -15752 2568 -15736 2632
rect -15672 2568 -15656 2632
rect -14340 2632 -14244 2668
rect -15752 2552 -15656 2568
rect -15752 2488 -15736 2552
rect -15672 2488 -15656 2552
rect -15752 2472 -15656 2488
rect -15752 2408 -15736 2472
rect -15672 2408 -15656 2472
rect -15752 2392 -15656 2408
rect -15752 2328 -15736 2392
rect -15672 2328 -15656 2392
rect -15752 2312 -15656 2328
rect -15752 2248 -15736 2312
rect -15672 2248 -15656 2312
rect -15752 2232 -15656 2248
rect -15752 2168 -15736 2232
rect -15672 2168 -15656 2232
rect -15752 2152 -15656 2168
rect -15752 2088 -15736 2152
rect -15672 2088 -15656 2152
rect -15752 2072 -15656 2088
rect -15752 2008 -15736 2072
rect -15672 2008 -15656 2072
rect -15752 1992 -15656 2008
rect -15752 1928 -15736 1992
rect -15672 1928 -15656 1992
rect -15752 1912 -15656 1928
rect -17164 1812 -17068 1848
rect -15752 1848 -15736 1912
rect -15672 1848 -15656 1912
rect -15333 2592 -14611 2601
rect -15333 1888 -15324 2592
rect -14620 1888 -14611 2592
rect -15333 1879 -14611 1888
rect -14340 2568 -14324 2632
rect -14260 2568 -14244 2632
rect -12928 2632 -12832 2668
rect -14340 2552 -14244 2568
rect -14340 2488 -14324 2552
rect -14260 2488 -14244 2552
rect -14340 2472 -14244 2488
rect -14340 2408 -14324 2472
rect -14260 2408 -14244 2472
rect -14340 2392 -14244 2408
rect -14340 2328 -14324 2392
rect -14260 2328 -14244 2392
rect -14340 2312 -14244 2328
rect -14340 2248 -14324 2312
rect -14260 2248 -14244 2312
rect -14340 2232 -14244 2248
rect -14340 2168 -14324 2232
rect -14260 2168 -14244 2232
rect -14340 2152 -14244 2168
rect -14340 2088 -14324 2152
rect -14260 2088 -14244 2152
rect -14340 2072 -14244 2088
rect -14340 2008 -14324 2072
rect -14260 2008 -14244 2072
rect -14340 1992 -14244 2008
rect -14340 1928 -14324 1992
rect -14260 1928 -14244 1992
rect -14340 1912 -14244 1928
rect -15752 1812 -15656 1848
rect -14340 1848 -14324 1912
rect -14260 1848 -14244 1912
rect -13921 2592 -13199 2601
rect -13921 1888 -13912 2592
rect -13208 1888 -13199 2592
rect -13921 1879 -13199 1888
rect -12928 2568 -12912 2632
rect -12848 2568 -12832 2632
rect -11516 2632 -11420 2668
rect -12928 2552 -12832 2568
rect -12928 2488 -12912 2552
rect -12848 2488 -12832 2552
rect -12928 2472 -12832 2488
rect -12928 2408 -12912 2472
rect -12848 2408 -12832 2472
rect -12928 2392 -12832 2408
rect -12928 2328 -12912 2392
rect -12848 2328 -12832 2392
rect -12928 2312 -12832 2328
rect -12928 2248 -12912 2312
rect -12848 2248 -12832 2312
rect -12928 2232 -12832 2248
rect -12928 2168 -12912 2232
rect -12848 2168 -12832 2232
rect -12928 2152 -12832 2168
rect -12928 2088 -12912 2152
rect -12848 2088 -12832 2152
rect -12928 2072 -12832 2088
rect -12928 2008 -12912 2072
rect -12848 2008 -12832 2072
rect -12928 1992 -12832 2008
rect -12928 1928 -12912 1992
rect -12848 1928 -12832 1992
rect -12928 1912 -12832 1928
rect -14340 1812 -14244 1848
rect -12928 1848 -12912 1912
rect -12848 1848 -12832 1912
rect -12509 2592 -11787 2601
rect -12509 1888 -12500 2592
rect -11796 1888 -11787 2592
rect -12509 1879 -11787 1888
rect -11516 2568 -11500 2632
rect -11436 2568 -11420 2632
rect -10104 2632 -10008 2668
rect -11516 2552 -11420 2568
rect -11516 2488 -11500 2552
rect -11436 2488 -11420 2552
rect -11516 2472 -11420 2488
rect -11516 2408 -11500 2472
rect -11436 2408 -11420 2472
rect -11516 2392 -11420 2408
rect -11516 2328 -11500 2392
rect -11436 2328 -11420 2392
rect -11516 2312 -11420 2328
rect -11516 2248 -11500 2312
rect -11436 2248 -11420 2312
rect -11516 2232 -11420 2248
rect -11516 2168 -11500 2232
rect -11436 2168 -11420 2232
rect -11516 2152 -11420 2168
rect -11516 2088 -11500 2152
rect -11436 2088 -11420 2152
rect -11516 2072 -11420 2088
rect -11516 2008 -11500 2072
rect -11436 2008 -11420 2072
rect -11516 1992 -11420 2008
rect -11516 1928 -11500 1992
rect -11436 1928 -11420 1992
rect -11516 1912 -11420 1928
rect -12928 1812 -12832 1848
rect -11516 1848 -11500 1912
rect -11436 1848 -11420 1912
rect -11097 2592 -10375 2601
rect -11097 1888 -11088 2592
rect -10384 1888 -10375 2592
rect -11097 1879 -10375 1888
rect -10104 2568 -10088 2632
rect -10024 2568 -10008 2632
rect -8692 2632 -8596 2668
rect -10104 2552 -10008 2568
rect -10104 2488 -10088 2552
rect -10024 2488 -10008 2552
rect -10104 2472 -10008 2488
rect -10104 2408 -10088 2472
rect -10024 2408 -10008 2472
rect -10104 2392 -10008 2408
rect -10104 2328 -10088 2392
rect -10024 2328 -10008 2392
rect -10104 2312 -10008 2328
rect -10104 2248 -10088 2312
rect -10024 2248 -10008 2312
rect -10104 2232 -10008 2248
rect -10104 2168 -10088 2232
rect -10024 2168 -10008 2232
rect -10104 2152 -10008 2168
rect -10104 2088 -10088 2152
rect -10024 2088 -10008 2152
rect -10104 2072 -10008 2088
rect -10104 2008 -10088 2072
rect -10024 2008 -10008 2072
rect -10104 1992 -10008 2008
rect -10104 1928 -10088 1992
rect -10024 1928 -10008 1992
rect -10104 1912 -10008 1928
rect -11516 1812 -11420 1848
rect -10104 1848 -10088 1912
rect -10024 1848 -10008 1912
rect -9685 2592 -8963 2601
rect -9685 1888 -9676 2592
rect -8972 1888 -8963 2592
rect -9685 1879 -8963 1888
rect -8692 2568 -8676 2632
rect -8612 2568 -8596 2632
rect -7280 2632 -7184 2668
rect -8692 2552 -8596 2568
rect -8692 2488 -8676 2552
rect -8612 2488 -8596 2552
rect -8692 2472 -8596 2488
rect -8692 2408 -8676 2472
rect -8612 2408 -8596 2472
rect -8692 2392 -8596 2408
rect -8692 2328 -8676 2392
rect -8612 2328 -8596 2392
rect -8692 2312 -8596 2328
rect -8692 2248 -8676 2312
rect -8612 2248 -8596 2312
rect -8692 2232 -8596 2248
rect -8692 2168 -8676 2232
rect -8612 2168 -8596 2232
rect -8692 2152 -8596 2168
rect -8692 2088 -8676 2152
rect -8612 2088 -8596 2152
rect -8692 2072 -8596 2088
rect -8692 2008 -8676 2072
rect -8612 2008 -8596 2072
rect -8692 1992 -8596 2008
rect -8692 1928 -8676 1992
rect -8612 1928 -8596 1992
rect -8692 1912 -8596 1928
rect -10104 1812 -10008 1848
rect -8692 1848 -8676 1912
rect -8612 1848 -8596 1912
rect -8273 2592 -7551 2601
rect -8273 1888 -8264 2592
rect -7560 1888 -7551 2592
rect -8273 1879 -7551 1888
rect -7280 2568 -7264 2632
rect -7200 2568 -7184 2632
rect -5868 2632 -5772 2668
rect -7280 2552 -7184 2568
rect -7280 2488 -7264 2552
rect -7200 2488 -7184 2552
rect -7280 2472 -7184 2488
rect -7280 2408 -7264 2472
rect -7200 2408 -7184 2472
rect -7280 2392 -7184 2408
rect -7280 2328 -7264 2392
rect -7200 2328 -7184 2392
rect -7280 2312 -7184 2328
rect -7280 2248 -7264 2312
rect -7200 2248 -7184 2312
rect -7280 2232 -7184 2248
rect -7280 2168 -7264 2232
rect -7200 2168 -7184 2232
rect -7280 2152 -7184 2168
rect -7280 2088 -7264 2152
rect -7200 2088 -7184 2152
rect -7280 2072 -7184 2088
rect -7280 2008 -7264 2072
rect -7200 2008 -7184 2072
rect -7280 1992 -7184 2008
rect -7280 1928 -7264 1992
rect -7200 1928 -7184 1992
rect -7280 1912 -7184 1928
rect -8692 1812 -8596 1848
rect -7280 1848 -7264 1912
rect -7200 1848 -7184 1912
rect -6861 2592 -6139 2601
rect -6861 1888 -6852 2592
rect -6148 1888 -6139 2592
rect -6861 1879 -6139 1888
rect -5868 2568 -5852 2632
rect -5788 2568 -5772 2632
rect -4456 2632 -4360 2668
rect -5868 2552 -5772 2568
rect -5868 2488 -5852 2552
rect -5788 2488 -5772 2552
rect -5868 2472 -5772 2488
rect -5868 2408 -5852 2472
rect -5788 2408 -5772 2472
rect -5868 2392 -5772 2408
rect -5868 2328 -5852 2392
rect -5788 2328 -5772 2392
rect -5868 2312 -5772 2328
rect -5868 2248 -5852 2312
rect -5788 2248 -5772 2312
rect -5868 2232 -5772 2248
rect -5868 2168 -5852 2232
rect -5788 2168 -5772 2232
rect -5868 2152 -5772 2168
rect -5868 2088 -5852 2152
rect -5788 2088 -5772 2152
rect -5868 2072 -5772 2088
rect -5868 2008 -5852 2072
rect -5788 2008 -5772 2072
rect -5868 1992 -5772 2008
rect -5868 1928 -5852 1992
rect -5788 1928 -5772 1992
rect -5868 1912 -5772 1928
rect -7280 1812 -7184 1848
rect -5868 1848 -5852 1912
rect -5788 1848 -5772 1912
rect -5449 2592 -4727 2601
rect -5449 1888 -5440 2592
rect -4736 1888 -4727 2592
rect -5449 1879 -4727 1888
rect -4456 2568 -4440 2632
rect -4376 2568 -4360 2632
rect -3044 2632 -2948 2668
rect -4456 2552 -4360 2568
rect -4456 2488 -4440 2552
rect -4376 2488 -4360 2552
rect -4456 2472 -4360 2488
rect -4456 2408 -4440 2472
rect -4376 2408 -4360 2472
rect -4456 2392 -4360 2408
rect -4456 2328 -4440 2392
rect -4376 2328 -4360 2392
rect -4456 2312 -4360 2328
rect -4456 2248 -4440 2312
rect -4376 2248 -4360 2312
rect -4456 2232 -4360 2248
rect -4456 2168 -4440 2232
rect -4376 2168 -4360 2232
rect -4456 2152 -4360 2168
rect -4456 2088 -4440 2152
rect -4376 2088 -4360 2152
rect -4456 2072 -4360 2088
rect -4456 2008 -4440 2072
rect -4376 2008 -4360 2072
rect -4456 1992 -4360 2008
rect -4456 1928 -4440 1992
rect -4376 1928 -4360 1992
rect -4456 1912 -4360 1928
rect -5868 1812 -5772 1848
rect -4456 1848 -4440 1912
rect -4376 1848 -4360 1912
rect -4037 2592 -3315 2601
rect -4037 1888 -4028 2592
rect -3324 1888 -3315 2592
rect -4037 1879 -3315 1888
rect -3044 2568 -3028 2632
rect -2964 2568 -2948 2632
rect -1632 2632 -1536 2668
rect -3044 2552 -2948 2568
rect -3044 2488 -3028 2552
rect -2964 2488 -2948 2552
rect -3044 2472 -2948 2488
rect -3044 2408 -3028 2472
rect -2964 2408 -2948 2472
rect -3044 2392 -2948 2408
rect -3044 2328 -3028 2392
rect -2964 2328 -2948 2392
rect -3044 2312 -2948 2328
rect -3044 2248 -3028 2312
rect -2964 2248 -2948 2312
rect -3044 2232 -2948 2248
rect -3044 2168 -3028 2232
rect -2964 2168 -2948 2232
rect -3044 2152 -2948 2168
rect -3044 2088 -3028 2152
rect -2964 2088 -2948 2152
rect -3044 2072 -2948 2088
rect -3044 2008 -3028 2072
rect -2964 2008 -2948 2072
rect -3044 1992 -2948 2008
rect -3044 1928 -3028 1992
rect -2964 1928 -2948 1992
rect -3044 1912 -2948 1928
rect -4456 1812 -4360 1848
rect -3044 1848 -3028 1912
rect -2964 1848 -2948 1912
rect -2625 2592 -1903 2601
rect -2625 1888 -2616 2592
rect -1912 1888 -1903 2592
rect -2625 1879 -1903 1888
rect -1632 2568 -1616 2632
rect -1552 2568 -1536 2632
rect -220 2632 -124 2668
rect -1632 2552 -1536 2568
rect -1632 2488 -1616 2552
rect -1552 2488 -1536 2552
rect -1632 2472 -1536 2488
rect -1632 2408 -1616 2472
rect -1552 2408 -1536 2472
rect -1632 2392 -1536 2408
rect -1632 2328 -1616 2392
rect -1552 2328 -1536 2392
rect -1632 2312 -1536 2328
rect -1632 2248 -1616 2312
rect -1552 2248 -1536 2312
rect -1632 2232 -1536 2248
rect -1632 2168 -1616 2232
rect -1552 2168 -1536 2232
rect -1632 2152 -1536 2168
rect -1632 2088 -1616 2152
rect -1552 2088 -1536 2152
rect -1632 2072 -1536 2088
rect -1632 2008 -1616 2072
rect -1552 2008 -1536 2072
rect -1632 1992 -1536 2008
rect -1632 1928 -1616 1992
rect -1552 1928 -1536 1992
rect -1632 1912 -1536 1928
rect -3044 1812 -2948 1848
rect -1632 1848 -1616 1912
rect -1552 1848 -1536 1912
rect -1213 2592 -491 2601
rect -1213 1888 -1204 2592
rect -500 1888 -491 2592
rect -1213 1879 -491 1888
rect -220 2568 -204 2632
rect -140 2568 -124 2632
rect 1192 2632 1288 2668
rect -220 2552 -124 2568
rect -220 2488 -204 2552
rect -140 2488 -124 2552
rect -220 2472 -124 2488
rect -220 2408 -204 2472
rect -140 2408 -124 2472
rect -220 2392 -124 2408
rect -220 2328 -204 2392
rect -140 2328 -124 2392
rect -220 2312 -124 2328
rect -220 2248 -204 2312
rect -140 2248 -124 2312
rect -220 2232 -124 2248
rect -220 2168 -204 2232
rect -140 2168 -124 2232
rect -220 2152 -124 2168
rect -220 2088 -204 2152
rect -140 2088 -124 2152
rect -220 2072 -124 2088
rect -220 2008 -204 2072
rect -140 2008 -124 2072
rect -220 1992 -124 2008
rect -220 1928 -204 1992
rect -140 1928 -124 1992
rect -220 1912 -124 1928
rect -1632 1812 -1536 1848
rect -220 1848 -204 1912
rect -140 1848 -124 1912
rect 199 2592 921 2601
rect 199 1888 208 2592
rect 912 1888 921 2592
rect 199 1879 921 1888
rect 1192 2568 1208 2632
rect 1272 2568 1288 2632
rect 2604 2632 2700 2668
rect 1192 2552 1288 2568
rect 1192 2488 1208 2552
rect 1272 2488 1288 2552
rect 1192 2472 1288 2488
rect 1192 2408 1208 2472
rect 1272 2408 1288 2472
rect 1192 2392 1288 2408
rect 1192 2328 1208 2392
rect 1272 2328 1288 2392
rect 1192 2312 1288 2328
rect 1192 2248 1208 2312
rect 1272 2248 1288 2312
rect 1192 2232 1288 2248
rect 1192 2168 1208 2232
rect 1272 2168 1288 2232
rect 1192 2152 1288 2168
rect 1192 2088 1208 2152
rect 1272 2088 1288 2152
rect 1192 2072 1288 2088
rect 1192 2008 1208 2072
rect 1272 2008 1288 2072
rect 1192 1992 1288 2008
rect 1192 1928 1208 1992
rect 1272 1928 1288 1992
rect 1192 1912 1288 1928
rect -220 1812 -124 1848
rect 1192 1848 1208 1912
rect 1272 1848 1288 1912
rect 1611 2592 2333 2601
rect 1611 1888 1620 2592
rect 2324 1888 2333 2592
rect 1611 1879 2333 1888
rect 2604 2568 2620 2632
rect 2684 2568 2700 2632
rect 4016 2632 4112 2668
rect 2604 2552 2700 2568
rect 2604 2488 2620 2552
rect 2684 2488 2700 2552
rect 2604 2472 2700 2488
rect 2604 2408 2620 2472
rect 2684 2408 2700 2472
rect 2604 2392 2700 2408
rect 2604 2328 2620 2392
rect 2684 2328 2700 2392
rect 2604 2312 2700 2328
rect 2604 2248 2620 2312
rect 2684 2248 2700 2312
rect 2604 2232 2700 2248
rect 2604 2168 2620 2232
rect 2684 2168 2700 2232
rect 2604 2152 2700 2168
rect 2604 2088 2620 2152
rect 2684 2088 2700 2152
rect 2604 2072 2700 2088
rect 2604 2008 2620 2072
rect 2684 2008 2700 2072
rect 2604 1992 2700 2008
rect 2604 1928 2620 1992
rect 2684 1928 2700 1992
rect 2604 1912 2700 1928
rect 1192 1812 1288 1848
rect 2604 1848 2620 1912
rect 2684 1848 2700 1912
rect 3023 2592 3745 2601
rect 3023 1888 3032 2592
rect 3736 1888 3745 2592
rect 3023 1879 3745 1888
rect 4016 2568 4032 2632
rect 4096 2568 4112 2632
rect 5428 2632 5524 2668
rect 4016 2552 4112 2568
rect 4016 2488 4032 2552
rect 4096 2488 4112 2552
rect 4016 2472 4112 2488
rect 4016 2408 4032 2472
rect 4096 2408 4112 2472
rect 4016 2392 4112 2408
rect 4016 2328 4032 2392
rect 4096 2328 4112 2392
rect 4016 2312 4112 2328
rect 4016 2248 4032 2312
rect 4096 2248 4112 2312
rect 4016 2232 4112 2248
rect 4016 2168 4032 2232
rect 4096 2168 4112 2232
rect 4016 2152 4112 2168
rect 4016 2088 4032 2152
rect 4096 2088 4112 2152
rect 4016 2072 4112 2088
rect 4016 2008 4032 2072
rect 4096 2008 4112 2072
rect 4016 1992 4112 2008
rect 4016 1928 4032 1992
rect 4096 1928 4112 1992
rect 4016 1912 4112 1928
rect 2604 1812 2700 1848
rect 4016 1848 4032 1912
rect 4096 1848 4112 1912
rect 4435 2592 5157 2601
rect 4435 1888 4444 2592
rect 5148 1888 5157 2592
rect 4435 1879 5157 1888
rect 5428 2568 5444 2632
rect 5508 2568 5524 2632
rect 6840 2632 6936 2668
rect 5428 2552 5524 2568
rect 5428 2488 5444 2552
rect 5508 2488 5524 2552
rect 5428 2472 5524 2488
rect 5428 2408 5444 2472
rect 5508 2408 5524 2472
rect 5428 2392 5524 2408
rect 5428 2328 5444 2392
rect 5508 2328 5524 2392
rect 5428 2312 5524 2328
rect 5428 2248 5444 2312
rect 5508 2248 5524 2312
rect 5428 2232 5524 2248
rect 5428 2168 5444 2232
rect 5508 2168 5524 2232
rect 5428 2152 5524 2168
rect 5428 2088 5444 2152
rect 5508 2088 5524 2152
rect 5428 2072 5524 2088
rect 5428 2008 5444 2072
rect 5508 2008 5524 2072
rect 5428 1992 5524 2008
rect 5428 1928 5444 1992
rect 5508 1928 5524 1992
rect 5428 1912 5524 1928
rect 4016 1812 4112 1848
rect 5428 1848 5444 1912
rect 5508 1848 5524 1912
rect 5847 2592 6569 2601
rect 5847 1888 5856 2592
rect 6560 1888 6569 2592
rect 5847 1879 6569 1888
rect 6840 2568 6856 2632
rect 6920 2568 6936 2632
rect 8252 2632 8348 2668
rect 6840 2552 6936 2568
rect 6840 2488 6856 2552
rect 6920 2488 6936 2552
rect 6840 2472 6936 2488
rect 6840 2408 6856 2472
rect 6920 2408 6936 2472
rect 6840 2392 6936 2408
rect 6840 2328 6856 2392
rect 6920 2328 6936 2392
rect 6840 2312 6936 2328
rect 6840 2248 6856 2312
rect 6920 2248 6936 2312
rect 6840 2232 6936 2248
rect 6840 2168 6856 2232
rect 6920 2168 6936 2232
rect 6840 2152 6936 2168
rect 6840 2088 6856 2152
rect 6920 2088 6936 2152
rect 6840 2072 6936 2088
rect 6840 2008 6856 2072
rect 6920 2008 6936 2072
rect 6840 1992 6936 2008
rect 6840 1928 6856 1992
rect 6920 1928 6936 1992
rect 6840 1912 6936 1928
rect 5428 1812 5524 1848
rect 6840 1848 6856 1912
rect 6920 1848 6936 1912
rect 7259 2592 7981 2601
rect 7259 1888 7268 2592
rect 7972 1888 7981 2592
rect 7259 1879 7981 1888
rect 8252 2568 8268 2632
rect 8332 2568 8348 2632
rect 9664 2632 9760 2668
rect 8252 2552 8348 2568
rect 8252 2488 8268 2552
rect 8332 2488 8348 2552
rect 8252 2472 8348 2488
rect 8252 2408 8268 2472
rect 8332 2408 8348 2472
rect 8252 2392 8348 2408
rect 8252 2328 8268 2392
rect 8332 2328 8348 2392
rect 8252 2312 8348 2328
rect 8252 2248 8268 2312
rect 8332 2248 8348 2312
rect 8252 2232 8348 2248
rect 8252 2168 8268 2232
rect 8332 2168 8348 2232
rect 8252 2152 8348 2168
rect 8252 2088 8268 2152
rect 8332 2088 8348 2152
rect 8252 2072 8348 2088
rect 8252 2008 8268 2072
rect 8332 2008 8348 2072
rect 8252 1992 8348 2008
rect 8252 1928 8268 1992
rect 8332 1928 8348 1992
rect 8252 1912 8348 1928
rect 6840 1812 6936 1848
rect 8252 1848 8268 1912
rect 8332 1848 8348 1912
rect 8671 2592 9393 2601
rect 8671 1888 8680 2592
rect 9384 1888 9393 2592
rect 8671 1879 9393 1888
rect 9664 2568 9680 2632
rect 9744 2568 9760 2632
rect 11076 2632 11172 2668
rect 9664 2552 9760 2568
rect 9664 2488 9680 2552
rect 9744 2488 9760 2552
rect 9664 2472 9760 2488
rect 9664 2408 9680 2472
rect 9744 2408 9760 2472
rect 9664 2392 9760 2408
rect 9664 2328 9680 2392
rect 9744 2328 9760 2392
rect 9664 2312 9760 2328
rect 9664 2248 9680 2312
rect 9744 2248 9760 2312
rect 9664 2232 9760 2248
rect 9664 2168 9680 2232
rect 9744 2168 9760 2232
rect 9664 2152 9760 2168
rect 9664 2088 9680 2152
rect 9744 2088 9760 2152
rect 9664 2072 9760 2088
rect 9664 2008 9680 2072
rect 9744 2008 9760 2072
rect 9664 1992 9760 2008
rect 9664 1928 9680 1992
rect 9744 1928 9760 1992
rect 9664 1912 9760 1928
rect 8252 1812 8348 1848
rect 9664 1848 9680 1912
rect 9744 1848 9760 1912
rect 10083 2592 10805 2601
rect 10083 1888 10092 2592
rect 10796 1888 10805 2592
rect 10083 1879 10805 1888
rect 11076 2568 11092 2632
rect 11156 2568 11172 2632
rect 12488 2632 12584 2668
rect 11076 2552 11172 2568
rect 11076 2488 11092 2552
rect 11156 2488 11172 2552
rect 11076 2472 11172 2488
rect 11076 2408 11092 2472
rect 11156 2408 11172 2472
rect 11076 2392 11172 2408
rect 11076 2328 11092 2392
rect 11156 2328 11172 2392
rect 11076 2312 11172 2328
rect 11076 2248 11092 2312
rect 11156 2248 11172 2312
rect 11076 2232 11172 2248
rect 11076 2168 11092 2232
rect 11156 2168 11172 2232
rect 11076 2152 11172 2168
rect 11076 2088 11092 2152
rect 11156 2088 11172 2152
rect 11076 2072 11172 2088
rect 11076 2008 11092 2072
rect 11156 2008 11172 2072
rect 11076 1992 11172 2008
rect 11076 1928 11092 1992
rect 11156 1928 11172 1992
rect 11076 1912 11172 1928
rect 9664 1812 9760 1848
rect 11076 1848 11092 1912
rect 11156 1848 11172 1912
rect 11495 2592 12217 2601
rect 11495 1888 11504 2592
rect 12208 1888 12217 2592
rect 11495 1879 12217 1888
rect 12488 2568 12504 2632
rect 12568 2568 12584 2632
rect 13900 2632 13996 2668
rect 12488 2552 12584 2568
rect 12488 2488 12504 2552
rect 12568 2488 12584 2552
rect 12488 2472 12584 2488
rect 12488 2408 12504 2472
rect 12568 2408 12584 2472
rect 12488 2392 12584 2408
rect 12488 2328 12504 2392
rect 12568 2328 12584 2392
rect 12488 2312 12584 2328
rect 12488 2248 12504 2312
rect 12568 2248 12584 2312
rect 12488 2232 12584 2248
rect 12488 2168 12504 2232
rect 12568 2168 12584 2232
rect 12488 2152 12584 2168
rect 12488 2088 12504 2152
rect 12568 2088 12584 2152
rect 12488 2072 12584 2088
rect 12488 2008 12504 2072
rect 12568 2008 12584 2072
rect 12488 1992 12584 2008
rect 12488 1928 12504 1992
rect 12568 1928 12584 1992
rect 12488 1912 12584 1928
rect 11076 1812 11172 1848
rect 12488 1848 12504 1912
rect 12568 1848 12584 1912
rect 12907 2592 13629 2601
rect 12907 1888 12916 2592
rect 13620 1888 13629 2592
rect 12907 1879 13629 1888
rect 13900 2568 13916 2632
rect 13980 2568 13996 2632
rect 15312 2632 15408 2668
rect 13900 2552 13996 2568
rect 13900 2488 13916 2552
rect 13980 2488 13996 2552
rect 13900 2472 13996 2488
rect 13900 2408 13916 2472
rect 13980 2408 13996 2472
rect 13900 2392 13996 2408
rect 13900 2328 13916 2392
rect 13980 2328 13996 2392
rect 13900 2312 13996 2328
rect 13900 2248 13916 2312
rect 13980 2248 13996 2312
rect 13900 2232 13996 2248
rect 13900 2168 13916 2232
rect 13980 2168 13996 2232
rect 13900 2152 13996 2168
rect 13900 2088 13916 2152
rect 13980 2088 13996 2152
rect 13900 2072 13996 2088
rect 13900 2008 13916 2072
rect 13980 2008 13996 2072
rect 13900 1992 13996 2008
rect 13900 1928 13916 1992
rect 13980 1928 13996 1992
rect 13900 1912 13996 1928
rect 12488 1812 12584 1848
rect 13900 1848 13916 1912
rect 13980 1848 13996 1912
rect 14319 2592 15041 2601
rect 14319 1888 14328 2592
rect 15032 1888 15041 2592
rect 14319 1879 15041 1888
rect 15312 2568 15328 2632
rect 15392 2568 15408 2632
rect 16724 2632 16820 2668
rect 15312 2552 15408 2568
rect 15312 2488 15328 2552
rect 15392 2488 15408 2552
rect 15312 2472 15408 2488
rect 15312 2408 15328 2472
rect 15392 2408 15408 2472
rect 15312 2392 15408 2408
rect 15312 2328 15328 2392
rect 15392 2328 15408 2392
rect 15312 2312 15408 2328
rect 15312 2248 15328 2312
rect 15392 2248 15408 2312
rect 15312 2232 15408 2248
rect 15312 2168 15328 2232
rect 15392 2168 15408 2232
rect 15312 2152 15408 2168
rect 15312 2088 15328 2152
rect 15392 2088 15408 2152
rect 15312 2072 15408 2088
rect 15312 2008 15328 2072
rect 15392 2008 15408 2072
rect 15312 1992 15408 2008
rect 15312 1928 15328 1992
rect 15392 1928 15408 1992
rect 15312 1912 15408 1928
rect 13900 1812 13996 1848
rect 15312 1848 15328 1912
rect 15392 1848 15408 1912
rect 15731 2592 16453 2601
rect 15731 1888 15740 2592
rect 16444 1888 16453 2592
rect 15731 1879 16453 1888
rect 16724 2568 16740 2632
rect 16804 2568 16820 2632
rect 18136 2632 18232 2668
rect 16724 2552 16820 2568
rect 16724 2488 16740 2552
rect 16804 2488 16820 2552
rect 16724 2472 16820 2488
rect 16724 2408 16740 2472
rect 16804 2408 16820 2472
rect 16724 2392 16820 2408
rect 16724 2328 16740 2392
rect 16804 2328 16820 2392
rect 16724 2312 16820 2328
rect 16724 2248 16740 2312
rect 16804 2248 16820 2312
rect 16724 2232 16820 2248
rect 16724 2168 16740 2232
rect 16804 2168 16820 2232
rect 16724 2152 16820 2168
rect 16724 2088 16740 2152
rect 16804 2088 16820 2152
rect 16724 2072 16820 2088
rect 16724 2008 16740 2072
rect 16804 2008 16820 2072
rect 16724 1992 16820 2008
rect 16724 1928 16740 1992
rect 16804 1928 16820 1992
rect 16724 1912 16820 1928
rect 15312 1812 15408 1848
rect 16724 1848 16740 1912
rect 16804 1848 16820 1912
rect 17143 2592 17865 2601
rect 17143 1888 17152 2592
rect 17856 1888 17865 2592
rect 17143 1879 17865 1888
rect 18136 2568 18152 2632
rect 18216 2568 18232 2632
rect 19548 2632 19644 2668
rect 18136 2552 18232 2568
rect 18136 2488 18152 2552
rect 18216 2488 18232 2552
rect 18136 2472 18232 2488
rect 18136 2408 18152 2472
rect 18216 2408 18232 2472
rect 18136 2392 18232 2408
rect 18136 2328 18152 2392
rect 18216 2328 18232 2392
rect 18136 2312 18232 2328
rect 18136 2248 18152 2312
rect 18216 2248 18232 2312
rect 18136 2232 18232 2248
rect 18136 2168 18152 2232
rect 18216 2168 18232 2232
rect 18136 2152 18232 2168
rect 18136 2088 18152 2152
rect 18216 2088 18232 2152
rect 18136 2072 18232 2088
rect 18136 2008 18152 2072
rect 18216 2008 18232 2072
rect 18136 1992 18232 2008
rect 18136 1928 18152 1992
rect 18216 1928 18232 1992
rect 18136 1912 18232 1928
rect 16724 1812 16820 1848
rect 18136 1848 18152 1912
rect 18216 1848 18232 1912
rect 18555 2592 19277 2601
rect 18555 1888 18564 2592
rect 19268 1888 19277 2592
rect 18555 1879 19277 1888
rect 19548 2568 19564 2632
rect 19628 2568 19644 2632
rect 20960 2632 21056 2668
rect 19548 2552 19644 2568
rect 19548 2488 19564 2552
rect 19628 2488 19644 2552
rect 19548 2472 19644 2488
rect 19548 2408 19564 2472
rect 19628 2408 19644 2472
rect 19548 2392 19644 2408
rect 19548 2328 19564 2392
rect 19628 2328 19644 2392
rect 19548 2312 19644 2328
rect 19548 2248 19564 2312
rect 19628 2248 19644 2312
rect 19548 2232 19644 2248
rect 19548 2168 19564 2232
rect 19628 2168 19644 2232
rect 19548 2152 19644 2168
rect 19548 2088 19564 2152
rect 19628 2088 19644 2152
rect 19548 2072 19644 2088
rect 19548 2008 19564 2072
rect 19628 2008 19644 2072
rect 19548 1992 19644 2008
rect 19548 1928 19564 1992
rect 19628 1928 19644 1992
rect 19548 1912 19644 1928
rect 18136 1812 18232 1848
rect 19548 1848 19564 1912
rect 19628 1848 19644 1912
rect 19967 2592 20689 2601
rect 19967 1888 19976 2592
rect 20680 1888 20689 2592
rect 19967 1879 20689 1888
rect 20960 2568 20976 2632
rect 21040 2568 21056 2632
rect 22372 2632 22468 2668
rect 20960 2552 21056 2568
rect 20960 2488 20976 2552
rect 21040 2488 21056 2552
rect 20960 2472 21056 2488
rect 20960 2408 20976 2472
rect 21040 2408 21056 2472
rect 20960 2392 21056 2408
rect 20960 2328 20976 2392
rect 21040 2328 21056 2392
rect 20960 2312 21056 2328
rect 20960 2248 20976 2312
rect 21040 2248 21056 2312
rect 20960 2232 21056 2248
rect 20960 2168 20976 2232
rect 21040 2168 21056 2232
rect 20960 2152 21056 2168
rect 20960 2088 20976 2152
rect 21040 2088 21056 2152
rect 20960 2072 21056 2088
rect 20960 2008 20976 2072
rect 21040 2008 21056 2072
rect 20960 1992 21056 2008
rect 20960 1928 20976 1992
rect 21040 1928 21056 1992
rect 20960 1912 21056 1928
rect 19548 1812 19644 1848
rect 20960 1848 20976 1912
rect 21040 1848 21056 1912
rect 21379 2592 22101 2601
rect 21379 1888 21388 2592
rect 22092 1888 22101 2592
rect 21379 1879 22101 1888
rect 22372 2568 22388 2632
rect 22452 2568 22468 2632
rect 23784 2632 23880 2668
rect 22372 2552 22468 2568
rect 22372 2488 22388 2552
rect 22452 2488 22468 2552
rect 22372 2472 22468 2488
rect 22372 2408 22388 2472
rect 22452 2408 22468 2472
rect 22372 2392 22468 2408
rect 22372 2328 22388 2392
rect 22452 2328 22468 2392
rect 22372 2312 22468 2328
rect 22372 2248 22388 2312
rect 22452 2248 22468 2312
rect 22372 2232 22468 2248
rect 22372 2168 22388 2232
rect 22452 2168 22468 2232
rect 22372 2152 22468 2168
rect 22372 2088 22388 2152
rect 22452 2088 22468 2152
rect 22372 2072 22468 2088
rect 22372 2008 22388 2072
rect 22452 2008 22468 2072
rect 22372 1992 22468 2008
rect 22372 1928 22388 1992
rect 22452 1928 22468 1992
rect 22372 1912 22468 1928
rect 20960 1812 21056 1848
rect 22372 1848 22388 1912
rect 22452 1848 22468 1912
rect 22791 2592 23513 2601
rect 22791 1888 22800 2592
rect 23504 1888 23513 2592
rect 22791 1879 23513 1888
rect 23784 2568 23800 2632
rect 23864 2568 23880 2632
rect 23784 2552 23880 2568
rect 23784 2488 23800 2552
rect 23864 2488 23880 2552
rect 23784 2472 23880 2488
rect 23784 2408 23800 2472
rect 23864 2408 23880 2472
rect 23784 2392 23880 2408
rect 23784 2328 23800 2392
rect 23864 2328 23880 2392
rect 23784 2312 23880 2328
rect 23784 2248 23800 2312
rect 23864 2248 23880 2312
rect 23784 2232 23880 2248
rect 23784 2168 23800 2232
rect 23864 2168 23880 2232
rect 23784 2152 23880 2168
rect 23784 2088 23800 2152
rect 23864 2088 23880 2152
rect 23784 2072 23880 2088
rect 23784 2008 23800 2072
rect 23864 2008 23880 2072
rect 23784 1992 23880 2008
rect 23784 1928 23800 1992
rect 23864 1928 23880 1992
rect 23784 1912 23880 1928
rect 22372 1812 22468 1848
rect 23784 1848 23800 1912
rect 23864 1848 23880 1912
rect 23784 1812 23880 1848
rect -22812 1512 -22716 1548
rect -23805 1472 -23083 1481
rect -23805 768 -23796 1472
rect -23092 768 -23083 1472
rect -23805 759 -23083 768
rect -22812 1448 -22796 1512
rect -22732 1448 -22716 1512
rect -21400 1512 -21304 1548
rect -22812 1432 -22716 1448
rect -22812 1368 -22796 1432
rect -22732 1368 -22716 1432
rect -22812 1352 -22716 1368
rect -22812 1288 -22796 1352
rect -22732 1288 -22716 1352
rect -22812 1272 -22716 1288
rect -22812 1208 -22796 1272
rect -22732 1208 -22716 1272
rect -22812 1192 -22716 1208
rect -22812 1128 -22796 1192
rect -22732 1128 -22716 1192
rect -22812 1112 -22716 1128
rect -22812 1048 -22796 1112
rect -22732 1048 -22716 1112
rect -22812 1032 -22716 1048
rect -22812 968 -22796 1032
rect -22732 968 -22716 1032
rect -22812 952 -22716 968
rect -22812 888 -22796 952
rect -22732 888 -22716 952
rect -22812 872 -22716 888
rect -22812 808 -22796 872
rect -22732 808 -22716 872
rect -22812 792 -22716 808
rect -22812 728 -22796 792
rect -22732 728 -22716 792
rect -22393 1472 -21671 1481
rect -22393 768 -22384 1472
rect -21680 768 -21671 1472
rect -22393 759 -21671 768
rect -21400 1448 -21384 1512
rect -21320 1448 -21304 1512
rect -19988 1512 -19892 1548
rect -21400 1432 -21304 1448
rect -21400 1368 -21384 1432
rect -21320 1368 -21304 1432
rect -21400 1352 -21304 1368
rect -21400 1288 -21384 1352
rect -21320 1288 -21304 1352
rect -21400 1272 -21304 1288
rect -21400 1208 -21384 1272
rect -21320 1208 -21304 1272
rect -21400 1192 -21304 1208
rect -21400 1128 -21384 1192
rect -21320 1128 -21304 1192
rect -21400 1112 -21304 1128
rect -21400 1048 -21384 1112
rect -21320 1048 -21304 1112
rect -21400 1032 -21304 1048
rect -21400 968 -21384 1032
rect -21320 968 -21304 1032
rect -21400 952 -21304 968
rect -21400 888 -21384 952
rect -21320 888 -21304 952
rect -21400 872 -21304 888
rect -21400 808 -21384 872
rect -21320 808 -21304 872
rect -21400 792 -21304 808
rect -22812 692 -22716 728
rect -21400 728 -21384 792
rect -21320 728 -21304 792
rect -20981 1472 -20259 1481
rect -20981 768 -20972 1472
rect -20268 768 -20259 1472
rect -20981 759 -20259 768
rect -19988 1448 -19972 1512
rect -19908 1448 -19892 1512
rect -18576 1512 -18480 1548
rect -19988 1432 -19892 1448
rect -19988 1368 -19972 1432
rect -19908 1368 -19892 1432
rect -19988 1352 -19892 1368
rect -19988 1288 -19972 1352
rect -19908 1288 -19892 1352
rect -19988 1272 -19892 1288
rect -19988 1208 -19972 1272
rect -19908 1208 -19892 1272
rect -19988 1192 -19892 1208
rect -19988 1128 -19972 1192
rect -19908 1128 -19892 1192
rect -19988 1112 -19892 1128
rect -19988 1048 -19972 1112
rect -19908 1048 -19892 1112
rect -19988 1032 -19892 1048
rect -19988 968 -19972 1032
rect -19908 968 -19892 1032
rect -19988 952 -19892 968
rect -19988 888 -19972 952
rect -19908 888 -19892 952
rect -19988 872 -19892 888
rect -19988 808 -19972 872
rect -19908 808 -19892 872
rect -19988 792 -19892 808
rect -21400 692 -21304 728
rect -19988 728 -19972 792
rect -19908 728 -19892 792
rect -19569 1472 -18847 1481
rect -19569 768 -19560 1472
rect -18856 768 -18847 1472
rect -19569 759 -18847 768
rect -18576 1448 -18560 1512
rect -18496 1448 -18480 1512
rect -17164 1512 -17068 1548
rect -18576 1432 -18480 1448
rect -18576 1368 -18560 1432
rect -18496 1368 -18480 1432
rect -18576 1352 -18480 1368
rect -18576 1288 -18560 1352
rect -18496 1288 -18480 1352
rect -18576 1272 -18480 1288
rect -18576 1208 -18560 1272
rect -18496 1208 -18480 1272
rect -18576 1192 -18480 1208
rect -18576 1128 -18560 1192
rect -18496 1128 -18480 1192
rect -18576 1112 -18480 1128
rect -18576 1048 -18560 1112
rect -18496 1048 -18480 1112
rect -18576 1032 -18480 1048
rect -18576 968 -18560 1032
rect -18496 968 -18480 1032
rect -18576 952 -18480 968
rect -18576 888 -18560 952
rect -18496 888 -18480 952
rect -18576 872 -18480 888
rect -18576 808 -18560 872
rect -18496 808 -18480 872
rect -18576 792 -18480 808
rect -19988 692 -19892 728
rect -18576 728 -18560 792
rect -18496 728 -18480 792
rect -18157 1472 -17435 1481
rect -18157 768 -18148 1472
rect -17444 768 -17435 1472
rect -18157 759 -17435 768
rect -17164 1448 -17148 1512
rect -17084 1448 -17068 1512
rect -15752 1512 -15656 1548
rect -17164 1432 -17068 1448
rect -17164 1368 -17148 1432
rect -17084 1368 -17068 1432
rect -17164 1352 -17068 1368
rect -17164 1288 -17148 1352
rect -17084 1288 -17068 1352
rect -17164 1272 -17068 1288
rect -17164 1208 -17148 1272
rect -17084 1208 -17068 1272
rect -17164 1192 -17068 1208
rect -17164 1128 -17148 1192
rect -17084 1128 -17068 1192
rect -17164 1112 -17068 1128
rect -17164 1048 -17148 1112
rect -17084 1048 -17068 1112
rect -17164 1032 -17068 1048
rect -17164 968 -17148 1032
rect -17084 968 -17068 1032
rect -17164 952 -17068 968
rect -17164 888 -17148 952
rect -17084 888 -17068 952
rect -17164 872 -17068 888
rect -17164 808 -17148 872
rect -17084 808 -17068 872
rect -17164 792 -17068 808
rect -18576 692 -18480 728
rect -17164 728 -17148 792
rect -17084 728 -17068 792
rect -16745 1472 -16023 1481
rect -16745 768 -16736 1472
rect -16032 768 -16023 1472
rect -16745 759 -16023 768
rect -15752 1448 -15736 1512
rect -15672 1448 -15656 1512
rect -14340 1512 -14244 1548
rect -15752 1432 -15656 1448
rect -15752 1368 -15736 1432
rect -15672 1368 -15656 1432
rect -15752 1352 -15656 1368
rect -15752 1288 -15736 1352
rect -15672 1288 -15656 1352
rect -15752 1272 -15656 1288
rect -15752 1208 -15736 1272
rect -15672 1208 -15656 1272
rect -15752 1192 -15656 1208
rect -15752 1128 -15736 1192
rect -15672 1128 -15656 1192
rect -15752 1112 -15656 1128
rect -15752 1048 -15736 1112
rect -15672 1048 -15656 1112
rect -15752 1032 -15656 1048
rect -15752 968 -15736 1032
rect -15672 968 -15656 1032
rect -15752 952 -15656 968
rect -15752 888 -15736 952
rect -15672 888 -15656 952
rect -15752 872 -15656 888
rect -15752 808 -15736 872
rect -15672 808 -15656 872
rect -15752 792 -15656 808
rect -17164 692 -17068 728
rect -15752 728 -15736 792
rect -15672 728 -15656 792
rect -15333 1472 -14611 1481
rect -15333 768 -15324 1472
rect -14620 768 -14611 1472
rect -15333 759 -14611 768
rect -14340 1448 -14324 1512
rect -14260 1448 -14244 1512
rect -12928 1512 -12832 1548
rect -14340 1432 -14244 1448
rect -14340 1368 -14324 1432
rect -14260 1368 -14244 1432
rect -14340 1352 -14244 1368
rect -14340 1288 -14324 1352
rect -14260 1288 -14244 1352
rect -14340 1272 -14244 1288
rect -14340 1208 -14324 1272
rect -14260 1208 -14244 1272
rect -14340 1192 -14244 1208
rect -14340 1128 -14324 1192
rect -14260 1128 -14244 1192
rect -14340 1112 -14244 1128
rect -14340 1048 -14324 1112
rect -14260 1048 -14244 1112
rect -14340 1032 -14244 1048
rect -14340 968 -14324 1032
rect -14260 968 -14244 1032
rect -14340 952 -14244 968
rect -14340 888 -14324 952
rect -14260 888 -14244 952
rect -14340 872 -14244 888
rect -14340 808 -14324 872
rect -14260 808 -14244 872
rect -14340 792 -14244 808
rect -15752 692 -15656 728
rect -14340 728 -14324 792
rect -14260 728 -14244 792
rect -13921 1472 -13199 1481
rect -13921 768 -13912 1472
rect -13208 768 -13199 1472
rect -13921 759 -13199 768
rect -12928 1448 -12912 1512
rect -12848 1448 -12832 1512
rect -11516 1512 -11420 1548
rect -12928 1432 -12832 1448
rect -12928 1368 -12912 1432
rect -12848 1368 -12832 1432
rect -12928 1352 -12832 1368
rect -12928 1288 -12912 1352
rect -12848 1288 -12832 1352
rect -12928 1272 -12832 1288
rect -12928 1208 -12912 1272
rect -12848 1208 -12832 1272
rect -12928 1192 -12832 1208
rect -12928 1128 -12912 1192
rect -12848 1128 -12832 1192
rect -12928 1112 -12832 1128
rect -12928 1048 -12912 1112
rect -12848 1048 -12832 1112
rect -12928 1032 -12832 1048
rect -12928 968 -12912 1032
rect -12848 968 -12832 1032
rect -12928 952 -12832 968
rect -12928 888 -12912 952
rect -12848 888 -12832 952
rect -12928 872 -12832 888
rect -12928 808 -12912 872
rect -12848 808 -12832 872
rect -12928 792 -12832 808
rect -14340 692 -14244 728
rect -12928 728 -12912 792
rect -12848 728 -12832 792
rect -12509 1472 -11787 1481
rect -12509 768 -12500 1472
rect -11796 768 -11787 1472
rect -12509 759 -11787 768
rect -11516 1448 -11500 1512
rect -11436 1448 -11420 1512
rect -10104 1512 -10008 1548
rect -11516 1432 -11420 1448
rect -11516 1368 -11500 1432
rect -11436 1368 -11420 1432
rect -11516 1352 -11420 1368
rect -11516 1288 -11500 1352
rect -11436 1288 -11420 1352
rect -11516 1272 -11420 1288
rect -11516 1208 -11500 1272
rect -11436 1208 -11420 1272
rect -11516 1192 -11420 1208
rect -11516 1128 -11500 1192
rect -11436 1128 -11420 1192
rect -11516 1112 -11420 1128
rect -11516 1048 -11500 1112
rect -11436 1048 -11420 1112
rect -11516 1032 -11420 1048
rect -11516 968 -11500 1032
rect -11436 968 -11420 1032
rect -11516 952 -11420 968
rect -11516 888 -11500 952
rect -11436 888 -11420 952
rect -11516 872 -11420 888
rect -11516 808 -11500 872
rect -11436 808 -11420 872
rect -11516 792 -11420 808
rect -12928 692 -12832 728
rect -11516 728 -11500 792
rect -11436 728 -11420 792
rect -11097 1472 -10375 1481
rect -11097 768 -11088 1472
rect -10384 768 -10375 1472
rect -11097 759 -10375 768
rect -10104 1448 -10088 1512
rect -10024 1448 -10008 1512
rect -8692 1512 -8596 1548
rect -10104 1432 -10008 1448
rect -10104 1368 -10088 1432
rect -10024 1368 -10008 1432
rect -10104 1352 -10008 1368
rect -10104 1288 -10088 1352
rect -10024 1288 -10008 1352
rect -10104 1272 -10008 1288
rect -10104 1208 -10088 1272
rect -10024 1208 -10008 1272
rect -10104 1192 -10008 1208
rect -10104 1128 -10088 1192
rect -10024 1128 -10008 1192
rect -10104 1112 -10008 1128
rect -10104 1048 -10088 1112
rect -10024 1048 -10008 1112
rect -10104 1032 -10008 1048
rect -10104 968 -10088 1032
rect -10024 968 -10008 1032
rect -10104 952 -10008 968
rect -10104 888 -10088 952
rect -10024 888 -10008 952
rect -10104 872 -10008 888
rect -10104 808 -10088 872
rect -10024 808 -10008 872
rect -10104 792 -10008 808
rect -11516 692 -11420 728
rect -10104 728 -10088 792
rect -10024 728 -10008 792
rect -9685 1472 -8963 1481
rect -9685 768 -9676 1472
rect -8972 768 -8963 1472
rect -9685 759 -8963 768
rect -8692 1448 -8676 1512
rect -8612 1448 -8596 1512
rect -7280 1512 -7184 1548
rect -8692 1432 -8596 1448
rect -8692 1368 -8676 1432
rect -8612 1368 -8596 1432
rect -8692 1352 -8596 1368
rect -8692 1288 -8676 1352
rect -8612 1288 -8596 1352
rect -8692 1272 -8596 1288
rect -8692 1208 -8676 1272
rect -8612 1208 -8596 1272
rect -8692 1192 -8596 1208
rect -8692 1128 -8676 1192
rect -8612 1128 -8596 1192
rect -8692 1112 -8596 1128
rect -8692 1048 -8676 1112
rect -8612 1048 -8596 1112
rect -8692 1032 -8596 1048
rect -8692 968 -8676 1032
rect -8612 968 -8596 1032
rect -8692 952 -8596 968
rect -8692 888 -8676 952
rect -8612 888 -8596 952
rect -8692 872 -8596 888
rect -8692 808 -8676 872
rect -8612 808 -8596 872
rect -8692 792 -8596 808
rect -10104 692 -10008 728
rect -8692 728 -8676 792
rect -8612 728 -8596 792
rect -8273 1472 -7551 1481
rect -8273 768 -8264 1472
rect -7560 768 -7551 1472
rect -8273 759 -7551 768
rect -7280 1448 -7264 1512
rect -7200 1448 -7184 1512
rect -5868 1512 -5772 1548
rect -7280 1432 -7184 1448
rect -7280 1368 -7264 1432
rect -7200 1368 -7184 1432
rect -7280 1352 -7184 1368
rect -7280 1288 -7264 1352
rect -7200 1288 -7184 1352
rect -7280 1272 -7184 1288
rect -7280 1208 -7264 1272
rect -7200 1208 -7184 1272
rect -7280 1192 -7184 1208
rect -7280 1128 -7264 1192
rect -7200 1128 -7184 1192
rect -7280 1112 -7184 1128
rect -7280 1048 -7264 1112
rect -7200 1048 -7184 1112
rect -7280 1032 -7184 1048
rect -7280 968 -7264 1032
rect -7200 968 -7184 1032
rect -7280 952 -7184 968
rect -7280 888 -7264 952
rect -7200 888 -7184 952
rect -7280 872 -7184 888
rect -7280 808 -7264 872
rect -7200 808 -7184 872
rect -7280 792 -7184 808
rect -8692 692 -8596 728
rect -7280 728 -7264 792
rect -7200 728 -7184 792
rect -6861 1472 -6139 1481
rect -6861 768 -6852 1472
rect -6148 768 -6139 1472
rect -6861 759 -6139 768
rect -5868 1448 -5852 1512
rect -5788 1448 -5772 1512
rect -4456 1512 -4360 1548
rect -5868 1432 -5772 1448
rect -5868 1368 -5852 1432
rect -5788 1368 -5772 1432
rect -5868 1352 -5772 1368
rect -5868 1288 -5852 1352
rect -5788 1288 -5772 1352
rect -5868 1272 -5772 1288
rect -5868 1208 -5852 1272
rect -5788 1208 -5772 1272
rect -5868 1192 -5772 1208
rect -5868 1128 -5852 1192
rect -5788 1128 -5772 1192
rect -5868 1112 -5772 1128
rect -5868 1048 -5852 1112
rect -5788 1048 -5772 1112
rect -5868 1032 -5772 1048
rect -5868 968 -5852 1032
rect -5788 968 -5772 1032
rect -5868 952 -5772 968
rect -5868 888 -5852 952
rect -5788 888 -5772 952
rect -5868 872 -5772 888
rect -5868 808 -5852 872
rect -5788 808 -5772 872
rect -5868 792 -5772 808
rect -7280 692 -7184 728
rect -5868 728 -5852 792
rect -5788 728 -5772 792
rect -5449 1472 -4727 1481
rect -5449 768 -5440 1472
rect -4736 768 -4727 1472
rect -5449 759 -4727 768
rect -4456 1448 -4440 1512
rect -4376 1448 -4360 1512
rect -3044 1512 -2948 1548
rect -4456 1432 -4360 1448
rect -4456 1368 -4440 1432
rect -4376 1368 -4360 1432
rect -4456 1352 -4360 1368
rect -4456 1288 -4440 1352
rect -4376 1288 -4360 1352
rect -4456 1272 -4360 1288
rect -4456 1208 -4440 1272
rect -4376 1208 -4360 1272
rect -4456 1192 -4360 1208
rect -4456 1128 -4440 1192
rect -4376 1128 -4360 1192
rect -4456 1112 -4360 1128
rect -4456 1048 -4440 1112
rect -4376 1048 -4360 1112
rect -4456 1032 -4360 1048
rect -4456 968 -4440 1032
rect -4376 968 -4360 1032
rect -4456 952 -4360 968
rect -4456 888 -4440 952
rect -4376 888 -4360 952
rect -4456 872 -4360 888
rect -4456 808 -4440 872
rect -4376 808 -4360 872
rect -4456 792 -4360 808
rect -5868 692 -5772 728
rect -4456 728 -4440 792
rect -4376 728 -4360 792
rect -4037 1472 -3315 1481
rect -4037 768 -4028 1472
rect -3324 768 -3315 1472
rect -4037 759 -3315 768
rect -3044 1448 -3028 1512
rect -2964 1448 -2948 1512
rect -1632 1512 -1536 1548
rect -3044 1432 -2948 1448
rect -3044 1368 -3028 1432
rect -2964 1368 -2948 1432
rect -3044 1352 -2948 1368
rect -3044 1288 -3028 1352
rect -2964 1288 -2948 1352
rect -3044 1272 -2948 1288
rect -3044 1208 -3028 1272
rect -2964 1208 -2948 1272
rect -3044 1192 -2948 1208
rect -3044 1128 -3028 1192
rect -2964 1128 -2948 1192
rect -3044 1112 -2948 1128
rect -3044 1048 -3028 1112
rect -2964 1048 -2948 1112
rect -3044 1032 -2948 1048
rect -3044 968 -3028 1032
rect -2964 968 -2948 1032
rect -3044 952 -2948 968
rect -3044 888 -3028 952
rect -2964 888 -2948 952
rect -3044 872 -2948 888
rect -3044 808 -3028 872
rect -2964 808 -2948 872
rect -3044 792 -2948 808
rect -4456 692 -4360 728
rect -3044 728 -3028 792
rect -2964 728 -2948 792
rect -2625 1472 -1903 1481
rect -2625 768 -2616 1472
rect -1912 768 -1903 1472
rect -2625 759 -1903 768
rect -1632 1448 -1616 1512
rect -1552 1448 -1536 1512
rect -220 1512 -124 1548
rect -1632 1432 -1536 1448
rect -1632 1368 -1616 1432
rect -1552 1368 -1536 1432
rect -1632 1352 -1536 1368
rect -1632 1288 -1616 1352
rect -1552 1288 -1536 1352
rect -1632 1272 -1536 1288
rect -1632 1208 -1616 1272
rect -1552 1208 -1536 1272
rect -1632 1192 -1536 1208
rect -1632 1128 -1616 1192
rect -1552 1128 -1536 1192
rect -1632 1112 -1536 1128
rect -1632 1048 -1616 1112
rect -1552 1048 -1536 1112
rect -1632 1032 -1536 1048
rect -1632 968 -1616 1032
rect -1552 968 -1536 1032
rect -1632 952 -1536 968
rect -1632 888 -1616 952
rect -1552 888 -1536 952
rect -1632 872 -1536 888
rect -1632 808 -1616 872
rect -1552 808 -1536 872
rect -1632 792 -1536 808
rect -3044 692 -2948 728
rect -1632 728 -1616 792
rect -1552 728 -1536 792
rect -1213 1472 -491 1481
rect -1213 768 -1204 1472
rect -500 768 -491 1472
rect -1213 759 -491 768
rect -220 1448 -204 1512
rect -140 1448 -124 1512
rect 1192 1512 1288 1548
rect -220 1432 -124 1448
rect -220 1368 -204 1432
rect -140 1368 -124 1432
rect -220 1352 -124 1368
rect -220 1288 -204 1352
rect -140 1288 -124 1352
rect -220 1272 -124 1288
rect -220 1208 -204 1272
rect -140 1208 -124 1272
rect -220 1192 -124 1208
rect -220 1128 -204 1192
rect -140 1128 -124 1192
rect -220 1112 -124 1128
rect -220 1048 -204 1112
rect -140 1048 -124 1112
rect -220 1032 -124 1048
rect -220 968 -204 1032
rect -140 968 -124 1032
rect -220 952 -124 968
rect -220 888 -204 952
rect -140 888 -124 952
rect -220 872 -124 888
rect -220 808 -204 872
rect -140 808 -124 872
rect -220 792 -124 808
rect -1632 692 -1536 728
rect -220 728 -204 792
rect -140 728 -124 792
rect 199 1472 921 1481
rect 199 768 208 1472
rect 912 768 921 1472
rect 199 759 921 768
rect 1192 1448 1208 1512
rect 1272 1448 1288 1512
rect 2604 1512 2700 1548
rect 1192 1432 1288 1448
rect 1192 1368 1208 1432
rect 1272 1368 1288 1432
rect 1192 1352 1288 1368
rect 1192 1288 1208 1352
rect 1272 1288 1288 1352
rect 1192 1272 1288 1288
rect 1192 1208 1208 1272
rect 1272 1208 1288 1272
rect 1192 1192 1288 1208
rect 1192 1128 1208 1192
rect 1272 1128 1288 1192
rect 1192 1112 1288 1128
rect 1192 1048 1208 1112
rect 1272 1048 1288 1112
rect 1192 1032 1288 1048
rect 1192 968 1208 1032
rect 1272 968 1288 1032
rect 1192 952 1288 968
rect 1192 888 1208 952
rect 1272 888 1288 952
rect 1192 872 1288 888
rect 1192 808 1208 872
rect 1272 808 1288 872
rect 1192 792 1288 808
rect -220 692 -124 728
rect 1192 728 1208 792
rect 1272 728 1288 792
rect 1611 1472 2333 1481
rect 1611 768 1620 1472
rect 2324 768 2333 1472
rect 1611 759 2333 768
rect 2604 1448 2620 1512
rect 2684 1448 2700 1512
rect 4016 1512 4112 1548
rect 2604 1432 2700 1448
rect 2604 1368 2620 1432
rect 2684 1368 2700 1432
rect 2604 1352 2700 1368
rect 2604 1288 2620 1352
rect 2684 1288 2700 1352
rect 2604 1272 2700 1288
rect 2604 1208 2620 1272
rect 2684 1208 2700 1272
rect 2604 1192 2700 1208
rect 2604 1128 2620 1192
rect 2684 1128 2700 1192
rect 2604 1112 2700 1128
rect 2604 1048 2620 1112
rect 2684 1048 2700 1112
rect 2604 1032 2700 1048
rect 2604 968 2620 1032
rect 2684 968 2700 1032
rect 2604 952 2700 968
rect 2604 888 2620 952
rect 2684 888 2700 952
rect 2604 872 2700 888
rect 2604 808 2620 872
rect 2684 808 2700 872
rect 2604 792 2700 808
rect 1192 692 1288 728
rect 2604 728 2620 792
rect 2684 728 2700 792
rect 3023 1472 3745 1481
rect 3023 768 3032 1472
rect 3736 768 3745 1472
rect 3023 759 3745 768
rect 4016 1448 4032 1512
rect 4096 1448 4112 1512
rect 5428 1512 5524 1548
rect 4016 1432 4112 1448
rect 4016 1368 4032 1432
rect 4096 1368 4112 1432
rect 4016 1352 4112 1368
rect 4016 1288 4032 1352
rect 4096 1288 4112 1352
rect 4016 1272 4112 1288
rect 4016 1208 4032 1272
rect 4096 1208 4112 1272
rect 4016 1192 4112 1208
rect 4016 1128 4032 1192
rect 4096 1128 4112 1192
rect 4016 1112 4112 1128
rect 4016 1048 4032 1112
rect 4096 1048 4112 1112
rect 4016 1032 4112 1048
rect 4016 968 4032 1032
rect 4096 968 4112 1032
rect 4016 952 4112 968
rect 4016 888 4032 952
rect 4096 888 4112 952
rect 4016 872 4112 888
rect 4016 808 4032 872
rect 4096 808 4112 872
rect 4016 792 4112 808
rect 2604 692 2700 728
rect 4016 728 4032 792
rect 4096 728 4112 792
rect 4435 1472 5157 1481
rect 4435 768 4444 1472
rect 5148 768 5157 1472
rect 4435 759 5157 768
rect 5428 1448 5444 1512
rect 5508 1448 5524 1512
rect 6840 1512 6936 1548
rect 5428 1432 5524 1448
rect 5428 1368 5444 1432
rect 5508 1368 5524 1432
rect 5428 1352 5524 1368
rect 5428 1288 5444 1352
rect 5508 1288 5524 1352
rect 5428 1272 5524 1288
rect 5428 1208 5444 1272
rect 5508 1208 5524 1272
rect 5428 1192 5524 1208
rect 5428 1128 5444 1192
rect 5508 1128 5524 1192
rect 5428 1112 5524 1128
rect 5428 1048 5444 1112
rect 5508 1048 5524 1112
rect 5428 1032 5524 1048
rect 5428 968 5444 1032
rect 5508 968 5524 1032
rect 5428 952 5524 968
rect 5428 888 5444 952
rect 5508 888 5524 952
rect 5428 872 5524 888
rect 5428 808 5444 872
rect 5508 808 5524 872
rect 5428 792 5524 808
rect 4016 692 4112 728
rect 5428 728 5444 792
rect 5508 728 5524 792
rect 5847 1472 6569 1481
rect 5847 768 5856 1472
rect 6560 768 6569 1472
rect 5847 759 6569 768
rect 6840 1448 6856 1512
rect 6920 1448 6936 1512
rect 8252 1512 8348 1548
rect 6840 1432 6936 1448
rect 6840 1368 6856 1432
rect 6920 1368 6936 1432
rect 6840 1352 6936 1368
rect 6840 1288 6856 1352
rect 6920 1288 6936 1352
rect 6840 1272 6936 1288
rect 6840 1208 6856 1272
rect 6920 1208 6936 1272
rect 6840 1192 6936 1208
rect 6840 1128 6856 1192
rect 6920 1128 6936 1192
rect 6840 1112 6936 1128
rect 6840 1048 6856 1112
rect 6920 1048 6936 1112
rect 6840 1032 6936 1048
rect 6840 968 6856 1032
rect 6920 968 6936 1032
rect 6840 952 6936 968
rect 6840 888 6856 952
rect 6920 888 6936 952
rect 6840 872 6936 888
rect 6840 808 6856 872
rect 6920 808 6936 872
rect 6840 792 6936 808
rect 5428 692 5524 728
rect 6840 728 6856 792
rect 6920 728 6936 792
rect 7259 1472 7981 1481
rect 7259 768 7268 1472
rect 7972 768 7981 1472
rect 7259 759 7981 768
rect 8252 1448 8268 1512
rect 8332 1448 8348 1512
rect 9664 1512 9760 1548
rect 8252 1432 8348 1448
rect 8252 1368 8268 1432
rect 8332 1368 8348 1432
rect 8252 1352 8348 1368
rect 8252 1288 8268 1352
rect 8332 1288 8348 1352
rect 8252 1272 8348 1288
rect 8252 1208 8268 1272
rect 8332 1208 8348 1272
rect 8252 1192 8348 1208
rect 8252 1128 8268 1192
rect 8332 1128 8348 1192
rect 8252 1112 8348 1128
rect 8252 1048 8268 1112
rect 8332 1048 8348 1112
rect 8252 1032 8348 1048
rect 8252 968 8268 1032
rect 8332 968 8348 1032
rect 8252 952 8348 968
rect 8252 888 8268 952
rect 8332 888 8348 952
rect 8252 872 8348 888
rect 8252 808 8268 872
rect 8332 808 8348 872
rect 8252 792 8348 808
rect 6840 692 6936 728
rect 8252 728 8268 792
rect 8332 728 8348 792
rect 8671 1472 9393 1481
rect 8671 768 8680 1472
rect 9384 768 9393 1472
rect 8671 759 9393 768
rect 9664 1448 9680 1512
rect 9744 1448 9760 1512
rect 11076 1512 11172 1548
rect 9664 1432 9760 1448
rect 9664 1368 9680 1432
rect 9744 1368 9760 1432
rect 9664 1352 9760 1368
rect 9664 1288 9680 1352
rect 9744 1288 9760 1352
rect 9664 1272 9760 1288
rect 9664 1208 9680 1272
rect 9744 1208 9760 1272
rect 9664 1192 9760 1208
rect 9664 1128 9680 1192
rect 9744 1128 9760 1192
rect 9664 1112 9760 1128
rect 9664 1048 9680 1112
rect 9744 1048 9760 1112
rect 9664 1032 9760 1048
rect 9664 968 9680 1032
rect 9744 968 9760 1032
rect 9664 952 9760 968
rect 9664 888 9680 952
rect 9744 888 9760 952
rect 9664 872 9760 888
rect 9664 808 9680 872
rect 9744 808 9760 872
rect 9664 792 9760 808
rect 8252 692 8348 728
rect 9664 728 9680 792
rect 9744 728 9760 792
rect 10083 1472 10805 1481
rect 10083 768 10092 1472
rect 10796 768 10805 1472
rect 10083 759 10805 768
rect 11076 1448 11092 1512
rect 11156 1448 11172 1512
rect 12488 1512 12584 1548
rect 11076 1432 11172 1448
rect 11076 1368 11092 1432
rect 11156 1368 11172 1432
rect 11076 1352 11172 1368
rect 11076 1288 11092 1352
rect 11156 1288 11172 1352
rect 11076 1272 11172 1288
rect 11076 1208 11092 1272
rect 11156 1208 11172 1272
rect 11076 1192 11172 1208
rect 11076 1128 11092 1192
rect 11156 1128 11172 1192
rect 11076 1112 11172 1128
rect 11076 1048 11092 1112
rect 11156 1048 11172 1112
rect 11076 1032 11172 1048
rect 11076 968 11092 1032
rect 11156 968 11172 1032
rect 11076 952 11172 968
rect 11076 888 11092 952
rect 11156 888 11172 952
rect 11076 872 11172 888
rect 11076 808 11092 872
rect 11156 808 11172 872
rect 11076 792 11172 808
rect 9664 692 9760 728
rect 11076 728 11092 792
rect 11156 728 11172 792
rect 11495 1472 12217 1481
rect 11495 768 11504 1472
rect 12208 768 12217 1472
rect 11495 759 12217 768
rect 12488 1448 12504 1512
rect 12568 1448 12584 1512
rect 13900 1512 13996 1548
rect 12488 1432 12584 1448
rect 12488 1368 12504 1432
rect 12568 1368 12584 1432
rect 12488 1352 12584 1368
rect 12488 1288 12504 1352
rect 12568 1288 12584 1352
rect 12488 1272 12584 1288
rect 12488 1208 12504 1272
rect 12568 1208 12584 1272
rect 12488 1192 12584 1208
rect 12488 1128 12504 1192
rect 12568 1128 12584 1192
rect 12488 1112 12584 1128
rect 12488 1048 12504 1112
rect 12568 1048 12584 1112
rect 12488 1032 12584 1048
rect 12488 968 12504 1032
rect 12568 968 12584 1032
rect 12488 952 12584 968
rect 12488 888 12504 952
rect 12568 888 12584 952
rect 12488 872 12584 888
rect 12488 808 12504 872
rect 12568 808 12584 872
rect 12488 792 12584 808
rect 11076 692 11172 728
rect 12488 728 12504 792
rect 12568 728 12584 792
rect 12907 1472 13629 1481
rect 12907 768 12916 1472
rect 13620 768 13629 1472
rect 12907 759 13629 768
rect 13900 1448 13916 1512
rect 13980 1448 13996 1512
rect 15312 1512 15408 1548
rect 13900 1432 13996 1448
rect 13900 1368 13916 1432
rect 13980 1368 13996 1432
rect 13900 1352 13996 1368
rect 13900 1288 13916 1352
rect 13980 1288 13996 1352
rect 13900 1272 13996 1288
rect 13900 1208 13916 1272
rect 13980 1208 13996 1272
rect 13900 1192 13996 1208
rect 13900 1128 13916 1192
rect 13980 1128 13996 1192
rect 13900 1112 13996 1128
rect 13900 1048 13916 1112
rect 13980 1048 13996 1112
rect 13900 1032 13996 1048
rect 13900 968 13916 1032
rect 13980 968 13996 1032
rect 13900 952 13996 968
rect 13900 888 13916 952
rect 13980 888 13996 952
rect 13900 872 13996 888
rect 13900 808 13916 872
rect 13980 808 13996 872
rect 13900 792 13996 808
rect 12488 692 12584 728
rect 13900 728 13916 792
rect 13980 728 13996 792
rect 14319 1472 15041 1481
rect 14319 768 14328 1472
rect 15032 768 15041 1472
rect 14319 759 15041 768
rect 15312 1448 15328 1512
rect 15392 1448 15408 1512
rect 16724 1512 16820 1548
rect 15312 1432 15408 1448
rect 15312 1368 15328 1432
rect 15392 1368 15408 1432
rect 15312 1352 15408 1368
rect 15312 1288 15328 1352
rect 15392 1288 15408 1352
rect 15312 1272 15408 1288
rect 15312 1208 15328 1272
rect 15392 1208 15408 1272
rect 15312 1192 15408 1208
rect 15312 1128 15328 1192
rect 15392 1128 15408 1192
rect 15312 1112 15408 1128
rect 15312 1048 15328 1112
rect 15392 1048 15408 1112
rect 15312 1032 15408 1048
rect 15312 968 15328 1032
rect 15392 968 15408 1032
rect 15312 952 15408 968
rect 15312 888 15328 952
rect 15392 888 15408 952
rect 15312 872 15408 888
rect 15312 808 15328 872
rect 15392 808 15408 872
rect 15312 792 15408 808
rect 13900 692 13996 728
rect 15312 728 15328 792
rect 15392 728 15408 792
rect 15731 1472 16453 1481
rect 15731 768 15740 1472
rect 16444 768 16453 1472
rect 15731 759 16453 768
rect 16724 1448 16740 1512
rect 16804 1448 16820 1512
rect 18136 1512 18232 1548
rect 16724 1432 16820 1448
rect 16724 1368 16740 1432
rect 16804 1368 16820 1432
rect 16724 1352 16820 1368
rect 16724 1288 16740 1352
rect 16804 1288 16820 1352
rect 16724 1272 16820 1288
rect 16724 1208 16740 1272
rect 16804 1208 16820 1272
rect 16724 1192 16820 1208
rect 16724 1128 16740 1192
rect 16804 1128 16820 1192
rect 16724 1112 16820 1128
rect 16724 1048 16740 1112
rect 16804 1048 16820 1112
rect 16724 1032 16820 1048
rect 16724 968 16740 1032
rect 16804 968 16820 1032
rect 16724 952 16820 968
rect 16724 888 16740 952
rect 16804 888 16820 952
rect 16724 872 16820 888
rect 16724 808 16740 872
rect 16804 808 16820 872
rect 16724 792 16820 808
rect 15312 692 15408 728
rect 16724 728 16740 792
rect 16804 728 16820 792
rect 17143 1472 17865 1481
rect 17143 768 17152 1472
rect 17856 768 17865 1472
rect 17143 759 17865 768
rect 18136 1448 18152 1512
rect 18216 1448 18232 1512
rect 19548 1512 19644 1548
rect 18136 1432 18232 1448
rect 18136 1368 18152 1432
rect 18216 1368 18232 1432
rect 18136 1352 18232 1368
rect 18136 1288 18152 1352
rect 18216 1288 18232 1352
rect 18136 1272 18232 1288
rect 18136 1208 18152 1272
rect 18216 1208 18232 1272
rect 18136 1192 18232 1208
rect 18136 1128 18152 1192
rect 18216 1128 18232 1192
rect 18136 1112 18232 1128
rect 18136 1048 18152 1112
rect 18216 1048 18232 1112
rect 18136 1032 18232 1048
rect 18136 968 18152 1032
rect 18216 968 18232 1032
rect 18136 952 18232 968
rect 18136 888 18152 952
rect 18216 888 18232 952
rect 18136 872 18232 888
rect 18136 808 18152 872
rect 18216 808 18232 872
rect 18136 792 18232 808
rect 16724 692 16820 728
rect 18136 728 18152 792
rect 18216 728 18232 792
rect 18555 1472 19277 1481
rect 18555 768 18564 1472
rect 19268 768 19277 1472
rect 18555 759 19277 768
rect 19548 1448 19564 1512
rect 19628 1448 19644 1512
rect 20960 1512 21056 1548
rect 19548 1432 19644 1448
rect 19548 1368 19564 1432
rect 19628 1368 19644 1432
rect 19548 1352 19644 1368
rect 19548 1288 19564 1352
rect 19628 1288 19644 1352
rect 19548 1272 19644 1288
rect 19548 1208 19564 1272
rect 19628 1208 19644 1272
rect 19548 1192 19644 1208
rect 19548 1128 19564 1192
rect 19628 1128 19644 1192
rect 19548 1112 19644 1128
rect 19548 1048 19564 1112
rect 19628 1048 19644 1112
rect 19548 1032 19644 1048
rect 19548 968 19564 1032
rect 19628 968 19644 1032
rect 19548 952 19644 968
rect 19548 888 19564 952
rect 19628 888 19644 952
rect 19548 872 19644 888
rect 19548 808 19564 872
rect 19628 808 19644 872
rect 19548 792 19644 808
rect 18136 692 18232 728
rect 19548 728 19564 792
rect 19628 728 19644 792
rect 19967 1472 20689 1481
rect 19967 768 19976 1472
rect 20680 768 20689 1472
rect 19967 759 20689 768
rect 20960 1448 20976 1512
rect 21040 1448 21056 1512
rect 22372 1512 22468 1548
rect 20960 1432 21056 1448
rect 20960 1368 20976 1432
rect 21040 1368 21056 1432
rect 20960 1352 21056 1368
rect 20960 1288 20976 1352
rect 21040 1288 21056 1352
rect 20960 1272 21056 1288
rect 20960 1208 20976 1272
rect 21040 1208 21056 1272
rect 20960 1192 21056 1208
rect 20960 1128 20976 1192
rect 21040 1128 21056 1192
rect 20960 1112 21056 1128
rect 20960 1048 20976 1112
rect 21040 1048 21056 1112
rect 20960 1032 21056 1048
rect 20960 968 20976 1032
rect 21040 968 21056 1032
rect 20960 952 21056 968
rect 20960 888 20976 952
rect 21040 888 21056 952
rect 20960 872 21056 888
rect 20960 808 20976 872
rect 21040 808 21056 872
rect 20960 792 21056 808
rect 19548 692 19644 728
rect 20960 728 20976 792
rect 21040 728 21056 792
rect 21379 1472 22101 1481
rect 21379 768 21388 1472
rect 22092 768 22101 1472
rect 21379 759 22101 768
rect 22372 1448 22388 1512
rect 22452 1448 22468 1512
rect 23784 1512 23880 1548
rect 22372 1432 22468 1448
rect 22372 1368 22388 1432
rect 22452 1368 22468 1432
rect 22372 1352 22468 1368
rect 22372 1288 22388 1352
rect 22452 1288 22468 1352
rect 22372 1272 22468 1288
rect 22372 1208 22388 1272
rect 22452 1208 22468 1272
rect 22372 1192 22468 1208
rect 22372 1128 22388 1192
rect 22452 1128 22468 1192
rect 22372 1112 22468 1128
rect 22372 1048 22388 1112
rect 22452 1048 22468 1112
rect 22372 1032 22468 1048
rect 22372 968 22388 1032
rect 22452 968 22468 1032
rect 22372 952 22468 968
rect 22372 888 22388 952
rect 22452 888 22468 952
rect 22372 872 22468 888
rect 22372 808 22388 872
rect 22452 808 22468 872
rect 22372 792 22468 808
rect 20960 692 21056 728
rect 22372 728 22388 792
rect 22452 728 22468 792
rect 22791 1472 23513 1481
rect 22791 768 22800 1472
rect 23504 768 23513 1472
rect 22791 759 23513 768
rect 23784 1448 23800 1512
rect 23864 1448 23880 1512
rect 23784 1432 23880 1448
rect 23784 1368 23800 1432
rect 23864 1368 23880 1432
rect 23784 1352 23880 1368
rect 23784 1288 23800 1352
rect 23864 1288 23880 1352
rect 23784 1272 23880 1288
rect 23784 1208 23800 1272
rect 23864 1208 23880 1272
rect 23784 1192 23880 1208
rect 23784 1128 23800 1192
rect 23864 1128 23880 1192
rect 23784 1112 23880 1128
rect 23784 1048 23800 1112
rect 23864 1048 23880 1112
rect 23784 1032 23880 1048
rect 23784 968 23800 1032
rect 23864 968 23880 1032
rect 23784 952 23880 968
rect 23784 888 23800 952
rect 23864 888 23880 952
rect 23784 872 23880 888
rect 23784 808 23800 872
rect 23864 808 23880 872
rect 23784 792 23880 808
rect 22372 692 22468 728
rect 23784 728 23800 792
rect 23864 728 23880 792
rect 23784 692 23880 728
rect -22812 392 -22716 428
rect -23805 352 -23083 361
rect -23805 -352 -23796 352
rect -23092 -352 -23083 352
rect -23805 -361 -23083 -352
rect -22812 328 -22796 392
rect -22732 328 -22716 392
rect -21400 392 -21304 428
rect -22812 312 -22716 328
rect -22812 248 -22796 312
rect -22732 248 -22716 312
rect -22812 232 -22716 248
rect -22812 168 -22796 232
rect -22732 168 -22716 232
rect -22812 152 -22716 168
rect -22812 88 -22796 152
rect -22732 88 -22716 152
rect -22812 72 -22716 88
rect -22812 8 -22796 72
rect -22732 8 -22716 72
rect -22812 -8 -22716 8
rect -22812 -72 -22796 -8
rect -22732 -72 -22716 -8
rect -22812 -88 -22716 -72
rect -22812 -152 -22796 -88
rect -22732 -152 -22716 -88
rect -22812 -168 -22716 -152
rect -22812 -232 -22796 -168
rect -22732 -232 -22716 -168
rect -22812 -248 -22716 -232
rect -22812 -312 -22796 -248
rect -22732 -312 -22716 -248
rect -22812 -328 -22716 -312
rect -22812 -392 -22796 -328
rect -22732 -392 -22716 -328
rect -22393 352 -21671 361
rect -22393 -352 -22384 352
rect -21680 -352 -21671 352
rect -22393 -361 -21671 -352
rect -21400 328 -21384 392
rect -21320 328 -21304 392
rect -19988 392 -19892 428
rect -21400 312 -21304 328
rect -21400 248 -21384 312
rect -21320 248 -21304 312
rect -21400 232 -21304 248
rect -21400 168 -21384 232
rect -21320 168 -21304 232
rect -21400 152 -21304 168
rect -21400 88 -21384 152
rect -21320 88 -21304 152
rect -21400 72 -21304 88
rect -21400 8 -21384 72
rect -21320 8 -21304 72
rect -21400 -8 -21304 8
rect -21400 -72 -21384 -8
rect -21320 -72 -21304 -8
rect -21400 -88 -21304 -72
rect -21400 -152 -21384 -88
rect -21320 -152 -21304 -88
rect -21400 -168 -21304 -152
rect -21400 -232 -21384 -168
rect -21320 -232 -21304 -168
rect -21400 -248 -21304 -232
rect -21400 -312 -21384 -248
rect -21320 -312 -21304 -248
rect -21400 -328 -21304 -312
rect -22812 -428 -22716 -392
rect -21400 -392 -21384 -328
rect -21320 -392 -21304 -328
rect -20981 352 -20259 361
rect -20981 -352 -20972 352
rect -20268 -352 -20259 352
rect -20981 -361 -20259 -352
rect -19988 328 -19972 392
rect -19908 328 -19892 392
rect -18576 392 -18480 428
rect -19988 312 -19892 328
rect -19988 248 -19972 312
rect -19908 248 -19892 312
rect -19988 232 -19892 248
rect -19988 168 -19972 232
rect -19908 168 -19892 232
rect -19988 152 -19892 168
rect -19988 88 -19972 152
rect -19908 88 -19892 152
rect -19988 72 -19892 88
rect -19988 8 -19972 72
rect -19908 8 -19892 72
rect -19988 -8 -19892 8
rect -19988 -72 -19972 -8
rect -19908 -72 -19892 -8
rect -19988 -88 -19892 -72
rect -19988 -152 -19972 -88
rect -19908 -152 -19892 -88
rect -19988 -168 -19892 -152
rect -19988 -232 -19972 -168
rect -19908 -232 -19892 -168
rect -19988 -248 -19892 -232
rect -19988 -312 -19972 -248
rect -19908 -312 -19892 -248
rect -19988 -328 -19892 -312
rect -21400 -428 -21304 -392
rect -19988 -392 -19972 -328
rect -19908 -392 -19892 -328
rect -19569 352 -18847 361
rect -19569 -352 -19560 352
rect -18856 -352 -18847 352
rect -19569 -361 -18847 -352
rect -18576 328 -18560 392
rect -18496 328 -18480 392
rect -17164 392 -17068 428
rect -18576 312 -18480 328
rect -18576 248 -18560 312
rect -18496 248 -18480 312
rect -18576 232 -18480 248
rect -18576 168 -18560 232
rect -18496 168 -18480 232
rect -18576 152 -18480 168
rect -18576 88 -18560 152
rect -18496 88 -18480 152
rect -18576 72 -18480 88
rect -18576 8 -18560 72
rect -18496 8 -18480 72
rect -18576 -8 -18480 8
rect -18576 -72 -18560 -8
rect -18496 -72 -18480 -8
rect -18576 -88 -18480 -72
rect -18576 -152 -18560 -88
rect -18496 -152 -18480 -88
rect -18576 -168 -18480 -152
rect -18576 -232 -18560 -168
rect -18496 -232 -18480 -168
rect -18576 -248 -18480 -232
rect -18576 -312 -18560 -248
rect -18496 -312 -18480 -248
rect -18576 -328 -18480 -312
rect -19988 -428 -19892 -392
rect -18576 -392 -18560 -328
rect -18496 -392 -18480 -328
rect -18157 352 -17435 361
rect -18157 -352 -18148 352
rect -17444 -352 -17435 352
rect -18157 -361 -17435 -352
rect -17164 328 -17148 392
rect -17084 328 -17068 392
rect -15752 392 -15656 428
rect -17164 312 -17068 328
rect -17164 248 -17148 312
rect -17084 248 -17068 312
rect -17164 232 -17068 248
rect -17164 168 -17148 232
rect -17084 168 -17068 232
rect -17164 152 -17068 168
rect -17164 88 -17148 152
rect -17084 88 -17068 152
rect -17164 72 -17068 88
rect -17164 8 -17148 72
rect -17084 8 -17068 72
rect -17164 -8 -17068 8
rect -17164 -72 -17148 -8
rect -17084 -72 -17068 -8
rect -17164 -88 -17068 -72
rect -17164 -152 -17148 -88
rect -17084 -152 -17068 -88
rect -17164 -168 -17068 -152
rect -17164 -232 -17148 -168
rect -17084 -232 -17068 -168
rect -17164 -248 -17068 -232
rect -17164 -312 -17148 -248
rect -17084 -312 -17068 -248
rect -17164 -328 -17068 -312
rect -18576 -428 -18480 -392
rect -17164 -392 -17148 -328
rect -17084 -392 -17068 -328
rect -16745 352 -16023 361
rect -16745 -352 -16736 352
rect -16032 -352 -16023 352
rect -16745 -361 -16023 -352
rect -15752 328 -15736 392
rect -15672 328 -15656 392
rect -14340 392 -14244 428
rect -15752 312 -15656 328
rect -15752 248 -15736 312
rect -15672 248 -15656 312
rect -15752 232 -15656 248
rect -15752 168 -15736 232
rect -15672 168 -15656 232
rect -15752 152 -15656 168
rect -15752 88 -15736 152
rect -15672 88 -15656 152
rect -15752 72 -15656 88
rect -15752 8 -15736 72
rect -15672 8 -15656 72
rect -15752 -8 -15656 8
rect -15752 -72 -15736 -8
rect -15672 -72 -15656 -8
rect -15752 -88 -15656 -72
rect -15752 -152 -15736 -88
rect -15672 -152 -15656 -88
rect -15752 -168 -15656 -152
rect -15752 -232 -15736 -168
rect -15672 -232 -15656 -168
rect -15752 -248 -15656 -232
rect -15752 -312 -15736 -248
rect -15672 -312 -15656 -248
rect -15752 -328 -15656 -312
rect -17164 -428 -17068 -392
rect -15752 -392 -15736 -328
rect -15672 -392 -15656 -328
rect -15333 352 -14611 361
rect -15333 -352 -15324 352
rect -14620 -352 -14611 352
rect -15333 -361 -14611 -352
rect -14340 328 -14324 392
rect -14260 328 -14244 392
rect -12928 392 -12832 428
rect -14340 312 -14244 328
rect -14340 248 -14324 312
rect -14260 248 -14244 312
rect -14340 232 -14244 248
rect -14340 168 -14324 232
rect -14260 168 -14244 232
rect -14340 152 -14244 168
rect -14340 88 -14324 152
rect -14260 88 -14244 152
rect -14340 72 -14244 88
rect -14340 8 -14324 72
rect -14260 8 -14244 72
rect -14340 -8 -14244 8
rect -14340 -72 -14324 -8
rect -14260 -72 -14244 -8
rect -14340 -88 -14244 -72
rect -14340 -152 -14324 -88
rect -14260 -152 -14244 -88
rect -14340 -168 -14244 -152
rect -14340 -232 -14324 -168
rect -14260 -232 -14244 -168
rect -14340 -248 -14244 -232
rect -14340 -312 -14324 -248
rect -14260 -312 -14244 -248
rect -14340 -328 -14244 -312
rect -15752 -428 -15656 -392
rect -14340 -392 -14324 -328
rect -14260 -392 -14244 -328
rect -13921 352 -13199 361
rect -13921 -352 -13912 352
rect -13208 -352 -13199 352
rect -13921 -361 -13199 -352
rect -12928 328 -12912 392
rect -12848 328 -12832 392
rect -11516 392 -11420 428
rect -12928 312 -12832 328
rect -12928 248 -12912 312
rect -12848 248 -12832 312
rect -12928 232 -12832 248
rect -12928 168 -12912 232
rect -12848 168 -12832 232
rect -12928 152 -12832 168
rect -12928 88 -12912 152
rect -12848 88 -12832 152
rect -12928 72 -12832 88
rect -12928 8 -12912 72
rect -12848 8 -12832 72
rect -12928 -8 -12832 8
rect -12928 -72 -12912 -8
rect -12848 -72 -12832 -8
rect -12928 -88 -12832 -72
rect -12928 -152 -12912 -88
rect -12848 -152 -12832 -88
rect -12928 -168 -12832 -152
rect -12928 -232 -12912 -168
rect -12848 -232 -12832 -168
rect -12928 -248 -12832 -232
rect -12928 -312 -12912 -248
rect -12848 -312 -12832 -248
rect -12928 -328 -12832 -312
rect -14340 -428 -14244 -392
rect -12928 -392 -12912 -328
rect -12848 -392 -12832 -328
rect -12509 352 -11787 361
rect -12509 -352 -12500 352
rect -11796 -352 -11787 352
rect -12509 -361 -11787 -352
rect -11516 328 -11500 392
rect -11436 328 -11420 392
rect -10104 392 -10008 428
rect -11516 312 -11420 328
rect -11516 248 -11500 312
rect -11436 248 -11420 312
rect -11516 232 -11420 248
rect -11516 168 -11500 232
rect -11436 168 -11420 232
rect -11516 152 -11420 168
rect -11516 88 -11500 152
rect -11436 88 -11420 152
rect -11516 72 -11420 88
rect -11516 8 -11500 72
rect -11436 8 -11420 72
rect -11516 -8 -11420 8
rect -11516 -72 -11500 -8
rect -11436 -72 -11420 -8
rect -11516 -88 -11420 -72
rect -11516 -152 -11500 -88
rect -11436 -152 -11420 -88
rect -11516 -168 -11420 -152
rect -11516 -232 -11500 -168
rect -11436 -232 -11420 -168
rect -11516 -248 -11420 -232
rect -11516 -312 -11500 -248
rect -11436 -312 -11420 -248
rect -11516 -328 -11420 -312
rect -12928 -428 -12832 -392
rect -11516 -392 -11500 -328
rect -11436 -392 -11420 -328
rect -11097 352 -10375 361
rect -11097 -352 -11088 352
rect -10384 -352 -10375 352
rect -11097 -361 -10375 -352
rect -10104 328 -10088 392
rect -10024 328 -10008 392
rect -8692 392 -8596 428
rect -10104 312 -10008 328
rect -10104 248 -10088 312
rect -10024 248 -10008 312
rect -10104 232 -10008 248
rect -10104 168 -10088 232
rect -10024 168 -10008 232
rect -10104 152 -10008 168
rect -10104 88 -10088 152
rect -10024 88 -10008 152
rect -10104 72 -10008 88
rect -10104 8 -10088 72
rect -10024 8 -10008 72
rect -10104 -8 -10008 8
rect -10104 -72 -10088 -8
rect -10024 -72 -10008 -8
rect -10104 -88 -10008 -72
rect -10104 -152 -10088 -88
rect -10024 -152 -10008 -88
rect -10104 -168 -10008 -152
rect -10104 -232 -10088 -168
rect -10024 -232 -10008 -168
rect -10104 -248 -10008 -232
rect -10104 -312 -10088 -248
rect -10024 -312 -10008 -248
rect -10104 -328 -10008 -312
rect -11516 -428 -11420 -392
rect -10104 -392 -10088 -328
rect -10024 -392 -10008 -328
rect -9685 352 -8963 361
rect -9685 -352 -9676 352
rect -8972 -352 -8963 352
rect -9685 -361 -8963 -352
rect -8692 328 -8676 392
rect -8612 328 -8596 392
rect -7280 392 -7184 428
rect -8692 312 -8596 328
rect -8692 248 -8676 312
rect -8612 248 -8596 312
rect -8692 232 -8596 248
rect -8692 168 -8676 232
rect -8612 168 -8596 232
rect -8692 152 -8596 168
rect -8692 88 -8676 152
rect -8612 88 -8596 152
rect -8692 72 -8596 88
rect -8692 8 -8676 72
rect -8612 8 -8596 72
rect -8692 -8 -8596 8
rect -8692 -72 -8676 -8
rect -8612 -72 -8596 -8
rect -8692 -88 -8596 -72
rect -8692 -152 -8676 -88
rect -8612 -152 -8596 -88
rect -8692 -168 -8596 -152
rect -8692 -232 -8676 -168
rect -8612 -232 -8596 -168
rect -8692 -248 -8596 -232
rect -8692 -312 -8676 -248
rect -8612 -312 -8596 -248
rect -8692 -328 -8596 -312
rect -10104 -428 -10008 -392
rect -8692 -392 -8676 -328
rect -8612 -392 -8596 -328
rect -8273 352 -7551 361
rect -8273 -352 -8264 352
rect -7560 -352 -7551 352
rect -8273 -361 -7551 -352
rect -7280 328 -7264 392
rect -7200 328 -7184 392
rect -5868 392 -5772 428
rect -7280 312 -7184 328
rect -7280 248 -7264 312
rect -7200 248 -7184 312
rect -7280 232 -7184 248
rect -7280 168 -7264 232
rect -7200 168 -7184 232
rect -7280 152 -7184 168
rect -7280 88 -7264 152
rect -7200 88 -7184 152
rect -7280 72 -7184 88
rect -7280 8 -7264 72
rect -7200 8 -7184 72
rect -7280 -8 -7184 8
rect -7280 -72 -7264 -8
rect -7200 -72 -7184 -8
rect -7280 -88 -7184 -72
rect -7280 -152 -7264 -88
rect -7200 -152 -7184 -88
rect -7280 -168 -7184 -152
rect -7280 -232 -7264 -168
rect -7200 -232 -7184 -168
rect -7280 -248 -7184 -232
rect -7280 -312 -7264 -248
rect -7200 -312 -7184 -248
rect -7280 -328 -7184 -312
rect -8692 -428 -8596 -392
rect -7280 -392 -7264 -328
rect -7200 -392 -7184 -328
rect -6861 352 -6139 361
rect -6861 -352 -6852 352
rect -6148 -352 -6139 352
rect -6861 -361 -6139 -352
rect -5868 328 -5852 392
rect -5788 328 -5772 392
rect -4456 392 -4360 428
rect -5868 312 -5772 328
rect -5868 248 -5852 312
rect -5788 248 -5772 312
rect -5868 232 -5772 248
rect -5868 168 -5852 232
rect -5788 168 -5772 232
rect -5868 152 -5772 168
rect -5868 88 -5852 152
rect -5788 88 -5772 152
rect -5868 72 -5772 88
rect -5868 8 -5852 72
rect -5788 8 -5772 72
rect -5868 -8 -5772 8
rect -5868 -72 -5852 -8
rect -5788 -72 -5772 -8
rect -5868 -88 -5772 -72
rect -5868 -152 -5852 -88
rect -5788 -152 -5772 -88
rect -5868 -168 -5772 -152
rect -5868 -232 -5852 -168
rect -5788 -232 -5772 -168
rect -5868 -248 -5772 -232
rect -5868 -312 -5852 -248
rect -5788 -312 -5772 -248
rect -5868 -328 -5772 -312
rect -7280 -428 -7184 -392
rect -5868 -392 -5852 -328
rect -5788 -392 -5772 -328
rect -5449 352 -4727 361
rect -5449 -352 -5440 352
rect -4736 -352 -4727 352
rect -5449 -361 -4727 -352
rect -4456 328 -4440 392
rect -4376 328 -4360 392
rect -3044 392 -2948 428
rect -4456 312 -4360 328
rect -4456 248 -4440 312
rect -4376 248 -4360 312
rect -4456 232 -4360 248
rect -4456 168 -4440 232
rect -4376 168 -4360 232
rect -4456 152 -4360 168
rect -4456 88 -4440 152
rect -4376 88 -4360 152
rect -4456 72 -4360 88
rect -4456 8 -4440 72
rect -4376 8 -4360 72
rect -4456 -8 -4360 8
rect -4456 -72 -4440 -8
rect -4376 -72 -4360 -8
rect -4456 -88 -4360 -72
rect -4456 -152 -4440 -88
rect -4376 -152 -4360 -88
rect -4456 -168 -4360 -152
rect -4456 -232 -4440 -168
rect -4376 -232 -4360 -168
rect -4456 -248 -4360 -232
rect -4456 -312 -4440 -248
rect -4376 -312 -4360 -248
rect -4456 -328 -4360 -312
rect -5868 -428 -5772 -392
rect -4456 -392 -4440 -328
rect -4376 -392 -4360 -328
rect -4037 352 -3315 361
rect -4037 -352 -4028 352
rect -3324 -352 -3315 352
rect -4037 -361 -3315 -352
rect -3044 328 -3028 392
rect -2964 328 -2948 392
rect -1632 392 -1536 428
rect -3044 312 -2948 328
rect -3044 248 -3028 312
rect -2964 248 -2948 312
rect -3044 232 -2948 248
rect -3044 168 -3028 232
rect -2964 168 -2948 232
rect -3044 152 -2948 168
rect -3044 88 -3028 152
rect -2964 88 -2948 152
rect -3044 72 -2948 88
rect -3044 8 -3028 72
rect -2964 8 -2948 72
rect -3044 -8 -2948 8
rect -3044 -72 -3028 -8
rect -2964 -72 -2948 -8
rect -3044 -88 -2948 -72
rect -3044 -152 -3028 -88
rect -2964 -152 -2948 -88
rect -3044 -168 -2948 -152
rect -3044 -232 -3028 -168
rect -2964 -232 -2948 -168
rect -3044 -248 -2948 -232
rect -3044 -312 -3028 -248
rect -2964 -312 -2948 -248
rect -3044 -328 -2948 -312
rect -4456 -428 -4360 -392
rect -3044 -392 -3028 -328
rect -2964 -392 -2948 -328
rect -2625 352 -1903 361
rect -2625 -352 -2616 352
rect -1912 -352 -1903 352
rect -2625 -361 -1903 -352
rect -1632 328 -1616 392
rect -1552 328 -1536 392
rect -220 392 -124 428
rect -1632 312 -1536 328
rect -1632 248 -1616 312
rect -1552 248 -1536 312
rect -1632 232 -1536 248
rect -1632 168 -1616 232
rect -1552 168 -1536 232
rect -1632 152 -1536 168
rect -1632 88 -1616 152
rect -1552 88 -1536 152
rect -1632 72 -1536 88
rect -1632 8 -1616 72
rect -1552 8 -1536 72
rect -1632 -8 -1536 8
rect -1632 -72 -1616 -8
rect -1552 -72 -1536 -8
rect -1632 -88 -1536 -72
rect -1632 -152 -1616 -88
rect -1552 -152 -1536 -88
rect -1632 -168 -1536 -152
rect -1632 -232 -1616 -168
rect -1552 -232 -1536 -168
rect -1632 -248 -1536 -232
rect -1632 -312 -1616 -248
rect -1552 -312 -1536 -248
rect -1632 -328 -1536 -312
rect -3044 -428 -2948 -392
rect -1632 -392 -1616 -328
rect -1552 -392 -1536 -328
rect -1213 352 -491 361
rect -1213 -352 -1204 352
rect -500 -352 -491 352
rect -1213 -361 -491 -352
rect -220 328 -204 392
rect -140 328 -124 392
rect 1192 392 1288 428
rect -220 312 -124 328
rect -220 248 -204 312
rect -140 248 -124 312
rect -220 232 -124 248
rect -220 168 -204 232
rect -140 168 -124 232
rect -220 152 -124 168
rect -220 88 -204 152
rect -140 88 -124 152
rect -220 72 -124 88
rect -220 8 -204 72
rect -140 8 -124 72
rect -220 -8 -124 8
rect -220 -72 -204 -8
rect -140 -72 -124 -8
rect -220 -88 -124 -72
rect -220 -152 -204 -88
rect -140 -152 -124 -88
rect -220 -168 -124 -152
rect -220 -232 -204 -168
rect -140 -232 -124 -168
rect -220 -248 -124 -232
rect -220 -312 -204 -248
rect -140 -312 -124 -248
rect -220 -328 -124 -312
rect -1632 -428 -1536 -392
rect -220 -392 -204 -328
rect -140 -392 -124 -328
rect 199 352 921 361
rect 199 -352 208 352
rect 912 -352 921 352
rect 199 -361 921 -352
rect 1192 328 1208 392
rect 1272 328 1288 392
rect 2604 392 2700 428
rect 1192 312 1288 328
rect 1192 248 1208 312
rect 1272 248 1288 312
rect 1192 232 1288 248
rect 1192 168 1208 232
rect 1272 168 1288 232
rect 1192 152 1288 168
rect 1192 88 1208 152
rect 1272 88 1288 152
rect 1192 72 1288 88
rect 1192 8 1208 72
rect 1272 8 1288 72
rect 1192 -8 1288 8
rect 1192 -72 1208 -8
rect 1272 -72 1288 -8
rect 1192 -88 1288 -72
rect 1192 -152 1208 -88
rect 1272 -152 1288 -88
rect 1192 -168 1288 -152
rect 1192 -232 1208 -168
rect 1272 -232 1288 -168
rect 1192 -248 1288 -232
rect 1192 -312 1208 -248
rect 1272 -312 1288 -248
rect 1192 -328 1288 -312
rect -220 -428 -124 -392
rect 1192 -392 1208 -328
rect 1272 -392 1288 -328
rect 1611 352 2333 361
rect 1611 -352 1620 352
rect 2324 -352 2333 352
rect 1611 -361 2333 -352
rect 2604 328 2620 392
rect 2684 328 2700 392
rect 4016 392 4112 428
rect 2604 312 2700 328
rect 2604 248 2620 312
rect 2684 248 2700 312
rect 2604 232 2700 248
rect 2604 168 2620 232
rect 2684 168 2700 232
rect 2604 152 2700 168
rect 2604 88 2620 152
rect 2684 88 2700 152
rect 2604 72 2700 88
rect 2604 8 2620 72
rect 2684 8 2700 72
rect 2604 -8 2700 8
rect 2604 -72 2620 -8
rect 2684 -72 2700 -8
rect 2604 -88 2700 -72
rect 2604 -152 2620 -88
rect 2684 -152 2700 -88
rect 2604 -168 2700 -152
rect 2604 -232 2620 -168
rect 2684 -232 2700 -168
rect 2604 -248 2700 -232
rect 2604 -312 2620 -248
rect 2684 -312 2700 -248
rect 2604 -328 2700 -312
rect 1192 -428 1288 -392
rect 2604 -392 2620 -328
rect 2684 -392 2700 -328
rect 3023 352 3745 361
rect 3023 -352 3032 352
rect 3736 -352 3745 352
rect 3023 -361 3745 -352
rect 4016 328 4032 392
rect 4096 328 4112 392
rect 5428 392 5524 428
rect 4016 312 4112 328
rect 4016 248 4032 312
rect 4096 248 4112 312
rect 4016 232 4112 248
rect 4016 168 4032 232
rect 4096 168 4112 232
rect 4016 152 4112 168
rect 4016 88 4032 152
rect 4096 88 4112 152
rect 4016 72 4112 88
rect 4016 8 4032 72
rect 4096 8 4112 72
rect 4016 -8 4112 8
rect 4016 -72 4032 -8
rect 4096 -72 4112 -8
rect 4016 -88 4112 -72
rect 4016 -152 4032 -88
rect 4096 -152 4112 -88
rect 4016 -168 4112 -152
rect 4016 -232 4032 -168
rect 4096 -232 4112 -168
rect 4016 -248 4112 -232
rect 4016 -312 4032 -248
rect 4096 -312 4112 -248
rect 4016 -328 4112 -312
rect 2604 -428 2700 -392
rect 4016 -392 4032 -328
rect 4096 -392 4112 -328
rect 4435 352 5157 361
rect 4435 -352 4444 352
rect 5148 -352 5157 352
rect 4435 -361 5157 -352
rect 5428 328 5444 392
rect 5508 328 5524 392
rect 6840 392 6936 428
rect 5428 312 5524 328
rect 5428 248 5444 312
rect 5508 248 5524 312
rect 5428 232 5524 248
rect 5428 168 5444 232
rect 5508 168 5524 232
rect 5428 152 5524 168
rect 5428 88 5444 152
rect 5508 88 5524 152
rect 5428 72 5524 88
rect 5428 8 5444 72
rect 5508 8 5524 72
rect 5428 -8 5524 8
rect 5428 -72 5444 -8
rect 5508 -72 5524 -8
rect 5428 -88 5524 -72
rect 5428 -152 5444 -88
rect 5508 -152 5524 -88
rect 5428 -168 5524 -152
rect 5428 -232 5444 -168
rect 5508 -232 5524 -168
rect 5428 -248 5524 -232
rect 5428 -312 5444 -248
rect 5508 -312 5524 -248
rect 5428 -328 5524 -312
rect 4016 -428 4112 -392
rect 5428 -392 5444 -328
rect 5508 -392 5524 -328
rect 5847 352 6569 361
rect 5847 -352 5856 352
rect 6560 -352 6569 352
rect 5847 -361 6569 -352
rect 6840 328 6856 392
rect 6920 328 6936 392
rect 8252 392 8348 428
rect 6840 312 6936 328
rect 6840 248 6856 312
rect 6920 248 6936 312
rect 6840 232 6936 248
rect 6840 168 6856 232
rect 6920 168 6936 232
rect 6840 152 6936 168
rect 6840 88 6856 152
rect 6920 88 6936 152
rect 6840 72 6936 88
rect 6840 8 6856 72
rect 6920 8 6936 72
rect 6840 -8 6936 8
rect 6840 -72 6856 -8
rect 6920 -72 6936 -8
rect 6840 -88 6936 -72
rect 6840 -152 6856 -88
rect 6920 -152 6936 -88
rect 6840 -168 6936 -152
rect 6840 -232 6856 -168
rect 6920 -232 6936 -168
rect 6840 -248 6936 -232
rect 6840 -312 6856 -248
rect 6920 -312 6936 -248
rect 6840 -328 6936 -312
rect 5428 -428 5524 -392
rect 6840 -392 6856 -328
rect 6920 -392 6936 -328
rect 7259 352 7981 361
rect 7259 -352 7268 352
rect 7972 -352 7981 352
rect 7259 -361 7981 -352
rect 8252 328 8268 392
rect 8332 328 8348 392
rect 9664 392 9760 428
rect 8252 312 8348 328
rect 8252 248 8268 312
rect 8332 248 8348 312
rect 8252 232 8348 248
rect 8252 168 8268 232
rect 8332 168 8348 232
rect 8252 152 8348 168
rect 8252 88 8268 152
rect 8332 88 8348 152
rect 8252 72 8348 88
rect 8252 8 8268 72
rect 8332 8 8348 72
rect 8252 -8 8348 8
rect 8252 -72 8268 -8
rect 8332 -72 8348 -8
rect 8252 -88 8348 -72
rect 8252 -152 8268 -88
rect 8332 -152 8348 -88
rect 8252 -168 8348 -152
rect 8252 -232 8268 -168
rect 8332 -232 8348 -168
rect 8252 -248 8348 -232
rect 8252 -312 8268 -248
rect 8332 -312 8348 -248
rect 8252 -328 8348 -312
rect 6840 -428 6936 -392
rect 8252 -392 8268 -328
rect 8332 -392 8348 -328
rect 8671 352 9393 361
rect 8671 -352 8680 352
rect 9384 -352 9393 352
rect 8671 -361 9393 -352
rect 9664 328 9680 392
rect 9744 328 9760 392
rect 11076 392 11172 428
rect 9664 312 9760 328
rect 9664 248 9680 312
rect 9744 248 9760 312
rect 9664 232 9760 248
rect 9664 168 9680 232
rect 9744 168 9760 232
rect 9664 152 9760 168
rect 9664 88 9680 152
rect 9744 88 9760 152
rect 9664 72 9760 88
rect 9664 8 9680 72
rect 9744 8 9760 72
rect 9664 -8 9760 8
rect 9664 -72 9680 -8
rect 9744 -72 9760 -8
rect 9664 -88 9760 -72
rect 9664 -152 9680 -88
rect 9744 -152 9760 -88
rect 9664 -168 9760 -152
rect 9664 -232 9680 -168
rect 9744 -232 9760 -168
rect 9664 -248 9760 -232
rect 9664 -312 9680 -248
rect 9744 -312 9760 -248
rect 9664 -328 9760 -312
rect 8252 -428 8348 -392
rect 9664 -392 9680 -328
rect 9744 -392 9760 -328
rect 10083 352 10805 361
rect 10083 -352 10092 352
rect 10796 -352 10805 352
rect 10083 -361 10805 -352
rect 11076 328 11092 392
rect 11156 328 11172 392
rect 12488 392 12584 428
rect 11076 312 11172 328
rect 11076 248 11092 312
rect 11156 248 11172 312
rect 11076 232 11172 248
rect 11076 168 11092 232
rect 11156 168 11172 232
rect 11076 152 11172 168
rect 11076 88 11092 152
rect 11156 88 11172 152
rect 11076 72 11172 88
rect 11076 8 11092 72
rect 11156 8 11172 72
rect 11076 -8 11172 8
rect 11076 -72 11092 -8
rect 11156 -72 11172 -8
rect 11076 -88 11172 -72
rect 11076 -152 11092 -88
rect 11156 -152 11172 -88
rect 11076 -168 11172 -152
rect 11076 -232 11092 -168
rect 11156 -232 11172 -168
rect 11076 -248 11172 -232
rect 11076 -312 11092 -248
rect 11156 -312 11172 -248
rect 11076 -328 11172 -312
rect 9664 -428 9760 -392
rect 11076 -392 11092 -328
rect 11156 -392 11172 -328
rect 11495 352 12217 361
rect 11495 -352 11504 352
rect 12208 -352 12217 352
rect 11495 -361 12217 -352
rect 12488 328 12504 392
rect 12568 328 12584 392
rect 13900 392 13996 428
rect 12488 312 12584 328
rect 12488 248 12504 312
rect 12568 248 12584 312
rect 12488 232 12584 248
rect 12488 168 12504 232
rect 12568 168 12584 232
rect 12488 152 12584 168
rect 12488 88 12504 152
rect 12568 88 12584 152
rect 12488 72 12584 88
rect 12488 8 12504 72
rect 12568 8 12584 72
rect 12488 -8 12584 8
rect 12488 -72 12504 -8
rect 12568 -72 12584 -8
rect 12488 -88 12584 -72
rect 12488 -152 12504 -88
rect 12568 -152 12584 -88
rect 12488 -168 12584 -152
rect 12488 -232 12504 -168
rect 12568 -232 12584 -168
rect 12488 -248 12584 -232
rect 12488 -312 12504 -248
rect 12568 -312 12584 -248
rect 12488 -328 12584 -312
rect 11076 -428 11172 -392
rect 12488 -392 12504 -328
rect 12568 -392 12584 -328
rect 12907 352 13629 361
rect 12907 -352 12916 352
rect 13620 -352 13629 352
rect 12907 -361 13629 -352
rect 13900 328 13916 392
rect 13980 328 13996 392
rect 15312 392 15408 428
rect 13900 312 13996 328
rect 13900 248 13916 312
rect 13980 248 13996 312
rect 13900 232 13996 248
rect 13900 168 13916 232
rect 13980 168 13996 232
rect 13900 152 13996 168
rect 13900 88 13916 152
rect 13980 88 13996 152
rect 13900 72 13996 88
rect 13900 8 13916 72
rect 13980 8 13996 72
rect 13900 -8 13996 8
rect 13900 -72 13916 -8
rect 13980 -72 13996 -8
rect 13900 -88 13996 -72
rect 13900 -152 13916 -88
rect 13980 -152 13996 -88
rect 13900 -168 13996 -152
rect 13900 -232 13916 -168
rect 13980 -232 13996 -168
rect 13900 -248 13996 -232
rect 13900 -312 13916 -248
rect 13980 -312 13996 -248
rect 13900 -328 13996 -312
rect 12488 -428 12584 -392
rect 13900 -392 13916 -328
rect 13980 -392 13996 -328
rect 14319 352 15041 361
rect 14319 -352 14328 352
rect 15032 -352 15041 352
rect 14319 -361 15041 -352
rect 15312 328 15328 392
rect 15392 328 15408 392
rect 16724 392 16820 428
rect 15312 312 15408 328
rect 15312 248 15328 312
rect 15392 248 15408 312
rect 15312 232 15408 248
rect 15312 168 15328 232
rect 15392 168 15408 232
rect 15312 152 15408 168
rect 15312 88 15328 152
rect 15392 88 15408 152
rect 15312 72 15408 88
rect 15312 8 15328 72
rect 15392 8 15408 72
rect 15312 -8 15408 8
rect 15312 -72 15328 -8
rect 15392 -72 15408 -8
rect 15312 -88 15408 -72
rect 15312 -152 15328 -88
rect 15392 -152 15408 -88
rect 15312 -168 15408 -152
rect 15312 -232 15328 -168
rect 15392 -232 15408 -168
rect 15312 -248 15408 -232
rect 15312 -312 15328 -248
rect 15392 -312 15408 -248
rect 15312 -328 15408 -312
rect 13900 -428 13996 -392
rect 15312 -392 15328 -328
rect 15392 -392 15408 -328
rect 15731 352 16453 361
rect 15731 -352 15740 352
rect 16444 -352 16453 352
rect 15731 -361 16453 -352
rect 16724 328 16740 392
rect 16804 328 16820 392
rect 18136 392 18232 428
rect 16724 312 16820 328
rect 16724 248 16740 312
rect 16804 248 16820 312
rect 16724 232 16820 248
rect 16724 168 16740 232
rect 16804 168 16820 232
rect 16724 152 16820 168
rect 16724 88 16740 152
rect 16804 88 16820 152
rect 16724 72 16820 88
rect 16724 8 16740 72
rect 16804 8 16820 72
rect 16724 -8 16820 8
rect 16724 -72 16740 -8
rect 16804 -72 16820 -8
rect 16724 -88 16820 -72
rect 16724 -152 16740 -88
rect 16804 -152 16820 -88
rect 16724 -168 16820 -152
rect 16724 -232 16740 -168
rect 16804 -232 16820 -168
rect 16724 -248 16820 -232
rect 16724 -312 16740 -248
rect 16804 -312 16820 -248
rect 16724 -328 16820 -312
rect 15312 -428 15408 -392
rect 16724 -392 16740 -328
rect 16804 -392 16820 -328
rect 17143 352 17865 361
rect 17143 -352 17152 352
rect 17856 -352 17865 352
rect 17143 -361 17865 -352
rect 18136 328 18152 392
rect 18216 328 18232 392
rect 19548 392 19644 428
rect 18136 312 18232 328
rect 18136 248 18152 312
rect 18216 248 18232 312
rect 18136 232 18232 248
rect 18136 168 18152 232
rect 18216 168 18232 232
rect 18136 152 18232 168
rect 18136 88 18152 152
rect 18216 88 18232 152
rect 18136 72 18232 88
rect 18136 8 18152 72
rect 18216 8 18232 72
rect 18136 -8 18232 8
rect 18136 -72 18152 -8
rect 18216 -72 18232 -8
rect 18136 -88 18232 -72
rect 18136 -152 18152 -88
rect 18216 -152 18232 -88
rect 18136 -168 18232 -152
rect 18136 -232 18152 -168
rect 18216 -232 18232 -168
rect 18136 -248 18232 -232
rect 18136 -312 18152 -248
rect 18216 -312 18232 -248
rect 18136 -328 18232 -312
rect 16724 -428 16820 -392
rect 18136 -392 18152 -328
rect 18216 -392 18232 -328
rect 18555 352 19277 361
rect 18555 -352 18564 352
rect 19268 -352 19277 352
rect 18555 -361 19277 -352
rect 19548 328 19564 392
rect 19628 328 19644 392
rect 20960 392 21056 428
rect 19548 312 19644 328
rect 19548 248 19564 312
rect 19628 248 19644 312
rect 19548 232 19644 248
rect 19548 168 19564 232
rect 19628 168 19644 232
rect 19548 152 19644 168
rect 19548 88 19564 152
rect 19628 88 19644 152
rect 19548 72 19644 88
rect 19548 8 19564 72
rect 19628 8 19644 72
rect 19548 -8 19644 8
rect 19548 -72 19564 -8
rect 19628 -72 19644 -8
rect 19548 -88 19644 -72
rect 19548 -152 19564 -88
rect 19628 -152 19644 -88
rect 19548 -168 19644 -152
rect 19548 -232 19564 -168
rect 19628 -232 19644 -168
rect 19548 -248 19644 -232
rect 19548 -312 19564 -248
rect 19628 -312 19644 -248
rect 19548 -328 19644 -312
rect 18136 -428 18232 -392
rect 19548 -392 19564 -328
rect 19628 -392 19644 -328
rect 19967 352 20689 361
rect 19967 -352 19976 352
rect 20680 -352 20689 352
rect 19967 -361 20689 -352
rect 20960 328 20976 392
rect 21040 328 21056 392
rect 22372 392 22468 428
rect 20960 312 21056 328
rect 20960 248 20976 312
rect 21040 248 21056 312
rect 20960 232 21056 248
rect 20960 168 20976 232
rect 21040 168 21056 232
rect 20960 152 21056 168
rect 20960 88 20976 152
rect 21040 88 21056 152
rect 20960 72 21056 88
rect 20960 8 20976 72
rect 21040 8 21056 72
rect 20960 -8 21056 8
rect 20960 -72 20976 -8
rect 21040 -72 21056 -8
rect 20960 -88 21056 -72
rect 20960 -152 20976 -88
rect 21040 -152 21056 -88
rect 20960 -168 21056 -152
rect 20960 -232 20976 -168
rect 21040 -232 21056 -168
rect 20960 -248 21056 -232
rect 20960 -312 20976 -248
rect 21040 -312 21056 -248
rect 20960 -328 21056 -312
rect 19548 -428 19644 -392
rect 20960 -392 20976 -328
rect 21040 -392 21056 -328
rect 21379 352 22101 361
rect 21379 -352 21388 352
rect 22092 -352 22101 352
rect 21379 -361 22101 -352
rect 22372 328 22388 392
rect 22452 328 22468 392
rect 23784 392 23880 428
rect 22372 312 22468 328
rect 22372 248 22388 312
rect 22452 248 22468 312
rect 22372 232 22468 248
rect 22372 168 22388 232
rect 22452 168 22468 232
rect 22372 152 22468 168
rect 22372 88 22388 152
rect 22452 88 22468 152
rect 22372 72 22468 88
rect 22372 8 22388 72
rect 22452 8 22468 72
rect 22372 -8 22468 8
rect 22372 -72 22388 -8
rect 22452 -72 22468 -8
rect 22372 -88 22468 -72
rect 22372 -152 22388 -88
rect 22452 -152 22468 -88
rect 22372 -168 22468 -152
rect 22372 -232 22388 -168
rect 22452 -232 22468 -168
rect 22372 -248 22468 -232
rect 22372 -312 22388 -248
rect 22452 -312 22468 -248
rect 22372 -328 22468 -312
rect 20960 -428 21056 -392
rect 22372 -392 22388 -328
rect 22452 -392 22468 -328
rect 22791 352 23513 361
rect 22791 -352 22800 352
rect 23504 -352 23513 352
rect 22791 -361 23513 -352
rect 23784 328 23800 392
rect 23864 328 23880 392
rect 23784 312 23880 328
rect 23784 248 23800 312
rect 23864 248 23880 312
rect 23784 232 23880 248
rect 23784 168 23800 232
rect 23864 168 23880 232
rect 23784 152 23880 168
rect 23784 88 23800 152
rect 23864 88 23880 152
rect 23784 72 23880 88
rect 23784 8 23800 72
rect 23864 8 23880 72
rect 23784 -8 23880 8
rect 23784 -72 23800 -8
rect 23864 -72 23880 -8
rect 23784 -88 23880 -72
rect 23784 -152 23800 -88
rect 23864 -152 23880 -88
rect 23784 -168 23880 -152
rect 23784 -232 23800 -168
rect 23864 -232 23880 -168
rect 23784 -248 23880 -232
rect 23784 -312 23800 -248
rect 23864 -312 23880 -248
rect 23784 -328 23880 -312
rect 22372 -428 22468 -392
rect 23784 -392 23800 -328
rect 23864 -392 23880 -328
rect 23784 -428 23880 -392
rect -22812 -728 -22716 -692
rect -23805 -768 -23083 -759
rect -23805 -1472 -23796 -768
rect -23092 -1472 -23083 -768
rect -23805 -1481 -23083 -1472
rect -22812 -792 -22796 -728
rect -22732 -792 -22716 -728
rect -21400 -728 -21304 -692
rect -22812 -808 -22716 -792
rect -22812 -872 -22796 -808
rect -22732 -872 -22716 -808
rect -22812 -888 -22716 -872
rect -22812 -952 -22796 -888
rect -22732 -952 -22716 -888
rect -22812 -968 -22716 -952
rect -22812 -1032 -22796 -968
rect -22732 -1032 -22716 -968
rect -22812 -1048 -22716 -1032
rect -22812 -1112 -22796 -1048
rect -22732 -1112 -22716 -1048
rect -22812 -1128 -22716 -1112
rect -22812 -1192 -22796 -1128
rect -22732 -1192 -22716 -1128
rect -22812 -1208 -22716 -1192
rect -22812 -1272 -22796 -1208
rect -22732 -1272 -22716 -1208
rect -22812 -1288 -22716 -1272
rect -22812 -1352 -22796 -1288
rect -22732 -1352 -22716 -1288
rect -22812 -1368 -22716 -1352
rect -22812 -1432 -22796 -1368
rect -22732 -1432 -22716 -1368
rect -22812 -1448 -22716 -1432
rect -22812 -1512 -22796 -1448
rect -22732 -1512 -22716 -1448
rect -22393 -768 -21671 -759
rect -22393 -1472 -22384 -768
rect -21680 -1472 -21671 -768
rect -22393 -1481 -21671 -1472
rect -21400 -792 -21384 -728
rect -21320 -792 -21304 -728
rect -19988 -728 -19892 -692
rect -21400 -808 -21304 -792
rect -21400 -872 -21384 -808
rect -21320 -872 -21304 -808
rect -21400 -888 -21304 -872
rect -21400 -952 -21384 -888
rect -21320 -952 -21304 -888
rect -21400 -968 -21304 -952
rect -21400 -1032 -21384 -968
rect -21320 -1032 -21304 -968
rect -21400 -1048 -21304 -1032
rect -21400 -1112 -21384 -1048
rect -21320 -1112 -21304 -1048
rect -21400 -1128 -21304 -1112
rect -21400 -1192 -21384 -1128
rect -21320 -1192 -21304 -1128
rect -21400 -1208 -21304 -1192
rect -21400 -1272 -21384 -1208
rect -21320 -1272 -21304 -1208
rect -21400 -1288 -21304 -1272
rect -21400 -1352 -21384 -1288
rect -21320 -1352 -21304 -1288
rect -21400 -1368 -21304 -1352
rect -21400 -1432 -21384 -1368
rect -21320 -1432 -21304 -1368
rect -21400 -1448 -21304 -1432
rect -22812 -1548 -22716 -1512
rect -21400 -1512 -21384 -1448
rect -21320 -1512 -21304 -1448
rect -20981 -768 -20259 -759
rect -20981 -1472 -20972 -768
rect -20268 -1472 -20259 -768
rect -20981 -1481 -20259 -1472
rect -19988 -792 -19972 -728
rect -19908 -792 -19892 -728
rect -18576 -728 -18480 -692
rect -19988 -808 -19892 -792
rect -19988 -872 -19972 -808
rect -19908 -872 -19892 -808
rect -19988 -888 -19892 -872
rect -19988 -952 -19972 -888
rect -19908 -952 -19892 -888
rect -19988 -968 -19892 -952
rect -19988 -1032 -19972 -968
rect -19908 -1032 -19892 -968
rect -19988 -1048 -19892 -1032
rect -19988 -1112 -19972 -1048
rect -19908 -1112 -19892 -1048
rect -19988 -1128 -19892 -1112
rect -19988 -1192 -19972 -1128
rect -19908 -1192 -19892 -1128
rect -19988 -1208 -19892 -1192
rect -19988 -1272 -19972 -1208
rect -19908 -1272 -19892 -1208
rect -19988 -1288 -19892 -1272
rect -19988 -1352 -19972 -1288
rect -19908 -1352 -19892 -1288
rect -19988 -1368 -19892 -1352
rect -19988 -1432 -19972 -1368
rect -19908 -1432 -19892 -1368
rect -19988 -1448 -19892 -1432
rect -21400 -1548 -21304 -1512
rect -19988 -1512 -19972 -1448
rect -19908 -1512 -19892 -1448
rect -19569 -768 -18847 -759
rect -19569 -1472 -19560 -768
rect -18856 -1472 -18847 -768
rect -19569 -1481 -18847 -1472
rect -18576 -792 -18560 -728
rect -18496 -792 -18480 -728
rect -17164 -728 -17068 -692
rect -18576 -808 -18480 -792
rect -18576 -872 -18560 -808
rect -18496 -872 -18480 -808
rect -18576 -888 -18480 -872
rect -18576 -952 -18560 -888
rect -18496 -952 -18480 -888
rect -18576 -968 -18480 -952
rect -18576 -1032 -18560 -968
rect -18496 -1032 -18480 -968
rect -18576 -1048 -18480 -1032
rect -18576 -1112 -18560 -1048
rect -18496 -1112 -18480 -1048
rect -18576 -1128 -18480 -1112
rect -18576 -1192 -18560 -1128
rect -18496 -1192 -18480 -1128
rect -18576 -1208 -18480 -1192
rect -18576 -1272 -18560 -1208
rect -18496 -1272 -18480 -1208
rect -18576 -1288 -18480 -1272
rect -18576 -1352 -18560 -1288
rect -18496 -1352 -18480 -1288
rect -18576 -1368 -18480 -1352
rect -18576 -1432 -18560 -1368
rect -18496 -1432 -18480 -1368
rect -18576 -1448 -18480 -1432
rect -19988 -1548 -19892 -1512
rect -18576 -1512 -18560 -1448
rect -18496 -1512 -18480 -1448
rect -18157 -768 -17435 -759
rect -18157 -1472 -18148 -768
rect -17444 -1472 -17435 -768
rect -18157 -1481 -17435 -1472
rect -17164 -792 -17148 -728
rect -17084 -792 -17068 -728
rect -15752 -728 -15656 -692
rect -17164 -808 -17068 -792
rect -17164 -872 -17148 -808
rect -17084 -872 -17068 -808
rect -17164 -888 -17068 -872
rect -17164 -952 -17148 -888
rect -17084 -952 -17068 -888
rect -17164 -968 -17068 -952
rect -17164 -1032 -17148 -968
rect -17084 -1032 -17068 -968
rect -17164 -1048 -17068 -1032
rect -17164 -1112 -17148 -1048
rect -17084 -1112 -17068 -1048
rect -17164 -1128 -17068 -1112
rect -17164 -1192 -17148 -1128
rect -17084 -1192 -17068 -1128
rect -17164 -1208 -17068 -1192
rect -17164 -1272 -17148 -1208
rect -17084 -1272 -17068 -1208
rect -17164 -1288 -17068 -1272
rect -17164 -1352 -17148 -1288
rect -17084 -1352 -17068 -1288
rect -17164 -1368 -17068 -1352
rect -17164 -1432 -17148 -1368
rect -17084 -1432 -17068 -1368
rect -17164 -1448 -17068 -1432
rect -18576 -1548 -18480 -1512
rect -17164 -1512 -17148 -1448
rect -17084 -1512 -17068 -1448
rect -16745 -768 -16023 -759
rect -16745 -1472 -16736 -768
rect -16032 -1472 -16023 -768
rect -16745 -1481 -16023 -1472
rect -15752 -792 -15736 -728
rect -15672 -792 -15656 -728
rect -14340 -728 -14244 -692
rect -15752 -808 -15656 -792
rect -15752 -872 -15736 -808
rect -15672 -872 -15656 -808
rect -15752 -888 -15656 -872
rect -15752 -952 -15736 -888
rect -15672 -952 -15656 -888
rect -15752 -968 -15656 -952
rect -15752 -1032 -15736 -968
rect -15672 -1032 -15656 -968
rect -15752 -1048 -15656 -1032
rect -15752 -1112 -15736 -1048
rect -15672 -1112 -15656 -1048
rect -15752 -1128 -15656 -1112
rect -15752 -1192 -15736 -1128
rect -15672 -1192 -15656 -1128
rect -15752 -1208 -15656 -1192
rect -15752 -1272 -15736 -1208
rect -15672 -1272 -15656 -1208
rect -15752 -1288 -15656 -1272
rect -15752 -1352 -15736 -1288
rect -15672 -1352 -15656 -1288
rect -15752 -1368 -15656 -1352
rect -15752 -1432 -15736 -1368
rect -15672 -1432 -15656 -1368
rect -15752 -1448 -15656 -1432
rect -17164 -1548 -17068 -1512
rect -15752 -1512 -15736 -1448
rect -15672 -1512 -15656 -1448
rect -15333 -768 -14611 -759
rect -15333 -1472 -15324 -768
rect -14620 -1472 -14611 -768
rect -15333 -1481 -14611 -1472
rect -14340 -792 -14324 -728
rect -14260 -792 -14244 -728
rect -12928 -728 -12832 -692
rect -14340 -808 -14244 -792
rect -14340 -872 -14324 -808
rect -14260 -872 -14244 -808
rect -14340 -888 -14244 -872
rect -14340 -952 -14324 -888
rect -14260 -952 -14244 -888
rect -14340 -968 -14244 -952
rect -14340 -1032 -14324 -968
rect -14260 -1032 -14244 -968
rect -14340 -1048 -14244 -1032
rect -14340 -1112 -14324 -1048
rect -14260 -1112 -14244 -1048
rect -14340 -1128 -14244 -1112
rect -14340 -1192 -14324 -1128
rect -14260 -1192 -14244 -1128
rect -14340 -1208 -14244 -1192
rect -14340 -1272 -14324 -1208
rect -14260 -1272 -14244 -1208
rect -14340 -1288 -14244 -1272
rect -14340 -1352 -14324 -1288
rect -14260 -1352 -14244 -1288
rect -14340 -1368 -14244 -1352
rect -14340 -1432 -14324 -1368
rect -14260 -1432 -14244 -1368
rect -14340 -1448 -14244 -1432
rect -15752 -1548 -15656 -1512
rect -14340 -1512 -14324 -1448
rect -14260 -1512 -14244 -1448
rect -13921 -768 -13199 -759
rect -13921 -1472 -13912 -768
rect -13208 -1472 -13199 -768
rect -13921 -1481 -13199 -1472
rect -12928 -792 -12912 -728
rect -12848 -792 -12832 -728
rect -11516 -728 -11420 -692
rect -12928 -808 -12832 -792
rect -12928 -872 -12912 -808
rect -12848 -872 -12832 -808
rect -12928 -888 -12832 -872
rect -12928 -952 -12912 -888
rect -12848 -952 -12832 -888
rect -12928 -968 -12832 -952
rect -12928 -1032 -12912 -968
rect -12848 -1032 -12832 -968
rect -12928 -1048 -12832 -1032
rect -12928 -1112 -12912 -1048
rect -12848 -1112 -12832 -1048
rect -12928 -1128 -12832 -1112
rect -12928 -1192 -12912 -1128
rect -12848 -1192 -12832 -1128
rect -12928 -1208 -12832 -1192
rect -12928 -1272 -12912 -1208
rect -12848 -1272 -12832 -1208
rect -12928 -1288 -12832 -1272
rect -12928 -1352 -12912 -1288
rect -12848 -1352 -12832 -1288
rect -12928 -1368 -12832 -1352
rect -12928 -1432 -12912 -1368
rect -12848 -1432 -12832 -1368
rect -12928 -1448 -12832 -1432
rect -14340 -1548 -14244 -1512
rect -12928 -1512 -12912 -1448
rect -12848 -1512 -12832 -1448
rect -12509 -768 -11787 -759
rect -12509 -1472 -12500 -768
rect -11796 -1472 -11787 -768
rect -12509 -1481 -11787 -1472
rect -11516 -792 -11500 -728
rect -11436 -792 -11420 -728
rect -10104 -728 -10008 -692
rect -11516 -808 -11420 -792
rect -11516 -872 -11500 -808
rect -11436 -872 -11420 -808
rect -11516 -888 -11420 -872
rect -11516 -952 -11500 -888
rect -11436 -952 -11420 -888
rect -11516 -968 -11420 -952
rect -11516 -1032 -11500 -968
rect -11436 -1032 -11420 -968
rect -11516 -1048 -11420 -1032
rect -11516 -1112 -11500 -1048
rect -11436 -1112 -11420 -1048
rect -11516 -1128 -11420 -1112
rect -11516 -1192 -11500 -1128
rect -11436 -1192 -11420 -1128
rect -11516 -1208 -11420 -1192
rect -11516 -1272 -11500 -1208
rect -11436 -1272 -11420 -1208
rect -11516 -1288 -11420 -1272
rect -11516 -1352 -11500 -1288
rect -11436 -1352 -11420 -1288
rect -11516 -1368 -11420 -1352
rect -11516 -1432 -11500 -1368
rect -11436 -1432 -11420 -1368
rect -11516 -1448 -11420 -1432
rect -12928 -1548 -12832 -1512
rect -11516 -1512 -11500 -1448
rect -11436 -1512 -11420 -1448
rect -11097 -768 -10375 -759
rect -11097 -1472 -11088 -768
rect -10384 -1472 -10375 -768
rect -11097 -1481 -10375 -1472
rect -10104 -792 -10088 -728
rect -10024 -792 -10008 -728
rect -8692 -728 -8596 -692
rect -10104 -808 -10008 -792
rect -10104 -872 -10088 -808
rect -10024 -872 -10008 -808
rect -10104 -888 -10008 -872
rect -10104 -952 -10088 -888
rect -10024 -952 -10008 -888
rect -10104 -968 -10008 -952
rect -10104 -1032 -10088 -968
rect -10024 -1032 -10008 -968
rect -10104 -1048 -10008 -1032
rect -10104 -1112 -10088 -1048
rect -10024 -1112 -10008 -1048
rect -10104 -1128 -10008 -1112
rect -10104 -1192 -10088 -1128
rect -10024 -1192 -10008 -1128
rect -10104 -1208 -10008 -1192
rect -10104 -1272 -10088 -1208
rect -10024 -1272 -10008 -1208
rect -10104 -1288 -10008 -1272
rect -10104 -1352 -10088 -1288
rect -10024 -1352 -10008 -1288
rect -10104 -1368 -10008 -1352
rect -10104 -1432 -10088 -1368
rect -10024 -1432 -10008 -1368
rect -10104 -1448 -10008 -1432
rect -11516 -1548 -11420 -1512
rect -10104 -1512 -10088 -1448
rect -10024 -1512 -10008 -1448
rect -9685 -768 -8963 -759
rect -9685 -1472 -9676 -768
rect -8972 -1472 -8963 -768
rect -9685 -1481 -8963 -1472
rect -8692 -792 -8676 -728
rect -8612 -792 -8596 -728
rect -7280 -728 -7184 -692
rect -8692 -808 -8596 -792
rect -8692 -872 -8676 -808
rect -8612 -872 -8596 -808
rect -8692 -888 -8596 -872
rect -8692 -952 -8676 -888
rect -8612 -952 -8596 -888
rect -8692 -968 -8596 -952
rect -8692 -1032 -8676 -968
rect -8612 -1032 -8596 -968
rect -8692 -1048 -8596 -1032
rect -8692 -1112 -8676 -1048
rect -8612 -1112 -8596 -1048
rect -8692 -1128 -8596 -1112
rect -8692 -1192 -8676 -1128
rect -8612 -1192 -8596 -1128
rect -8692 -1208 -8596 -1192
rect -8692 -1272 -8676 -1208
rect -8612 -1272 -8596 -1208
rect -8692 -1288 -8596 -1272
rect -8692 -1352 -8676 -1288
rect -8612 -1352 -8596 -1288
rect -8692 -1368 -8596 -1352
rect -8692 -1432 -8676 -1368
rect -8612 -1432 -8596 -1368
rect -8692 -1448 -8596 -1432
rect -10104 -1548 -10008 -1512
rect -8692 -1512 -8676 -1448
rect -8612 -1512 -8596 -1448
rect -8273 -768 -7551 -759
rect -8273 -1472 -8264 -768
rect -7560 -1472 -7551 -768
rect -8273 -1481 -7551 -1472
rect -7280 -792 -7264 -728
rect -7200 -792 -7184 -728
rect -5868 -728 -5772 -692
rect -7280 -808 -7184 -792
rect -7280 -872 -7264 -808
rect -7200 -872 -7184 -808
rect -7280 -888 -7184 -872
rect -7280 -952 -7264 -888
rect -7200 -952 -7184 -888
rect -7280 -968 -7184 -952
rect -7280 -1032 -7264 -968
rect -7200 -1032 -7184 -968
rect -7280 -1048 -7184 -1032
rect -7280 -1112 -7264 -1048
rect -7200 -1112 -7184 -1048
rect -7280 -1128 -7184 -1112
rect -7280 -1192 -7264 -1128
rect -7200 -1192 -7184 -1128
rect -7280 -1208 -7184 -1192
rect -7280 -1272 -7264 -1208
rect -7200 -1272 -7184 -1208
rect -7280 -1288 -7184 -1272
rect -7280 -1352 -7264 -1288
rect -7200 -1352 -7184 -1288
rect -7280 -1368 -7184 -1352
rect -7280 -1432 -7264 -1368
rect -7200 -1432 -7184 -1368
rect -7280 -1448 -7184 -1432
rect -8692 -1548 -8596 -1512
rect -7280 -1512 -7264 -1448
rect -7200 -1512 -7184 -1448
rect -6861 -768 -6139 -759
rect -6861 -1472 -6852 -768
rect -6148 -1472 -6139 -768
rect -6861 -1481 -6139 -1472
rect -5868 -792 -5852 -728
rect -5788 -792 -5772 -728
rect -4456 -728 -4360 -692
rect -5868 -808 -5772 -792
rect -5868 -872 -5852 -808
rect -5788 -872 -5772 -808
rect -5868 -888 -5772 -872
rect -5868 -952 -5852 -888
rect -5788 -952 -5772 -888
rect -5868 -968 -5772 -952
rect -5868 -1032 -5852 -968
rect -5788 -1032 -5772 -968
rect -5868 -1048 -5772 -1032
rect -5868 -1112 -5852 -1048
rect -5788 -1112 -5772 -1048
rect -5868 -1128 -5772 -1112
rect -5868 -1192 -5852 -1128
rect -5788 -1192 -5772 -1128
rect -5868 -1208 -5772 -1192
rect -5868 -1272 -5852 -1208
rect -5788 -1272 -5772 -1208
rect -5868 -1288 -5772 -1272
rect -5868 -1352 -5852 -1288
rect -5788 -1352 -5772 -1288
rect -5868 -1368 -5772 -1352
rect -5868 -1432 -5852 -1368
rect -5788 -1432 -5772 -1368
rect -5868 -1448 -5772 -1432
rect -7280 -1548 -7184 -1512
rect -5868 -1512 -5852 -1448
rect -5788 -1512 -5772 -1448
rect -5449 -768 -4727 -759
rect -5449 -1472 -5440 -768
rect -4736 -1472 -4727 -768
rect -5449 -1481 -4727 -1472
rect -4456 -792 -4440 -728
rect -4376 -792 -4360 -728
rect -3044 -728 -2948 -692
rect -4456 -808 -4360 -792
rect -4456 -872 -4440 -808
rect -4376 -872 -4360 -808
rect -4456 -888 -4360 -872
rect -4456 -952 -4440 -888
rect -4376 -952 -4360 -888
rect -4456 -968 -4360 -952
rect -4456 -1032 -4440 -968
rect -4376 -1032 -4360 -968
rect -4456 -1048 -4360 -1032
rect -4456 -1112 -4440 -1048
rect -4376 -1112 -4360 -1048
rect -4456 -1128 -4360 -1112
rect -4456 -1192 -4440 -1128
rect -4376 -1192 -4360 -1128
rect -4456 -1208 -4360 -1192
rect -4456 -1272 -4440 -1208
rect -4376 -1272 -4360 -1208
rect -4456 -1288 -4360 -1272
rect -4456 -1352 -4440 -1288
rect -4376 -1352 -4360 -1288
rect -4456 -1368 -4360 -1352
rect -4456 -1432 -4440 -1368
rect -4376 -1432 -4360 -1368
rect -4456 -1448 -4360 -1432
rect -5868 -1548 -5772 -1512
rect -4456 -1512 -4440 -1448
rect -4376 -1512 -4360 -1448
rect -4037 -768 -3315 -759
rect -4037 -1472 -4028 -768
rect -3324 -1472 -3315 -768
rect -4037 -1481 -3315 -1472
rect -3044 -792 -3028 -728
rect -2964 -792 -2948 -728
rect -1632 -728 -1536 -692
rect -3044 -808 -2948 -792
rect -3044 -872 -3028 -808
rect -2964 -872 -2948 -808
rect -3044 -888 -2948 -872
rect -3044 -952 -3028 -888
rect -2964 -952 -2948 -888
rect -3044 -968 -2948 -952
rect -3044 -1032 -3028 -968
rect -2964 -1032 -2948 -968
rect -3044 -1048 -2948 -1032
rect -3044 -1112 -3028 -1048
rect -2964 -1112 -2948 -1048
rect -3044 -1128 -2948 -1112
rect -3044 -1192 -3028 -1128
rect -2964 -1192 -2948 -1128
rect -3044 -1208 -2948 -1192
rect -3044 -1272 -3028 -1208
rect -2964 -1272 -2948 -1208
rect -3044 -1288 -2948 -1272
rect -3044 -1352 -3028 -1288
rect -2964 -1352 -2948 -1288
rect -3044 -1368 -2948 -1352
rect -3044 -1432 -3028 -1368
rect -2964 -1432 -2948 -1368
rect -3044 -1448 -2948 -1432
rect -4456 -1548 -4360 -1512
rect -3044 -1512 -3028 -1448
rect -2964 -1512 -2948 -1448
rect -2625 -768 -1903 -759
rect -2625 -1472 -2616 -768
rect -1912 -1472 -1903 -768
rect -2625 -1481 -1903 -1472
rect -1632 -792 -1616 -728
rect -1552 -792 -1536 -728
rect -220 -728 -124 -692
rect -1632 -808 -1536 -792
rect -1632 -872 -1616 -808
rect -1552 -872 -1536 -808
rect -1632 -888 -1536 -872
rect -1632 -952 -1616 -888
rect -1552 -952 -1536 -888
rect -1632 -968 -1536 -952
rect -1632 -1032 -1616 -968
rect -1552 -1032 -1536 -968
rect -1632 -1048 -1536 -1032
rect -1632 -1112 -1616 -1048
rect -1552 -1112 -1536 -1048
rect -1632 -1128 -1536 -1112
rect -1632 -1192 -1616 -1128
rect -1552 -1192 -1536 -1128
rect -1632 -1208 -1536 -1192
rect -1632 -1272 -1616 -1208
rect -1552 -1272 -1536 -1208
rect -1632 -1288 -1536 -1272
rect -1632 -1352 -1616 -1288
rect -1552 -1352 -1536 -1288
rect -1632 -1368 -1536 -1352
rect -1632 -1432 -1616 -1368
rect -1552 -1432 -1536 -1368
rect -1632 -1448 -1536 -1432
rect -3044 -1548 -2948 -1512
rect -1632 -1512 -1616 -1448
rect -1552 -1512 -1536 -1448
rect -1213 -768 -491 -759
rect -1213 -1472 -1204 -768
rect -500 -1472 -491 -768
rect -1213 -1481 -491 -1472
rect -220 -792 -204 -728
rect -140 -792 -124 -728
rect 1192 -728 1288 -692
rect -220 -808 -124 -792
rect -220 -872 -204 -808
rect -140 -872 -124 -808
rect -220 -888 -124 -872
rect -220 -952 -204 -888
rect -140 -952 -124 -888
rect -220 -968 -124 -952
rect -220 -1032 -204 -968
rect -140 -1032 -124 -968
rect -220 -1048 -124 -1032
rect -220 -1112 -204 -1048
rect -140 -1112 -124 -1048
rect -220 -1128 -124 -1112
rect -220 -1192 -204 -1128
rect -140 -1192 -124 -1128
rect -220 -1208 -124 -1192
rect -220 -1272 -204 -1208
rect -140 -1272 -124 -1208
rect -220 -1288 -124 -1272
rect -220 -1352 -204 -1288
rect -140 -1352 -124 -1288
rect -220 -1368 -124 -1352
rect -220 -1432 -204 -1368
rect -140 -1432 -124 -1368
rect -220 -1448 -124 -1432
rect -1632 -1548 -1536 -1512
rect -220 -1512 -204 -1448
rect -140 -1512 -124 -1448
rect 199 -768 921 -759
rect 199 -1472 208 -768
rect 912 -1472 921 -768
rect 199 -1481 921 -1472
rect 1192 -792 1208 -728
rect 1272 -792 1288 -728
rect 2604 -728 2700 -692
rect 1192 -808 1288 -792
rect 1192 -872 1208 -808
rect 1272 -872 1288 -808
rect 1192 -888 1288 -872
rect 1192 -952 1208 -888
rect 1272 -952 1288 -888
rect 1192 -968 1288 -952
rect 1192 -1032 1208 -968
rect 1272 -1032 1288 -968
rect 1192 -1048 1288 -1032
rect 1192 -1112 1208 -1048
rect 1272 -1112 1288 -1048
rect 1192 -1128 1288 -1112
rect 1192 -1192 1208 -1128
rect 1272 -1192 1288 -1128
rect 1192 -1208 1288 -1192
rect 1192 -1272 1208 -1208
rect 1272 -1272 1288 -1208
rect 1192 -1288 1288 -1272
rect 1192 -1352 1208 -1288
rect 1272 -1352 1288 -1288
rect 1192 -1368 1288 -1352
rect 1192 -1432 1208 -1368
rect 1272 -1432 1288 -1368
rect 1192 -1448 1288 -1432
rect -220 -1548 -124 -1512
rect 1192 -1512 1208 -1448
rect 1272 -1512 1288 -1448
rect 1611 -768 2333 -759
rect 1611 -1472 1620 -768
rect 2324 -1472 2333 -768
rect 1611 -1481 2333 -1472
rect 2604 -792 2620 -728
rect 2684 -792 2700 -728
rect 4016 -728 4112 -692
rect 2604 -808 2700 -792
rect 2604 -872 2620 -808
rect 2684 -872 2700 -808
rect 2604 -888 2700 -872
rect 2604 -952 2620 -888
rect 2684 -952 2700 -888
rect 2604 -968 2700 -952
rect 2604 -1032 2620 -968
rect 2684 -1032 2700 -968
rect 2604 -1048 2700 -1032
rect 2604 -1112 2620 -1048
rect 2684 -1112 2700 -1048
rect 2604 -1128 2700 -1112
rect 2604 -1192 2620 -1128
rect 2684 -1192 2700 -1128
rect 2604 -1208 2700 -1192
rect 2604 -1272 2620 -1208
rect 2684 -1272 2700 -1208
rect 2604 -1288 2700 -1272
rect 2604 -1352 2620 -1288
rect 2684 -1352 2700 -1288
rect 2604 -1368 2700 -1352
rect 2604 -1432 2620 -1368
rect 2684 -1432 2700 -1368
rect 2604 -1448 2700 -1432
rect 1192 -1548 1288 -1512
rect 2604 -1512 2620 -1448
rect 2684 -1512 2700 -1448
rect 3023 -768 3745 -759
rect 3023 -1472 3032 -768
rect 3736 -1472 3745 -768
rect 3023 -1481 3745 -1472
rect 4016 -792 4032 -728
rect 4096 -792 4112 -728
rect 5428 -728 5524 -692
rect 4016 -808 4112 -792
rect 4016 -872 4032 -808
rect 4096 -872 4112 -808
rect 4016 -888 4112 -872
rect 4016 -952 4032 -888
rect 4096 -952 4112 -888
rect 4016 -968 4112 -952
rect 4016 -1032 4032 -968
rect 4096 -1032 4112 -968
rect 4016 -1048 4112 -1032
rect 4016 -1112 4032 -1048
rect 4096 -1112 4112 -1048
rect 4016 -1128 4112 -1112
rect 4016 -1192 4032 -1128
rect 4096 -1192 4112 -1128
rect 4016 -1208 4112 -1192
rect 4016 -1272 4032 -1208
rect 4096 -1272 4112 -1208
rect 4016 -1288 4112 -1272
rect 4016 -1352 4032 -1288
rect 4096 -1352 4112 -1288
rect 4016 -1368 4112 -1352
rect 4016 -1432 4032 -1368
rect 4096 -1432 4112 -1368
rect 4016 -1448 4112 -1432
rect 2604 -1548 2700 -1512
rect 4016 -1512 4032 -1448
rect 4096 -1512 4112 -1448
rect 4435 -768 5157 -759
rect 4435 -1472 4444 -768
rect 5148 -1472 5157 -768
rect 4435 -1481 5157 -1472
rect 5428 -792 5444 -728
rect 5508 -792 5524 -728
rect 6840 -728 6936 -692
rect 5428 -808 5524 -792
rect 5428 -872 5444 -808
rect 5508 -872 5524 -808
rect 5428 -888 5524 -872
rect 5428 -952 5444 -888
rect 5508 -952 5524 -888
rect 5428 -968 5524 -952
rect 5428 -1032 5444 -968
rect 5508 -1032 5524 -968
rect 5428 -1048 5524 -1032
rect 5428 -1112 5444 -1048
rect 5508 -1112 5524 -1048
rect 5428 -1128 5524 -1112
rect 5428 -1192 5444 -1128
rect 5508 -1192 5524 -1128
rect 5428 -1208 5524 -1192
rect 5428 -1272 5444 -1208
rect 5508 -1272 5524 -1208
rect 5428 -1288 5524 -1272
rect 5428 -1352 5444 -1288
rect 5508 -1352 5524 -1288
rect 5428 -1368 5524 -1352
rect 5428 -1432 5444 -1368
rect 5508 -1432 5524 -1368
rect 5428 -1448 5524 -1432
rect 4016 -1548 4112 -1512
rect 5428 -1512 5444 -1448
rect 5508 -1512 5524 -1448
rect 5847 -768 6569 -759
rect 5847 -1472 5856 -768
rect 6560 -1472 6569 -768
rect 5847 -1481 6569 -1472
rect 6840 -792 6856 -728
rect 6920 -792 6936 -728
rect 8252 -728 8348 -692
rect 6840 -808 6936 -792
rect 6840 -872 6856 -808
rect 6920 -872 6936 -808
rect 6840 -888 6936 -872
rect 6840 -952 6856 -888
rect 6920 -952 6936 -888
rect 6840 -968 6936 -952
rect 6840 -1032 6856 -968
rect 6920 -1032 6936 -968
rect 6840 -1048 6936 -1032
rect 6840 -1112 6856 -1048
rect 6920 -1112 6936 -1048
rect 6840 -1128 6936 -1112
rect 6840 -1192 6856 -1128
rect 6920 -1192 6936 -1128
rect 6840 -1208 6936 -1192
rect 6840 -1272 6856 -1208
rect 6920 -1272 6936 -1208
rect 6840 -1288 6936 -1272
rect 6840 -1352 6856 -1288
rect 6920 -1352 6936 -1288
rect 6840 -1368 6936 -1352
rect 6840 -1432 6856 -1368
rect 6920 -1432 6936 -1368
rect 6840 -1448 6936 -1432
rect 5428 -1548 5524 -1512
rect 6840 -1512 6856 -1448
rect 6920 -1512 6936 -1448
rect 7259 -768 7981 -759
rect 7259 -1472 7268 -768
rect 7972 -1472 7981 -768
rect 7259 -1481 7981 -1472
rect 8252 -792 8268 -728
rect 8332 -792 8348 -728
rect 9664 -728 9760 -692
rect 8252 -808 8348 -792
rect 8252 -872 8268 -808
rect 8332 -872 8348 -808
rect 8252 -888 8348 -872
rect 8252 -952 8268 -888
rect 8332 -952 8348 -888
rect 8252 -968 8348 -952
rect 8252 -1032 8268 -968
rect 8332 -1032 8348 -968
rect 8252 -1048 8348 -1032
rect 8252 -1112 8268 -1048
rect 8332 -1112 8348 -1048
rect 8252 -1128 8348 -1112
rect 8252 -1192 8268 -1128
rect 8332 -1192 8348 -1128
rect 8252 -1208 8348 -1192
rect 8252 -1272 8268 -1208
rect 8332 -1272 8348 -1208
rect 8252 -1288 8348 -1272
rect 8252 -1352 8268 -1288
rect 8332 -1352 8348 -1288
rect 8252 -1368 8348 -1352
rect 8252 -1432 8268 -1368
rect 8332 -1432 8348 -1368
rect 8252 -1448 8348 -1432
rect 6840 -1548 6936 -1512
rect 8252 -1512 8268 -1448
rect 8332 -1512 8348 -1448
rect 8671 -768 9393 -759
rect 8671 -1472 8680 -768
rect 9384 -1472 9393 -768
rect 8671 -1481 9393 -1472
rect 9664 -792 9680 -728
rect 9744 -792 9760 -728
rect 11076 -728 11172 -692
rect 9664 -808 9760 -792
rect 9664 -872 9680 -808
rect 9744 -872 9760 -808
rect 9664 -888 9760 -872
rect 9664 -952 9680 -888
rect 9744 -952 9760 -888
rect 9664 -968 9760 -952
rect 9664 -1032 9680 -968
rect 9744 -1032 9760 -968
rect 9664 -1048 9760 -1032
rect 9664 -1112 9680 -1048
rect 9744 -1112 9760 -1048
rect 9664 -1128 9760 -1112
rect 9664 -1192 9680 -1128
rect 9744 -1192 9760 -1128
rect 9664 -1208 9760 -1192
rect 9664 -1272 9680 -1208
rect 9744 -1272 9760 -1208
rect 9664 -1288 9760 -1272
rect 9664 -1352 9680 -1288
rect 9744 -1352 9760 -1288
rect 9664 -1368 9760 -1352
rect 9664 -1432 9680 -1368
rect 9744 -1432 9760 -1368
rect 9664 -1448 9760 -1432
rect 8252 -1548 8348 -1512
rect 9664 -1512 9680 -1448
rect 9744 -1512 9760 -1448
rect 10083 -768 10805 -759
rect 10083 -1472 10092 -768
rect 10796 -1472 10805 -768
rect 10083 -1481 10805 -1472
rect 11076 -792 11092 -728
rect 11156 -792 11172 -728
rect 12488 -728 12584 -692
rect 11076 -808 11172 -792
rect 11076 -872 11092 -808
rect 11156 -872 11172 -808
rect 11076 -888 11172 -872
rect 11076 -952 11092 -888
rect 11156 -952 11172 -888
rect 11076 -968 11172 -952
rect 11076 -1032 11092 -968
rect 11156 -1032 11172 -968
rect 11076 -1048 11172 -1032
rect 11076 -1112 11092 -1048
rect 11156 -1112 11172 -1048
rect 11076 -1128 11172 -1112
rect 11076 -1192 11092 -1128
rect 11156 -1192 11172 -1128
rect 11076 -1208 11172 -1192
rect 11076 -1272 11092 -1208
rect 11156 -1272 11172 -1208
rect 11076 -1288 11172 -1272
rect 11076 -1352 11092 -1288
rect 11156 -1352 11172 -1288
rect 11076 -1368 11172 -1352
rect 11076 -1432 11092 -1368
rect 11156 -1432 11172 -1368
rect 11076 -1448 11172 -1432
rect 9664 -1548 9760 -1512
rect 11076 -1512 11092 -1448
rect 11156 -1512 11172 -1448
rect 11495 -768 12217 -759
rect 11495 -1472 11504 -768
rect 12208 -1472 12217 -768
rect 11495 -1481 12217 -1472
rect 12488 -792 12504 -728
rect 12568 -792 12584 -728
rect 13900 -728 13996 -692
rect 12488 -808 12584 -792
rect 12488 -872 12504 -808
rect 12568 -872 12584 -808
rect 12488 -888 12584 -872
rect 12488 -952 12504 -888
rect 12568 -952 12584 -888
rect 12488 -968 12584 -952
rect 12488 -1032 12504 -968
rect 12568 -1032 12584 -968
rect 12488 -1048 12584 -1032
rect 12488 -1112 12504 -1048
rect 12568 -1112 12584 -1048
rect 12488 -1128 12584 -1112
rect 12488 -1192 12504 -1128
rect 12568 -1192 12584 -1128
rect 12488 -1208 12584 -1192
rect 12488 -1272 12504 -1208
rect 12568 -1272 12584 -1208
rect 12488 -1288 12584 -1272
rect 12488 -1352 12504 -1288
rect 12568 -1352 12584 -1288
rect 12488 -1368 12584 -1352
rect 12488 -1432 12504 -1368
rect 12568 -1432 12584 -1368
rect 12488 -1448 12584 -1432
rect 11076 -1548 11172 -1512
rect 12488 -1512 12504 -1448
rect 12568 -1512 12584 -1448
rect 12907 -768 13629 -759
rect 12907 -1472 12916 -768
rect 13620 -1472 13629 -768
rect 12907 -1481 13629 -1472
rect 13900 -792 13916 -728
rect 13980 -792 13996 -728
rect 15312 -728 15408 -692
rect 13900 -808 13996 -792
rect 13900 -872 13916 -808
rect 13980 -872 13996 -808
rect 13900 -888 13996 -872
rect 13900 -952 13916 -888
rect 13980 -952 13996 -888
rect 13900 -968 13996 -952
rect 13900 -1032 13916 -968
rect 13980 -1032 13996 -968
rect 13900 -1048 13996 -1032
rect 13900 -1112 13916 -1048
rect 13980 -1112 13996 -1048
rect 13900 -1128 13996 -1112
rect 13900 -1192 13916 -1128
rect 13980 -1192 13996 -1128
rect 13900 -1208 13996 -1192
rect 13900 -1272 13916 -1208
rect 13980 -1272 13996 -1208
rect 13900 -1288 13996 -1272
rect 13900 -1352 13916 -1288
rect 13980 -1352 13996 -1288
rect 13900 -1368 13996 -1352
rect 13900 -1432 13916 -1368
rect 13980 -1432 13996 -1368
rect 13900 -1448 13996 -1432
rect 12488 -1548 12584 -1512
rect 13900 -1512 13916 -1448
rect 13980 -1512 13996 -1448
rect 14319 -768 15041 -759
rect 14319 -1472 14328 -768
rect 15032 -1472 15041 -768
rect 14319 -1481 15041 -1472
rect 15312 -792 15328 -728
rect 15392 -792 15408 -728
rect 16724 -728 16820 -692
rect 15312 -808 15408 -792
rect 15312 -872 15328 -808
rect 15392 -872 15408 -808
rect 15312 -888 15408 -872
rect 15312 -952 15328 -888
rect 15392 -952 15408 -888
rect 15312 -968 15408 -952
rect 15312 -1032 15328 -968
rect 15392 -1032 15408 -968
rect 15312 -1048 15408 -1032
rect 15312 -1112 15328 -1048
rect 15392 -1112 15408 -1048
rect 15312 -1128 15408 -1112
rect 15312 -1192 15328 -1128
rect 15392 -1192 15408 -1128
rect 15312 -1208 15408 -1192
rect 15312 -1272 15328 -1208
rect 15392 -1272 15408 -1208
rect 15312 -1288 15408 -1272
rect 15312 -1352 15328 -1288
rect 15392 -1352 15408 -1288
rect 15312 -1368 15408 -1352
rect 15312 -1432 15328 -1368
rect 15392 -1432 15408 -1368
rect 15312 -1448 15408 -1432
rect 13900 -1548 13996 -1512
rect 15312 -1512 15328 -1448
rect 15392 -1512 15408 -1448
rect 15731 -768 16453 -759
rect 15731 -1472 15740 -768
rect 16444 -1472 16453 -768
rect 15731 -1481 16453 -1472
rect 16724 -792 16740 -728
rect 16804 -792 16820 -728
rect 18136 -728 18232 -692
rect 16724 -808 16820 -792
rect 16724 -872 16740 -808
rect 16804 -872 16820 -808
rect 16724 -888 16820 -872
rect 16724 -952 16740 -888
rect 16804 -952 16820 -888
rect 16724 -968 16820 -952
rect 16724 -1032 16740 -968
rect 16804 -1032 16820 -968
rect 16724 -1048 16820 -1032
rect 16724 -1112 16740 -1048
rect 16804 -1112 16820 -1048
rect 16724 -1128 16820 -1112
rect 16724 -1192 16740 -1128
rect 16804 -1192 16820 -1128
rect 16724 -1208 16820 -1192
rect 16724 -1272 16740 -1208
rect 16804 -1272 16820 -1208
rect 16724 -1288 16820 -1272
rect 16724 -1352 16740 -1288
rect 16804 -1352 16820 -1288
rect 16724 -1368 16820 -1352
rect 16724 -1432 16740 -1368
rect 16804 -1432 16820 -1368
rect 16724 -1448 16820 -1432
rect 15312 -1548 15408 -1512
rect 16724 -1512 16740 -1448
rect 16804 -1512 16820 -1448
rect 17143 -768 17865 -759
rect 17143 -1472 17152 -768
rect 17856 -1472 17865 -768
rect 17143 -1481 17865 -1472
rect 18136 -792 18152 -728
rect 18216 -792 18232 -728
rect 19548 -728 19644 -692
rect 18136 -808 18232 -792
rect 18136 -872 18152 -808
rect 18216 -872 18232 -808
rect 18136 -888 18232 -872
rect 18136 -952 18152 -888
rect 18216 -952 18232 -888
rect 18136 -968 18232 -952
rect 18136 -1032 18152 -968
rect 18216 -1032 18232 -968
rect 18136 -1048 18232 -1032
rect 18136 -1112 18152 -1048
rect 18216 -1112 18232 -1048
rect 18136 -1128 18232 -1112
rect 18136 -1192 18152 -1128
rect 18216 -1192 18232 -1128
rect 18136 -1208 18232 -1192
rect 18136 -1272 18152 -1208
rect 18216 -1272 18232 -1208
rect 18136 -1288 18232 -1272
rect 18136 -1352 18152 -1288
rect 18216 -1352 18232 -1288
rect 18136 -1368 18232 -1352
rect 18136 -1432 18152 -1368
rect 18216 -1432 18232 -1368
rect 18136 -1448 18232 -1432
rect 16724 -1548 16820 -1512
rect 18136 -1512 18152 -1448
rect 18216 -1512 18232 -1448
rect 18555 -768 19277 -759
rect 18555 -1472 18564 -768
rect 19268 -1472 19277 -768
rect 18555 -1481 19277 -1472
rect 19548 -792 19564 -728
rect 19628 -792 19644 -728
rect 20960 -728 21056 -692
rect 19548 -808 19644 -792
rect 19548 -872 19564 -808
rect 19628 -872 19644 -808
rect 19548 -888 19644 -872
rect 19548 -952 19564 -888
rect 19628 -952 19644 -888
rect 19548 -968 19644 -952
rect 19548 -1032 19564 -968
rect 19628 -1032 19644 -968
rect 19548 -1048 19644 -1032
rect 19548 -1112 19564 -1048
rect 19628 -1112 19644 -1048
rect 19548 -1128 19644 -1112
rect 19548 -1192 19564 -1128
rect 19628 -1192 19644 -1128
rect 19548 -1208 19644 -1192
rect 19548 -1272 19564 -1208
rect 19628 -1272 19644 -1208
rect 19548 -1288 19644 -1272
rect 19548 -1352 19564 -1288
rect 19628 -1352 19644 -1288
rect 19548 -1368 19644 -1352
rect 19548 -1432 19564 -1368
rect 19628 -1432 19644 -1368
rect 19548 -1448 19644 -1432
rect 18136 -1548 18232 -1512
rect 19548 -1512 19564 -1448
rect 19628 -1512 19644 -1448
rect 19967 -768 20689 -759
rect 19967 -1472 19976 -768
rect 20680 -1472 20689 -768
rect 19967 -1481 20689 -1472
rect 20960 -792 20976 -728
rect 21040 -792 21056 -728
rect 22372 -728 22468 -692
rect 20960 -808 21056 -792
rect 20960 -872 20976 -808
rect 21040 -872 21056 -808
rect 20960 -888 21056 -872
rect 20960 -952 20976 -888
rect 21040 -952 21056 -888
rect 20960 -968 21056 -952
rect 20960 -1032 20976 -968
rect 21040 -1032 21056 -968
rect 20960 -1048 21056 -1032
rect 20960 -1112 20976 -1048
rect 21040 -1112 21056 -1048
rect 20960 -1128 21056 -1112
rect 20960 -1192 20976 -1128
rect 21040 -1192 21056 -1128
rect 20960 -1208 21056 -1192
rect 20960 -1272 20976 -1208
rect 21040 -1272 21056 -1208
rect 20960 -1288 21056 -1272
rect 20960 -1352 20976 -1288
rect 21040 -1352 21056 -1288
rect 20960 -1368 21056 -1352
rect 20960 -1432 20976 -1368
rect 21040 -1432 21056 -1368
rect 20960 -1448 21056 -1432
rect 19548 -1548 19644 -1512
rect 20960 -1512 20976 -1448
rect 21040 -1512 21056 -1448
rect 21379 -768 22101 -759
rect 21379 -1472 21388 -768
rect 22092 -1472 22101 -768
rect 21379 -1481 22101 -1472
rect 22372 -792 22388 -728
rect 22452 -792 22468 -728
rect 23784 -728 23880 -692
rect 22372 -808 22468 -792
rect 22372 -872 22388 -808
rect 22452 -872 22468 -808
rect 22372 -888 22468 -872
rect 22372 -952 22388 -888
rect 22452 -952 22468 -888
rect 22372 -968 22468 -952
rect 22372 -1032 22388 -968
rect 22452 -1032 22468 -968
rect 22372 -1048 22468 -1032
rect 22372 -1112 22388 -1048
rect 22452 -1112 22468 -1048
rect 22372 -1128 22468 -1112
rect 22372 -1192 22388 -1128
rect 22452 -1192 22468 -1128
rect 22372 -1208 22468 -1192
rect 22372 -1272 22388 -1208
rect 22452 -1272 22468 -1208
rect 22372 -1288 22468 -1272
rect 22372 -1352 22388 -1288
rect 22452 -1352 22468 -1288
rect 22372 -1368 22468 -1352
rect 22372 -1432 22388 -1368
rect 22452 -1432 22468 -1368
rect 22372 -1448 22468 -1432
rect 20960 -1548 21056 -1512
rect 22372 -1512 22388 -1448
rect 22452 -1512 22468 -1448
rect 22791 -768 23513 -759
rect 22791 -1472 22800 -768
rect 23504 -1472 23513 -768
rect 22791 -1481 23513 -1472
rect 23784 -792 23800 -728
rect 23864 -792 23880 -728
rect 23784 -808 23880 -792
rect 23784 -872 23800 -808
rect 23864 -872 23880 -808
rect 23784 -888 23880 -872
rect 23784 -952 23800 -888
rect 23864 -952 23880 -888
rect 23784 -968 23880 -952
rect 23784 -1032 23800 -968
rect 23864 -1032 23880 -968
rect 23784 -1048 23880 -1032
rect 23784 -1112 23800 -1048
rect 23864 -1112 23880 -1048
rect 23784 -1128 23880 -1112
rect 23784 -1192 23800 -1128
rect 23864 -1192 23880 -1128
rect 23784 -1208 23880 -1192
rect 23784 -1272 23800 -1208
rect 23864 -1272 23880 -1208
rect 23784 -1288 23880 -1272
rect 23784 -1352 23800 -1288
rect 23864 -1352 23880 -1288
rect 23784 -1368 23880 -1352
rect 23784 -1432 23800 -1368
rect 23864 -1432 23880 -1368
rect 23784 -1448 23880 -1432
rect 22372 -1548 22468 -1512
rect 23784 -1512 23800 -1448
rect 23864 -1512 23880 -1448
rect 23784 -1548 23880 -1512
rect -22812 -1848 -22716 -1812
rect -23805 -1888 -23083 -1879
rect -23805 -2592 -23796 -1888
rect -23092 -2592 -23083 -1888
rect -23805 -2601 -23083 -2592
rect -22812 -1912 -22796 -1848
rect -22732 -1912 -22716 -1848
rect -21400 -1848 -21304 -1812
rect -22812 -1928 -22716 -1912
rect -22812 -1992 -22796 -1928
rect -22732 -1992 -22716 -1928
rect -22812 -2008 -22716 -1992
rect -22812 -2072 -22796 -2008
rect -22732 -2072 -22716 -2008
rect -22812 -2088 -22716 -2072
rect -22812 -2152 -22796 -2088
rect -22732 -2152 -22716 -2088
rect -22812 -2168 -22716 -2152
rect -22812 -2232 -22796 -2168
rect -22732 -2232 -22716 -2168
rect -22812 -2248 -22716 -2232
rect -22812 -2312 -22796 -2248
rect -22732 -2312 -22716 -2248
rect -22812 -2328 -22716 -2312
rect -22812 -2392 -22796 -2328
rect -22732 -2392 -22716 -2328
rect -22812 -2408 -22716 -2392
rect -22812 -2472 -22796 -2408
rect -22732 -2472 -22716 -2408
rect -22812 -2488 -22716 -2472
rect -22812 -2552 -22796 -2488
rect -22732 -2552 -22716 -2488
rect -22812 -2568 -22716 -2552
rect -22812 -2632 -22796 -2568
rect -22732 -2632 -22716 -2568
rect -22393 -1888 -21671 -1879
rect -22393 -2592 -22384 -1888
rect -21680 -2592 -21671 -1888
rect -22393 -2601 -21671 -2592
rect -21400 -1912 -21384 -1848
rect -21320 -1912 -21304 -1848
rect -19988 -1848 -19892 -1812
rect -21400 -1928 -21304 -1912
rect -21400 -1992 -21384 -1928
rect -21320 -1992 -21304 -1928
rect -21400 -2008 -21304 -1992
rect -21400 -2072 -21384 -2008
rect -21320 -2072 -21304 -2008
rect -21400 -2088 -21304 -2072
rect -21400 -2152 -21384 -2088
rect -21320 -2152 -21304 -2088
rect -21400 -2168 -21304 -2152
rect -21400 -2232 -21384 -2168
rect -21320 -2232 -21304 -2168
rect -21400 -2248 -21304 -2232
rect -21400 -2312 -21384 -2248
rect -21320 -2312 -21304 -2248
rect -21400 -2328 -21304 -2312
rect -21400 -2392 -21384 -2328
rect -21320 -2392 -21304 -2328
rect -21400 -2408 -21304 -2392
rect -21400 -2472 -21384 -2408
rect -21320 -2472 -21304 -2408
rect -21400 -2488 -21304 -2472
rect -21400 -2552 -21384 -2488
rect -21320 -2552 -21304 -2488
rect -21400 -2568 -21304 -2552
rect -22812 -2668 -22716 -2632
rect -21400 -2632 -21384 -2568
rect -21320 -2632 -21304 -2568
rect -20981 -1888 -20259 -1879
rect -20981 -2592 -20972 -1888
rect -20268 -2592 -20259 -1888
rect -20981 -2601 -20259 -2592
rect -19988 -1912 -19972 -1848
rect -19908 -1912 -19892 -1848
rect -18576 -1848 -18480 -1812
rect -19988 -1928 -19892 -1912
rect -19988 -1992 -19972 -1928
rect -19908 -1992 -19892 -1928
rect -19988 -2008 -19892 -1992
rect -19988 -2072 -19972 -2008
rect -19908 -2072 -19892 -2008
rect -19988 -2088 -19892 -2072
rect -19988 -2152 -19972 -2088
rect -19908 -2152 -19892 -2088
rect -19988 -2168 -19892 -2152
rect -19988 -2232 -19972 -2168
rect -19908 -2232 -19892 -2168
rect -19988 -2248 -19892 -2232
rect -19988 -2312 -19972 -2248
rect -19908 -2312 -19892 -2248
rect -19988 -2328 -19892 -2312
rect -19988 -2392 -19972 -2328
rect -19908 -2392 -19892 -2328
rect -19988 -2408 -19892 -2392
rect -19988 -2472 -19972 -2408
rect -19908 -2472 -19892 -2408
rect -19988 -2488 -19892 -2472
rect -19988 -2552 -19972 -2488
rect -19908 -2552 -19892 -2488
rect -19988 -2568 -19892 -2552
rect -21400 -2668 -21304 -2632
rect -19988 -2632 -19972 -2568
rect -19908 -2632 -19892 -2568
rect -19569 -1888 -18847 -1879
rect -19569 -2592 -19560 -1888
rect -18856 -2592 -18847 -1888
rect -19569 -2601 -18847 -2592
rect -18576 -1912 -18560 -1848
rect -18496 -1912 -18480 -1848
rect -17164 -1848 -17068 -1812
rect -18576 -1928 -18480 -1912
rect -18576 -1992 -18560 -1928
rect -18496 -1992 -18480 -1928
rect -18576 -2008 -18480 -1992
rect -18576 -2072 -18560 -2008
rect -18496 -2072 -18480 -2008
rect -18576 -2088 -18480 -2072
rect -18576 -2152 -18560 -2088
rect -18496 -2152 -18480 -2088
rect -18576 -2168 -18480 -2152
rect -18576 -2232 -18560 -2168
rect -18496 -2232 -18480 -2168
rect -18576 -2248 -18480 -2232
rect -18576 -2312 -18560 -2248
rect -18496 -2312 -18480 -2248
rect -18576 -2328 -18480 -2312
rect -18576 -2392 -18560 -2328
rect -18496 -2392 -18480 -2328
rect -18576 -2408 -18480 -2392
rect -18576 -2472 -18560 -2408
rect -18496 -2472 -18480 -2408
rect -18576 -2488 -18480 -2472
rect -18576 -2552 -18560 -2488
rect -18496 -2552 -18480 -2488
rect -18576 -2568 -18480 -2552
rect -19988 -2668 -19892 -2632
rect -18576 -2632 -18560 -2568
rect -18496 -2632 -18480 -2568
rect -18157 -1888 -17435 -1879
rect -18157 -2592 -18148 -1888
rect -17444 -2592 -17435 -1888
rect -18157 -2601 -17435 -2592
rect -17164 -1912 -17148 -1848
rect -17084 -1912 -17068 -1848
rect -15752 -1848 -15656 -1812
rect -17164 -1928 -17068 -1912
rect -17164 -1992 -17148 -1928
rect -17084 -1992 -17068 -1928
rect -17164 -2008 -17068 -1992
rect -17164 -2072 -17148 -2008
rect -17084 -2072 -17068 -2008
rect -17164 -2088 -17068 -2072
rect -17164 -2152 -17148 -2088
rect -17084 -2152 -17068 -2088
rect -17164 -2168 -17068 -2152
rect -17164 -2232 -17148 -2168
rect -17084 -2232 -17068 -2168
rect -17164 -2248 -17068 -2232
rect -17164 -2312 -17148 -2248
rect -17084 -2312 -17068 -2248
rect -17164 -2328 -17068 -2312
rect -17164 -2392 -17148 -2328
rect -17084 -2392 -17068 -2328
rect -17164 -2408 -17068 -2392
rect -17164 -2472 -17148 -2408
rect -17084 -2472 -17068 -2408
rect -17164 -2488 -17068 -2472
rect -17164 -2552 -17148 -2488
rect -17084 -2552 -17068 -2488
rect -17164 -2568 -17068 -2552
rect -18576 -2668 -18480 -2632
rect -17164 -2632 -17148 -2568
rect -17084 -2632 -17068 -2568
rect -16745 -1888 -16023 -1879
rect -16745 -2592 -16736 -1888
rect -16032 -2592 -16023 -1888
rect -16745 -2601 -16023 -2592
rect -15752 -1912 -15736 -1848
rect -15672 -1912 -15656 -1848
rect -14340 -1848 -14244 -1812
rect -15752 -1928 -15656 -1912
rect -15752 -1992 -15736 -1928
rect -15672 -1992 -15656 -1928
rect -15752 -2008 -15656 -1992
rect -15752 -2072 -15736 -2008
rect -15672 -2072 -15656 -2008
rect -15752 -2088 -15656 -2072
rect -15752 -2152 -15736 -2088
rect -15672 -2152 -15656 -2088
rect -15752 -2168 -15656 -2152
rect -15752 -2232 -15736 -2168
rect -15672 -2232 -15656 -2168
rect -15752 -2248 -15656 -2232
rect -15752 -2312 -15736 -2248
rect -15672 -2312 -15656 -2248
rect -15752 -2328 -15656 -2312
rect -15752 -2392 -15736 -2328
rect -15672 -2392 -15656 -2328
rect -15752 -2408 -15656 -2392
rect -15752 -2472 -15736 -2408
rect -15672 -2472 -15656 -2408
rect -15752 -2488 -15656 -2472
rect -15752 -2552 -15736 -2488
rect -15672 -2552 -15656 -2488
rect -15752 -2568 -15656 -2552
rect -17164 -2668 -17068 -2632
rect -15752 -2632 -15736 -2568
rect -15672 -2632 -15656 -2568
rect -15333 -1888 -14611 -1879
rect -15333 -2592 -15324 -1888
rect -14620 -2592 -14611 -1888
rect -15333 -2601 -14611 -2592
rect -14340 -1912 -14324 -1848
rect -14260 -1912 -14244 -1848
rect -12928 -1848 -12832 -1812
rect -14340 -1928 -14244 -1912
rect -14340 -1992 -14324 -1928
rect -14260 -1992 -14244 -1928
rect -14340 -2008 -14244 -1992
rect -14340 -2072 -14324 -2008
rect -14260 -2072 -14244 -2008
rect -14340 -2088 -14244 -2072
rect -14340 -2152 -14324 -2088
rect -14260 -2152 -14244 -2088
rect -14340 -2168 -14244 -2152
rect -14340 -2232 -14324 -2168
rect -14260 -2232 -14244 -2168
rect -14340 -2248 -14244 -2232
rect -14340 -2312 -14324 -2248
rect -14260 -2312 -14244 -2248
rect -14340 -2328 -14244 -2312
rect -14340 -2392 -14324 -2328
rect -14260 -2392 -14244 -2328
rect -14340 -2408 -14244 -2392
rect -14340 -2472 -14324 -2408
rect -14260 -2472 -14244 -2408
rect -14340 -2488 -14244 -2472
rect -14340 -2552 -14324 -2488
rect -14260 -2552 -14244 -2488
rect -14340 -2568 -14244 -2552
rect -15752 -2668 -15656 -2632
rect -14340 -2632 -14324 -2568
rect -14260 -2632 -14244 -2568
rect -13921 -1888 -13199 -1879
rect -13921 -2592 -13912 -1888
rect -13208 -2592 -13199 -1888
rect -13921 -2601 -13199 -2592
rect -12928 -1912 -12912 -1848
rect -12848 -1912 -12832 -1848
rect -11516 -1848 -11420 -1812
rect -12928 -1928 -12832 -1912
rect -12928 -1992 -12912 -1928
rect -12848 -1992 -12832 -1928
rect -12928 -2008 -12832 -1992
rect -12928 -2072 -12912 -2008
rect -12848 -2072 -12832 -2008
rect -12928 -2088 -12832 -2072
rect -12928 -2152 -12912 -2088
rect -12848 -2152 -12832 -2088
rect -12928 -2168 -12832 -2152
rect -12928 -2232 -12912 -2168
rect -12848 -2232 -12832 -2168
rect -12928 -2248 -12832 -2232
rect -12928 -2312 -12912 -2248
rect -12848 -2312 -12832 -2248
rect -12928 -2328 -12832 -2312
rect -12928 -2392 -12912 -2328
rect -12848 -2392 -12832 -2328
rect -12928 -2408 -12832 -2392
rect -12928 -2472 -12912 -2408
rect -12848 -2472 -12832 -2408
rect -12928 -2488 -12832 -2472
rect -12928 -2552 -12912 -2488
rect -12848 -2552 -12832 -2488
rect -12928 -2568 -12832 -2552
rect -14340 -2668 -14244 -2632
rect -12928 -2632 -12912 -2568
rect -12848 -2632 -12832 -2568
rect -12509 -1888 -11787 -1879
rect -12509 -2592 -12500 -1888
rect -11796 -2592 -11787 -1888
rect -12509 -2601 -11787 -2592
rect -11516 -1912 -11500 -1848
rect -11436 -1912 -11420 -1848
rect -10104 -1848 -10008 -1812
rect -11516 -1928 -11420 -1912
rect -11516 -1992 -11500 -1928
rect -11436 -1992 -11420 -1928
rect -11516 -2008 -11420 -1992
rect -11516 -2072 -11500 -2008
rect -11436 -2072 -11420 -2008
rect -11516 -2088 -11420 -2072
rect -11516 -2152 -11500 -2088
rect -11436 -2152 -11420 -2088
rect -11516 -2168 -11420 -2152
rect -11516 -2232 -11500 -2168
rect -11436 -2232 -11420 -2168
rect -11516 -2248 -11420 -2232
rect -11516 -2312 -11500 -2248
rect -11436 -2312 -11420 -2248
rect -11516 -2328 -11420 -2312
rect -11516 -2392 -11500 -2328
rect -11436 -2392 -11420 -2328
rect -11516 -2408 -11420 -2392
rect -11516 -2472 -11500 -2408
rect -11436 -2472 -11420 -2408
rect -11516 -2488 -11420 -2472
rect -11516 -2552 -11500 -2488
rect -11436 -2552 -11420 -2488
rect -11516 -2568 -11420 -2552
rect -12928 -2668 -12832 -2632
rect -11516 -2632 -11500 -2568
rect -11436 -2632 -11420 -2568
rect -11097 -1888 -10375 -1879
rect -11097 -2592 -11088 -1888
rect -10384 -2592 -10375 -1888
rect -11097 -2601 -10375 -2592
rect -10104 -1912 -10088 -1848
rect -10024 -1912 -10008 -1848
rect -8692 -1848 -8596 -1812
rect -10104 -1928 -10008 -1912
rect -10104 -1992 -10088 -1928
rect -10024 -1992 -10008 -1928
rect -10104 -2008 -10008 -1992
rect -10104 -2072 -10088 -2008
rect -10024 -2072 -10008 -2008
rect -10104 -2088 -10008 -2072
rect -10104 -2152 -10088 -2088
rect -10024 -2152 -10008 -2088
rect -10104 -2168 -10008 -2152
rect -10104 -2232 -10088 -2168
rect -10024 -2232 -10008 -2168
rect -10104 -2248 -10008 -2232
rect -10104 -2312 -10088 -2248
rect -10024 -2312 -10008 -2248
rect -10104 -2328 -10008 -2312
rect -10104 -2392 -10088 -2328
rect -10024 -2392 -10008 -2328
rect -10104 -2408 -10008 -2392
rect -10104 -2472 -10088 -2408
rect -10024 -2472 -10008 -2408
rect -10104 -2488 -10008 -2472
rect -10104 -2552 -10088 -2488
rect -10024 -2552 -10008 -2488
rect -10104 -2568 -10008 -2552
rect -11516 -2668 -11420 -2632
rect -10104 -2632 -10088 -2568
rect -10024 -2632 -10008 -2568
rect -9685 -1888 -8963 -1879
rect -9685 -2592 -9676 -1888
rect -8972 -2592 -8963 -1888
rect -9685 -2601 -8963 -2592
rect -8692 -1912 -8676 -1848
rect -8612 -1912 -8596 -1848
rect -7280 -1848 -7184 -1812
rect -8692 -1928 -8596 -1912
rect -8692 -1992 -8676 -1928
rect -8612 -1992 -8596 -1928
rect -8692 -2008 -8596 -1992
rect -8692 -2072 -8676 -2008
rect -8612 -2072 -8596 -2008
rect -8692 -2088 -8596 -2072
rect -8692 -2152 -8676 -2088
rect -8612 -2152 -8596 -2088
rect -8692 -2168 -8596 -2152
rect -8692 -2232 -8676 -2168
rect -8612 -2232 -8596 -2168
rect -8692 -2248 -8596 -2232
rect -8692 -2312 -8676 -2248
rect -8612 -2312 -8596 -2248
rect -8692 -2328 -8596 -2312
rect -8692 -2392 -8676 -2328
rect -8612 -2392 -8596 -2328
rect -8692 -2408 -8596 -2392
rect -8692 -2472 -8676 -2408
rect -8612 -2472 -8596 -2408
rect -8692 -2488 -8596 -2472
rect -8692 -2552 -8676 -2488
rect -8612 -2552 -8596 -2488
rect -8692 -2568 -8596 -2552
rect -10104 -2668 -10008 -2632
rect -8692 -2632 -8676 -2568
rect -8612 -2632 -8596 -2568
rect -8273 -1888 -7551 -1879
rect -8273 -2592 -8264 -1888
rect -7560 -2592 -7551 -1888
rect -8273 -2601 -7551 -2592
rect -7280 -1912 -7264 -1848
rect -7200 -1912 -7184 -1848
rect -5868 -1848 -5772 -1812
rect -7280 -1928 -7184 -1912
rect -7280 -1992 -7264 -1928
rect -7200 -1992 -7184 -1928
rect -7280 -2008 -7184 -1992
rect -7280 -2072 -7264 -2008
rect -7200 -2072 -7184 -2008
rect -7280 -2088 -7184 -2072
rect -7280 -2152 -7264 -2088
rect -7200 -2152 -7184 -2088
rect -7280 -2168 -7184 -2152
rect -7280 -2232 -7264 -2168
rect -7200 -2232 -7184 -2168
rect -7280 -2248 -7184 -2232
rect -7280 -2312 -7264 -2248
rect -7200 -2312 -7184 -2248
rect -7280 -2328 -7184 -2312
rect -7280 -2392 -7264 -2328
rect -7200 -2392 -7184 -2328
rect -7280 -2408 -7184 -2392
rect -7280 -2472 -7264 -2408
rect -7200 -2472 -7184 -2408
rect -7280 -2488 -7184 -2472
rect -7280 -2552 -7264 -2488
rect -7200 -2552 -7184 -2488
rect -7280 -2568 -7184 -2552
rect -8692 -2668 -8596 -2632
rect -7280 -2632 -7264 -2568
rect -7200 -2632 -7184 -2568
rect -6861 -1888 -6139 -1879
rect -6861 -2592 -6852 -1888
rect -6148 -2592 -6139 -1888
rect -6861 -2601 -6139 -2592
rect -5868 -1912 -5852 -1848
rect -5788 -1912 -5772 -1848
rect -4456 -1848 -4360 -1812
rect -5868 -1928 -5772 -1912
rect -5868 -1992 -5852 -1928
rect -5788 -1992 -5772 -1928
rect -5868 -2008 -5772 -1992
rect -5868 -2072 -5852 -2008
rect -5788 -2072 -5772 -2008
rect -5868 -2088 -5772 -2072
rect -5868 -2152 -5852 -2088
rect -5788 -2152 -5772 -2088
rect -5868 -2168 -5772 -2152
rect -5868 -2232 -5852 -2168
rect -5788 -2232 -5772 -2168
rect -5868 -2248 -5772 -2232
rect -5868 -2312 -5852 -2248
rect -5788 -2312 -5772 -2248
rect -5868 -2328 -5772 -2312
rect -5868 -2392 -5852 -2328
rect -5788 -2392 -5772 -2328
rect -5868 -2408 -5772 -2392
rect -5868 -2472 -5852 -2408
rect -5788 -2472 -5772 -2408
rect -5868 -2488 -5772 -2472
rect -5868 -2552 -5852 -2488
rect -5788 -2552 -5772 -2488
rect -5868 -2568 -5772 -2552
rect -7280 -2668 -7184 -2632
rect -5868 -2632 -5852 -2568
rect -5788 -2632 -5772 -2568
rect -5449 -1888 -4727 -1879
rect -5449 -2592 -5440 -1888
rect -4736 -2592 -4727 -1888
rect -5449 -2601 -4727 -2592
rect -4456 -1912 -4440 -1848
rect -4376 -1912 -4360 -1848
rect -3044 -1848 -2948 -1812
rect -4456 -1928 -4360 -1912
rect -4456 -1992 -4440 -1928
rect -4376 -1992 -4360 -1928
rect -4456 -2008 -4360 -1992
rect -4456 -2072 -4440 -2008
rect -4376 -2072 -4360 -2008
rect -4456 -2088 -4360 -2072
rect -4456 -2152 -4440 -2088
rect -4376 -2152 -4360 -2088
rect -4456 -2168 -4360 -2152
rect -4456 -2232 -4440 -2168
rect -4376 -2232 -4360 -2168
rect -4456 -2248 -4360 -2232
rect -4456 -2312 -4440 -2248
rect -4376 -2312 -4360 -2248
rect -4456 -2328 -4360 -2312
rect -4456 -2392 -4440 -2328
rect -4376 -2392 -4360 -2328
rect -4456 -2408 -4360 -2392
rect -4456 -2472 -4440 -2408
rect -4376 -2472 -4360 -2408
rect -4456 -2488 -4360 -2472
rect -4456 -2552 -4440 -2488
rect -4376 -2552 -4360 -2488
rect -4456 -2568 -4360 -2552
rect -5868 -2668 -5772 -2632
rect -4456 -2632 -4440 -2568
rect -4376 -2632 -4360 -2568
rect -4037 -1888 -3315 -1879
rect -4037 -2592 -4028 -1888
rect -3324 -2592 -3315 -1888
rect -4037 -2601 -3315 -2592
rect -3044 -1912 -3028 -1848
rect -2964 -1912 -2948 -1848
rect -1632 -1848 -1536 -1812
rect -3044 -1928 -2948 -1912
rect -3044 -1992 -3028 -1928
rect -2964 -1992 -2948 -1928
rect -3044 -2008 -2948 -1992
rect -3044 -2072 -3028 -2008
rect -2964 -2072 -2948 -2008
rect -3044 -2088 -2948 -2072
rect -3044 -2152 -3028 -2088
rect -2964 -2152 -2948 -2088
rect -3044 -2168 -2948 -2152
rect -3044 -2232 -3028 -2168
rect -2964 -2232 -2948 -2168
rect -3044 -2248 -2948 -2232
rect -3044 -2312 -3028 -2248
rect -2964 -2312 -2948 -2248
rect -3044 -2328 -2948 -2312
rect -3044 -2392 -3028 -2328
rect -2964 -2392 -2948 -2328
rect -3044 -2408 -2948 -2392
rect -3044 -2472 -3028 -2408
rect -2964 -2472 -2948 -2408
rect -3044 -2488 -2948 -2472
rect -3044 -2552 -3028 -2488
rect -2964 -2552 -2948 -2488
rect -3044 -2568 -2948 -2552
rect -4456 -2668 -4360 -2632
rect -3044 -2632 -3028 -2568
rect -2964 -2632 -2948 -2568
rect -2625 -1888 -1903 -1879
rect -2625 -2592 -2616 -1888
rect -1912 -2592 -1903 -1888
rect -2625 -2601 -1903 -2592
rect -1632 -1912 -1616 -1848
rect -1552 -1912 -1536 -1848
rect -220 -1848 -124 -1812
rect -1632 -1928 -1536 -1912
rect -1632 -1992 -1616 -1928
rect -1552 -1992 -1536 -1928
rect -1632 -2008 -1536 -1992
rect -1632 -2072 -1616 -2008
rect -1552 -2072 -1536 -2008
rect -1632 -2088 -1536 -2072
rect -1632 -2152 -1616 -2088
rect -1552 -2152 -1536 -2088
rect -1632 -2168 -1536 -2152
rect -1632 -2232 -1616 -2168
rect -1552 -2232 -1536 -2168
rect -1632 -2248 -1536 -2232
rect -1632 -2312 -1616 -2248
rect -1552 -2312 -1536 -2248
rect -1632 -2328 -1536 -2312
rect -1632 -2392 -1616 -2328
rect -1552 -2392 -1536 -2328
rect -1632 -2408 -1536 -2392
rect -1632 -2472 -1616 -2408
rect -1552 -2472 -1536 -2408
rect -1632 -2488 -1536 -2472
rect -1632 -2552 -1616 -2488
rect -1552 -2552 -1536 -2488
rect -1632 -2568 -1536 -2552
rect -3044 -2668 -2948 -2632
rect -1632 -2632 -1616 -2568
rect -1552 -2632 -1536 -2568
rect -1213 -1888 -491 -1879
rect -1213 -2592 -1204 -1888
rect -500 -2592 -491 -1888
rect -1213 -2601 -491 -2592
rect -220 -1912 -204 -1848
rect -140 -1912 -124 -1848
rect 1192 -1848 1288 -1812
rect -220 -1928 -124 -1912
rect -220 -1992 -204 -1928
rect -140 -1992 -124 -1928
rect -220 -2008 -124 -1992
rect -220 -2072 -204 -2008
rect -140 -2072 -124 -2008
rect -220 -2088 -124 -2072
rect -220 -2152 -204 -2088
rect -140 -2152 -124 -2088
rect -220 -2168 -124 -2152
rect -220 -2232 -204 -2168
rect -140 -2232 -124 -2168
rect -220 -2248 -124 -2232
rect -220 -2312 -204 -2248
rect -140 -2312 -124 -2248
rect -220 -2328 -124 -2312
rect -220 -2392 -204 -2328
rect -140 -2392 -124 -2328
rect -220 -2408 -124 -2392
rect -220 -2472 -204 -2408
rect -140 -2472 -124 -2408
rect -220 -2488 -124 -2472
rect -220 -2552 -204 -2488
rect -140 -2552 -124 -2488
rect -220 -2568 -124 -2552
rect -1632 -2668 -1536 -2632
rect -220 -2632 -204 -2568
rect -140 -2632 -124 -2568
rect 199 -1888 921 -1879
rect 199 -2592 208 -1888
rect 912 -2592 921 -1888
rect 199 -2601 921 -2592
rect 1192 -1912 1208 -1848
rect 1272 -1912 1288 -1848
rect 2604 -1848 2700 -1812
rect 1192 -1928 1288 -1912
rect 1192 -1992 1208 -1928
rect 1272 -1992 1288 -1928
rect 1192 -2008 1288 -1992
rect 1192 -2072 1208 -2008
rect 1272 -2072 1288 -2008
rect 1192 -2088 1288 -2072
rect 1192 -2152 1208 -2088
rect 1272 -2152 1288 -2088
rect 1192 -2168 1288 -2152
rect 1192 -2232 1208 -2168
rect 1272 -2232 1288 -2168
rect 1192 -2248 1288 -2232
rect 1192 -2312 1208 -2248
rect 1272 -2312 1288 -2248
rect 1192 -2328 1288 -2312
rect 1192 -2392 1208 -2328
rect 1272 -2392 1288 -2328
rect 1192 -2408 1288 -2392
rect 1192 -2472 1208 -2408
rect 1272 -2472 1288 -2408
rect 1192 -2488 1288 -2472
rect 1192 -2552 1208 -2488
rect 1272 -2552 1288 -2488
rect 1192 -2568 1288 -2552
rect -220 -2668 -124 -2632
rect 1192 -2632 1208 -2568
rect 1272 -2632 1288 -2568
rect 1611 -1888 2333 -1879
rect 1611 -2592 1620 -1888
rect 2324 -2592 2333 -1888
rect 1611 -2601 2333 -2592
rect 2604 -1912 2620 -1848
rect 2684 -1912 2700 -1848
rect 4016 -1848 4112 -1812
rect 2604 -1928 2700 -1912
rect 2604 -1992 2620 -1928
rect 2684 -1992 2700 -1928
rect 2604 -2008 2700 -1992
rect 2604 -2072 2620 -2008
rect 2684 -2072 2700 -2008
rect 2604 -2088 2700 -2072
rect 2604 -2152 2620 -2088
rect 2684 -2152 2700 -2088
rect 2604 -2168 2700 -2152
rect 2604 -2232 2620 -2168
rect 2684 -2232 2700 -2168
rect 2604 -2248 2700 -2232
rect 2604 -2312 2620 -2248
rect 2684 -2312 2700 -2248
rect 2604 -2328 2700 -2312
rect 2604 -2392 2620 -2328
rect 2684 -2392 2700 -2328
rect 2604 -2408 2700 -2392
rect 2604 -2472 2620 -2408
rect 2684 -2472 2700 -2408
rect 2604 -2488 2700 -2472
rect 2604 -2552 2620 -2488
rect 2684 -2552 2700 -2488
rect 2604 -2568 2700 -2552
rect 1192 -2668 1288 -2632
rect 2604 -2632 2620 -2568
rect 2684 -2632 2700 -2568
rect 3023 -1888 3745 -1879
rect 3023 -2592 3032 -1888
rect 3736 -2592 3745 -1888
rect 3023 -2601 3745 -2592
rect 4016 -1912 4032 -1848
rect 4096 -1912 4112 -1848
rect 5428 -1848 5524 -1812
rect 4016 -1928 4112 -1912
rect 4016 -1992 4032 -1928
rect 4096 -1992 4112 -1928
rect 4016 -2008 4112 -1992
rect 4016 -2072 4032 -2008
rect 4096 -2072 4112 -2008
rect 4016 -2088 4112 -2072
rect 4016 -2152 4032 -2088
rect 4096 -2152 4112 -2088
rect 4016 -2168 4112 -2152
rect 4016 -2232 4032 -2168
rect 4096 -2232 4112 -2168
rect 4016 -2248 4112 -2232
rect 4016 -2312 4032 -2248
rect 4096 -2312 4112 -2248
rect 4016 -2328 4112 -2312
rect 4016 -2392 4032 -2328
rect 4096 -2392 4112 -2328
rect 4016 -2408 4112 -2392
rect 4016 -2472 4032 -2408
rect 4096 -2472 4112 -2408
rect 4016 -2488 4112 -2472
rect 4016 -2552 4032 -2488
rect 4096 -2552 4112 -2488
rect 4016 -2568 4112 -2552
rect 2604 -2668 2700 -2632
rect 4016 -2632 4032 -2568
rect 4096 -2632 4112 -2568
rect 4435 -1888 5157 -1879
rect 4435 -2592 4444 -1888
rect 5148 -2592 5157 -1888
rect 4435 -2601 5157 -2592
rect 5428 -1912 5444 -1848
rect 5508 -1912 5524 -1848
rect 6840 -1848 6936 -1812
rect 5428 -1928 5524 -1912
rect 5428 -1992 5444 -1928
rect 5508 -1992 5524 -1928
rect 5428 -2008 5524 -1992
rect 5428 -2072 5444 -2008
rect 5508 -2072 5524 -2008
rect 5428 -2088 5524 -2072
rect 5428 -2152 5444 -2088
rect 5508 -2152 5524 -2088
rect 5428 -2168 5524 -2152
rect 5428 -2232 5444 -2168
rect 5508 -2232 5524 -2168
rect 5428 -2248 5524 -2232
rect 5428 -2312 5444 -2248
rect 5508 -2312 5524 -2248
rect 5428 -2328 5524 -2312
rect 5428 -2392 5444 -2328
rect 5508 -2392 5524 -2328
rect 5428 -2408 5524 -2392
rect 5428 -2472 5444 -2408
rect 5508 -2472 5524 -2408
rect 5428 -2488 5524 -2472
rect 5428 -2552 5444 -2488
rect 5508 -2552 5524 -2488
rect 5428 -2568 5524 -2552
rect 4016 -2668 4112 -2632
rect 5428 -2632 5444 -2568
rect 5508 -2632 5524 -2568
rect 5847 -1888 6569 -1879
rect 5847 -2592 5856 -1888
rect 6560 -2592 6569 -1888
rect 5847 -2601 6569 -2592
rect 6840 -1912 6856 -1848
rect 6920 -1912 6936 -1848
rect 8252 -1848 8348 -1812
rect 6840 -1928 6936 -1912
rect 6840 -1992 6856 -1928
rect 6920 -1992 6936 -1928
rect 6840 -2008 6936 -1992
rect 6840 -2072 6856 -2008
rect 6920 -2072 6936 -2008
rect 6840 -2088 6936 -2072
rect 6840 -2152 6856 -2088
rect 6920 -2152 6936 -2088
rect 6840 -2168 6936 -2152
rect 6840 -2232 6856 -2168
rect 6920 -2232 6936 -2168
rect 6840 -2248 6936 -2232
rect 6840 -2312 6856 -2248
rect 6920 -2312 6936 -2248
rect 6840 -2328 6936 -2312
rect 6840 -2392 6856 -2328
rect 6920 -2392 6936 -2328
rect 6840 -2408 6936 -2392
rect 6840 -2472 6856 -2408
rect 6920 -2472 6936 -2408
rect 6840 -2488 6936 -2472
rect 6840 -2552 6856 -2488
rect 6920 -2552 6936 -2488
rect 6840 -2568 6936 -2552
rect 5428 -2668 5524 -2632
rect 6840 -2632 6856 -2568
rect 6920 -2632 6936 -2568
rect 7259 -1888 7981 -1879
rect 7259 -2592 7268 -1888
rect 7972 -2592 7981 -1888
rect 7259 -2601 7981 -2592
rect 8252 -1912 8268 -1848
rect 8332 -1912 8348 -1848
rect 9664 -1848 9760 -1812
rect 8252 -1928 8348 -1912
rect 8252 -1992 8268 -1928
rect 8332 -1992 8348 -1928
rect 8252 -2008 8348 -1992
rect 8252 -2072 8268 -2008
rect 8332 -2072 8348 -2008
rect 8252 -2088 8348 -2072
rect 8252 -2152 8268 -2088
rect 8332 -2152 8348 -2088
rect 8252 -2168 8348 -2152
rect 8252 -2232 8268 -2168
rect 8332 -2232 8348 -2168
rect 8252 -2248 8348 -2232
rect 8252 -2312 8268 -2248
rect 8332 -2312 8348 -2248
rect 8252 -2328 8348 -2312
rect 8252 -2392 8268 -2328
rect 8332 -2392 8348 -2328
rect 8252 -2408 8348 -2392
rect 8252 -2472 8268 -2408
rect 8332 -2472 8348 -2408
rect 8252 -2488 8348 -2472
rect 8252 -2552 8268 -2488
rect 8332 -2552 8348 -2488
rect 8252 -2568 8348 -2552
rect 6840 -2668 6936 -2632
rect 8252 -2632 8268 -2568
rect 8332 -2632 8348 -2568
rect 8671 -1888 9393 -1879
rect 8671 -2592 8680 -1888
rect 9384 -2592 9393 -1888
rect 8671 -2601 9393 -2592
rect 9664 -1912 9680 -1848
rect 9744 -1912 9760 -1848
rect 11076 -1848 11172 -1812
rect 9664 -1928 9760 -1912
rect 9664 -1992 9680 -1928
rect 9744 -1992 9760 -1928
rect 9664 -2008 9760 -1992
rect 9664 -2072 9680 -2008
rect 9744 -2072 9760 -2008
rect 9664 -2088 9760 -2072
rect 9664 -2152 9680 -2088
rect 9744 -2152 9760 -2088
rect 9664 -2168 9760 -2152
rect 9664 -2232 9680 -2168
rect 9744 -2232 9760 -2168
rect 9664 -2248 9760 -2232
rect 9664 -2312 9680 -2248
rect 9744 -2312 9760 -2248
rect 9664 -2328 9760 -2312
rect 9664 -2392 9680 -2328
rect 9744 -2392 9760 -2328
rect 9664 -2408 9760 -2392
rect 9664 -2472 9680 -2408
rect 9744 -2472 9760 -2408
rect 9664 -2488 9760 -2472
rect 9664 -2552 9680 -2488
rect 9744 -2552 9760 -2488
rect 9664 -2568 9760 -2552
rect 8252 -2668 8348 -2632
rect 9664 -2632 9680 -2568
rect 9744 -2632 9760 -2568
rect 10083 -1888 10805 -1879
rect 10083 -2592 10092 -1888
rect 10796 -2592 10805 -1888
rect 10083 -2601 10805 -2592
rect 11076 -1912 11092 -1848
rect 11156 -1912 11172 -1848
rect 12488 -1848 12584 -1812
rect 11076 -1928 11172 -1912
rect 11076 -1992 11092 -1928
rect 11156 -1992 11172 -1928
rect 11076 -2008 11172 -1992
rect 11076 -2072 11092 -2008
rect 11156 -2072 11172 -2008
rect 11076 -2088 11172 -2072
rect 11076 -2152 11092 -2088
rect 11156 -2152 11172 -2088
rect 11076 -2168 11172 -2152
rect 11076 -2232 11092 -2168
rect 11156 -2232 11172 -2168
rect 11076 -2248 11172 -2232
rect 11076 -2312 11092 -2248
rect 11156 -2312 11172 -2248
rect 11076 -2328 11172 -2312
rect 11076 -2392 11092 -2328
rect 11156 -2392 11172 -2328
rect 11076 -2408 11172 -2392
rect 11076 -2472 11092 -2408
rect 11156 -2472 11172 -2408
rect 11076 -2488 11172 -2472
rect 11076 -2552 11092 -2488
rect 11156 -2552 11172 -2488
rect 11076 -2568 11172 -2552
rect 9664 -2668 9760 -2632
rect 11076 -2632 11092 -2568
rect 11156 -2632 11172 -2568
rect 11495 -1888 12217 -1879
rect 11495 -2592 11504 -1888
rect 12208 -2592 12217 -1888
rect 11495 -2601 12217 -2592
rect 12488 -1912 12504 -1848
rect 12568 -1912 12584 -1848
rect 13900 -1848 13996 -1812
rect 12488 -1928 12584 -1912
rect 12488 -1992 12504 -1928
rect 12568 -1992 12584 -1928
rect 12488 -2008 12584 -1992
rect 12488 -2072 12504 -2008
rect 12568 -2072 12584 -2008
rect 12488 -2088 12584 -2072
rect 12488 -2152 12504 -2088
rect 12568 -2152 12584 -2088
rect 12488 -2168 12584 -2152
rect 12488 -2232 12504 -2168
rect 12568 -2232 12584 -2168
rect 12488 -2248 12584 -2232
rect 12488 -2312 12504 -2248
rect 12568 -2312 12584 -2248
rect 12488 -2328 12584 -2312
rect 12488 -2392 12504 -2328
rect 12568 -2392 12584 -2328
rect 12488 -2408 12584 -2392
rect 12488 -2472 12504 -2408
rect 12568 -2472 12584 -2408
rect 12488 -2488 12584 -2472
rect 12488 -2552 12504 -2488
rect 12568 -2552 12584 -2488
rect 12488 -2568 12584 -2552
rect 11076 -2668 11172 -2632
rect 12488 -2632 12504 -2568
rect 12568 -2632 12584 -2568
rect 12907 -1888 13629 -1879
rect 12907 -2592 12916 -1888
rect 13620 -2592 13629 -1888
rect 12907 -2601 13629 -2592
rect 13900 -1912 13916 -1848
rect 13980 -1912 13996 -1848
rect 15312 -1848 15408 -1812
rect 13900 -1928 13996 -1912
rect 13900 -1992 13916 -1928
rect 13980 -1992 13996 -1928
rect 13900 -2008 13996 -1992
rect 13900 -2072 13916 -2008
rect 13980 -2072 13996 -2008
rect 13900 -2088 13996 -2072
rect 13900 -2152 13916 -2088
rect 13980 -2152 13996 -2088
rect 13900 -2168 13996 -2152
rect 13900 -2232 13916 -2168
rect 13980 -2232 13996 -2168
rect 13900 -2248 13996 -2232
rect 13900 -2312 13916 -2248
rect 13980 -2312 13996 -2248
rect 13900 -2328 13996 -2312
rect 13900 -2392 13916 -2328
rect 13980 -2392 13996 -2328
rect 13900 -2408 13996 -2392
rect 13900 -2472 13916 -2408
rect 13980 -2472 13996 -2408
rect 13900 -2488 13996 -2472
rect 13900 -2552 13916 -2488
rect 13980 -2552 13996 -2488
rect 13900 -2568 13996 -2552
rect 12488 -2668 12584 -2632
rect 13900 -2632 13916 -2568
rect 13980 -2632 13996 -2568
rect 14319 -1888 15041 -1879
rect 14319 -2592 14328 -1888
rect 15032 -2592 15041 -1888
rect 14319 -2601 15041 -2592
rect 15312 -1912 15328 -1848
rect 15392 -1912 15408 -1848
rect 16724 -1848 16820 -1812
rect 15312 -1928 15408 -1912
rect 15312 -1992 15328 -1928
rect 15392 -1992 15408 -1928
rect 15312 -2008 15408 -1992
rect 15312 -2072 15328 -2008
rect 15392 -2072 15408 -2008
rect 15312 -2088 15408 -2072
rect 15312 -2152 15328 -2088
rect 15392 -2152 15408 -2088
rect 15312 -2168 15408 -2152
rect 15312 -2232 15328 -2168
rect 15392 -2232 15408 -2168
rect 15312 -2248 15408 -2232
rect 15312 -2312 15328 -2248
rect 15392 -2312 15408 -2248
rect 15312 -2328 15408 -2312
rect 15312 -2392 15328 -2328
rect 15392 -2392 15408 -2328
rect 15312 -2408 15408 -2392
rect 15312 -2472 15328 -2408
rect 15392 -2472 15408 -2408
rect 15312 -2488 15408 -2472
rect 15312 -2552 15328 -2488
rect 15392 -2552 15408 -2488
rect 15312 -2568 15408 -2552
rect 13900 -2668 13996 -2632
rect 15312 -2632 15328 -2568
rect 15392 -2632 15408 -2568
rect 15731 -1888 16453 -1879
rect 15731 -2592 15740 -1888
rect 16444 -2592 16453 -1888
rect 15731 -2601 16453 -2592
rect 16724 -1912 16740 -1848
rect 16804 -1912 16820 -1848
rect 18136 -1848 18232 -1812
rect 16724 -1928 16820 -1912
rect 16724 -1992 16740 -1928
rect 16804 -1992 16820 -1928
rect 16724 -2008 16820 -1992
rect 16724 -2072 16740 -2008
rect 16804 -2072 16820 -2008
rect 16724 -2088 16820 -2072
rect 16724 -2152 16740 -2088
rect 16804 -2152 16820 -2088
rect 16724 -2168 16820 -2152
rect 16724 -2232 16740 -2168
rect 16804 -2232 16820 -2168
rect 16724 -2248 16820 -2232
rect 16724 -2312 16740 -2248
rect 16804 -2312 16820 -2248
rect 16724 -2328 16820 -2312
rect 16724 -2392 16740 -2328
rect 16804 -2392 16820 -2328
rect 16724 -2408 16820 -2392
rect 16724 -2472 16740 -2408
rect 16804 -2472 16820 -2408
rect 16724 -2488 16820 -2472
rect 16724 -2552 16740 -2488
rect 16804 -2552 16820 -2488
rect 16724 -2568 16820 -2552
rect 15312 -2668 15408 -2632
rect 16724 -2632 16740 -2568
rect 16804 -2632 16820 -2568
rect 17143 -1888 17865 -1879
rect 17143 -2592 17152 -1888
rect 17856 -2592 17865 -1888
rect 17143 -2601 17865 -2592
rect 18136 -1912 18152 -1848
rect 18216 -1912 18232 -1848
rect 19548 -1848 19644 -1812
rect 18136 -1928 18232 -1912
rect 18136 -1992 18152 -1928
rect 18216 -1992 18232 -1928
rect 18136 -2008 18232 -1992
rect 18136 -2072 18152 -2008
rect 18216 -2072 18232 -2008
rect 18136 -2088 18232 -2072
rect 18136 -2152 18152 -2088
rect 18216 -2152 18232 -2088
rect 18136 -2168 18232 -2152
rect 18136 -2232 18152 -2168
rect 18216 -2232 18232 -2168
rect 18136 -2248 18232 -2232
rect 18136 -2312 18152 -2248
rect 18216 -2312 18232 -2248
rect 18136 -2328 18232 -2312
rect 18136 -2392 18152 -2328
rect 18216 -2392 18232 -2328
rect 18136 -2408 18232 -2392
rect 18136 -2472 18152 -2408
rect 18216 -2472 18232 -2408
rect 18136 -2488 18232 -2472
rect 18136 -2552 18152 -2488
rect 18216 -2552 18232 -2488
rect 18136 -2568 18232 -2552
rect 16724 -2668 16820 -2632
rect 18136 -2632 18152 -2568
rect 18216 -2632 18232 -2568
rect 18555 -1888 19277 -1879
rect 18555 -2592 18564 -1888
rect 19268 -2592 19277 -1888
rect 18555 -2601 19277 -2592
rect 19548 -1912 19564 -1848
rect 19628 -1912 19644 -1848
rect 20960 -1848 21056 -1812
rect 19548 -1928 19644 -1912
rect 19548 -1992 19564 -1928
rect 19628 -1992 19644 -1928
rect 19548 -2008 19644 -1992
rect 19548 -2072 19564 -2008
rect 19628 -2072 19644 -2008
rect 19548 -2088 19644 -2072
rect 19548 -2152 19564 -2088
rect 19628 -2152 19644 -2088
rect 19548 -2168 19644 -2152
rect 19548 -2232 19564 -2168
rect 19628 -2232 19644 -2168
rect 19548 -2248 19644 -2232
rect 19548 -2312 19564 -2248
rect 19628 -2312 19644 -2248
rect 19548 -2328 19644 -2312
rect 19548 -2392 19564 -2328
rect 19628 -2392 19644 -2328
rect 19548 -2408 19644 -2392
rect 19548 -2472 19564 -2408
rect 19628 -2472 19644 -2408
rect 19548 -2488 19644 -2472
rect 19548 -2552 19564 -2488
rect 19628 -2552 19644 -2488
rect 19548 -2568 19644 -2552
rect 18136 -2668 18232 -2632
rect 19548 -2632 19564 -2568
rect 19628 -2632 19644 -2568
rect 19967 -1888 20689 -1879
rect 19967 -2592 19976 -1888
rect 20680 -2592 20689 -1888
rect 19967 -2601 20689 -2592
rect 20960 -1912 20976 -1848
rect 21040 -1912 21056 -1848
rect 22372 -1848 22468 -1812
rect 20960 -1928 21056 -1912
rect 20960 -1992 20976 -1928
rect 21040 -1992 21056 -1928
rect 20960 -2008 21056 -1992
rect 20960 -2072 20976 -2008
rect 21040 -2072 21056 -2008
rect 20960 -2088 21056 -2072
rect 20960 -2152 20976 -2088
rect 21040 -2152 21056 -2088
rect 20960 -2168 21056 -2152
rect 20960 -2232 20976 -2168
rect 21040 -2232 21056 -2168
rect 20960 -2248 21056 -2232
rect 20960 -2312 20976 -2248
rect 21040 -2312 21056 -2248
rect 20960 -2328 21056 -2312
rect 20960 -2392 20976 -2328
rect 21040 -2392 21056 -2328
rect 20960 -2408 21056 -2392
rect 20960 -2472 20976 -2408
rect 21040 -2472 21056 -2408
rect 20960 -2488 21056 -2472
rect 20960 -2552 20976 -2488
rect 21040 -2552 21056 -2488
rect 20960 -2568 21056 -2552
rect 19548 -2668 19644 -2632
rect 20960 -2632 20976 -2568
rect 21040 -2632 21056 -2568
rect 21379 -1888 22101 -1879
rect 21379 -2592 21388 -1888
rect 22092 -2592 22101 -1888
rect 21379 -2601 22101 -2592
rect 22372 -1912 22388 -1848
rect 22452 -1912 22468 -1848
rect 23784 -1848 23880 -1812
rect 22372 -1928 22468 -1912
rect 22372 -1992 22388 -1928
rect 22452 -1992 22468 -1928
rect 22372 -2008 22468 -1992
rect 22372 -2072 22388 -2008
rect 22452 -2072 22468 -2008
rect 22372 -2088 22468 -2072
rect 22372 -2152 22388 -2088
rect 22452 -2152 22468 -2088
rect 22372 -2168 22468 -2152
rect 22372 -2232 22388 -2168
rect 22452 -2232 22468 -2168
rect 22372 -2248 22468 -2232
rect 22372 -2312 22388 -2248
rect 22452 -2312 22468 -2248
rect 22372 -2328 22468 -2312
rect 22372 -2392 22388 -2328
rect 22452 -2392 22468 -2328
rect 22372 -2408 22468 -2392
rect 22372 -2472 22388 -2408
rect 22452 -2472 22468 -2408
rect 22372 -2488 22468 -2472
rect 22372 -2552 22388 -2488
rect 22452 -2552 22468 -2488
rect 22372 -2568 22468 -2552
rect 20960 -2668 21056 -2632
rect 22372 -2632 22388 -2568
rect 22452 -2632 22468 -2568
rect 22791 -1888 23513 -1879
rect 22791 -2592 22800 -1888
rect 23504 -2592 23513 -1888
rect 22791 -2601 23513 -2592
rect 23784 -1912 23800 -1848
rect 23864 -1912 23880 -1848
rect 23784 -1928 23880 -1912
rect 23784 -1992 23800 -1928
rect 23864 -1992 23880 -1928
rect 23784 -2008 23880 -1992
rect 23784 -2072 23800 -2008
rect 23864 -2072 23880 -2008
rect 23784 -2088 23880 -2072
rect 23784 -2152 23800 -2088
rect 23864 -2152 23880 -2088
rect 23784 -2168 23880 -2152
rect 23784 -2232 23800 -2168
rect 23864 -2232 23880 -2168
rect 23784 -2248 23880 -2232
rect 23784 -2312 23800 -2248
rect 23864 -2312 23880 -2248
rect 23784 -2328 23880 -2312
rect 23784 -2392 23800 -2328
rect 23864 -2392 23880 -2328
rect 23784 -2408 23880 -2392
rect 23784 -2472 23800 -2408
rect 23864 -2472 23880 -2408
rect 23784 -2488 23880 -2472
rect 23784 -2552 23800 -2488
rect 23864 -2552 23880 -2488
rect 23784 -2568 23880 -2552
rect 22372 -2668 22468 -2632
rect 23784 -2632 23800 -2568
rect 23864 -2632 23880 -2568
rect 23784 -2668 23880 -2632
rect -22812 -2968 -22716 -2932
rect -23805 -3008 -23083 -2999
rect -23805 -3712 -23796 -3008
rect -23092 -3712 -23083 -3008
rect -23805 -3721 -23083 -3712
rect -22812 -3032 -22796 -2968
rect -22732 -3032 -22716 -2968
rect -21400 -2968 -21304 -2932
rect -22812 -3048 -22716 -3032
rect -22812 -3112 -22796 -3048
rect -22732 -3112 -22716 -3048
rect -22812 -3128 -22716 -3112
rect -22812 -3192 -22796 -3128
rect -22732 -3192 -22716 -3128
rect -22812 -3208 -22716 -3192
rect -22812 -3272 -22796 -3208
rect -22732 -3272 -22716 -3208
rect -22812 -3288 -22716 -3272
rect -22812 -3352 -22796 -3288
rect -22732 -3352 -22716 -3288
rect -22812 -3368 -22716 -3352
rect -22812 -3432 -22796 -3368
rect -22732 -3432 -22716 -3368
rect -22812 -3448 -22716 -3432
rect -22812 -3512 -22796 -3448
rect -22732 -3512 -22716 -3448
rect -22812 -3528 -22716 -3512
rect -22812 -3592 -22796 -3528
rect -22732 -3592 -22716 -3528
rect -22812 -3608 -22716 -3592
rect -22812 -3672 -22796 -3608
rect -22732 -3672 -22716 -3608
rect -22812 -3688 -22716 -3672
rect -22812 -3752 -22796 -3688
rect -22732 -3752 -22716 -3688
rect -22393 -3008 -21671 -2999
rect -22393 -3712 -22384 -3008
rect -21680 -3712 -21671 -3008
rect -22393 -3721 -21671 -3712
rect -21400 -3032 -21384 -2968
rect -21320 -3032 -21304 -2968
rect -19988 -2968 -19892 -2932
rect -21400 -3048 -21304 -3032
rect -21400 -3112 -21384 -3048
rect -21320 -3112 -21304 -3048
rect -21400 -3128 -21304 -3112
rect -21400 -3192 -21384 -3128
rect -21320 -3192 -21304 -3128
rect -21400 -3208 -21304 -3192
rect -21400 -3272 -21384 -3208
rect -21320 -3272 -21304 -3208
rect -21400 -3288 -21304 -3272
rect -21400 -3352 -21384 -3288
rect -21320 -3352 -21304 -3288
rect -21400 -3368 -21304 -3352
rect -21400 -3432 -21384 -3368
rect -21320 -3432 -21304 -3368
rect -21400 -3448 -21304 -3432
rect -21400 -3512 -21384 -3448
rect -21320 -3512 -21304 -3448
rect -21400 -3528 -21304 -3512
rect -21400 -3592 -21384 -3528
rect -21320 -3592 -21304 -3528
rect -21400 -3608 -21304 -3592
rect -21400 -3672 -21384 -3608
rect -21320 -3672 -21304 -3608
rect -21400 -3688 -21304 -3672
rect -22812 -3788 -22716 -3752
rect -21400 -3752 -21384 -3688
rect -21320 -3752 -21304 -3688
rect -20981 -3008 -20259 -2999
rect -20981 -3712 -20972 -3008
rect -20268 -3712 -20259 -3008
rect -20981 -3721 -20259 -3712
rect -19988 -3032 -19972 -2968
rect -19908 -3032 -19892 -2968
rect -18576 -2968 -18480 -2932
rect -19988 -3048 -19892 -3032
rect -19988 -3112 -19972 -3048
rect -19908 -3112 -19892 -3048
rect -19988 -3128 -19892 -3112
rect -19988 -3192 -19972 -3128
rect -19908 -3192 -19892 -3128
rect -19988 -3208 -19892 -3192
rect -19988 -3272 -19972 -3208
rect -19908 -3272 -19892 -3208
rect -19988 -3288 -19892 -3272
rect -19988 -3352 -19972 -3288
rect -19908 -3352 -19892 -3288
rect -19988 -3368 -19892 -3352
rect -19988 -3432 -19972 -3368
rect -19908 -3432 -19892 -3368
rect -19988 -3448 -19892 -3432
rect -19988 -3512 -19972 -3448
rect -19908 -3512 -19892 -3448
rect -19988 -3528 -19892 -3512
rect -19988 -3592 -19972 -3528
rect -19908 -3592 -19892 -3528
rect -19988 -3608 -19892 -3592
rect -19988 -3672 -19972 -3608
rect -19908 -3672 -19892 -3608
rect -19988 -3688 -19892 -3672
rect -21400 -3788 -21304 -3752
rect -19988 -3752 -19972 -3688
rect -19908 -3752 -19892 -3688
rect -19569 -3008 -18847 -2999
rect -19569 -3712 -19560 -3008
rect -18856 -3712 -18847 -3008
rect -19569 -3721 -18847 -3712
rect -18576 -3032 -18560 -2968
rect -18496 -3032 -18480 -2968
rect -17164 -2968 -17068 -2932
rect -18576 -3048 -18480 -3032
rect -18576 -3112 -18560 -3048
rect -18496 -3112 -18480 -3048
rect -18576 -3128 -18480 -3112
rect -18576 -3192 -18560 -3128
rect -18496 -3192 -18480 -3128
rect -18576 -3208 -18480 -3192
rect -18576 -3272 -18560 -3208
rect -18496 -3272 -18480 -3208
rect -18576 -3288 -18480 -3272
rect -18576 -3352 -18560 -3288
rect -18496 -3352 -18480 -3288
rect -18576 -3368 -18480 -3352
rect -18576 -3432 -18560 -3368
rect -18496 -3432 -18480 -3368
rect -18576 -3448 -18480 -3432
rect -18576 -3512 -18560 -3448
rect -18496 -3512 -18480 -3448
rect -18576 -3528 -18480 -3512
rect -18576 -3592 -18560 -3528
rect -18496 -3592 -18480 -3528
rect -18576 -3608 -18480 -3592
rect -18576 -3672 -18560 -3608
rect -18496 -3672 -18480 -3608
rect -18576 -3688 -18480 -3672
rect -19988 -3788 -19892 -3752
rect -18576 -3752 -18560 -3688
rect -18496 -3752 -18480 -3688
rect -18157 -3008 -17435 -2999
rect -18157 -3712 -18148 -3008
rect -17444 -3712 -17435 -3008
rect -18157 -3721 -17435 -3712
rect -17164 -3032 -17148 -2968
rect -17084 -3032 -17068 -2968
rect -15752 -2968 -15656 -2932
rect -17164 -3048 -17068 -3032
rect -17164 -3112 -17148 -3048
rect -17084 -3112 -17068 -3048
rect -17164 -3128 -17068 -3112
rect -17164 -3192 -17148 -3128
rect -17084 -3192 -17068 -3128
rect -17164 -3208 -17068 -3192
rect -17164 -3272 -17148 -3208
rect -17084 -3272 -17068 -3208
rect -17164 -3288 -17068 -3272
rect -17164 -3352 -17148 -3288
rect -17084 -3352 -17068 -3288
rect -17164 -3368 -17068 -3352
rect -17164 -3432 -17148 -3368
rect -17084 -3432 -17068 -3368
rect -17164 -3448 -17068 -3432
rect -17164 -3512 -17148 -3448
rect -17084 -3512 -17068 -3448
rect -17164 -3528 -17068 -3512
rect -17164 -3592 -17148 -3528
rect -17084 -3592 -17068 -3528
rect -17164 -3608 -17068 -3592
rect -17164 -3672 -17148 -3608
rect -17084 -3672 -17068 -3608
rect -17164 -3688 -17068 -3672
rect -18576 -3788 -18480 -3752
rect -17164 -3752 -17148 -3688
rect -17084 -3752 -17068 -3688
rect -16745 -3008 -16023 -2999
rect -16745 -3712 -16736 -3008
rect -16032 -3712 -16023 -3008
rect -16745 -3721 -16023 -3712
rect -15752 -3032 -15736 -2968
rect -15672 -3032 -15656 -2968
rect -14340 -2968 -14244 -2932
rect -15752 -3048 -15656 -3032
rect -15752 -3112 -15736 -3048
rect -15672 -3112 -15656 -3048
rect -15752 -3128 -15656 -3112
rect -15752 -3192 -15736 -3128
rect -15672 -3192 -15656 -3128
rect -15752 -3208 -15656 -3192
rect -15752 -3272 -15736 -3208
rect -15672 -3272 -15656 -3208
rect -15752 -3288 -15656 -3272
rect -15752 -3352 -15736 -3288
rect -15672 -3352 -15656 -3288
rect -15752 -3368 -15656 -3352
rect -15752 -3432 -15736 -3368
rect -15672 -3432 -15656 -3368
rect -15752 -3448 -15656 -3432
rect -15752 -3512 -15736 -3448
rect -15672 -3512 -15656 -3448
rect -15752 -3528 -15656 -3512
rect -15752 -3592 -15736 -3528
rect -15672 -3592 -15656 -3528
rect -15752 -3608 -15656 -3592
rect -15752 -3672 -15736 -3608
rect -15672 -3672 -15656 -3608
rect -15752 -3688 -15656 -3672
rect -17164 -3788 -17068 -3752
rect -15752 -3752 -15736 -3688
rect -15672 -3752 -15656 -3688
rect -15333 -3008 -14611 -2999
rect -15333 -3712 -15324 -3008
rect -14620 -3712 -14611 -3008
rect -15333 -3721 -14611 -3712
rect -14340 -3032 -14324 -2968
rect -14260 -3032 -14244 -2968
rect -12928 -2968 -12832 -2932
rect -14340 -3048 -14244 -3032
rect -14340 -3112 -14324 -3048
rect -14260 -3112 -14244 -3048
rect -14340 -3128 -14244 -3112
rect -14340 -3192 -14324 -3128
rect -14260 -3192 -14244 -3128
rect -14340 -3208 -14244 -3192
rect -14340 -3272 -14324 -3208
rect -14260 -3272 -14244 -3208
rect -14340 -3288 -14244 -3272
rect -14340 -3352 -14324 -3288
rect -14260 -3352 -14244 -3288
rect -14340 -3368 -14244 -3352
rect -14340 -3432 -14324 -3368
rect -14260 -3432 -14244 -3368
rect -14340 -3448 -14244 -3432
rect -14340 -3512 -14324 -3448
rect -14260 -3512 -14244 -3448
rect -14340 -3528 -14244 -3512
rect -14340 -3592 -14324 -3528
rect -14260 -3592 -14244 -3528
rect -14340 -3608 -14244 -3592
rect -14340 -3672 -14324 -3608
rect -14260 -3672 -14244 -3608
rect -14340 -3688 -14244 -3672
rect -15752 -3788 -15656 -3752
rect -14340 -3752 -14324 -3688
rect -14260 -3752 -14244 -3688
rect -13921 -3008 -13199 -2999
rect -13921 -3712 -13912 -3008
rect -13208 -3712 -13199 -3008
rect -13921 -3721 -13199 -3712
rect -12928 -3032 -12912 -2968
rect -12848 -3032 -12832 -2968
rect -11516 -2968 -11420 -2932
rect -12928 -3048 -12832 -3032
rect -12928 -3112 -12912 -3048
rect -12848 -3112 -12832 -3048
rect -12928 -3128 -12832 -3112
rect -12928 -3192 -12912 -3128
rect -12848 -3192 -12832 -3128
rect -12928 -3208 -12832 -3192
rect -12928 -3272 -12912 -3208
rect -12848 -3272 -12832 -3208
rect -12928 -3288 -12832 -3272
rect -12928 -3352 -12912 -3288
rect -12848 -3352 -12832 -3288
rect -12928 -3368 -12832 -3352
rect -12928 -3432 -12912 -3368
rect -12848 -3432 -12832 -3368
rect -12928 -3448 -12832 -3432
rect -12928 -3512 -12912 -3448
rect -12848 -3512 -12832 -3448
rect -12928 -3528 -12832 -3512
rect -12928 -3592 -12912 -3528
rect -12848 -3592 -12832 -3528
rect -12928 -3608 -12832 -3592
rect -12928 -3672 -12912 -3608
rect -12848 -3672 -12832 -3608
rect -12928 -3688 -12832 -3672
rect -14340 -3788 -14244 -3752
rect -12928 -3752 -12912 -3688
rect -12848 -3752 -12832 -3688
rect -12509 -3008 -11787 -2999
rect -12509 -3712 -12500 -3008
rect -11796 -3712 -11787 -3008
rect -12509 -3721 -11787 -3712
rect -11516 -3032 -11500 -2968
rect -11436 -3032 -11420 -2968
rect -10104 -2968 -10008 -2932
rect -11516 -3048 -11420 -3032
rect -11516 -3112 -11500 -3048
rect -11436 -3112 -11420 -3048
rect -11516 -3128 -11420 -3112
rect -11516 -3192 -11500 -3128
rect -11436 -3192 -11420 -3128
rect -11516 -3208 -11420 -3192
rect -11516 -3272 -11500 -3208
rect -11436 -3272 -11420 -3208
rect -11516 -3288 -11420 -3272
rect -11516 -3352 -11500 -3288
rect -11436 -3352 -11420 -3288
rect -11516 -3368 -11420 -3352
rect -11516 -3432 -11500 -3368
rect -11436 -3432 -11420 -3368
rect -11516 -3448 -11420 -3432
rect -11516 -3512 -11500 -3448
rect -11436 -3512 -11420 -3448
rect -11516 -3528 -11420 -3512
rect -11516 -3592 -11500 -3528
rect -11436 -3592 -11420 -3528
rect -11516 -3608 -11420 -3592
rect -11516 -3672 -11500 -3608
rect -11436 -3672 -11420 -3608
rect -11516 -3688 -11420 -3672
rect -12928 -3788 -12832 -3752
rect -11516 -3752 -11500 -3688
rect -11436 -3752 -11420 -3688
rect -11097 -3008 -10375 -2999
rect -11097 -3712 -11088 -3008
rect -10384 -3712 -10375 -3008
rect -11097 -3721 -10375 -3712
rect -10104 -3032 -10088 -2968
rect -10024 -3032 -10008 -2968
rect -8692 -2968 -8596 -2932
rect -10104 -3048 -10008 -3032
rect -10104 -3112 -10088 -3048
rect -10024 -3112 -10008 -3048
rect -10104 -3128 -10008 -3112
rect -10104 -3192 -10088 -3128
rect -10024 -3192 -10008 -3128
rect -10104 -3208 -10008 -3192
rect -10104 -3272 -10088 -3208
rect -10024 -3272 -10008 -3208
rect -10104 -3288 -10008 -3272
rect -10104 -3352 -10088 -3288
rect -10024 -3352 -10008 -3288
rect -10104 -3368 -10008 -3352
rect -10104 -3432 -10088 -3368
rect -10024 -3432 -10008 -3368
rect -10104 -3448 -10008 -3432
rect -10104 -3512 -10088 -3448
rect -10024 -3512 -10008 -3448
rect -10104 -3528 -10008 -3512
rect -10104 -3592 -10088 -3528
rect -10024 -3592 -10008 -3528
rect -10104 -3608 -10008 -3592
rect -10104 -3672 -10088 -3608
rect -10024 -3672 -10008 -3608
rect -10104 -3688 -10008 -3672
rect -11516 -3788 -11420 -3752
rect -10104 -3752 -10088 -3688
rect -10024 -3752 -10008 -3688
rect -9685 -3008 -8963 -2999
rect -9685 -3712 -9676 -3008
rect -8972 -3712 -8963 -3008
rect -9685 -3721 -8963 -3712
rect -8692 -3032 -8676 -2968
rect -8612 -3032 -8596 -2968
rect -7280 -2968 -7184 -2932
rect -8692 -3048 -8596 -3032
rect -8692 -3112 -8676 -3048
rect -8612 -3112 -8596 -3048
rect -8692 -3128 -8596 -3112
rect -8692 -3192 -8676 -3128
rect -8612 -3192 -8596 -3128
rect -8692 -3208 -8596 -3192
rect -8692 -3272 -8676 -3208
rect -8612 -3272 -8596 -3208
rect -8692 -3288 -8596 -3272
rect -8692 -3352 -8676 -3288
rect -8612 -3352 -8596 -3288
rect -8692 -3368 -8596 -3352
rect -8692 -3432 -8676 -3368
rect -8612 -3432 -8596 -3368
rect -8692 -3448 -8596 -3432
rect -8692 -3512 -8676 -3448
rect -8612 -3512 -8596 -3448
rect -8692 -3528 -8596 -3512
rect -8692 -3592 -8676 -3528
rect -8612 -3592 -8596 -3528
rect -8692 -3608 -8596 -3592
rect -8692 -3672 -8676 -3608
rect -8612 -3672 -8596 -3608
rect -8692 -3688 -8596 -3672
rect -10104 -3788 -10008 -3752
rect -8692 -3752 -8676 -3688
rect -8612 -3752 -8596 -3688
rect -8273 -3008 -7551 -2999
rect -8273 -3712 -8264 -3008
rect -7560 -3712 -7551 -3008
rect -8273 -3721 -7551 -3712
rect -7280 -3032 -7264 -2968
rect -7200 -3032 -7184 -2968
rect -5868 -2968 -5772 -2932
rect -7280 -3048 -7184 -3032
rect -7280 -3112 -7264 -3048
rect -7200 -3112 -7184 -3048
rect -7280 -3128 -7184 -3112
rect -7280 -3192 -7264 -3128
rect -7200 -3192 -7184 -3128
rect -7280 -3208 -7184 -3192
rect -7280 -3272 -7264 -3208
rect -7200 -3272 -7184 -3208
rect -7280 -3288 -7184 -3272
rect -7280 -3352 -7264 -3288
rect -7200 -3352 -7184 -3288
rect -7280 -3368 -7184 -3352
rect -7280 -3432 -7264 -3368
rect -7200 -3432 -7184 -3368
rect -7280 -3448 -7184 -3432
rect -7280 -3512 -7264 -3448
rect -7200 -3512 -7184 -3448
rect -7280 -3528 -7184 -3512
rect -7280 -3592 -7264 -3528
rect -7200 -3592 -7184 -3528
rect -7280 -3608 -7184 -3592
rect -7280 -3672 -7264 -3608
rect -7200 -3672 -7184 -3608
rect -7280 -3688 -7184 -3672
rect -8692 -3788 -8596 -3752
rect -7280 -3752 -7264 -3688
rect -7200 -3752 -7184 -3688
rect -6861 -3008 -6139 -2999
rect -6861 -3712 -6852 -3008
rect -6148 -3712 -6139 -3008
rect -6861 -3721 -6139 -3712
rect -5868 -3032 -5852 -2968
rect -5788 -3032 -5772 -2968
rect -4456 -2968 -4360 -2932
rect -5868 -3048 -5772 -3032
rect -5868 -3112 -5852 -3048
rect -5788 -3112 -5772 -3048
rect -5868 -3128 -5772 -3112
rect -5868 -3192 -5852 -3128
rect -5788 -3192 -5772 -3128
rect -5868 -3208 -5772 -3192
rect -5868 -3272 -5852 -3208
rect -5788 -3272 -5772 -3208
rect -5868 -3288 -5772 -3272
rect -5868 -3352 -5852 -3288
rect -5788 -3352 -5772 -3288
rect -5868 -3368 -5772 -3352
rect -5868 -3432 -5852 -3368
rect -5788 -3432 -5772 -3368
rect -5868 -3448 -5772 -3432
rect -5868 -3512 -5852 -3448
rect -5788 -3512 -5772 -3448
rect -5868 -3528 -5772 -3512
rect -5868 -3592 -5852 -3528
rect -5788 -3592 -5772 -3528
rect -5868 -3608 -5772 -3592
rect -5868 -3672 -5852 -3608
rect -5788 -3672 -5772 -3608
rect -5868 -3688 -5772 -3672
rect -7280 -3788 -7184 -3752
rect -5868 -3752 -5852 -3688
rect -5788 -3752 -5772 -3688
rect -5449 -3008 -4727 -2999
rect -5449 -3712 -5440 -3008
rect -4736 -3712 -4727 -3008
rect -5449 -3721 -4727 -3712
rect -4456 -3032 -4440 -2968
rect -4376 -3032 -4360 -2968
rect -3044 -2968 -2948 -2932
rect -4456 -3048 -4360 -3032
rect -4456 -3112 -4440 -3048
rect -4376 -3112 -4360 -3048
rect -4456 -3128 -4360 -3112
rect -4456 -3192 -4440 -3128
rect -4376 -3192 -4360 -3128
rect -4456 -3208 -4360 -3192
rect -4456 -3272 -4440 -3208
rect -4376 -3272 -4360 -3208
rect -4456 -3288 -4360 -3272
rect -4456 -3352 -4440 -3288
rect -4376 -3352 -4360 -3288
rect -4456 -3368 -4360 -3352
rect -4456 -3432 -4440 -3368
rect -4376 -3432 -4360 -3368
rect -4456 -3448 -4360 -3432
rect -4456 -3512 -4440 -3448
rect -4376 -3512 -4360 -3448
rect -4456 -3528 -4360 -3512
rect -4456 -3592 -4440 -3528
rect -4376 -3592 -4360 -3528
rect -4456 -3608 -4360 -3592
rect -4456 -3672 -4440 -3608
rect -4376 -3672 -4360 -3608
rect -4456 -3688 -4360 -3672
rect -5868 -3788 -5772 -3752
rect -4456 -3752 -4440 -3688
rect -4376 -3752 -4360 -3688
rect -4037 -3008 -3315 -2999
rect -4037 -3712 -4028 -3008
rect -3324 -3712 -3315 -3008
rect -4037 -3721 -3315 -3712
rect -3044 -3032 -3028 -2968
rect -2964 -3032 -2948 -2968
rect -1632 -2968 -1536 -2932
rect -3044 -3048 -2948 -3032
rect -3044 -3112 -3028 -3048
rect -2964 -3112 -2948 -3048
rect -3044 -3128 -2948 -3112
rect -3044 -3192 -3028 -3128
rect -2964 -3192 -2948 -3128
rect -3044 -3208 -2948 -3192
rect -3044 -3272 -3028 -3208
rect -2964 -3272 -2948 -3208
rect -3044 -3288 -2948 -3272
rect -3044 -3352 -3028 -3288
rect -2964 -3352 -2948 -3288
rect -3044 -3368 -2948 -3352
rect -3044 -3432 -3028 -3368
rect -2964 -3432 -2948 -3368
rect -3044 -3448 -2948 -3432
rect -3044 -3512 -3028 -3448
rect -2964 -3512 -2948 -3448
rect -3044 -3528 -2948 -3512
rect -3044 -3592 -3028 -3528
rect -2964 -3592 -2948 -3528
rect -3044 -3608 -2948 -3592
rect -3044 -3672 -3028 -3608
rect -2964 -3672 -2948 -3608
rect -3044 -3688 -2948 -3672
rect -4456 -3788 -4360 -3752
rect -3044 -3752 -3028 -3688
rect -2964 -3752 -2948 -3688
rect -2625 -3008 -1903 -2999
rect -2625 -3712 -2616 -3008
rect -1912 -3712 -1903 -3008
rect -2625 -3721 -1903 -3712
rect -1632 -3032 -1616 -2968
rect -1552 -3032 -1536 -2968
rect -220 -2968 -124 -2932
rect -1632 -3048 -1536 -3032
rect -1632 -3112 -1616 -3048
rect -1552 -3112 -1536 -3048
rect -1632 -3128 -1536 -3112
rect -1632 -3192 -1616 -3128
rect -1552 -3192 -1536 -3128
rect -1632 -3208 -1536 -3192
rect -1632 -3272 -1616 -3208
rect -1552 -3272 -1536 -3208
rect -1632 -3288 -1536 -3272
rect -1632 -3352 -1616 -3288
rect -1552 -3352 -1536 -3288
rect -1632 -3368 -1536 -3352
rect -1632 -3432 -1616 -3368
rect -1552 -3432 -1536 -3368
rect -1632 -3448 -1536 -3432
rect -1632 -3512 -1616 -3448
rect -1552 -3512 -1536 -3448
rect -1632 -3528 -1536 -3512
rect -1632 -3592 -1616 -3528
rect -1552 -3592 -1536 -3528
rect -1632 -3608 -1536 -3592
rect -1632 -3672 -1616 -3608
rect -1552 -3672 -1536 -3608
rect -1632 -3688 -1536 -3672
rect -3044 -3788 -2948 -3752
rect -1632 -3752 -1616 -3688
rect -1552 -3752 -1536 -3688
rect -1213 -3008 -491 -2999
rect -1213 -3712 -1204 -3008
rect -500 -3712 -491 -3008
rect -1213 -3721 -491 -3712
rect -220 -3032 -204 -2968
rect -140 -3032 -124 -2968
rect 1192 -2968 1288 -2932
rect -220 -3048 -124 -3032
rect -220 -3112 -204 -3048
rect -140 -3112 -124 -3048
rect -220 -3128 -124 -3112
rect -220 -3192 -204 -3128
rect -140 -3192 -124 -3128
rect -220 -3208 -124 -3192
rect -220 -3272 -204 -3208
rect -140 -3272 -124 -3208
rect -220 -3288 -124 -3272
rect -220 -3352 -204 -3288
rect -140 -3352 -124 -3288
rect -220 -3368 -124 -3352
rect -220 -3432 -204 -3368
rect -140 -3432 -124 -3368
rect -220 -3448 -124 -3432
rect -220 -3512 -204 -3448
rect -140 -3512 -124 -3448
rect -220 -3528 -124 -3512
rect -220 -3592 -204 -3528
rect -140 -3592 -124 -3528
rect -220 -3608 -124 -3592
rect -220 -3672 -204 -3608
rect -140 -3672 -124 -3608
rect -220 -3688 -124 -3672
rect -1632 -3788 -1536 -3752
rect -220 -3752 -204 -3688
rect -140 -3752 -124 -3688
rect 199 -3008 921 -2999
rect 199 -3712 208 -3008
rect 912 -3712 921 -3008
rect 199 -3721 921 -3712
rect 1192 -3032 1208 -2968
rect 1272 -3032 1288 -2968
rect 2604 -2968 2700 -2932
rect 1192 -3048 1288 -3032
rect 1192 -3112 1208 -3048
rect 1272 -3112 1288 -3048
rect 1192 -3128 1288 -3112
rect 1192 -3192 1208 -3128
rect 1272 -3192 1288 -3128
rect 1192 -3208 1288 -3192
rect 1192 -3272 1208 -3208
rect 1272 -3272 1288 -3208
rect 1192 -3288 1288 -3272
rect 1192 -3352 1208 -3288
rect 1272 -3352 1288 -3288
rect 1192 -3368 1288 -3352
rect 1192 -3432 1208 -3368
rect 1272 -3432 1288 -3368
rect 1192 -3448 1288 -3432
rect 1192 -3512 1208 -3448
rect 1272 -3512 1288 -3448
rect 1192 -3528 1288 -3512
rect 1192 -3592 1208 -3528
rect 1272 -3592 1288 -3528
rect 1192 -3608 1288 -3592
rect 1192 -3672 1208 -3608
rect 1272 -3672 1288 -3608
rect 1192 -3688 1288 -3672
rect -220 -3788 -124 -3752
rect 1192 -3752 1208 -3688
rect 1272 -3752 1288 -3688
rect 1611 -3008 2333 -2999
rect 1611 -3712 1620 -3008
rect 2324 -3712 2333 -3008
rect 1611 -3721 2333 -3712
rect 2604 -3032 2620 -2968
rect 2684 -3032 2700 -2968
rect 4016 -2968 4112 -2932
rect 2604 -3048 2700 -3032
rect 2604 -3112 2620 -3048
rect 2684 -3112 2700 -3048
rect 2604 -3128 2700 -3112
rect 2604 -3192 2620 -3128
rect 2684 -3192 2700 -3128
rect 2604 -3208 2700 -3192
rect 2604 -3272 2620 -3208
rect 2684 -3272 2700 -3208
rect 2604 -3288 2700 -3272
rect 2604 -3352 2620 -3288
rect 2684 -3352 2700 -3288
rect 2604 -3368 2700 -3352
rect 2604 -3432 2620 -3368
rect 2684 -3432 2700 -3368
rect 2604 -3448 2700 -3432
rect 2604 -3512 2620 -3448
rect 2684 -3512 2700 -3448
rect 2604 -3528 2700 -3512
rect 2604 -3592 2620 -3528
rect 2684 -3592 2700 -3528
rect 2604 -3608 2700 -3592
rect 2604 -3672 2620 -3608
rect 2684 -3672 2700 -3608
rect 2604 -3688 2700 -3672
rect 1192 -3788 1288 -3752
rect 2604 -3752 2620 -3688
rect 2684 -3752 2700 -3688
rect 3023 -3008 3745 -2999
rect 3023 -3712 3032 -3008
rect 3736 -3712 3745 -3008
rect 3023 -3721 3745 -3712
rect 4016 -3032 4032 -2968
rect 4096 -3032 4112 -2968
rect 5428 -2968 5524 -2932
rect 4016 -3048 4112 -3032
rect 4016 -3112 4032 -3048
rect 4096 -3112 4112 -3048
rect 4016 -3128 4112 -3112
rect 4016 -3192 4032 -3128
rect 4096 -3192 4112 -3128
rect 4016 -3208 4112 -3192
rect 4016 -3272 4032 -3208
rect 4096 -3272 4112 -3208
rect 4016 -3288 4112 -3272
rect 4016 -3352 4032 -3288
rect 4096 -3352 4112 -3288
rect 4016 -3368 4112 -3352
rect 4016 -3432 4032 -3368
rect 4096 -3432 4112 -3368
rect 4016 -3448 4112 -3432
rect 4016 -3512 4032 -3448
rect 4096 -3512 4112 -3448
rect 4016 -3528 4112 -3512
rect 4016 -3592 4032 -3528
rect 4096 -3592 4112 -3528
rect 4016 -3608 4112 -3592
rect 4016 -3672 4032 -3608
rect 4096 -3672 4112 -3608
rect 4016 -3688 4112 -3672
rect 2604 -3788 2700 -3752
rect 4016 -3752 4032 -3688
rect 4096 -3752 4112 -3688
rect 4435 -3008 5157 -2999
rect 4435 -3712 4444 -3008
rect 5148 -3712 5157 -3008
rect 4435 -3721 5157 -3712
rect 5428 -3032 5444 -2968
rect 5508 -3032 5524 -2968
rect 6840 -2968 6936 -2932
rect 5428 -3048 5524 -3032
rect 5428 -3112 5444 -3048
rect 5508 -3112 5524 -3048
rect 5428 -3128 5524 -3112
rect 5428 -3192 5444 -3128
rect 5508 -3192 5524 -3128
rect 5428 -3208 5524 -3192
rect 5428 -3272 5444 -3208
rect 5508 -3272 5524 -3208
rect 5428 -3288 5524 -3272
rect 5428 -3352 5444 -3288
rect 5508 -3352 5524 -3288
rect 5428 -3368 5524 -3352
rect 5428 -3432 5444 -3368
rect 5508 -3432 5524 -3368
rect 5428 -3448 5524 -3432
rect 5428 -3512 5444 -3448
rect 5508 -3512 5524 -3448
rect 5428 -3528 5524 -3512
rect 5428 -3592 5444 -3528
rect 5508 -3592 5524 -3528
rect 5428 -3608 5524 -3592
rect 5428 -3672 5444 -3608
rect 5508 -3672 5524 -3608
rect 5428 -3688 5524 -3672
rect 4016 -3788 4112 -3752
rect 5428 -3752 5444 -3688
rect 5508 -3752 5524 -3688
rect 5847 -3008 6569 -2999
rect 5847 -3712 5856 -3008
rect 6560 -3712 6569 -3008
rect 5847 -3721 6569 -3712
rect 6840 -3032 6856 -2968
rect 6920 -3032 6936 -2968
rect 8252 -2968 8348 -2932
rect 6840 -3048 6936 -3032
rect 6840 -3112 6856 -3048
rect 6920 -3112 6936 -3048
rect 6840 -3128 6936 -3112
rect 6840 -3192 6856 -3128
rect 6920 -3192 6936 -3128
rect 6840 -3208 6936 -3192
rect 6840 -3272 6856 -3208
rect 6920 -3272 6936 -3208
rect 6840 -3288 6936 -3272
rect 6840 -3352 6856 -3288
rect 6920 -3352 6936 -3288
rect 6840 -3368 6936 -3352
rect 6840 -3432 6856 -3368
rect 6920 -3432 6936 -3368
rect 6840 -3448 6936 -3432
rect 6840 -3512 6856 -3448
rect 6920 -3512 6936 -3448
rect 6840 -3528 6936 -3512
rect 6840 -3592 6856 -3528
rect 6920 -3592 6936 -3528
rect 6840 -3608 6936 -3592
rect 6840 -3672 6856 -3608
rect 6920 -3672 6936 -3608
rect 6840 -3688 6936 -3672
rect 5428 -3788 5524 -3752
rect 6840 -3752 6856 -3688
rect 6920 -3752 6936 -3688
rect 7259 -3008 7981 -2999
rect 7259 -3712 7268 -3008
rect 7972 -3712 7981 -3008
rect 7259 -3721 7981 -3712
rect 8252 -3032 8268 -2968
rect 8332 -3032 8348 -2968
rect 9664 -2968 9760 -2932
rect 8252 -3048 8348 -3032
rect 8252 -3112 8268 -3048
rect 8332 -3112 8348 -3048
rect 8252 -3128 8348 -3112
rect 8252 -3192 8268 -3128
rect 8332 -3192 8348 -3128
rect 8252 -3208 8348 -3192
rect 8252 -3272 8268 -3208
rect 8332 -3272 8348 -3208
rect 8252 -3288 8348 -3272
rect 8252 -3352 8268 -3288
rect 8332 -3352 8348 -3288
rect 8252 -3368 8348 -3352
rect 8252 -3432 8268 -3368
rect 8332 -3432 8348 -3368
rect 8252 -3448 8348 -3432
rect 8252 -3512 8268 -3448
rect 8332 -3512 8348 -3448
rect 8252 -3528 8348 -3512
rect 8252 -3592 8268 -3528
rect 8332 -3592 8348 -3528
rect 8252 -3608 8348 -3592
rect 8252 -3672 8268 -3608
rect 8332 -3672 8348 -3608
rect 8252 -3688 8348 -3672
rect 6840 -3788 6936 -3752
rect 8252 -3752 8268 -3688
rect 8332 -3752 8348 -3688
rect 8671 -3008 9393 -2999
rect 8671 -3712 8680 -3008
rect 9384 -3712 9393 -3008
rect 8671 -3721 9393 -3712
rect 9664 -3032 9680 -2968
rect 9744 -3032 9760 -2968
rect 11076 -2968 11172 -2932
rect 9664 -3048 9760 -3032
rect 9664 -3112 9680 -3048
rect 9744 -3112 9760 -3048
rect 9664 -3128 9760 -3112
rect 9664 -3192 9680 -3128
rect 9744 -3192 9760 -3128
rect 9664 -3208 9760 -3192
rect 9664 -3272 9680 -3208
rect 9744 -3272 9760 -3208
rect 9664 -3288 9760 -3272
rect 9664 -3352 9680 -3288
rect 9744 -3352 9760 -3288
rect 9664 -3368 9760 -3352
rect 9664 -3432 9680 -3368
rect 9744 -3432 9760 -3368
rect 9664 -3448 9760 -3432
rect 9664 -3512 9680 -3448
rect 9744 -3512 9760 -3448
rect 9664 -3528 9760 -3512
rect 9664 -3592 9680 -3528
rect 9744 -3592 9760 -3528
rect 9664 -3608 9760 -3592
rect 9664 -3672 9680 -3608
rect 9744 -3672 9760 -3608
rect 9664 -3688 9760 -3672
rect 8252 -3788 8348 -3752
rect 9664 -3752 9680 -3688
rect 9744 -3752 9760 -3688
rect 10083 -3008 10805 -2999
rect 10083 -3712 10092 -3008
rect 10796 -3712 10805 -3008
rect 10083 -3721 10805 -3712
rect 11076 -3032 11092 -2968
rect 11156 -3032 11172 -2968
rect 12488 -2968 12584 -2932
rect 11076 -3048 11172 -3032
rect 11076 -3112 11092 -3048
rect 11156 -3112 11172 -3048
rect 11076 -3128 11172 -3112
rect 11076 -3192 11092 -3128
rect 11156 -3192 11172 -3128
rect 11076 -3208 11172 -3192
rect 11076 -3272 11092 -3208
rect 11156 -3272 11172 -3208
rect 11076 -3288 11172 -3272
rect 11076 -3352 11092 -3288
rect 11156 -3352 11172 -3288
rect 11076 -3368 11172 -3352
rect 11076 -3432 11092 -3368
rect 11156 -3432 11172 -3368
rect 11076 -3448 11172 -3432
rect 11076 -3512 11092 -3448
rect 11156 -3512 11172 -3448
rect 11076 -3528 11172 -3512
rect 11076 -3592 11092 -3528
rect 11156 -3592 11172 -3528
rect 11076 -3608 11172 -3592
rect 11076 -3672 11092 -3608
rect 11156 -3672 11172 -3608
rect 11076 -3688 11172 -3672
rect 9664 -3788 9760 -3752
rect 11076 -3752 11092 -3688
rect 11156 -3752 11172 -3688
rect 11495 -3008 12217 -2999
rect 11495 -3712 11504 -3008
rect 12208 -3712 12217 -3008
rect 11495 -3721 12217 -3712
rect 12488 -3032 12504 -2968
rect 12568 -3032 12584 -2968
rect 13900 -2968 13996 -2932
rect 12488 -3048 12584 -3032
rect 12488 -3112 12504 -3048
rect 12568 -3112 12584 -3048
rect 12488 -3128 12584 -3112
rect 12488 -3192 12504 -3128
rect 12568 -3192 12584 -3128
rect 12488 -3208 12584 -3192
rect 12488 -3272 12504 -3208
rect 12568 -3272 12584 -3208
rect 12488 -3288 12584 -3272
rect 12488 -3352 12504 -3288
rect 12568 -3352 12584 -3288
rect 12488 -3368 12584 -3352
rect 12488 -3432 12504 -3368
rect 12568 -3432 12584 -3368
rect 12488 -3448 12584 -3432
rect 12488 -3512 12504 -3448
rect 12568 -3512 12584 -3448
rect 12488 -3528 12584 -3512
rect 12488 -3592 12504 -3528
rect 12568 -3592 12584 -3528
rect 12488 -3608 12584 -3592
rect 12488 -3672 12504 -3608
rect 12568 -3672 12584 -3608
rect 12488 -3688 12584 -3672
rect 11076 -3788 11172 -3752
rect 12488 -3752 12504 -3688
rect 12568 -3752 12584 -3688
rect 12907 -3008 13629 -2999
rect 12907 -3712 12916 -3008
rect 13620 -3712 13629 -3008
rect 12907 -3721 13629 -3712
rect 13900 -3032 13916 -2968
rect 13980 -3032 13996 -2968
rect 15312 -2968 15408 -2932
rect 13900 -3048 13996 -3032
rect 13900 -3112 13916 -3048
rect 13980 -3112 13996 -3048
rect 13900 -3128 13996 -3112
rect 13900 -3192 13916 -3128
rect 13980 -3192 13996 -3128
rect 13900 -3208 13996 -3192
rect 13900 -3272 13916 -3208
rect 13980 -3272 13996 -3208
rect 13900 -3288 13996 -3272
rect 13900 -3352 13916 -3288
rect 13980 -3352 13996 -3288
rect 13900 -3368 13996 -3352
rect 13900 -3432 13916 -3368
rect 13980 -3432 13996 -3368
rect 13900 -3448 13996 -3432
rect 13900 -3512 13916 -3448
rect 13980 -3512 13996 -3448
rect 13900 -3528 13996 -3512
rect 13900 -3592 13916 -3528
rect 13980 -3592 13996 -3528
rect 13900 -3608 13996 -3592
rect 13900 -3672 13916 -3608
rect 13980 -3672 13996 -3608
rect 13900 -3688 13996 -3672
rect 12488 -3788 12584 -3752
rect 13900 -3752 13916 -3688
rect 13980 -3752 13996 -3688
rect 14319 -3008 15041 -2999
rect 14319 -3712 14328 -3008
rect 15032 -3712 15041 -3008
rect 14319 -3721 15041 -3712
rect 15312 -3032 15328 -2968
rect 15392 -3032 15408 -2968
rect 16724 -2968 16820 -2932
rect 15312 -3048 15408 -3032
rect 15312 -3112 15328 -3048
rect 15392 -3112 15408 -3048
rect 15312 -3128 15408 -3112
rect 15312 -3192 15328 -3128
rect 15392 -3192 15408 -3128
rect 15312 -3208 15408 -3192
rect 15312 -3272 15328 -3208
rect 15392 -3272 15408 -3208
rect 15312 -3288 15408 -3272
rect 15312 -3352 15328 -3288
rect 15392 -3352 15408 -3288
rect 15312 -3368 15408 -3352
rect 15312 -3432 15328 -3368
rect 15392 -3432 15408 -3368
rect 15312 -3448 15408 -3432
rect 15312 -3512 15328 -3448
rect 15392 -3512 15408 -3448
rect 15312 -3528 15408 -3512
rect 15312 -3592 15328 -3528
rect 15392 -3592 15408 -3528
rect 15312 -3608 15408 -3592
rect 15312 -3672 15328 -3608
rect 15392 -3672 15408 -3608
rect 15312 -3688 15408 -3672
rect 13900 -3788 13996 -3752
rect 15312 -3752 15328 -3688
rect 15392 -3752 15408 -3688
rect 15731 -3008 16453 -2999
rect 15731 -3712 15740 -3008
rect 16444 -3712 16453 -3008
rect 15731 -3721 16453 -3712
rect 16724 -3032 16740 -2968
rect 16804 -3032 16820 -2968
rect 18136 -2968 18232 -2932
rect 16724 -3048 16820 -3032
rect 16724 -3112 16740 -3048
rect 16804 -3112 16820 -3048
rect 16724 -3128 16820 -3112
rect 16724 -3192 16740 -3128
rect 16804 -3192 16820 -3128
rect 16724 -3208 16820 -3192
rect 16724 -3272 16740 -3208
rect 16804 -3272 16820 -3208
rect 16724 -3288 16820 -3272
rect 16724 -3352 16740 -3288
rect 16804 -3352 16820 -3288
rect 16724 -3368 16820 -3352
rect 16724 -3432 16740 -3368
rect 16804 -3432 16820 -3368
rect 16724 -3448 16820 -3432
rect 16724 -3512 16740 -3448
rect 16804 -3512 16820 -3448
rect 16724 -3528 16820 -3512
rect 16724 -3592 16740 -3528
rect 16804 -3592 16820 -3528
rect 16724 -3608 16820 -3592
rect 16724 -3672 16740 -3608
rect 16804 -3672 16820 -3608
rect 16724 -3688 16820 -3672
rect 15312 -3788 15408 -3752
rect 16724 -3752 16740 -3688
rect 16804 -3752 16820 -3688
rect 17143 -3008 17865 -2999
rect 17143 -3712 17152 -3008
rect 17856 -3712 17865 -3008
rect 17143 -3721 17865 -3712
rect 18136 -3032 18152 -2968
rect 18216 -3032 18232 -2968
rect 19548 -2968 19644 -2932
rect 18136 -3048 18232 -3032
rect 18136 -3112 18152 -3048
rect 18216 -3112 18232 -3048
rect 18136 -3128 18232 -3112
rect 18136 -3192 18152 -3128
rect 18216 -3192 18232 -3128
rect 18136 -3208 18232 -3192
rect 18136 -3272 18152 -3208
rect 18216 -3272 18232 -3208
rect 18136 -3288 18232 -3272
rect 18136 -3352 18152 -3288
rect 18216 -3352 18232 -3288
rect 18136 -3368 18232 -3352
rect 18136 -3432 18152 -3368
rect 18216 -3432 18232 -3368
rect 18136 -3448 18232 -3432
rect 18136 -3512 18152 -3448
rect 18216 -3512 18232 -3448
rect 18136 -3528 18232 -3512
rect 18136 -3592 18152 -3528
rect 18216 -3592 18232 -3528
rect 18136 -3608 18232 -3592
rect 18136 -3672 18152 -3608
rect 18216 -3672 18232 -3608
rect 18136 -3688 18232 -3672
rect 16724 -3788 16820 -3752
rect 18136 -3752 18152 -3688
rect 18216 -3752 18232 -3688
rect 18555 -3008 19277 -2999
rect 18555 -3712 18564 -3008
rect 19268 -3712 19277 -3008
rect 18555 -3721 19277 -3712
rect 19548 -3032 19564 -2968
rect 19628 -3032 19644 -2968
rect 20960 -2968 21056 -2932
rect 19548 -3048 19644 -3032
rect 19548 -3112 19564 -3048
rect 19628 -3112 19644 -3048
rect 19548 -3128 19644 -3112
rect 19548 -3192 19564 -3128
rect 19628 -3192 19644 -3128
rect 19548 -3208 19644 -3192
rect 19548 -3272 19564 -3208
rect 19628 -3272 19644 -3208
rect 19548 -3288 19644 -3272
rect 19548 -3352 19564 -3288
rect 19628 -3352 19644 -3288
rect 19548 -3368 19644 -3352
rect 19548 -3432 19564 -3368
rect 19628 -3432 19644 -3368
rect 19548 -3448 19644 -3432
rect 19548 -3512 19564 -3448
rect 19628 -3512 19644 -3448
rect 19548 -3528 19644 -3512
rect 19548 -3592 19564 -3528
rect 19628 -3592 19644 -3528
rect 19548 -3608 19644 -3592
rect 19548 -3672 19564 -3608
rect 19628 -3672 19644 -3608
rect 19548 -3688 19644 -3672
rect 18136 -3788 18232 -3752
rect 19548 -3752 19564 -3688
rect 19628 -3752 19644 -3688
rect 19967 -3008 20689 -2999
rect 19967 -3712 19976 -3008
rect 20680 -3712 20689 -3008
rect 19967 -3721 20689 -3712
rect 20960 -3032 20976 -2968
rect 21040 -3032 21056 -2968
rect 22372 -2968 22468 -2932
rect 20960 -3048 21056 -3032
rect 20960 -3112 20976 -3048
rect 21040 -3112 21056 -3048
rect 20960 -3128 21056 -3112
rect 20960 -3192 20976 -3128
rect 21040 -3192 21056 -3128
rect 20960 -3208 21056 -3192
rect 20960 -3272 20976 -3208
rect 21040 -3272 21056 -3208
rect 20960 -3288 21056 -3272
rect 20960 -3352 20976 -3288
rect 21040 -3352 21056 -3288
rect 20960 -3368 21056 -3352
rect 20960 -3432 20976 -3368
rect 21040 -3432 21056 -3368
rect 20960 -3448 21056 -3432
rect 20960 -3512 20976 -3448
rect 21040 -3512 21056 -3448
rect 20960 -3528 21056 -3512
rect 20960 -3592 20976 -3528
rect 21040 -3592 21056 -3528
rect 20960 -3608 21056 -3592
rect 20960 -3672 20976 -3608
rect 21040 -3672 21056 -3608
rect 20960 -3688 21056 -3672
rect 19548 -3788 19644 -3752
rect 20960 -3752 20976 -3688
rect 21040 -3752 21056 -3688
rect 21379 -3008 22101 -2999
rect 21379 -3712 21388 -3008
rect 22092 -3712 22101 -3008
rect 21379 -3721 22101 -3712
rect 22372 -3032 22388 -2968
rect 22452 -3032 22468 -2968
rect 23784 -2968 23880 -2932
rect 22372 -3048 22468 -3032
rect 22372 -3112 22388 -3048
rect 22452 -3112 22468 -3048
rect 22372 -3128 22468 -3112
rect 22372 -3192 22388 -3128
rect 22452 -3192 22468 -3128
rect 22372 -3208 22468 -3192
rect 22372 -3272 22388 -3208
rect 22452 -3272 22468 -3208
rect 22372 -3288 22468 -3272
rect 22372 -3352 22388 -3288
rect 22452 -3352 22468 -3288
rect 22372 -3368 22468 -3352
rect 22372 -3432 22388 -3368
rect 22452 -3432 22468 -3368
rect 22372 -3448 22468 -3432
rect 22372 -3512 22388 -3448
rect 22452 -3512 22468 -3448
rect 22372 -3528 22468 -3512
rect 22372 -3592 22388 -3528
rect 22452 -3592 22468 -3528
rect 22372 -3608 22468 -3592
rect 22372 -3672 22388 -3608
rect 22452 -3672 22468 -3608
rect 22372 -3688 22468 -3672
rect 20960 -3788 21056 -3752
rect 22372 -3752 22388 -3688
rect 22452 -3752 22468 -3688
rect 22791 -3008 23513 -2999
rect 22791 -3712 22800 -3008
rect 23504 -3712 23513 -3008
rect 22791 -3721 23513 -3712
rect 23784 -3032 23800 -2968
rect 23864 -3032 23880 -2968
rect 23784 -3048 23880 -3032
rect 23784 -3112 23800 -3048
rect 23864 -3112 23880 -3048
rect 23784 -3128 23880 -3112
rect 23784 -3192 23800 -3128
rect 23864 -3192 23880 -3128
rect 23784 -3208 23880 -3192
rect 23784 -3272 23800 -3208
rect 23864 -3272 23880 -3208
rect 23784 -3288 23880 -3272
rect 23784 -3352 23800 -3288
rect 23864 -3352 23880 -3288
rect 23784 -3368 23880 -3352
rect 23784 -3432 23800 -3368
rect 23864 -3432 23880 -3368
rect 23784 -3448 23880 -3432
rect 23784 -3512 23800 -3448
rect 23864 -3512 23880 -3448
rect 23784 -3528 23880 -3512
rect 23784 -3592 23800 -3528
rect 23864 -3592 23880 -3528
rect 23784 -3608 23880 -3592
rect 23784 -3672 23800 -3608
rect 23864 -3672 23880 -3608
rect 23784 -3688 23880 -3672
rect 22372 -3788 22468 -3752
rect 23784 -3752 23800 -3688
rect 23864 -3752 23880 -3688
rect 23784 -3788 23880 -3752
rect -22812 -4088 -22716 -4052
rect -23805 -4128 -23083 -4119
rect -23805 -4832 -23796 -4128
rect -23092 -4832 -23083 -4128
rect -23805 -4841 -23083 -4832
rect -22812 -4152 -22796 -4088
rect -22732 -4152 -22716 -4088
rect -21400 -4088 -21304 -4052
rect -22812 -4168 -22716 -4152
rect -22812 -4232 -22796 -4168
rect -22732 -4232 -22716 -4168
rect -22812 -4248 -22716 -4232
rect -22812 -4312 -22796 -4248
rect -22732 -4312 -22716 -4248
rect -22812 -4328 -22716 -4312
rect -22812 -4392 -22796 -4328
rect -22732 -4392 -22716 -4328
rect -22812 -4408 -22716 -4392
rect -22812 -4472 -22796 -4408
rect -22732 -4472 -22716 -4408
rect -22812 -4488 -22716 -4472
rect -22812 -4552 -22796 -4488
rect -22732 -4552 -22716 -4488
rect -22812 -4568 -22716 -4552
rect -22812 -4632 -22796 -4568
rect -22732 -4632 -22716 -4568
rect -22812 -4648 -22716 -4632
rect -22812 -4712 -22796 -4648
rect -22732 -4712 -22716 -4648
rect -22812 -4728 -22716 -4712
rect -22812 -4792 -22796 -4728
rect -22732 -4792 -22716 -4728
rect -22812 -4808 -22716 -4792
rect -22812 -4872 -22796 -4808
rect -22732 -4872 -22716 -4808
rect -22393 -4128 -21671 -4119
rect -22393 -4832 -22384 -4128
rect -21680 -4832 -21671 -4128
rect -22393 -4841 -21671 -4832
rect -21400 -4152 -21384 -4088
rect -21320 -4152 -21304 -4088
rect -19988 -4088 -19892 -4052
rect -21400 -4168 -21304 -4152
rect -21400 -4232 -21384 -4168
rect -21320 -4232 -21304 -4168
rect -21400 -4248 -21304 -4232
rect -21400 -4312 -21384 -4248
rect -21320 -4312 -21304 -4248
rect -21400 -4328 -21304 -4312
rect -21400 -4392 -21384 -4328
rect -21320 -4392 -21304 -4328
rect -21400 -4408 -21304 -4392
rect -21400 -4472 -21384 -4408
rect -21320 -4472 -21304 -4408
rect -21400 -4488 -21304 -4472
rect -21400 -4552 -21384 -4488
rect -21320 -4552 -21304 -4488
rect -21400 -4568 -21304 -4552
rect -21400 -4632 -21384 -4568
rect -21320 -4632 -21304 -4568
rect -21400 -4648 -21304 -4632
rect -21400 -4712 -21384 -4648
rect -21320 -4712 -21304 -4648
rect -21400 -4728 -21304 -4712
rect -21400 -4792 -21384 -4728
rect -21320 -4792 -21304 -4728
rect -21400 -4808 -21304 -4792
rect -22812 -4908 -22716 -4872
rect -21400 -4872 -21384 -4808
rect -21320 -4872 -21304 -4808
rect -20981 -4128 -20259 -4119
rect -20981 -4832 -20972 -4128
rect -20268 -4832 -20259 -4128
rect -20981 -4841 -20259 -4832
rect -19988 -4152 -19972 -4088
rect -19908 -4152 -19892 -4088
rect -18576 -4088 -18480 -4052
rect -19988 -4168 -19892 -4152
rect -19988 -4232 -19972 -4168
rect -19908 -4232 -19892 -4168
rect -19988 -4248 -19892 -4232
rect -19988 -4312 -19972 -4248
rect -19908 -4312 -19892 -4248
rect -19988 -4328 -19892 -4312
rect -19988 -4392 -19972 -4328
rect -19908 -4392 -19892 -4328
rect -19988 -4408 -19892 -4392
rect -19988 -4472 -19972 -4408
rect -19908 -4472 -19892 -4408
rect -19988 -4488 -19892 -4472
rect -19988 -4552 -19972 -4488
rect -19908 -4552 -19892 -4488
rect -19988 -4568 -19892 -4552
rect -19988 -4632 -19972 -4568
rect -19908 -4632 -19892 -4568
rect -19988 -4648 -19892 -4632
rect -19988 -4712 -19972 -4648
rect -19908 -4712 -19892 -4648
rect -19988 -4728 -19892 -4712
rect -19988 -4792 -19972 -4728
rect -19908 -4792 -19892 -4728
rect -19988 -4808 -19892 -4792
rect -21400 -4908 -21304 -4872
rect -19988 -4872 -19972 -4808
rect -19908 -4872 -19892 -4808
rect -19569 -4128 -18847 -4119
rect -19569 -4832 -19560 -4128
rect -18856 -4832 -18847 -4128
rect -19569 -4841 -18847 -4832
rect -18576 -4152 -18560 -4088
rect -18496 -4152 -18480 -4088
rect -17164 -4088 -17068 -4052
rect -18576 -4168 -18480 -4152
rect -18576 -4232 -18560 -4168
rect -18496 -4232 -18480 -4168
rect -18576 -4248 -18480 -4232
rect -18576 -4312 -18560 -4248
rect -18496 -4312 -18480 -4248
rect -18576 -4328 -18480 -4312
rect -18576 -4392 -18560 -4328
rect -18496 -4392 -18480 -4328
rect -18576 -4408 -18480 -4392
rect -18576 -4472 -18560 -4408
rect -18496 -4472 -18480 -4408
rect -18576 -4488 -18480 -4472
rect -18576 -4552 -18560 -4488
rect -18496 -4552 -18480 -4488
rect -18576 -4568 -18480 -4552
rect -18576 -4632 -18560 -4568
rect -18496 -4632 -18480 -4568
rect -18576 -4648 -18480 -4632
rect -18576 -4712 -18560 -4648
rect -18496 -4712 -18480 -4648
rect -18576 -4728 -18480 -4712
rect -18576 -4792 -18560 -4728
rect -18496 -4792 -18480 -4728
rect -18576 -4808 -18480 -4792
rect -19988 -4908 -19892 -4872
rect -18576 -4872 -18560 -4808
rect -18496 -4872 -18480 -4808
rect -18157 -4128 -17435 -4119
rect -18157 -4832 -18148 -4128
rect -17444 -4832 -17435 -4128
rect -18157 -4841 -17435 -4832
rect -17164 -4152 -17148 -4088
rect -17084 -4152 -17068 -4088
rect -15752 -4088 -15656 -4052
rect -17164 -4168 -17068 -4152
rect -17164 -4232 -17148 -4168
rect -17084 -4232 -17068 -4168
rect -17164 -4248 -17068 -4232
rect -17164 -4312 -17148 -4248
rect -17084 -4312 -17068 -4248
rect -17164 -4328 -17068 -4312
rect -17164 -4392 -17148 -4328
rect -17084 -4392 -17068 -4328
rect -17164 -4408 -17068 -4392
rect -17164 -4472 -17148 -4408
rect -17084 -4472 -17068 -4408
rect -17164 -4488 -17068 -4472
rect -17164 -4552 -17148 -4488
rect -17084 -4552 -17068 -4488
rect -17164 -4568 -17068 -4552
rect -17164 -4632 -17148 -4568
rect -17084 -4632 -17068 -4568
rect -17164 -4648 -17068 -4632
rect -17164 -4712 -17148 -4648
rect -17084 -4712 -17068 -4648
rect -17164 -4728 -17068 -4712
rect -17164 -4792 -17148 -4728
rect -17084 -4792 -17068 -4728
rect -17164 -4808 -17068 -4792
rect -18576 -4908 -18480 -4872
rect -17164 -4872 -17148 -4808
rect -17084 -4872 -17068 -4808
rect -16745 -4128 -16023 -4119
rect -16745 -4832 -16736 -4128
rect -16032 -4832 -16023 -4128
rect -16745 -4841 -16023 -4832
rect -15752 -4152 -15736 -4088
rect -15672 -4152 -15656 -4088
rect -14340 -4088 -14244 -4052
rect -15752 -4168 -15656 -4152
rect -15752 -4232 -15736 -4168
rect -15672 -4232 -15656 -4168
rect -15752 -4248 -15656 -4232
rect -15752 -4312 -15736 -4248
rect -15672 -4312 -15656 -4248
rect -15752 -4328 -15656 -4312
rect -15752 -4392 -15736 -4328
rect -15672 -4392 -15656 -4328
rect -15752 -4408 -15656 -4392
rect -15752 -4472 -15736 -4408
rect -15672 -4472 -15656 -4408
rect -15752 -4488 -15656 -4472
rect -15752 -4552 -15736 -4488
rect -15672 -4552 -15656 -4488
rect -15752 -4568 -15656 -4552
rect -15752 -4632 -15736 -4568
rect -15672 -4632 -15656 -4568
rect -15752 -4648 -15656 -4632
rect -15752 -4712 -15736 -4648
rect -15672 -4712 -15656 -4648
rect -15752 -4728 -15656 -4712
rect -15752 -4792 -15736 -4728
rect -15672 -4792 -15656 -4728
rect -15752 -4808 -15656 -4792
rect -17164 -4908 -17068 -4872
rect -15752 -4872 -15736 -4808
rect -15672 -4872 -15656 -4808
rect -15333 -4128 -14611 -4119
rect -15333 -4832 -15324 -4128
rect -14620 -4832 -14611 -4128
rect -15333 -4841 -14611 -4832
rect -14340 -4152 -14324 -4088
rect -14260 -4152 -14244 -4088
rect -12928 -4088 -12832 -4052
rect -14340 -4168 -14244 -4152
rect -14340 -4232 -14324 -4168
rect -14260 -4232 -14244 -4168
rect -14340 -4248 -14244 -4232
rect -14340 -4312 -14324 -4248
rect -14260 -4312 -14244 -4248
rect -14340 -4328 -14244 -4312
rect -14340 -4392 -14324 -4328
rect -14260 -4392 -14244 -4328
rect -14340 -4408 -14244 -4392
rect -14340 -4472 -14324 -4408
rect -14260 -4472 -14244 -4408
rect -14340 -4488 -14244 -4472
rect -14340 -4552 -14324 -4488
rect -14260 -4552 -14244 -4488
rect -14340 -4568 -14244 -4552
rect -14340 -4632 -14324 -4568
rect -14260 -4632 -14244 -4568
rect -14340 -4648 -14244 -4632
rect -14340 -4712 -14324 -4648
rect -14260 -4712 -14244 -4648
rect -14340 -4728 -14244 -4712
rect -14340 -4792 -14324 -4728
rect -14260 -4792 -14244 -4728
rect -14340 -4808 -14244 -4792
rect -15752 -4908 -15656 -4872
rect -14340 -4872 -14324 -4808
rect -14260 -4872 -14244 -4808
rect -13921 -4128 -13199 -4119
rect -13921 -4832 -13912 -4128
rect -13208 -4832 -13199 -4128
rect -13921 -4841 -13199 -4832
rect -12928 -4152 -12912 -4088
rect -12848 -4152 -12832 -4088
rect -11516 -4088 -11420 -4052
rect -12928 -4168 -12832 -4152
rect -12928 -4232 -12912 -4168
rect -12848 -4232 -12832 -4168
rect -12928 -4248 -12832 -4232
rect -12928 -4312 -12912 -4248
rect -12848 -4312 -12832 -4248
rect -12928 -4328 -12832 -4312
rect -12928 -4392 -12912 -4328
rect -12848 -4392 -12832 -4328
rect -12928 -4408 -12832 -4392
rect -12928 -4472 -12912 -4408
rect -12848 -4472 -12832 -4408
rect -12928 -4488 -12832 -4472
rect -12928 -4552 -12912 -4488
rect -12848 -4552 -12832 -4488
rect -12928 -4568 -12832 -4552
rect -12928 -4632 -12912 -4568
rect -12848 -4632 -12832 -4568
rect -12928 -4648 -12832 -4632
rect -12928 -4712 -12912 -4648
rect -12848 -4712 -12832 -4648
rect -12928 -4728 -12832 -4712
rect -12928 -4792 -12912 -4728
rect -12848 -4792 -12832 -4728
rect -12928 -4808 -12832 -4792
rect -14340 -4908 -14244 -4872
rect -12928 -4872 -12912 -4808
rect -12848 -4872 -12832 -4808
rect -12509 -4128 -11787 -4119
rect -12509 -4832 -12500 -4128
rect -11796 -4832 -11787 -4128
rect -12509 -4841 -11787 -4832
rect -11516 -4152 -11500 -4088
rect -11436 -4152 -11420 -4088
rect -10104 -4088 -10008 -4052
rect -11516 -4168 -11420 -4152
rect -11516 -4232 -11500 -4168
rect -11436 -4232 -11420 -4168
rect -11516 -4248 -11420 -4232
rect -11516 -4312 -11500 -4248
rect -11436 -4312 -11420 -4248
rect -11516 -4328 -11420 -4312
rect -11516 -4392 -11500 -4328
rect -11436 -4392 -11420 -4328
rect -11516 -4408 -11420 -4392
rect -11516 -4472 -11500 -4408
rect -11436 -4472 -11420 -4408
rect -11516 -4488 -11420 -4472
rect -11516 -4552 -11500 -4488
rect -11436 -4552 -11420 -4488
rect -11516 -4568 -11420 -4552
rect -11516 -4632 -11500 -4568
rect -11436 -4632 -11420 -4568
rect -11516 -4648 -11420 -4632
rect -11516 -4712 -11500 -4648
rect -11436 -4712 -11420 -4648
rect -11516 -4728 -11420 -4712
rect -11516 -4792 -11500 -4728
rect -11436 -4792 -11420 -4728
rect -11516 -4808 -11420 -4792
rect -12928 -4908 -12832 -4872
rect -11516 -4872 -11500 -4808
rect -11436 -4872 -11420 -4808
rect -11097 -4128 -10375 -4119
rect -11097 -4832 -11088 -4128
rect -10384 -4832 -10375 -4128
rect -11097 -4841 -10375 -4832
rect -10104 -4152 -10088 -4088
rect -10024 -4152 -10008 -4088
rect -8692 -4088 -8596 -4052
rect -10104 -4168 -10008 -4152
rect -10104 -4232 -10088 -4168
rect -10024 -4232 -10008 -4168
rect -10104 -4248 -10008 -4232
rect -10104 -4312 -10088 -4248
rect -10024 -4312 -10008 -4248
rect -10104 -4328 -10008 -4312
rect -10104 -4392 -10088 -4328
rect -10024 -4392 -10008 -4328
rect -10104 -4408 -10008 -4392
rect -10104 -4472 -10088 -4408
rect -10024 -4472 -10008 -4408
rect -10104 -4488 -10008 -4472
rect -10104 -4552 -10088 -4488
rect -10024 -4552 -10008 -4488
rect -10104 -4568 -10008 -4552
rect -10104 -4632 -10088 -4568
rect -10024 -4632 -10008 -4568
rect -10104 -4648 -10008 -4632
rect -10104 -4712 -10088 -4648
rect -10024 -4712 -10008 -4648
rect -10104 -4728 -10008 -4712
rect -10104 -4792 -10088 -4728
rect -10024 -4792 -10008 -4728
rect -10104 -4808 -10008 -4792
rect -11516 -4908 -11420 -4872
rect -10104 -4872 -10088 -4808
rect -10024 -4872 -10008 -4808
rect -9685 -4128 -8963 -4119
rect -9685 -4832 -9676 -4128
rect -8972 -4832 -8963 -4128
rect -9685 -4841 -8963 -4832
rect -8692 -4152 -8676 -4088
rect -8612 -4152 -8596 -4088
rect -7280 -4088 -7184 -4052
rect -8692 -4168 -8596 -4152
rect -8692 -4232 -8676 -4168
rect -8612 -4232 -8596 -4168
rect -8692 -4248 -8596 -4232
rect -8692 -4312 -8676 -4248
rect -8612 -4312 -8596 -4248
rect -8692 -4328 -8596 -4312
rect -8692 -4392 -8676 -4328
rect -8612 -4392 -8596 -4328
rect -8692 -4408 -8596 -4392
rect -8692 -4472 -8676 -4408
rect -8612 -4472 -8596 -4408
rect -8692 -4488 -8596 -4472
rect -8692 -4552 -8676 -4488
rect -8612 -4552 -8596 -4488
rect -8692 -4568 -8596 -4552
rect -8692 -4632 -8676 -4568
rect -8612 -4632 -8596 -4568
rect -8692 -4648 -8596 -4632
rect -8692 -4712 -8676 -4648
rect -8612 -4712 -8596 -4648
rect -8692 -4728 -8596 -4712
rect -8692 -4792 -8676 -4728
rect -8612 -4792 -8596 -4728
rect -8692 -4808 -8596 -4792
rect -10104 -4908 -10008 -4872
rect -8692 -4872 -8676 -4808
rect -8612 -4872 -8596 -4808
rect -8273 -4128 -7551 -4119
rect -8273 -4832 -8264 -4128
rect -7560 -4832 -7551 -4128
rect -8273 -4841 -7551 -4832
rect -7280 -4152 -7264 -4088
rect -7200 -4152 -7184 -4088
rect -5868 -4088 -5772 -4052
rect -7280 -4168 -7184 -4152
rect -7280 -4232 -7264 -4168
rect -7200 -4232 -7184 -4168
rect -7280 -4248 -7184 -4232
rect -7280 -4312 -7264 -4248
rect -7200 -4312 -7184 -4248
rect -7280 -4328 -7184 -4312
rect -7280 -4392 -7264 -4328
rect -7200 -4392 -7184 -4328
rect -7280 -4408 -7184 -4392
rect -7280 -4472 -7264 -4408
rect -7200 -4472 -7184 -4408
rect -7280 -4488 -7184 -4472
rect -7280 -4552 -7264 -4488
rect -7200 -4552 -7184 -4488
rect -7280 -4568 -7184 -4552
rect -7280 -4632 -7264 -4568
rect -7200 -4632 -7184 -4568
rect -7280 -4648 -7184 -4632
rect -7280 -4712 -7264 -4648
rect -7200 -4712 -7184 -4648
rect -7280 -4728 -7184 -4712
rect -7280 -4792 -7264 -4728
rect -7200 -4792 -7184 -4728
rect -7280 -4808 -7184 -4792
rect -8692 -4908 -8596 -4872
rect -7280 -4872 -7264 -4808
rect -7200 -4872 -7184 -4808
rect -6861 -4128 -6139 -4119
rect -6861 -4832 -6852 -4128
rect -6148 -4832 -6139 -4128
rect -6861 -4841 -6139 -4832
rect -5868 -4152 -5852 -4088
rect -5788 -4152 -5772 -4088
rect -4456 -4088 -4360 -4052
rect -5868 -4168 -5772 -4152
rect -5868 -4232 -5852 -4168
rect -5788 -4232 -5772 -4168
rect -5868 -4248 -5772 -4232
rect -5868 -4312 -5852 -4248
rect -5788 -4312 -5772 -4248
rect -5868 -4328 -5772 -4312
rect -5868 -4392 -5852 -4328
rect -5788 -4392 -5772 -4328
rect -5868 -4408 -5772 -4392
rect -5868 -4472 -5852 -4408
rect -5788 -4472 -5772 -4408
rect -5868 -4488 -5772 -4472
rect -5868 -4552 -5852 -4488
rect -5788 -4552 -5772 -4488
rect -5868 -4568 -5772 -4552
rect -5868 -4632 -5852 -4568
rect -5788 -4632 -5772 -4568
rect -5868 -4648 -5772 -4632
rect -5868 -4712 -5852 -4648
rect -5788 -4712 -5772 -4648
rect -5868 -4728 -5772 -4712
rect -5868 -4792 -5852 -4728
rect -5788 -4792 -5772 -4728
rect -5868 -4808 -5772 -4792
rect -7280 -4908 -7184 -4872
rect -5868 -4872 -5852 -4808
rect -5788 -4872 -5772 -4808
rect -5449 -4128 -4727 -4119
rect -5449 -4832 -5440 -4128
rect -4736 -4832 -4727 -4128
rect -5449 -4841 -4727 -4832
rect -4456 -4152 -4440 -4088
rect -4376 -4152 -4360 -4088
rect -3044 -4088 -2948 -4052
rect -4456 -4168 -4360 -4152
rect -4456 -4232 -4440 -4168
rect -4376 -4232 -4360 -4168
rect -4456 -4248 -4360 -4232
rect -4456 -4312 -4440 -4248
rect -4376 -4312 -4360 -4248
rect -4456 -4328 -4360 -4312
rect -4456 -4392 -4440 -4328
rect -4376 -4392 -4360 -4328
rect -4456 -4408 -4360 -4392
rect -4456 -4472 -4440 -4408
rect -4376 -4472 -4360 -4408
rect -4456 -4488 -4360 -4472
rect -4456 -4552 -4440 -4488
rect -4376 -4552 -4360 -4488
rect -4456 -4568 -4360 -4552
rect -4456 -4632 -4440 -4568
rect -4376 -4632 -4360 -4568
rect -4456 -4648 -4360 -4632
rect -4456 -4712 -4440 -4648
rect -4376 -4712 -4360 -4648
rect -4456 -4728 -4360 -4712
rect -4456 -4792 -4440 -4728
rect -4376 -4792 -4360 -4728
rect -4456 -4808 -4360 -4792
rect -5868 -4908 -5772 -4872
rect -4456 -4872 -4440 -4808
rect -4376 -4872 -4360 -4808
rect -4037 -4128 -3315 -4119
rect -4037 -4832 -4028 -4128
rect -3324 -4832 -3315 -4128
rect -4037 -4841 -3315 -4832
rect -3044 -4152 -3028 -4088
rect -2964 -4152 -2948 -4088
rect -1632 -4088 -1536 -4052
rect -3044 -4168 -2948 -4152
rect -3044 -4232 -3028 -4168
rect -2964 -4232 -2948 -4168
rect -3044 -4248 -2948 -4232
rect -3044 -4312 -3028 -4248
rect -2964 -4312 -2948 -4248
rect -3044 -4328 -2948 -4312
rect -3044 -4392 -3028 -4328
rect -2964 -4392 -2948 -4328
rect -3044 -4408 -2948 -4392
rect -3044 -4472 -3028 -4408
rect -2964 -4472 -2948 -4408
rect -3044 -4488 -2948 -4472
rect -3044 -4552 -3028 -4488
rect -2964 -4552 -2948 -4488
rect -3044 -4568 -2948 -4552
rect -3044 -4632 -3028 -4568
rect -2964 -4632 -2948 -4568
rect -3044 -4648 -2948 -4632
rect -3044 -4712 -3028 -4648
rect -2964 -4712 -2948 -4648
rect -3044 -4728 -2948 -4712
rect -3044 -4792 -3028 -4728
rect -2964 -4792 -2948 -4728
rect -3044 -4808 -2948 -4792
rect -4456 -4908 -4360 -4872
rect -3044 -4872 -3028 -4808
rect -2964 -4872 -2948 -4808
rect -2625 -4128 -1903 -4119
rect -2625 -4832 -2616 -4128
rect -1912 -4832 -1903 -4128
rect -2625 -4841 -1903 -4832
rect -1632 -4152 -1616 -4088
rect -1552 -4152 -1536 -4088
rect -220 -4088 -124 -4052
rect -1632 -4168 -1536 -4152
rect -1632 -4232 -1616 -4168
rect -1552 -4232 -1536 -4168
rect -1632 -4248 -1536 -4232
rect -1632 -4312 -1616 -4248
rect -1552 -4312 -1536 -4248
rect -1632 -4328 -1536 -4312
rect -1632 -4392 -1616 -4328
rect -1552 -4392 -1536 -4328
rect -1632 -4408 -1536 -4392
rect -1632 -4472 -1616 -4408
rect -1552 -4472 -1536 -4408
rect -1632 -4488 -1536 -4472
rect -1632 -4552 -1616 -4488
rect -1552 -4552 -1536 -4488
rect -1632 -4568 -1536 -4552
rect -1632 -4632 -1616 -4568
rect -1552 -4632 -1536 -4568
rect -1632 -4648 -1536 -4632
rect -1632 -4712 -1616 -4648
rect -1552 -4712 -1536 -4648
rect -1632 -4728 -1536 -4712
rect -1632 -4792 -1616 -4728
rect -1552 -4792 -1536 -4728
rect -1632 -4808 -1536 -4792
rect -3044 -4908 -2948 -4872
rect -1632 -4872 -1616 -4808
rect -1552 -4872 -1536 -4808
rect -1213 -4128 -491 -4119
rect -1213 -4832 -1204 -4128
rect -500 -4832 -491 -4128
rect -1213 -4841 -491 -4832
rect -220 -4152 -204 -4088
rect -140 -4152 -124 -4088
rect 1192 -4088 1288 -4052
rect -220 -4168 -124 -4152
rect -220 -4232 -204 -4168
rect -140 -4232 -124 -4168
rect -220 -4248 -124 -4232
rect -220 -4312 -204 -4248
rect -140 -4312 -124 -4248
rect -220 -4328 -124 -4312
rect -220 -4392 -204 -4328
rect -140 -4392 -124 -4328
rect -220 -4408 -124 -4392
rect -220 -4472 -204 -4408
rect -140 -4472 -124 -4408
rect -220 -4488 -124 -4472
rect -220 -4552 -204 -4488
rect -140 -4552 -124 -4488
rect -220 -4568 -124 -4552
rect -220 -4632 -204 -4568
rect -140 -4632 -124 -4568
rect -220 -4648 -124 -4632
rect -220 -4712 -204 -4648
rect -140 -4712 -124 -4648
rect -220 -4728 -124 -4712
rect -220 -4792 -204 -4728
rect -140 -4792 -124 -4728
rect -220 -4808 -124 -4792
rect -1632 -4908 -1536 -4872
rect -220 -4872 -204 -4808
rect -140 -4872 -124 -4808
rect 199 -4128 921 -4119
rect 199 -4832 208 -4128
rect 912 -4832 921 -4128
rect 199 -4841 921 -4832
rect 1192 -4152 1208 -4088
rect 1272 -4152 1288 -4088
rect 2604 -4088 2700 -4052
rect 1192 -4168 1288 -4152
rect 1192 -4232 1208 -4168
rect 1272 -4232 1288 -4168
rect 1192 -4248 1288 -4232
rect 1192 -4312 1208 -4248
rect 1272 -4312 1288 -4248
rect 1192 -4328 1288 -4312
rect 1192 -4392 1208 -4328
rect 1272 -4392 1288 -4328
rect 1192 -4408 1288 -4392
rect 1192 -4472 1208 -4408
rect 1272 -4472 1288 -4408
rect 1192 -4488 1288 -4472
rect 1192 -4552 1208 -4488
rect 1272 -4552 1288 -4488
rect 1192 -4568 1288 -4552
rect 1192 -4632 1208 -4568
rect 1272 -4632 1288 -4568
rect 1192 -4648 1288 -4632
rect 1192 -4712 1208 -4648
rect 1272 -4712 1288 -4648
rect 1192 -4728 1288 -4712
rect 1192 -4792 1208 -4728
rect 1272 -4792 1288 -4728
rect 1192 -4808 1288 -4792
rect -220 -4908 -124 -4872
rect 1192 -4872 1208 -4808
rect 1272 -4872 1288 -4808
rect 1611 -4128 2333 -4119
rect 1611 -4832 1620 -4128
rect 2324 -4832 2333 -4128
rect 1611 -4841 2333 -4832
rect 2604 -4152 2620 -4088
rect 2684 -4152 2700 -4088
rect 4016 -4088 4112 -4052
rect 2604 -4168 2700 -4152
rect 2604 -4232 2620 -4168
rect 2684 -4232 2700 -4168
rect 2604 -4248 2700 -4232
rect 2604 -4312 2620 -4248
rect 2684 -4312 2700 -4248
rect 2604 -4328 2700 -4312
rect 2604 -4392 2620 -4328
rect 2684 -4392 2700 -4328
rect 2604 -4408 2700 -4392
rect 2604 -4472 2620 -4408
rect 2684 -4472 2700 -4408
rect 2604 -4488 2700 -4472
rect 2604 -4552 2620 -4488
rect 2684 -4552 2700 -4488
rect 2604 -4568 2700 -4552
rect 2604 -4632 2620 -4568
rect 2684 -4632 2700 -4568
rect 2604 -4648 2700 -4632
rect 2604 -4712 2620 -4648
rect 2684 -4712 2700 -4648
rect 2604 -4728 2700 -4712
rect 2604 -4792 2620 -4728
rect 2684 -4792 2700 -4728
rect 2604 -4808 2700 -4792
rect 1192 -4908 1288 -4872
rect 2604 -4872 2620 -4808
rect 2684 -4872 2700 -4808
rect 3023 -4128 3745 -4119
rect 3023 -4832 3032 -4128
rect 3736 -4832 3745 -4128
rect 3023 -4841 3745 -4832
rect 4016 -4152 4032 -4088
rect 4096 -4152 4112 -4088
rect 5428 -4088 5524 -4052
rect 4016 -4168 4112 -4152
rect 4016 -4232 4032 -4168
rect 4096 -4232 4112 -4168
rect 4016 -4248 4112 -4232
rect 4016 -4312 4032 -4248
rect 4096 -4312 4112 -4248
rect 4016 -4328 4112 -4312
rect 4016 -4392 4032 -4328
rect 4096 -4392 4112 -4328
rect 4016 -4408 4112 -4392
rect 4016 -4472 4032 -4408
rect 4096 -4472 4112 -4408
rect 4016 -4488 4112 -4472
rect 4016 -4552 4032 -4488
rect 4096 -4552 4112 -4488
rect 4016 -4568 4112 -4552
rect 4016 -4632 4032 -4568
rect 4096 -4632 4112 -4568
rect 4016 -4648 4112 -4632
rect 4016 -4712 4032 -4648
rect 4096 -4712 4112 -4648
rect 4016 -4728 4112 -4712
rect 4016 -4792 4032 -4728
rect 4096 -4792 4112 -4728
rect 4016 -4808 4112 -4792
rect 2604 -4908 2700 -4872
rect 4016 -4872 4032 -4808
rect 4096 -4872 4112 -4808
rect 4435 -4128 5157 -4119
rect 4435 -4832 4444 -4128
rect 5148 -4832 5157 -4128
rect 4435 -4841 5157 -4832
rect 5428 -4152 5444 -4088
rect 5508 -4152 5524 -4088
rect 6840 -4088 6936 -4052
rect 5428 -4168 5524 -4152
rect 5428 -4232 5444 -4168
rect 5508 -4232 5524 -4168
rect 5428 -4248 5524 -4232
rect 5428 -4312 5444 -4248
rect 5508 -4312 5524 -4248
rect 5428 -4328 5524 -4312
rect 5428 -4392 5444 -4328
rect 5508 -4392 5524 -4328
rect 5428 -4408 5524 -4392
rect 5428 -4472 5444 -4408
rect 5508 -4472 5524 -4408
rect 5428 -4488 5524 -4472
rect 5428 -4552 5444 -4488
rect 5508 -4552 5524 -4488
rect 5428 -4568 5524 -4552
rect 5428 -4632 5444 -4568
rect 5508 -4632 5524 -4568
rect 5428 -4648 5524 -4632
rect 5428 -4712 5444 -4648
rect 5508 -4712 5524 -4648
rect 5428 -4728 5524 -4712
rect 5428 -4792 5444 -4728
rect 5508 -4792 5524 -4728
rect 5428 -4808 5524 -4792
rect 4016 -4908 4112 -4872
rect 5428 -4872 5444 -4808
rect 5508 -4872 5524 -4808
rect 5847 -4128 6569 -4119
rect 5847 -4832 5856 -4128
rect 6560 -4832 6569 -4128
rect 5847 -4841 6569 -4832
rect 6840 -4152 6856 -4088
rect 6920 -4152 6936 -4088
rect 8252 -4088 8348 -4052
rect 6840 -4168 6936 -4152
rect 6840 -4232 6856 -4168
rect 6920 -4232 6936 -4168
rect 6840 -4248 6936 -4232
rect 6840 -4312 6856 -4248
rect 6920 -4312 6936 -4248
rect 6840 -4328 6936 -4312
rect 6840 -4392 6856 -4328
rect 6920 -4392 6936 -4328
rect 6840 -4408 6936 -4392
rect 6840 -4472 6856 -4408
rect 6920 -4472 6936 -4408
rect 6840 -4488 6936 -4472
rect 6840 -4552 6856 -4488
rect 6920 -4552 6936 -4488
rect 6840 -4568 6936 -4552
rect 6840 -4632 6856 -4568
rect 6920 -4632 6936 -4568
rect 6840 -4648 6936 -4632
rect 6840 -4712 6856 -4648
rect 6920 -4712 6936 -4648
rect 6840 -4728 6936 -4712
rect 6840 -4792 6856 -4728
rect 6920 -4792 6936 -4728
rect 6840 -4808 6936 -4792
rect 5428 -4908 5524 -4872
rect 6840 -4872 6856 -4808
rect 6920 -4872 6936 -4808
rect 7259 -4128 7981 -4119
rect 7259 -4832 7268 -4128
rect 7972 -4832 7981 -4128
rect 7259 -4841 7981 -4832
rect 8252 -4152 8268 -4088
rect 8332 -4152 8348 -4088
rect 9664 -4088 9760 -4052
rect 8252 -4168 8348 -4152
rect 8252 -4232 8268 -4168
rect 8332 -4232 8348 -4168
rect 8252 -4248 8348 -4232
rect 8252 -4312 8268 -4248
rect 8332 -4312 8348 -4248
rect 8252 -4328 8348 -4312
rect 8252 -4392 8268 -4328
rect 8332 -4392 8348 -4328
rect 8252 -4408 8348 -4392
rect 8252 -4472 8268 -4408
rect 8332 -4472 8348 -4408
rect 8252 -4488 8348 -4472
rect 8252 -4552 8268 -4488
rect 8332 -4552 8348 -4488
rect 8252 -4568 8348 -4552
rect 8252 -4632 8268 -4568
rect 8332 -4632 8348 -4568
rect 8252 -4648 8348 -4632
rect 8252 -4712 8268 -4648
rect 8332 -4712 8348 -4648
rect 8252 -4728 8348 -4712
rect 8252 -4792 8268 -4728
rect 8332 -4792 8348 -4728
rect 8252 -4808 8348 -4792
rect 6840 -4908 6936 -4872
rect 8252 -4872 8268 -4808
rect 8332 -4872 8348 -4808
rect 8671 -4128 9393 -4119
rect 8671 -4832 8680 -4128
rect 9384 -4832 9393 -4128
rect 8671 -4841 9393 -4832
rect 9664 -4152 9680 -4088
rect 9744 -4152 9760 -4088
rect 11076 -4088 11172 -4052
rect 9664 -4168 9760 -4152
rect 9664 -4232 9680 -4168
rect 9744 -4232 9760 -4168
rect 9664 -4248 9760 -4232
rect 9664 -4312 9680 -4248
rect 9744 -4312 9760 -4248
rect 9664 -4328 9760 -4312
rect 9664 -4392 9680 -4328
rect 9744 -4392 9760 -4328
rect 9664 -4408 9760 -4392
rect 9664 -4472 9680 -4408
rect 9744 -4472 9760 -4408
rect 9664 -4488 9760 -4472
rect 9664 -4552 9680 -4488
rect 9744 -4552 9760 -4488
rect 9664 -4568 9760 -4552
rect 9664 -4632 9680 -4568
rect 9744 -4632 9760 -4568
rect 9664 -4648 9760 -4632
rect 9664 -4712 9680 -4648
rect 9744 -4712 9760 -4648
rect 9664 -4728 9760 -4712
rect 9664 -4792 9680 -4728
rect 9744 -4792 9760 -4728
rect 9664 -4808 9760 -4792
rect 8252 -4908 8348 -4872
rect 9664 -4872 9680 -4808
rect 9744 -4872 9760 -4808
rect 10083 -4128 10805 -4119
rect 10083 -4832 10092 -4128
rect 10796 -4832 10805 -4128
rect 10083 -4841 10805 -4832
rect 11076 -4152 11092 -4088
rect 11156 -4152 11172 -4088
rect 12488 -4088 12584 -4052
rect 11076 -4168 11172 -4152
rect 11076 -4232 11092 -4168
rect 11156 -4232 11172 -4168
rect 11076 -4248 11172 -4232
rect 11076 -4312 11092 -4248
rect 11156 -4312 11172 -4248
rect 11076 -4328 11172 -4312
rect 11076 -4392 11092 -4328
rect 11156 -4392 11172 -4328
rect 11076 -4408 11172 -4392
rect 11076 -4472 11092 -4408
rect 11156 -4472 11172 -4408
rect 11076 -4488 11172 -4472
rect 11076 -4552 11092 -4488
rect 11156 -4552 11172 -4488
rect 11076 -4568 11172 -4552
rect 11076 -4632 11092 -4568
rect 11156 -4632 11172 -4568
rect 11076 -4648 11172 -4632
rect 11076 -4712 11092 -4648
rect 11156 -4712 11172 -4648
rect 11076 -4728 11172 -4712
rect 11076 -4792 11092 -4728
rect 11156 -4792 11172 -4728
rect 11076 -4808 11172 -4792
rect 9664 -4908 9760 -4872
rect 11076 -4872 11092 -4808
rect 11156 -4872 11172 -4808
rect 11495 -4128 12217 -4119
rect 11495 -4832 11504 -4128
rect 12208 -4832 12217 -4128
rect 11495 -4841 12217 -4832
rect 12488 -4152 12504 -4088
rect 12568 -4152 12584 -4088
rect 13900 -4088 13996 -4052
rect 12488 -4168 12584 -4152
rect 12488 -4232 12504 -4168
rect 12568 -4232 12584 -4168
rect 12488 -4248 12584 -4232
rect 12488 -4312 12504 -4248
rect 12568 -4312 12584 -4248
rect 12488 -4328 12584 -4312
rect 12488 -4392 12504 -4328
rect 12568 -4392 12584 -4328
rect 12488 -4408 12584 -4392
rect 12488 -4472 12504 -4408
rect 12568 -4472 12584 -4408
rect 12488 -4488 12584 -4472
rect 12488 -4552 12504 -4488
rect 12568 -4552 12584 -4488
rect 12488 -4568 12584 -4552
rect 12488 -4632 12504 -4568
rect 12568 -4632 12584 -4568
rect 12488 -4648 12584 -4632
rect 12488 -4712 12504 -4648
rect 12568 -4712 12584 -4648
rect 12488 -4728 12584 -4712
rect 12488 -4792 12504 -4728
rect 12568 -4792 12584 -4728
rect 12488 -4808 12584 -4792
rect 11076 -4908 11172 -4872
rect 12488 -4872 12504 -4808
rect 12568 -4872 12584 -4808
rect 12907 -4128 13629 -4119
rect 12907 -4832 12916 -4128
rect 13620 -4832 13629 -4128
rect 12907 -4841 13629 -4832
rect 13900 -4152 13916 -4088
rect 13980 -4152 13996 -4088
rect 15312 -4088 15408 -4052
rect 13900 -4168 13996 -4152
rect 13900 -4232 13916 -4168
rect 13980 -4232 13996 -4168
rect 13900 -4248 13996 -4232
rect 13900 -4312 13916 -4248
rect 13980 -4312 13996 -4248
rect 13900 -4328 13996 -4312
rect 13900 -4392 13916 -4328
rect 13980 -4392 13996 -4328
rect 13900 -4408 13996 -4392
rect 13900 -4472 13916 -4408
rect 13980 -4472 13996 -4408
rect 13900 -4488 13996 -4472
rect 13900 -4552 13916 -4488
rect 13980 -4552 13996 -4488
rect 13900 -4568 13996 -4552
rect 13900 -4632 13916 -4568
rect 13980 -4632 13996 -4568
rect 13900 -4648 13996 -4632
rect 13900 -4712 13916 -4648
rect 13980 -4712 13996 -4648
rect 13900 -4728 13996 -4712
rect 13900 -4792 13916 -4728
rect 13980 -4792 13996 -4728
rect 13900 -4808 13996 -4792
rect 12488 -4908 12584 -4872
rect 13900 -4872 13916 -4808
rect 13980 -4872 13996 -4808
rect 14319 -4128 15041 -4119
rect 14319 -4832 14328 -4128
rect 15032 -4832 15041 -4128
rect 14319 -4841 15041 -4832
rect 15312 -4152 15328 -4088
rect 15392 -4152 15408 -4088
rect 16724 -4088 16820 -4052
rect 15312 -4168 15408 -4152
rect 15312 -4232 15328 -4168
rect 15392 -4232 15408 -4168
rect 15312 -4248 15408 -4232
rect 15312 -4312 15328 -4248
rect 15392 -4312 15408 -4248
rect 15312 -4328 15408 -4312
rect 15312 -4392 15328 -4328
rect 15392 -4392 15408 -4328
rect 15312 -4408 15408 -4392
rect 15312 -4472 15328 -4408
rect 15392 -4472 15408 -4408
rect 15312 -4488 15408 -4472
rect 15312 -4552 15328 -4488
rect 15392 -4552 15408 -4488
rect 15312 -4568 15408 -4552
rect 15312 -4632 15328 -4568
rect 15392 -4632 15408 -4568
rect 15312 -4648 15408 -4632
rect 15312 -4712 15328 -4648
rect 15392 -4712 15408 -4648
rect 15312 -4728 15408 -4712
rect 15312 -4792 15328 -4728
rect 15392 -4792 15408 -4728
rect 15312 -4808 15408 -4792
rect 13900 -4908 13996 -4872
rect 15312 -4872 15328 -4808
rect 15392 -4872 15408 -4808
rect 15731 -4128 16453 -4119
rect 15731 -4832 15740 -4128
rect 16444 -4832 16453 -4128
rect 15731 -4841 16453 -4832
rect 16724 -4152 16740 -4088
rect 16804 -4152 16820 -4088
rect 18136 -4088 18232 -4052
rect 16724 -4168 16820 -4152
rect 16724 -4232 16740 -4168
rect 16804 -4232 16820 -4168
rect 16724 -4248 16820 -4232
rect 16724 -4312 16740 -4248
rect 16804 -4312 16820 -4248
rect 16724 -4328 16820 -4312
rect 16724 -4392 16740 -4328
rect 16804 -4392 16820 -4328
rect 16724 -4408 16820 -4392
rect 16724 -4472 16740 -4408
rect 16804 -4472 16820 -4408
rect 16724 -4488 16820 -4472
rect 16724 -4552 16740 -4488
rect 16804 -4552 16820 -4488
rect 16724 -4568 16820 -4552
rect 16724 -4632 16740 -4568
rect 16804 -4632 16820 -4568
rect 16724 -4648 16820 -4632
rect 16724 -4712 16740 -4648
rect 16804 -4712 16820 -4648
rect 16724 -4728 16820 -4712
rect 16724 -4792 16740 -4728
rect 16804 -4792 16820 -4728
rect 16724 -4808 16820 -4792
rect 15312 -4908 15408 -4872
rect 16724 -4872 16740 -4808
rect 16804 -4872 16820 -4808
rect 17143 -4128 17865 -4119
rect 17143 -4832 17152 -4128
rect 17856 -4832 17865 -4128
rect 17143 -4841 17865 -4832
rect 18136 -4152 18152 -4088
rect 18216 -4152 18232 -4088
rect 19548 -4088 19644 -4052
rect 18136 -4168 18232 -4152
rect 18136 -4232 18152 -4168
rect 18216 -4232 18232 -4168
rect 18136 -4248 18232 -4232
rect 18136 -4312 18152 -4248
rect 18216 -4312 18232 -4248
rect 18136 -4328 18232 -4312
rect 18136 -4392 18152 -4328
rect 18216 -4392 18232 -4328
rect 18136 -4408 18232 -4392
rect 18136 -4472 18152 -4408
rect 18216 -4472 18232 -4408
rect 18136 -4488 18232 -4472
rect 18136 -4552 18152 -4488
rect 18216 -4552 18232 -4488
rect 18136 -4568 18232 -4552
rect 18136 -4632 18152 -4568
rect 18216 -4632 18232 -4568
rect 18136 -4648 18232 -4632
rect 18136 -4712 18152 -4648
rect 18216 -4712 18232 -4648
rect 18136 -4728 18232 -4712
rect 18136 -4792 18152 -4728
rect 18216 -4792 18232 -4728
rect 18136 -4808 18232 -4792
rect 16724 -4908 16820 -4872
rect 18136 -4872 18152 -4808
rect 18216 -4872 18232 -4808
rect 18555 -4128 19277 -4119
rect 18555 -4832 18564 -4128
rect 19268 -4832 19277 -4128
rect 18555 -4841 19277 -4832
rect 19548 -4152 19564 -4088
rect 19628 -4152 19644 -4088
rect 20960 -4088 21056 -4052
rect 19548 -4168 19644 -4152
rect 19548 -4232 19564 -4168
rect 19628 -4232 19644 -4168
rect 19548 -4248 19644 -4232
rect 19548 -4312 19564 -4248
rect 19628 -4312 19644 -4248
rect 19548 -4328 19644 -4312
rect 19548 -4392 19564 -4328
rect 19628 -4392 19644 -4328
rect 19548 -4408 19644 -4392
rect 19548 -4472 19564 -4408
rect 19628 -4472 19644 -4408
rect 19548 -4488 19644 -4472
rect 19548 -4552 19564 -4488
rect 19628 -4552 19644 -4488
rect 19548 -4568 19644 -4552
rect 19548 -4632 19564 -4568
rect 19628 -4632 19644 -4568
rect 19548 -4648 19644 -4632
rect 19548 -4712 19564 -4648
rect 19628 -4712 19644 -4648
rect 19548 -4728 19644 -4712
rect 19548 -4792 19564 -4728
rect 19628 -4792 19644 -4728
rect 19548 -4808 19644 -4792
rect 18136 -4908 18232 -4872
rect 19548 -4872 19564 -4808
rect 19628 -4872 19644 -4808
rect 19967 -4128 20689 -4119
rect 19967 -4832 19976 -4128
rect 20680 -4832 20689 -4128
rect 19967 -4841 20689 -4832
rect 20960 -4152 20976 -4088
rect 21040 -4152 21056 -4088
rect 22372 -4088 22468 -4052
rect 20960 -4168 21056 -4152
rect 20960 -4232 20976 -4168
rect 21040 -4232 21056 -4168
rect 20960 -4248 21056 -4232
rect 20960 -4312 20976 -4248
rect 21040 -4312 21056 -4248
rect 20960 -4328 21056 -4312
rect 20960 -4392 20976 -4328
rect 21040 -4392 21056 -4328
rect 20960 -4408 21056 -4392
rect 20960 -4472 20976 -4408
rect 21040 -4472 21056 -4408
rect 20960 -4488 21056 -4472
rect 20960 -4552 20976 -4488
rect 21040 -4552 21056 -4488
rect 20960 -4568 21056 -4552
rect 20960 -4632 20976 -4568
rect 21040 -4632 21056 -4568
rect 20960 -4648 21056 -4632
rect 20960 -4712 20976 -4648
rect 21040 -4712 21056 -4648
rect 20960 -4728 21056 -4712
rect 20960 -4792 20976 -4728
rect 21040 -4792 21056 -4728
rect 20960 -4808 21056 -4792
rect 19548 -4908 19644 -4872
rect 20960 -4872 20976 -4808
rect 21040 -4872 21056 -4808
rect 21379 -4128 22101 -4119
rect 21379 -4832 21388 -4128
rect 22092 -4832 22101 -4128
rect 21379 -4841 22101 -4832
rect 22372 -4152 22388 -4088
rect 22452 -4152 22468 -4088
rect 23784 -4088 23880 -4052
rect 22372 -4168 22468 -4152
rect 22372 -4232 22388 -4168
rect 22452 -4232 22468 -4168
rect 22372 -4248 22468 -4232
rect 22372 -4312 22388 -4248
rect 22452 -4312 22468 -4248
rect 22372 -4328 22468 -4312
rect 22372 -4392 22388 -4328
rect 22452 -4392 22468 -4328
rect 22372 -4408 22468 -4392
rect 22372 -4472 22388 -4408
rect 22452 -4472 22468 -4408
rect 22372 -4488 22468 -4472
rect 22372 -4552 22388 -4488
rect 22452 -4552 22468 -4488
rect 22372 -4568 22468 -4552
rect 22372 -4632 22388 -4568
rect 22452 -4632 22468 -4568
rect 22372 -4648 22468 -4632
rect 22372 -4712 22388 -4648
rect 22452 -4712 22468 -4648
rect 22372 -4728 22468 -4712
rect 22372 -4792 22388 -4728
rect 22452 -4792 22468 -4728
rect 22372 -4808 22468 -4792
rect 20960 -4908 21056 -4872
rect 22372 -4872 22388 -4808
rect 22452 -4872 22468 -4808
rect 22791 -4128 23513 -4119
rect 22791 -4832 22800 -4128
rect 23504 -4832 23513 -4128
rect 22791 -4841 23513 -4832
rect 23784 -4152 23800 -4088
rect 23864 -4152 23880 -4088
rect 23784 -4168 23880 -4152
rect 23784 -4232 23800 -4168
rect 23864 -4232 23880 -4168
rect 23784 -4248 23880 -4232
rect 23784 -4312 23800 -4248
rect 23864 -4312 23880 -4248
rect 23784 -4328 23880 -4312
rect 23784 -4392 23800 -4328
rect 23864 -4392 23880 -4328
rect 23784 -4408 23880 -4392
rect 23784 -4472 23800 -4408
rect 23864 -4472 23880 -4408
rect 23784 -4488 23880 -4472
rect 23784 -4552 23800 -4488
rect 23864 -4552 23880 -4488
rect 23784 -4568 23880 -4552
rect 23784 -4632 23800 -4568
rect 23864 -4632 23880 -4568
rect 23784 -4648 23880 -4632
rect 23784 -4712 23800 -4648
rect 23864 -4712 23880 -4648
rect 23784 -4728 23880 -4712
rect 23784 -4792 23800 -4728
rect 23864 -4792 23880 -4728
rect 23784 -4808 23880 -4792
rect 22372 -4908 22468 -4872
rect 23784 -4872 23800 -4808
rect 23864 -4872 23880 -4808
rect 23784 -4908 23880 -4872
rect -22812 -5208 -22716 -5172
rect -23805 -5248 -23083 -5239
rect -23805 -5952 -23796 -5248
rect -23092 -5952 -23083 -5248
rect -23805 -5961 -23083 -5952
rect -22812 -5272 -22796 -5208
rect -22732 -5272 -22716 -5208
rect -21400 -5208 -21304 -5172
rect -22812 -5288 -22716 -5272
rect -22812 -5352 -22796 -5288
rect -22732 -5352 -22716 -5288
rect -22812 -5368 -22716 -5352
rect -22812 -5432 -22796 -5368
rect -22732 -5432 -22716 -5368
rect -22812 -5448 -22716 -5432
rect -22812 -5512 -22796 -5448
rect -22732 -5512 -22716 -5448
rect -22812 -5528 -22716 -5512
rect -22812 -5592 -22796 -5528
rect -22732 -5592 -22716 -5528
rect -22812 -5608 -22716 -5592
rect -22812 -5672 -22796 -5608
rect -22732 -5672 -22716 -5608
rect -22812 -5688 -22716 -5672
rect -22812 -5752 -22796 -5688
rect -22732 -5752 -22716 -5688
rect -22812 -5768 -22716 -5752
rect -22812 -5832 -22796 -5768
rect -22732 -5832 -22716 -5768
rect -22812 -5848 -22716 -5832
rect -22812 -5912 -22796 -5848
rect -22732 -5912 -22716 -5848
rect -22812 -5928 -22716 -5912
rect -22812 -5992 -22796 -5928
rect -22732 -5992 -22716 -5928
rect -22393 -5248 -21671 -5239
rect -22393 -5952 -22384 -5248
rect -21680 -5952 -21671 -5248
rect -22393 -5961 -21671 -5952
rect -21400 -5272 -21384 -5208
rect -21320 -5272 -21304 -5208
rect -19988 -5208 -19892 -5172
rect -21400 -5288 -21304 -5272
rect -21400 -5352 -21384 -5288
rect -21320 -5352 -21304 -5288
rect -21400 -5368 -21304 -5352
rect -21400 -5432 -21384 -5368
rect -21320 -5432 -21304 -5368
rect -21400 -5448 -21304 -5432
rect -21400 -5512 -21384 -5448
rect -21320 -5512 -21304 -5448
rect -21400 -5528 -21304 -5512
rect -21400 -5592 -21384 -5528
rect -21320 -5592 -21304 -5528
rect -21400 -5608 -21304 -5592
rect -21400 -5672 -21384 -5608
rect -21320 -5672 -21304 -5608
rect -21400 -5688 -21304 -5672
rect -21400 -5752 -21384 -5688
rect -21320 -5752 -21304 -5688
rect -21400 -5768 -21304 -5752
rect -21400 -5832 -21384 -5768
rect -21320 -5832 -21304 -5768
rect -21400 -5848 -21304 -5832
rect -21400 -5912 -21384 -5848
rect -21320 -5912 -21304 -5848
rect -21400 -5928 -21304 -5912
rect -22812 -6028 -22716 -5992
rect -21400 -5992 -21384 -5928
rect -21320 -5992 -21304 -5928
rect -20981 -5248 -20259 -5239
rect -20981 -5952 -20972 -5248
rect -20268 -5952 -20259 -5248
rect -20981 -5961 -20259 -5952
rect -19988 -5272 -19972 -5208
rect -19908 -5272 -19892 -5208
rect -18576 -5208 -18480 -5172
rect -19988 -5288 -19892 -5272
rect -19988 -5352 -19972 -5288
rect -19908 -5352 -19892 -5288
rect -19988 -5368 -19892 -5352
rect -19988 -5432 -19972 -5368
rect -19908 -5432 -19892 -5368
rect -19988 -5448 -19892 -5432
rect -19988 -5512 -19972 -5448
rect -19908 -5512 -19892 -5448
rect -19988 -5528 -19892 -5512
rect -19988 -5592 -19972 -5528
rect -19908 -5592 -19892 -5528
rect -19988 -5608 -19892 -5592
rect -19988 -5672 -19972 -5608
rect -19908 -5672 -19892 -5608
rect -19988 -5688 -19892 -5672
rect -19988 -5752 -19972 -5688
rect -19908 -5752 -19892 -5688
rect -19988 -5768 -19892 -5752
rect -19988 -5832 -19972 -5768
rect -19908 -5832 -19892 -5768
rect -19988 -5848 -19892 -5832
rect -19988 -5912 -19972 -5848
rect -19908 -5912 -19892 -5848
rect -19988 -5928 -19892 -5912
rect -21400 -6028 -21304 -5992
rect -19988 -5992 -19972 -5928
rect -19908 -5992 -19892 -5928
rect -19569 -5248 -18847 -5239
rect -19569 -5952 -19560 -5248
rect -18856 -5952 -18847 -5248
rect -19569 -5961 -18847 -5952
rect -18576 -5272 -18560 -5208
rect -18496 -5272 -18480 -5208
rect -17164 -5208 -17068 -5172
rect -18576 -5288 -18480 -5272
rect -18576 -5352 -18560 -5288
rect -18496 -5352 -18480 -5288
rect -18576 -5368 -18480 -5352
rect -18576 -5432 -18560 -5368
rect -18496 -5432 -18480 -5368
rect -18576 -5448 -18480 -5432
rect -18576 -5512 -18560 -5448
rect -18496 -5512 -18480 -5448
rect -18576 -5528 -18480 -5512
rect -18576 -5592 -18560 -5528
rect -18496 -5592 -18480 -5528
rect -18576 -5608 -18480 -5592
rect -18576 -5672 -18560 -5608
rect -18496 -5672 -18480 -5608
rect -18576 -5688 -18480 -5672
rect -18576 -5752 -18560 -5688
rect -18496 -5752 -18480 -5688
rect -18576 -5768 -18480 -5752
rect -18576 -5832 -18560 -5768
rect -18496 -5832 -18480 -5768
rect -18576 -5848 -18480 -5832
rect -18576 -5912 -18560 -5848
rect -18496 -5912 -18480 -5848
rect -18576 -5928 -18480 -5912
rect -19988 -6028 -19892 -5992
rect -18576 -5992 -18560 -5928
rect -18496 -5992 -18480 -5928
rect -18157 -5248 -17435 -5239
rect -18157 -5952 -18148 -5248
rect -17444 -5952 -17435 -5248
rect -18157 -5961 -17435 -5952
rect -17164 -5272 -17148 -5208
rect -17084 -5272 -17068 -5208
rect -15752 -5208 -15656 -5172
rect -17164 -5288 -17068 -5272
rect -17164 -5352 -17148 -5288
rect -17084 -5352 -17068 -5288
rect -17164 -5368 -17068 -5352
rect -17164 -5432 -17148 -5368
rect -17084 -5432 -17068 -5368
rect -17164 -5448 -17068 -5432
rect -17164 -5512 -17148 -5448
rect -17084 -5512 -17068 -5448
rect -17164 -5528 -17068 -5512
rect -17164 -5592 -17148 -5528
rect -17084 -5592 -17068 -5528
rect -17164 -5608 -17068 -5592
rect -17164 -5672 -17148 -5608
rect -17084 -5672 -17068 -5608
rect -17164 -5688 -17068 -5672
rect -17164 -5752 -17148 -5688
rect -17084 -5752 -17068 -5688
rect -17164 -5768 -17068 -5752
rect -17164 -5832 -17148 -5768
rect -17084 -5832 -17068 -5768
rect -17164 -5848 -17068 -5832
rect -17164 -5912 -17148 -5848
rect -17084 -5912 -17068 -5848
rect -17164 -5928 -17068 -5912
rect -18576 -6028 -18480 -5992
rect -17164 -5992 -17148 -5928
rect -17084 -5992 -17068 -5928
rect -16745 -5248 -16023 -5239
rect -16745 -5952 -16736 -5248
rect -16032 -5952 -16023 -5248
rect -16745 -5961 -16023 -5952
rect -15752 -5272 -15736 -5208
rect -15672 -5272 -15656 -5208
rect -14340 -5208 -14244 -5172
rect -15752 -5288 -15656 -5272
rect -15752 -5352 -15736 -5288
rect -15672 -5352 -15656 -5288
rect -15752 -5368 -15656 -5352
rect -15752 -5432 -15736 -5368
rect -15672 -5432 -15656 -5368
rect -15752 -5448 -15656 -5432
rect -15752 -5512 -15736 -5448
rect -15672 -5512 -15656 -5448
rect -15752 -5528 -15656 -5512
rect -15752 -5592 -15736 -5528
rect -15672 -5592 -15656 -5528
rect -15752 -5608 -15656 -5592
rect -15752 -5672 -15736 -5608
rect -15672 -5672 -15656 -5608
rect -15752 -5688 -15656 -5672
rect -15752 -5752 -15736 -5688
rect -15672 -5752 -15656 -5688
rect -15752 -5768 -15656 -5752
rect -15752 -5832 -15736 -5768
rect -15672 -5832 -15656 -5768
rect -15752 -5848 -15656 -5832
rect -15752 -5912 -15736 -5848
rect -15672 -5912 -15656 -5848
rect -15752 -5928 -15656 -5912
rect -17164 -6028 -17068 -5992
rect -15752 -5992 -15736 -5928
rect -15672 -5992 -15656 -5928
rect -15333 -5248 -14611 -5239
rect -15333 -5952 -15324 -5248
rect -14620 -5952 -14611 -5248
rect -15333 -5961 -14611 -5952
rect -14340 -5272 -14324 -5208
rect -14260 -5272 -14244 -5208
rect -12928 -5208 -12832 -5172
rect -14340 -5288 -14244 -5272
rect -14340 -5352 -14324 -5288
rect -14260 -5352 -14244 -5288
rect -14340 -5368 -14244 -5352
rect -14340 -5432 -14324 -5368
rect -14260 -5432 -14244 -5368
rect -14340 -5448 -14244 -5432
rect -14340 -5512 -14324 -5448
rect -14260 -5512 -14244 -5448
rect -14340 -5528 -14244 -5512
rect -14340 -5592 -14324 -5528
rect -14260 -5592 -14244 -5528
rect -14340 -5608 -14244 -5592
rect -14340 -5672 -14324 -5608
rect -14260 -5672 -14244 -5608
rect -14340 -5688 -14244 -5672
rect -14340 -5752 -14324 -5688
rect -14260 -5752 -14244 -5688
rect -14340 -5768 -14244 -5752
rect -14340 -5832 -14324 -5768
rect -14260 -5832 -14244 -5768
rect -14340 -5848 -14244 -5832
rect -14340 -5912 -14324 -5848
rect -14260 -5912 -14244 -5848
rect -14340 -5928 -14244 -5912
rect -15752 -6028 -15656 -5992
rect -14340 -5992 -14324 -5928
rect -14260 -5992 -14244 -5928
rect -13921 -5248 -13199 -5239
rect -13921 -5952 -13912 -5248
rect -13208 -5952 -13199 -5248
rect -13921 -5961 -13199 -5952
rect -12928 -5272 -12912 -5208
rect -12848 -5272 -12832 -5208
rect -11516 -5208 -11420 -5172
rect -12928 -5288 -12832 -5272
rect -12928 -5352 -12912 -5288
rect -12848 -5352 -12832 -5288
rect -12928 -5368 -12832 -5352
rect -12928 -5432 -12912 -5368
rect -12848 -5432 -12832 -5368
rect -12928 -5448 -12832 -5432
rect -12928 -5512 -12912 -5448
rect -12848 -5512 -12832 -5448
rect -12928 -5528 -12832 -5512
rect -12928 -5592 -12912 -5528
rect -12848 -5592 -12832 -5528
rect -12928 -5608 -12832 -5592
rect -12928 -5672 -12912 -5608
rect -12848 -5672 -12832 -5608
rect -12928 -5688 -12832 -5672
rect -12928 -5752 -12912 -5688
rect -12848 -5752 -12832 -5688
rect -12928 -5768 -12832 -5752
rect -12928 -5832 -12912 -5768
rect -12848 -5832 -12832 -5768
rect -12928 -5848 -12832 -5832
rect -12928 -5912 -12912 -5848
rect -12848 -5912 -12832 -5848
rect -12928 -5928 -12832 -5912
rect -14340 -6028 -14244 -5992
rect -12928 -5992 -12912 -5928
rect -12848 -5992 -12832 -5928
rect -12509 -5248 -11787 -5239
rect -12509 -5952 -12500 -5248
rect -11796 -5952 -11787 -5248
rect -12509 -5961 -11787 -5952
rect -11516 -5272 -11500 -5208
rect -11436 -5272 -11420 -5208
rect -10104 -5208 -10008 -5172
rect -11516 -5288 -11420 -5272
rect -11516 -5352 -11500 -5288
rect -11436 -5352 -11420 -5288
rect -11516 -5368 -11420 -5352
rect -11516 -5432 -11500 -5368
rect -11436 -5432 -11420 -5368
rect -11516 -5448 -11420 -5432
rect -11516 -5512 -11500 -5448
rect -11436 -5512 -11420 -5448
rect -11516 -5528 -11420 -5512
rect -11516 -5592 -11500 -5528
rect -11436 -5592 -11420 -5528
rect -11516 -5608 -11420 -5592
rect -11516 -5672 -11500 -5608
rect -11436 -5672 -11420 -5608
rect -11516 -5688 -11420 -5672
rect -11516 -5752 -11500 -5688
rect -11436 -5752 -11420 -5688
rect -11516 -5768 -11420 -5752
rect -11516 -5832 -11500 -5768
rect -11436 -5832 -11420 -5768
rect -11516 -5848 -11420 -5832
rect -11516 -5912 -11500 -5848
rect -11436 -5912 -11420 -5848
rect -11516 -5928 -11420 -5912
rect -12928 -6028 -12832 -5992
rect -11516 -5992 -11500 -5928
rect -11436 -5992 -11420 -5928
rect -11097 -5248 -10375 -5239
rect -11097 -5952 -11088 -5248
rect -10384 -5952 -10375 -5248
rect -11097 -5961 -10375 -5952
rect -10104 -5272 -10088 -5208
rect -10024 -5272 -10008 -5208
rect -8692 -5208 -8596 -5172
rect -10104 -5288 -10008 -5272
rect -10104 -5352 -10088 -5288
rect -10024 -5352 -10008 -5288
rect -10104 -5368 -10008 -5352
rect -10104 -5432 -10088 -5368
rect -10024 -5432 -10008 -5368
rect -10104 -5448 -10008 -5432
rect -10104 -5512 -10088 -5448
rect -10024 -5512 -10008 -5448
rect -10104 -5528 -10008 -5512
rect -10104 -5592 -10088 -5528
rect -10024 -5592 -10008 -5528
rect -10104 -5608 -10008 -5592
rect -10104 -5672 -10088 -5608
rect -10024 -5672 -10008 -5608
rect -10104 -5688 -10008 -5672
rect -10104 -5752 -10088 -5688
rect -10024 -5752 -10008 -5688
rect -10104 -5768 -10008 -5752
rect -10104 -5832 -10088 -5768
rect -10024 -5832 -10008 -5768
rect -10104 -5848 -10008 -5832
rect -10104 -5912 -10088 -5848
rect -10024 -5912 -10008 -5848
rect -10104 -5928 -10008 -5912
rect -11516 -6028 -11420 -5992
rect -10104 -5992 -10088 -5928
rect -10024 -5992 -10008 -5928
rect -9685 -5248 -8963 -5239
rect -9685 -5952 -9676 -5248
rect -8972 -5952 -8963 -5248
rect -9685 -5961 -8963 -5952
rect -8692 -5272 -8676 -5208
rect -8612 -5272 -8596 -5208
rect -7280 -5208 -7184 -5172
rect -8692 -5288 -8596 -5272
rect -8692 -5352 -8676 -5288
rect -8612 -5352 -8596 -5288
rect -8692 -5368 -8596 -5352
rect -8692 -5432 -8676 -5368
rect -8612 -5432 -8596 -5368
rect -8692 -5448 -8596 -5432
rect -8692 -5512 -8676 -5448
rect -8612 -5512 -8596 -5448
rect -8692 -5528 -8596 -5512
rect -8692 -5592 -8676 -5528
rect -8612 -5592 -8596 -5528
rect -8692 -5608 -8596 -5592
rect -8692 -5672 -8676 -5608
rect -8612 -5672 -8596 -5608
rect -8692 -5688 -8596 -5672
rect -8692 -5752 -8676 -5688
rect -8612 -5752 -8596 -5688
rect -8692 -5768 -8596 -5752
rect -8692 -5832 -8676 -5768
rect -8612 -5832 -8596 -5768
rect -8692 -5848 -8596 -5832
rect -8692 -5912 -8676 -5848
rect -8612 -5912 -8596 -5848
rect -8692 -5928 -8596 -5912
rect -10104 -6028 -10008 -5992
rect -8692 -5992 -8676 -5928
rect -8612 -5992 -8596 -5928
rect -8273 -5248 -7551 -5239
rect -8273 -5952 -8264 -5248
rect -7560 -5952 -7551 -5248
rect -8273 -5961 -7551 -5952
rect -7280 -5272 -7264 -5208
rect -7200 -5272 -7184 -5208
rect -5868 -5208 -5772 -5172
rect -7280 -5288 -7184 -5272
rect -7280 -5352 -7264 -5288
rect -7200 -5352 -7184 -5288
rect -7280 -5368 -7184 -5352
rect -7280 -5432 -7264 -5368
rect -7200 -5432 -7184 -5368
rect -7280 -5448 -7184 -5432
rect -7280 -5512 -7264 -5448
rect -7200 -5512 -7184 -5448
rect -7280 -5528 -7184 -5512
rect -7280 -5592 -7264 -5528
rect -7200 -5592 -7184 -5528
rect -7280 -5608 -7184 -5592
rect -7280 -5672 -7264 -5608
rect -7200 -5672 -7184 -5608
rect -7280 -5688 -7184 -5672
rect -7280 -5752 -7264 -5688
rect -7200 -5752 -7184 -5688
rect -7280 -5768 -7184 -5752
rect -7280 -5832 -7264 -5768
rect -7200 -5832 -7184 -5768
rect -7280 -5848 -7184 -5832
rect -7280 -5912 -7264 -5848
rect -7200 -5912 -7184 -5848
rect -7280 -5928 -7184 -5912
rect -8692 -6028 -8596 -5992
rect -7280 -5992 -7264 -5928
rect -7200 -5992 -7184 -5928
rect -6861 -5248 -6139 -5239
rect -6861 -5952 -6852 -5248
rect -6148 -5952 -6139 -5248
rect -6861 -5961 -6139 -5952
rect -5868 -5272 -5852 -5208
rect -5788 -5272 -5772 -5208
rect -4456 -5208 -4360 -5172
rect -5868 -5288 -5772 -5272
rect -5868 -5352 -5852 -5288
rect -5788 -5352 -5772 -5288
rect -5868 -5368 -5772 -5352
rect -5868 -5432 -5852 -5368
rect -5788 -5432 -5772 -5368
rect -5868 -5448 -5772 -5432
rect -5868 -5512 -5852 -5448
rect -5788 -5512 -5772 -5448
rect -5868 -5528 -5772 -5512
rect -5868 -5592 -5852 -5528
rect -5788 -5592 -5772 -5528
rect -5868 -5608 -5772 -5592
rect -5868 -5672 -5852 -5608
rect -5788 -5672 -5772 -5608
rect -5868 -5688 -5772 -5672
rect -5868 -5752 -5852 -5688
rect -5788 -5752 -5772 -5688
rect -5868 -5768 -5772 -5752
rect -5868 -5832 -5852 -5768
rect -5788 -5832 -5772 -5768
rect -5868 -5848 -5772 -5832
rect -5868 -5912 -5852 -5848
rect -5788 -5912 -5772 -5848
rect -5868 -5928 -5772 -5912
rect -7280 -6028 -7184 -5992
rect -5868 -5992 -5852 -5928
rect -5788 -5992 -5772 -5928
rect -5449 -5248 -4727 -5239
rect -5449 -5952 -5440 -5248
rect -4736 -5952 -4727 -5248
rect -5449 -5961 -4727 -5952
rect -4456 -5272 -4440 -5208
rect -4376 -5272 -4360 -5208
rect -3044 -5208 -2948 -5172
rect -4456 -5288 -4360 -5272
rect -4456 -5352 -4440 -5288
rect -4376 -5352 -4360 -5288
rect -4456 -5368 -4360 -5352
rect -4456 -5432 -4440 -5368
rect -4376 -5432 -4360 -5368
rect -4456 -5448 -4360 -5432
rect -4456 -5512 -4440 -5448
rect -4376 -5512 -4360 -5448
rect -4456 -5528 -4360 -5512
rect -4456 -5592 -4440 -5528
rect -4376 -5592 -4360 -5528
rect -4456 -5608 -4360 -5592
rect -4456 -5672 -4440 -5608
rect -4376 -5672 -4360 -5608
rect -4456 -5688 -4360 -5672
rect -4456 -5752 -4440 -5688
rect -4376 -5752 -4360 -5688
rect -4456 -5768 -4360 -5752
rect -4456 -5832 -4440 -5768
rect -4376 -5832 -4360 -5768
rect -4456 -5848 -4360 -5832
rect -4456 -5912 -4440 -5848
rect -4376 -5912 -4360 -5848
rect -4456 -5928 -4360 -5912
rect -5868 -6028 -5772 -5992
rect -4456 -5992 -4440 -5928
rect -4376 -5992 -4360 -5928
rect -4037 -5248 -3315 -5239
rect -4037 -5952 -4028 -5248
rect -3324 -5952 -3315 -5248
rect -4037 -5961 -3315 -5952
rect -3044 -5272 -3028 -5208
rect -2964 -5272 -2948 -5208
rect -1632 -5208 -1536 -5172
rect -3044 -5288 -2948 -5272
rect -3044 -5352 -3028 -5288
rect -2964 -5352 -2948 -5288
rect -3044 -5368 -2948 -5352
rect -3044 -5432 -3028 -5368
rect -2964 -5432 -2948 -5368
rect -3044 -5448 -2948 -5432
rect -3044 -5512 -3028 -5448
rect -2964 -5512 -2948 -5448
rect -3044 -5528 -2948 -5512
rect -3044 -5592 -3028 -5528
rect -2964 -5592 -2948 -5528
rect -3044 -5608 -2948 -5592
rect -3044 -5672 -3028 -5608
rect -2964 -5672 -2948 -5608
rect -3044 -5688 -2948 -5672
rect -3044 -5752 -3028 -5688
rect -2964 -5752 -2948 -5688
rect -3044 -5768 -2948 -5752
rect -3044 -5832 -3028 -5768
rect -2964 -5832 -2948 -5768
rect -3044 -5848 -2948 -5832
rect -3044 -5912 -3028 -5848
rect -2964 -5912 -2948 -5848
rect -3044 -5928 -2948 -5912
rect -4456 -6028 -4360 -5992
rect -3044 -5992 -3028 -5928
rect -2964 -5992 -2948 -5928
rect -2625 -5248 -1903 -5239
rect -2625 -5952 -2616 -5248
rect -1912 -5952 -1903 -5248
rect -2625 -5961 -1903 -5952
rect -1632 -5272 -1616 -5208
rect -1552 -5272 -1536 -5208
rect -220 -5208 -124 -5172
rect -1632 -5288 -1536 -5272
rect -1632 -5352 -1616 -5288
rect -1552 -5352 -1536 -5288
rect -1632 -5368 -1536 -5352
rect -1632 -5432 -1616 -5368
rect -1552 -5432 -1536 -5368
rect -1632 -5448 -1536 -5432
rect -1632 -5512 -1616 -5448
rect -1552 -5512 -1536 -5448
rect -1632 -5528 -1536 -5512
rect -1632 -5592 -1616 -5528
rect -1552 -5592 -1536 -5528
rect -1632 -5608 -1536 -5592
rect -1632 -5672 -1616 -5608
rect -1552 -5672 -1536 -5608
rect -1632 -5688 -1536 -5672
rect -1632 -5752 -1616 -5688
rect -1552 -5752 -1536 -5688
rect -1632 -5768 -1536 -5752
rect -1632 -5832 -1616 -5768
rect -1552 -5832 -1536 -5768
rect -1632 -5848 -1536 -5832
rect -1632 -5912 -1616 -5848
rect -1552 -5912 -1536 -5848
rect -1632 -5928 -1536 -5912
rect -3044 -6028 -2948 -5992
rect -1632 -5992 -1616 -5928
rect -1552 -5992 -1536 -5928
rect -1213 -5248 -491 -5239
rect -1213 -5952 -1204 -5248
rect -500 -5952 -491 -5248
rect -1213 -5961 -491 -5952
rect -220 -5272 -204 -5208
rect -140 -5272 -124 -5208
rect 1192 -5208 1288 -5172
rect -220 -5288 -124 -5272
rect -220 -5352 -204 -5288
rect -140 -5352 -124 -5288
rect -220 -5368 -124 -5352
rect -220 -5432 -204 -5368
rect -140 -5432 -124 -5368
rect -220 -5448 -124 -5432
rect -220 -5512 -204 -5448
rect -140 -5512 -124 -5448
rect -220 -5528 -124 -5512
rect -220 -5592 -204 -5528
rect -140 -5592 -124 -5528
rect -220 -5608 -124 -5592
rect -220 -5672 -204 -5608
rect -140 -5672 -124 -5608
rect -220 -5688 -124 -5672
rect -220 -5752 -204 -5688
rect -140 -5752 -124 -5688
rect -220 -5768 -124 -5752
rect -220 -5832 -204 -5768
rect -140 -5832 -124 -5768
rect -220 -5848 -124 -5832
rect -220 -5912 -204 -5848
rect -140 -5912 -124 -5848
rect -220 -5928 -124 -5912
rect -1632 -6028 -1536 -5992
rect -220 -5992 -204 -5928
rect -140 -5992 -124 -5928
rect 199 -5248 921 -5239
rect 199 -5952 208 -5248
rect 912 -5952 921 -5248
rect 199 -5961 921 -5952
rect 1192 -5272 1208 -5208
rect 1272 -5272 1288 -5208
rect 2604 -5208 2700 -5172
rect 1192 -5288 1288 -5272
rect 1192 -5352 1208 -5288
rect 1272 -5352 1288 -5288
rect 1192 -5368 1288 -5352
rect 1192 -5432 1208 -5368
rect 1272 -5432 1288 -5368
rect 1192 -5448 1288 -5432
rect 1192 -5512 1208 -5448
rect 1272 -5512 1288 -5448
rect 1192 -5528 1288 -5512
rect 1192 -5592 1208 -5528
rect 1272 -5592 1288 -5528
rect 1192 -5608 1288 -5592
rect 1192 -5672 1208 -5608
rect 1272 -5672 1288 -5608
rect 1192 -5688 1288 -5672
rect 1192 -5752 1208 -5688
rect 1272 -5752 1288 -5688
rect 1192 -5768 1288 -5752
rect 1192 -5832 1208 -5768
rect 1272 -5832 1288 -5768
rect 1192 -5848 1288 -5832
rect 1192 -5912 1208 -5848
rect 1272 -5912 1288 -5848
rect 1192 -5928 1288 -5912
rect -220 -6028 -124 -5992
rect 1192 -5992 1208 -5928
rect 1272 -5992 1288 -5928
rect 1611 -5248 2333 -5239
rect 1611 -5952 1620 -5248
rect 2324 -5952 2333 -5248
rect 1611 -5961 2333 -5952
rect 2604 -5272 2620 -5208
rect 2684 -5272 2700 -5208
rect 4016 -5208 4112 -5172
rect 2604 -5288 2700 -5272
rect 2604 -5352 2620 -5288
rect 2684 -5352 2700 -5288
rect 2604 -5368 2700 -5352
rect 2604 -5432 2620 -5368
rect 2684 -5432 2700 -5368
rect 2604 -5448 2700 -5432
rect 2604 -5512 2620 -5448
rect 2684 -5512 2700 -5448
rect 2604 -5528 2700 -5512
rect 2604 -5592 2620 -5528
rect 2684 -5592 2700 -5528
rect 2604 -5608 2700 -5592
rect 2604 -5672 2620 -5608
rect 2684 -5672 2700 -5608
rect 2604 -5688 2700 -5672
rect 2604 -5752 2620 -5688
rect 2684 -5752 2700 -5688
rect 2604 -5768 2700 -5752
rect 2604 -5832 2620 -5768
rect 2684 -5832 2700 -5768
rect 2604 -5848 2700 -5832
rect 2604 -5912 2620 -5848
rect 2684 -5912 2700 -5848
rect 2604 -5928 2700 -5912
rect 1192 -6028 1288 -5992
rect 2604 -5992 2620 -5928
rect 2684 -5992 2700 -5928
rect 3023 -5248 3745 -5239
rect 3023 -5952 3032 -5248
rect 3736 -5952 3745 -5248
rect 3023 -5961 3745 -5952
rect 4016 -5272 4032 -5208
rect 4096 -5272 4112 -5208
rect 5428 -5208 5524 -5172
rect 4016 -5288 4112 -5272
rect 4016 -5352 4032 -5288
rect 4096 -5352 4112 -5288
rect 4016 -5368 4112 -5352
rect 4016 -5432 4032 -5368
rect 4096 -5432 4112 -5368
rect 4016 -5448 4112 -5432
rect 4016 -5512 4032 -5448
rect 4096 -5512 4112 -5448
rect 4016 -5528 4112 -5512
rect 4016 -5592 4032 -5528
rect 4096 -5592 4112 -5528
rect 4016 -5608 4112 -5592
rect 4016 -5672 4032 -5608
rect 4096 -5672 4112 -5608
rect 4016 -5688 4112 -5672
rect 4016 -5752 4032 -5688
rect 4096 -5752 4112 -5688
rect 4016 -5768 4112 -5752
rect 4016 -5832 4032 -5768
rect 4096 -5832 4112 -5768
rect 4016 -5848 4112 -5832
rect 4016 -5912 4032 -5848
rect 4096 -5912 4112 -5848
rect 4016 -5928 4112 -5912
rect 2604 -6028 2700 -5992
rect 4016 -5992 4032 -5928
rect 4096 -5992 4112 -5928
rect 4435 -5248 5157 -5239
rect 4435 -5952 4444 -5248
rect 5148 -5952 5157 -5248
rect 4435 -5961 5157 -5952
rect 5428 -5272 5444 -5208
rect 5508 -5272 5524 -5208
rect 6840 -5208 6936 -5172
rect 5428 -5288 5524 -5272
rect 5428 -5352 5444 -5288
rect 5508 -5352 5524 -5288
rect 5428 -5368 5524 -5352
rect 5428 -5432 5444 -5368
rect 5508 -5432 5524 -5368
rect 5428 -5448 5524 -5432
rect 5428 -5512 5444 -5448
rect 5508 -5512 5524 -5448
rect 5428 -5528 5524 -5512
rect 5428 -5592 5444 -5528
rect 5508 -5592 5524 -5528
rect 5428 -5608 5524 -5592
rect 5428 -5672 5444 -5608
rect 5508 -5672 5524 -5608
rect 5428 -5688 5524 -5672
rect 5428 -5752 5444 -5688
rect 5508 -5752 5524 -5688
rect 5428 -5768 5524 -5752
rect 5428 -5832 5444 -5768
rect 5508 -5832 5524 -5768
rect 5428 -5848 5524 -5832
rect 5428 -5912 5444 -5848
rect 5508 -5912 5524 -5848
rect 5428 -5928 5524 -5912
rect 4016 -6028 4112 -5992
rect 5428 -5992 5444 -5928
rect 5508 -5992 5524 -5928
rect 5847 -5248 6569 -5239
rect 5847 -5952 5856 -5248
rect 6560 -5952 6569 -5248
rect 5847 -5961 6569 -5952
rect 6840 -5272 6856 -5208
rect 6920 -5272 6936 -5208
rect 8252 -5208 8348 -5172
rect 6840 -5288 6936 -5272
rect 6840 -5352 6856 -5288
rect 6920 -5352 6936 -5288
rect 6840 -5368 6936 -5352
rect 6840 -5432 6856 -5368
rect 6920 -5432 6936 -5368
rect 6840 -5448 6936 -5432
rect 6840 -5512 6856 -5448
rect 6920 -5512 6936 -5448
rect 6840 -5528 6936 -5512
rect 6840 -5592 6856 -5528
rect 6920 -5592 6936 -5528
rect 6840 -5608 6936 -5592
rect 6840 -5672 6856 -5608
rect 6920 -5672 6936 -5608
rect 6840 -5688 6936 -5672
rect 6840 -5752 6856 -5688
rect 6920 -5752 6936 -5688
rect 6840 -5768 6936 -5752
rect 6840 -5832 6856 -5768
rect 6920 -5832 6936 -5768
rect 6840 -5848 6936 -5832
rect 6840 -5912 6856 -5848
rect 6920 -5912 6936 -5848
rect 6840 -5928 6936 -5912
rect 5428 -6028 5524 -5992
rect 6840 -5992 6856 -5928
rect 6920 -5992 6936 -5928
rect 7259 -5248 7981 -5239
rect 7259 -5952 7268 -5248
rect 7972 -5952 7981 -5248
rect 7259 -5961 7981 -5952
rect 8252 -5272 8268 -5208
rect 8332 -5272 8348 -5208
rect 9664 -5208 9760 -5172
rect 8252 -5288 8348 -5272
rect 8252 -5352 8268 -5288
rect 8332 -5352 8348 -5288
rect 8252 -5368 8348 -5352
rect 8252 -5432 8268 -5368
rect 8332 -5432 8348 -5368
rect 8252 -5448 8348 -5432
rect 8252 -5512 8268 -5448
rect 8332 -5512 8348 -5448
rect 8252 -5528 8348 -5512
rect 8252 -5592 8268 -5528
rect 8332 -5592 8348 -5528
rect 8252 -5608 8348 -5592
rect 8252 -5672 8268 -5608
rect 8332 -5672 8348 -5608
rect 8252 -5688 8348 -5672
rect 8252 -5752 8268 -5688
rect 8332 -5752 8348 -5688
rect 8252 -5768 8348 -5752
rect 8252 -5832 8268 -5768
rect 8332 -5832 8348 -5768
rect 8252 -5848 8348 -5832
rect 8252 -5912 8268 -5848
rect 8332 -5912 8348 -5848
rect 8252 -5928 8348 -5912
rect 6840 -6028 6936 -5992
rect 8252 -5992 8268 -5928
rect 8332 -5992 8348 -5928
rect 8671 -5248 9393 -5239
rect 8671 -5952 8680 -5248
rect 9384 -5952 9393 -5248
rect 8671 -5961 9393 -5952
rect 9664 -5272 9680 -5208
rect 9744 -5272 9760 -5208
rect 11076 -5208 11172 -5172
rect 9664 -5288 9760 -5272
rect 9664 -5352 9680 -5288
rect 9744 -5352 9760 -5288
rect 9664 -5368 9760 -5352
rect 9664 -5432 9680 -5368
rect 9744 -5432 9760 -5368
rect 9664 -5448 9760 -5432
rect 9664 -5512 9680 -5448
rect 9744 -5512 9760 -5448
rect 9664 -5528 9760 -5512
rect 9664 -5592 9680 -5528
rect 9744 -5592 9760 -5528
rect 9664 -5608 9760 -5592
rect 9664 -5672 9680 -5608
rect 9744 -5672 9760 -5608
rect 9664 -5688 9760 -5672
rect 9664 -5752 9680 -5688
rect 9744 -5752 9760 -5688
rect 9664 -5768 9760 -5752
rect 9664 -5832 9680 -5768
rect 9744 -5832 9760 -5768
rect 9664 -5848 9760 -5832
rect 9664 -5912 9680 -5848
rect 9744 -5912 9760 -5848
rect 9664 -5928 9760 -5912
rect 8252 -6028 8348 -5992
rect 9664 -5992 9680 -5928
rect 9744 -5992 9760 -5928
rect 10083 -5248 10805 -5239
rect 10083 -5952 10092 -5248
rect 10796 -5952 10805 -5248
rect 10083 -5961 10805 -5952
rect 11076 -5272 11092 -5208
rect 11156 -5272 11172 -5208
rect 12488 -5208 12584 -5172
rect 11076 -5288 11172 -5272
rect 11076 -5352 11092 -5288
rect 11156 -5352 11172 -5288
rect 11076 -5368 11172 -5352
rect 11076 -5432 11092 -5368
rect 11156 -5432 11172 -5368
rect 11076 -5448 11172 -5432
rect 11076 -5512 11092 -5448
rect 11156 -5512 11172 -5448
rect 11076 -5528 11172 -5512
rect 11076 -5592 11092 -5528
rect 11156 -5592 11172 -5528
rect 11076 -5608 11172 -5592
rect 11076 -5672 11092 -5608
rect 11156 -5672 11172 -5608
rect 11076 -5688 11172 -5672
rect 11076 -5752 11092 -5688
rect 11156 -5752 11172 -5688
rect 11076 -5768 11172 -5752
rect 11076 -5832 11092 -5768
rect 11156 -5832 11172 -5768
rect 11076 -5848 11172 -5832
rect 11076 -5912 11092 -5848
rect 11156 -5912 11172 -5848
rect 11076 -5928 11172 -5912
rect 9664 -6028 9760 -5992
rect 11076 -5992 11092 -5928
rect 11156 -5992 11172 -5928
rect 11495 -5248 12217 -5239
rect 11495 -5952 11504 -5248
rect 12208 -5952 12217 -5248
rect 11495 -5961 12217 -5952
rect 12488 -5272 12504 -5208
rect 12568 -5272 12584 -5208
rect 13900 -5208 13996 -5172
rect 12488 -5288 12584 -5272
rect 12488 -5352 12504 -5288
rect 12568 -5352 12584 -5288
rect 12488 -5368 12584 -5352
rect 12488 -5432 12504 -5368
rect 12568 -5432 12584 -5368
rect 12488 -5448 12584 -5432
rect 12488 -5512 12504 -5448
rect 12568 -5512 12584 -5448
rect 12488 -5528 12584 -5512
rect 12488 -5592 12504 -5528
rect 12568 -5592 12584 -5528
rect 12488 -5608 12584 -5592
rect 12488 -5672 12504 -5608
rect 12568 -5672 12584 -5608
rect 12488 -5688 12584 -5672
rect 12488 -5752 12504 -5688
rect 12568 -5752 12584 -5688
rect 12488 -5768 12584 -5752
rect 12488 -5832 12504 -5768
rect 12568 -5832 12584 -5768
rect 12488 -5848 12584 -5832
rect 12488 -5912 12504 -5848
rect 12568 -5912 12584 -5848
rect 12488 -5928 12584 -5912
rect 11076 -6028 11172 -5992
rect 12488 -5992 12504 -5928
rect 12568 -5992 12584 -5928
rect 12907 -5248 13629 -5239
rect 12907 -5952 12916 -5248
rect 13620 -5952 13629 -5248
rect 12907 -5961 13629 -5952
rect 13900 -5272 13916 -5208
rect 13980 -5272 13996 -5208
rect 15312 -5208 15408 -5172
rect 13900 -5288 13996 -5272
rect 13900 -5352 13916 -5288
rect 13980 -5352 13996 -5288
rect 13900 -5368 13996 -5352
rect 13900 -5432 13916 -5368
rect 13980 -5432 13996 -5368
rect 13900 -5448 13996 -5432
rect 13900 -5512 13916 -5448
rect 13980 -5512 13996 -5448
rect 13900 -5528 13996 -5512
rect 13900 -5592 13916 -5528
rect 13980 -5592 13996 -5528
rect 13900 -5608 13996 -5592
rect 13900 -5672 13916 -5608
rect 13980 -5672 13996 -5608
rect 13900 -5688 13996 -5672
rect 13900 -5752 13916 -5688
rect 13980 -5752 13996 -5688
rect 13900 -5768 13996 -5752
rect 13900 -5832 13916 -5768
rect 13980 -5832 13996 -5768
rect 13900 -5848 13996 -5832
rect 13900 -5912 13916 -5848
rect 13980 -5912 13996 -5848
rect 13900 -5928 13996 -5912
rect 12488 -6028 12584 -5992
rect 13900 -5992 13916 -5928
rect 13980 -5992 13996 -5928
rect 14319 -5248 15041 -5239
rect 14319 -5952 14328 -5248
rect 15032 -5952 15041 -5248
rect 14319 -5961 15041 -5952
rect 15312 -5272 15328 -5208
rect 15392 -5272 15408 -5208
rect 16724 -5208 16820 -5172
rect 15312 -5288 15408 -5272
rect 15312 -5352 15328 -5288
rect 15392 -5352 15408 -5288
rect 15312 -5368 15408 -5352
rect 15312 -5432 15328 -5368
rect 15392 -5432 15408 -5368
rect 15312 -5448 15408 -5432
rect 15312 -5512 15328 -5448
rect 15392 -5512 15408 -5448
rect 15312 -5528 15408 -5512
rect 15312 -5592 15328 -5528
rect 15392 -5592 15408 -5528
rect 15312 -5608 15408 -5592
rect 15312 -5672 15328 -5608
rect 15392 -5672 15408 -5608
rect 15312 -5688 15408 -5672
rect 15312 -5752 15328 -5688
rect 15392 -5752 15408 -5688
rect 15312 -5768 15408 -5752
rect 15312 -5832 15328 -5768
rect 15392 -5832 15408 -5768
rect 15312 -5848 15408 -5832
rect 15312 -5912 15328 -5848
rect 15392 -5912 15408 -5848
rect 15312 -5928 15408 -5912
rect 13900 -6028 13996 -5992
rect 15312 -5992 15328 -5928
rect 15392 -5992 15408 -5928
rect 15731 -5248 16453 -5239
rect 15731 -5952 15740 -5248
rect 16444 -5952 16453 -5248
rect 15731 -5961 16453 -5952
rect 16724 -5272 16740 -5208
rect 16804 -5272 16820 -5208
rect 18136 -5208 18232 -5172
rect 16724 -5288 16820 -5272
rect 16724 -5352 16740 -5288
rect 16804 -5352 16820 -5288
rect 16724 -5368 16820 -5352
rect 16724 -5432 16740 -5368
rect 16804 -5432 16820 -5368
rect 16724 -5448 16820 -5432
rect 16724 -5512 16740 -5448
rect 16804 -5512 16820 -5448
rect 16724 -5528 16820 -5512
rect 16724 -5592 16740 -5528
rect 16804 -5592 16820 -5528
rect 16724 -5608 16820 -5592
rect 16724 -5672 16740 -5608
rect 16804 -5672 16820 -5608
rect 16724 -5688 16820 -5672
rect 16724 -5752 16740 -5688
rect 16804 -5752 16820 -5688
rect 16724 -5768 16820 -5752
rect 16724 -5832 16740 -5768
rect 16804 -5832 16820 -5768
rect 16724 -5848 16820 -5832
rect 16724 -5912 16740 -5848
rect 16804 -5912 16820 -5848
rect 16724 -5928 16820 -5912
rect 15312 -6028 15408 -5992
rect 16724 -5992 16740 -5928
rect 16804 -5992 16820 -5928
rect 17143 -5248 17865 -5239
rect 17143 -5952 17152 -5248
rect 17856 -5952 17865 -5248
rect 17143 -5961 17865 -5952
rect 18136 -5272 18152 -5208
rect 18216 -5272 18232 -5208
rect 19548 -5208 19644 -5172
rect 18136 -5288 18232 -5272
rect 18136 -5352 18152 -5288
rect 18216 -5352 18232 -5288
rect 18136 -5368 18232 -5352
rect 18136 -5432 18152 -5368
rect 18216 -5432 18232 -5368
rect 18136 -5448 18232 -5432
rect 18136 -5512 18152 -5448
rect 18216 -5512 18232 -5448
rect 18136 -5528 18232 -5512
rect 18136 -5592 18152 -5528
rect 18216 -5592 18232 -5528
rect 18136 -5608 18232 -5592
rect 18136 -5672 18152 -5608
rect 18216 -5672 18232 -5608
rect 18136 -5688 18232 -5672
rect 18136 -5752 18152 -5688
rect 18216 -5752 18232 -5688
rect 18136 -5768 18232 -5752
rect 18136 -5832 18152 -5768
rect 18216 -5832 18232 -5768
rect 18136 -5848 18232 -5832
rect 18136 -5912 18152 -5848
rect 18216 -5912 18232 -5848
rect 18136 -5928 18232 -5912
rect 16724 -6028 16820 -5992
rect 18136 -5992 18152 -5928
rect 18216 -5992 18232 -5928
rect 18555 -5248 19277 -5239
rect 18555 -5952 18564 -5248
rect 19268 -5952 19277 -5248
rect 18555 -5961 19277 -5952
rect 19548 -5272 19564 -5208
rect 19628 -5272 19644 -5208
rect 20960 -5208 21056 -5172
rect 19548 -5288 19644 -5272
rect 19548 -5352 19564 -5288
rect 19628 -5352 19644 -5288
rect 19548 -5368 19644 -5352
rect 19548 -5432 19564 -5368
rect 19628 -5432 19644 -5368
rect 19548 -5448 19644 -5432
rect 19548 -5512 19564 -5448
rect 19628 -5512 19644 -5448
rect 19548 -5528 19644 -5512
rect 19548 -5592 19564 -5528
rect 19628 -5592 19644 -5528
rect 19548 -5608 19644 -5592
rect 19548 -5672 19564 -5608
rect 19628 -5672 19644 -5608
rect 19548 -5688 19644 -5672
rect 19548 -5752 19564 -5688
rect 19628 -5752 19644 -5688
rect 19548 -5768 19644 -5752
rect 19548 -5832 19564 -5768
rect 19628 -5832 19644 -5768
rect 19548 -5848 19644 -5832
rect 19548 -5912 19564 -5848
rect 19628 -5912 19644 -5848
rect 19548 -5928 19644 -5912
rect 18136 -6028 18232 -5992
rect 19548 -5992 19564 -5928
rect 19628 -5992 19644 -5928
rect 19967 -5248 20689 -5239
rect 19967 -5952 19976 -5248
rect 20680 -5952 20689 -5248
rect 19967 -5961 20689 -5952
rect 20960 -5272 20976 -5208
rect 21040 -5272 21056 -5208
rect 22372 -5208 22468 -5172
rect 20960 -5288 21056 -5272
rect 20960 -5352 20976 -5288
rect 21040 -5352 21056 -5288
rect 20960 -5368 21056 -5352
rect 20960 -5432 20976 -5368
rect 21040 -5432 21056 -5368
rect 20960 -5448 21056 -5432
rect 20960 -5512 20976 -5448
rect 21040 -5512 21056 -5448
rect 20960 -5528 21056 -5512
rect 20960 -5592 20976 -5528
rect 21040 -5592 21056 -5528
rect 20960 -5608 21056 -5592
rect 20960 -5672 20976 -5608
rect 21040 -5672 21056 -5608
rect 20960 -5688 21056 -5672
rect 20960 -5752 20976 -5688
rect 21040 -5752 21056 -5688
rect 20960 -5768 21056 -5752
rect 20960 -5832 20976 -5768
rect 21040 -5832 21056 -5768
rect 20960 -5848 21056 -5832
rect 20960 -5912 20976 -5848
rect 21040 -5912 21056 -5848
rect 20960 -5928 21056 -5912
rect 19548 -6028 19644 -5992
rect 20960 -5992 20976 -5928
rect 21040 -5992 21056 -5928
rect 21379 -5248 22101 -5239
rect 21379 -5952 21388 -5248
rect 22092 -5952 22101 -5248
rect 21379 -5961 22101 -5952
rect 22372 -5272 22388 -5208
rect 22452 -5272 22468 -5208
rect 23784 -5208 23880 -5172
rect 22372 -5288 22468 -5272
rect 22372 -5352 22388 -5288
rect 22452 -5352 22468 -5288
rect 22372 -5368 22468 -5352
rect 22372 -5432 22388 -5368
rect 22452 -5432 22468 -5368
rect 22372 -5448 22468 -5432
rect 22372 -5512 22388 -5448
rect 22452 -5512 22468 -5448
rect 22372 -5528 22468 -5512
rect 22372 -5592 22388 -5528
rect 22452 -5592 22468 -5528
rect 22372 -5608 22468 -5592
rect 22372 -5672 22388 -5608
rect 22452 -5672 22468 -5608
rect 22372 -5688 22468 -5672
rect 22372 -5752 22388 -5688
rect 22452 -5752 22468 -5688
rect 22372 -5768 22468 -5752
rect 22372 -5832 22388 -5768
rect 22452 -5832 22468 -5768
rect 22372 -5848 22468 -5832
rect 22372 -5912 22388 -5848
rect 22452 -5912 22468 -5848
rect 22372 -5928 22468 -5912
rect 20960 -6028 21056 -5992
rect 22372 -5992 22388 -5928
rect 22452 -5992 22468 -5928
rect 22791 -5248 23513 -5239
rect 22791 -5952 22800 -5248
rect 23504 -5952 23513 -5248
rect 22791 -5961 23513 -5952
rect 23784 -5272 23800 -5208
rect 23864 -5272 23880 -5208
rect 23784 -5288 23880 -5272
rect 23784 -5352 23800 -5288
rect 23864 -5352 23880 -5288
rect 23784 -5368 23880 -5352
rect 23784 -5432 23800 -5368
rect 23864 -5432 23880 -5368
rect 23784 -5448 23880 -5432
rect 23784 -5512 23800 -5448
rect 23864 -5512 23880 -5448
rect 23784 -5528 23880 -5512
rect 23784 -5592 23800 -5528
rect 23864 -5592 23880 -5528
rect 23784 -5608 23880 -5592
rect 23784 -5672 23800 -5608
rect 23864 -5672 23880 -5608
rect 23784 -5688 23880 -5672
rect 23784 -5752 23800 -5688
rect 23864 -5752 23880 -5688
rect 23784 -5768 23880 -5752
rect 23784 -5832 23800 -5768
rect 23864 -5832 23880 -5768
rect 23784 -5848 23880 -5832
rect 23784 -5912 23800 -5848
rect 23864 -5912 23880 -5848
rect 23784 -5928 23880 -5912
rect 22372 -6028 22468 -5992
rect 23784 -5992 23800 -5928
rect 23864 -5992 23880 -5928
rect 23784 -6028 23880 -5992
rect -22812 -6328 -22716 -6292
rect -23805 -6368 -23083 -6359
rect -23805 -7072 -23796 -6368
rect -23092 -7072 -23083 -6368
rect -23805 -7081 -23083 -7072
rect -22812 -6392 -22796 -6328
rect -22732 -6392 -22716 -6328
rect -21400 -6328 -21304 -6292
rect -22812 -6408 -22716 -6392
rect -22812 -6472 -22796 -6408
rect -22732 -6472 -22716 -6408
rect -22812 -6488 -22716 -6472
rect -22812 -6552 -22796 -6488
rect -22732 -6552 -22716 -6488
rect -22812 -6568 -22716 -6552
rect -22812 -6632 -22796 -6568
rect -22732 -6632 -22716 -6568
rect -22812 -6648 -22716 -6632
rect -22812 -6712 -22796 -6648
rect -22732 -6712 -22716 -6648
rect -22812 -6728 -22716 -6712
rect -22812 -6792 -22796 -6728
rect -22732 -6792 -22716 -6728
rect -22812 -6808 -22716 -6792
rect -22812 -6872 -22796 -6808
rect -22732 -6872 -22716 -6808
rect -22812 -6888 -22716 -6872
rect -22812 -6952 -22796 -6888
rect -22732 -6952 -22716 -6888
rect -22812 -6968 -22716 -6952
rect -22812 -7032 -22796 -6968
rect -22732 -7032 -22716 -6968
rect -22812 -7048 -22716 -7032
rect -22812 -7112 -22796 -7048
rect -22732 -7112 -22716 -7048
rect -22393 -6368 -21671 -6359
rect -22393 -7072 -22384 -6368
rect -21680 -7072 -21671 -6368
rect -22393 -7081 -21671 -7072
rect -21400 -6392 -21384 -6328
rect -21320 -6392 -21304 -6328
rect -19988 -6328 -19892 -6292
rect -21400 -6408 -21304 -6392
rect -21400 -6472 -21384 -6408
rect -21320 -6472 -21304 -6408
rect -21400 -6488 -21304 -6472
rect -21400 -6552 -21384 -6488
rect -21320 -6552 -21304 -6488
rect -21400 -6568 -21304 -6552
rect -21400 -6632 -21384 -6568
rect -21320 -6632 -21304 -6568
rect -21400 -6648 -21304 -6632
rect -21400 -6712 -21384 -6648
rect -21320 -6712 -21304 -6648
rect -21400 -6728 -21304 -6712
rect -21400 -6792 -21384 -6728
rect -21320 -6792 -21304 -6728
rect -21400 -6808 -21304 -6792
rect -21400 -6872 -21384 -6808
rect -21320 -6872 -21304 -6808
rect -21400 -6888 -21304 -6872
rect -21400 -6952 -21384 -6888
rect -21320 -6952 -21304 -6888
rect -21400 -6968 -21304 -6952
rect -21400 -7032 -21384 -6968
rect -21320 -7032 -21304 -6968
rect -21400 -7048 -21304 -7032
rect -22812 -7148 -22716 -7112
rect -21400 -7112 -21384 -7048
rect -21320 -7112 -21304 -7048
rect -20981 -6368 -20259 -6359
rect -20981 -7072 -20972 -6368
rect -20268 -7072 -20259 -6368
rect -20981 -7081 -20259 -7072
rect -19988 -6392 -19972 -6328
rect -19908 -6392 -19892 -6328
rect -18576 -6328 -18480 -6292
rect -19988 -6408 -19892 -6392
rect -19988 -6472 -19972 -6408
rect -19908 -6472 -19892 -6408
rect -19988 -6488 -19892 -6472
rect -19988 -6552 -19972 -6488
rect -19908 -6552 -19892 -6488
rect -19988 -6568 -19892 -6552
rect -19988 -6632 -19972 -6568
rect -19908 -6632 -19892 -6568
rect -19988 -6648 -19892 -6632
rect -19988 -6712 -19972 -6648
rect -19908 -6712 -19892 -6648
rect -19988 -6728 -19892 -6712
rect -19988 -6792 -19972 -6728
rect -19908 -6792 -19892 -6728
rect -19988 -6808 -19892 -6792
rect -19988 -6872 -19972 -6808
rect -19908 -6872 -19892 -6808
rect -19988 -6888 -19892 -6872
rect -19988 -6952 -19972 -6888
rect -19908 -6952 -19892 -6888
rect -19988 -6968 -19892 -6952
rect -19988 -7032 -19972 -6968
rect -19908 -7032 -19892 -6968
rect -19988 -7048 -19892 -7032
rect -21400 -7148 -21304 -7112
rect -19988 -7112 -19972 -7048
rect -19908 -7112 -19892 -7048
rect -19569 -6368 -18847 -6359
rect -19569 -7072 -19560 -6368
rect -18856 -7072 -18847 -6368
rect -19569 -7081 -18847 -7072
rect -18576 -6392 -18560 -6328
rect -18496 -6392 -18480 -6328
rect -17164 -6328 -17068 -6292
rect -18576 -6408 -18480 -6392
rect -18576 -6472 -18560 -6408
rect -18496 -6472 -18480 -6408
rect -18576 -6488 -18480 -6472
rect -18576 -6552 -18560 -6488
rect -18496 -6552 -18480 -6488
rect -18576 -6568 -18480 -6552
rect -18576 -6632 -18560 -6568
rect -18496 -6632 -18480 -6568
rect -18576 -6648 -18480 -6632
rect -18576 -6712 -18560 -6648
rect -18496 -6712 -18480 -6648
rect -18576 -6728 -18480 -6712
rect -18576 -6792 -18560 -6728
rect -18496 -6792 -18480 -6728
rect -18576 -6808 -18480 -6792
rect -18576 -6872 -18560 -6808
rect -18496 -6872 -18480 -6808
rect -18576 -6888 -18480 -6872
rect -18576 -6952 -18560 -6888
rect -18496 -6952 -18480 -6888
rect -18576 -6968 -18480 -6952
rect -18576 -7032 -18560 -6968
rect -18496 -7032 -18480 -6968
rect -18576 -7048 -18480 -7032
rect -19988 -7148 -19892 -7112
rect -18576 -7112 -18560 -7048
rect -18496 -7112 -18480 -7048
rect -18157 -6368 -17435 -6359
rect -18157 -7072 -18148 -6368
rect -17444 -7072 -17435 -6368
rect -18157 -7081 -17435 -7072
rect -17164 -6392 -17148 -6328
rect -17084 -6392 -17068 -6328
rect -15752 -6328 -15656 -6292
rect -17164 -6408 -17068 -6392
rect -17164 -6472 -17148 -6408
rect -17084 -6472 -17068 -6408
rect -17164 -6488 -17068 -6472
rect -17164 -6552 -17148 -6488
rect -17084 -6552 -17068 -6488
rect -17164 -6568 -17068 -6552
rect -17164 -6632 -17148 -6568
rect -17084 -6632 -17068 -6568
rect -17164 -6648 -17068 -6632
rect -17164 -6712 -17148 -6648
rect -17084 -6712 -17068 -6648
rect -17164 -6728 -17068 -6712
rect -17164 -6792 -17148 -6728
rect -17084 -6792 -17068 -6728
rect -17164 -6808 -17068 -6792
rect -17164 -6872 -17148 -6808
rect -17084 -6872 -17068 -6808
rect -17164 -6888 -17068 -6872
rect -17164 -6952 -17148 -6888
rect -17084 -6952 -17068 -6888
rect -17164 -6968 -17068 -6952
rect -17164 -7032 -17148 -6968
rect -17084 -7032 -17068 -6968
rect -17164 -7048 -17068 -7032
rect -18576 -7148 -18480 -7112
rect -17164 -7112 -17148 -7048
rect -17084 -7112 -17068 -7048
rect -16745 -6368 -16023 -6359
rect -16745 -7072 -16736 -6368
rect -16032 -7072 -16023 -6368
rect -16745 -7081 -16023 -7072
rect -15752 -6392 -15736 -6328
rect -15672 -6392 -15656 -6328
rect -14340 -6328 -14244 -6292
rect -15752 -6408 -15656 -6392
rect -15752 -6472 -15736 -6408
rect -15672 -6472 -15656 -6408
rect -15752 -6488 -15656 -6472
rect -15752 -6552 -15736 -6488
rect -15672 -6552 -15656 -6488
rect -15752 -6568 -15656 -6552
rect -15752 -6632 -15736 -6568
rect -15672 -6632 -15656 -6568
rect -15752 -6648 -15656 -6632
rect -15752 -6712 -15736 -6648
rect -15672 -6712 -15656 -6648
rect -15752 -6728 -15656 -6712
rect -15752 -6792 -15736 -6728
rect -15672 -6792 -15656 -6728
rect -15752 -6808 -15656 -6792
rect -15752 -6872 -15736 -6808
rect -15672 -6872 -15656 -6808
rect -15752 -6888 -15656 -6872
rect -15752 -6952 -15736 -6888
rect -15672 -6952 -15656 -6888
rect -15752 -6968 -15656 -6952
rect -15752 -7032 -15736 -6968
rect -15672 -7032 -15656 -6968
rect -15752 -7048 -15656 -7032
rect -17164 -7148 -17068 -7112
rect -15752 -7112 -15736 -7048
rect -15672 -7112 -15656 -7048
rect -15333 -6368 -14611 -6359
rect -15333 -7072 -15324 -6368
rect -14620 -7072 -14611 -6368
rect -15333 -7081 -14611 -7072
rect -14340 -6392 -14324 -6328
rect -14260 -6392 -14244 -6328
rect -12928 -6328 -12832 -6292
rect -14340 -6408 -14244 -6392
rect -14340 -6472 -14324 -6408
rect -14260 -6472 -14244 -6408
rect -14340 -6488 -14244 -6472
rect -14340 -6552 -14324 -6488
rect -14260 -6552 -14244 -6488
rect -14340 -6568 -14244 -6552
rect -14340 -6632 -14324 -6568
rect -14260 -6632 -14244 -6568
rect -14340 -6648 -14244 -6632
rect -14340 -6712 -14324 -6648
rect -14260 -6712 -14244 -6648
rect -14340 -6728 -14244 -6712
rect -14340 -6792 -14324 -6728
rect -14260 -6792 -14244 -6728
rect -14340 -6808 -14244 -6792
rect -14340 -6872 -14324 -6808
rect -14260 -6872 -14244 -6808
rect -14340 -6888 -14244 -6872
rect -14340 -6952 -14324 -6888
rect -14260 -6952 -14244 -6888
rect -14340 -6968 -14244 -6952
rect -14340 -7032 -14324 -6968
rect -14260 -7032 -14244 -6968
rect -14340 -7048 -14244 -7032
rect -15752 -7148 -15656 -7112
rect -14340 -7112 -14324 -7048
rect -14260 -7112 -14244 -7048
rect -13921 -6368 -13199 -6359
rect -13921 -7072 -13912 -6368
rect -13208 -7072 -13199 -6368
rect -13921 -7081 -13199 -7072
rect -12928 -6392 -12912 -6328
rect -12848 -6392 -12832 -6328
rect -11516 -6328 -11420 -6292
rect -12928 -6408 -12832 -6392
rect -12928 -6472 -12912 -6408
rect -12848 -6472 -12832 -6408
rect -12928 -6488 -12832 -6472
rect -12928 -6552 -12912 -6488
rect -12848 -6552 -12832 -6488
rect -12928 -6568 -12832 -6552
rect -12928 -6632 -12912 -6568
rect -12848 -6632 -12832 -6568
rect -12928 -6648 -12832 -6632
rect -12928 -6712 -12912 -6648
rect -12848 -6712 -12832 -6648
rect -12928 -6728 -12832 -6712
rect -12928 -6792 -12912 -6728
rect -12848 -6792 -12832 -6728
rect -12928 -6808 -12832 -6792
rect -12928 -6872 -12912 -6808
rect -12848 -6872 -12832 -6808
rect -12928 -6888 -12832 -6872
rect -12928 -6952 -12912 -6888
rect -12848 -6952 -12832 -6888
rect -12928 -6968 -12832 -6952
rect -12928 -7032 -12912 -6968
rect -12848 -7032 -12832 -6968
rect -12928 -7048 -12832 -7032
rect -14340 -7148 -14244 -7112
rect -12928 -7112 -12912 -7048
rect -12848 -7112 -12832 -7048
rect -12509 -6368 -11787 -6359
rect -12509 -7072 -12500 -6368
rect -11796 -7072 -11787 -6368
rect -12509 -7081 -11787 -7072
rect -11516 -6392 -11500 -6328
rect -11436 -6392 -11420 -6328
rect -10104 -6328 -10008 -6292
rect -11516 -6408 -11420 -6392
rect -11516 -6472 -11500 -6408
rect -11436 -6472 -11420 -6408
rect -11516 -6488 -11420 -6472
rect -11516 -6552 -11500 -6488
rect -11436 -6552 -11420 -6488
rect -11516 -6568 -11420 -6552
rect -11516 -6632 -11500 -6568
rect -11436 -6632 -11420 -6568
rect -11516 -6648 -11420 -6632
rect -11516 -6712 -11500 -6648
rect -11436 -6712 -11420 -6648
rect -11516 -6728 -11420 -6712
rect -11516 -6792 -11500 -6728
rect -11436 -6792 -11420 -6728
rect -11516 -6808 -11420 -6792
rect -11516 -6872 -11500 -6808
rect -11436 -6872 -11420 -6808
rect -11516 -6888 -11420 -6872
rect -11516 -6952 -11500 -6888
rect -11436 -6952 -11420 -6888
rect -11516 -6968 -11420 -6952
rect -11516 -7032 -11500 -6968
rect -11436 -7032 -11420 -6968
rect -11516 -7048 -11420 -7032
rect -12928 -7148 -12832 -7112
rect -11516 -7112 -11500 -7048
rect -11436 -7112 -11420 -7048
rect -11097 -6368 -10375 -6359
rect -11097 -7072 -11088 -6368
rect -10384 -7072 -10375 -6368
rect -11097 -7081 -10375 -7072
rect -10104 -6392 -10088 -6328
rect -10024 -6392 -10008 -6328
rect -8692 -6328 -8596 -6292
rect -10104 -6408 -10008 -6392
rect -10104 -6472 -10088 -6408
rect -10024 -6472 -10008 -6408
rect -10104 -6488 -10008 -6472
rect -10104 -6552 -10088 -6488
rect -10024 -6552 -10008 -6488
rect -10104 -6568 -10008 -6552
rect -10104 -6632 -10088 -6568
rect -10024 -6632 -10008 -6568
rect -10104 -6648 -10008 -6632
rect -10104 -6712 -10088 -6648
rect -10024 -6712 -10008 -6648
rect -10104 -6728 -10008 -6712
rect -10104 -6792 -10088 -6728
rect -10024 -6792 -10008 -6728
rect -10104 -6808 -10008 -6792
rect -10104 -6872 -10088 -6808
rect -10024 -6872 -10008 -6808
rect -10104 -6888 -10008 -6872
rect -10104 -6952 -10088 -6888
rect -10024 -6952 -10008 -6888
rect -10104 -6968 -10008 -6952
rect -10104 -7032 -10088 -6968
rect -10024 -7032 -10008 -6968
rect -10104 -7048 -10008 -7032
rect -11516 -7148 -11420 -7112
rect -10104 -7112 -10088 -7048
rect -10024 -7112 -10008 -7048
rect -9685 -6368 -8963 -6359
rect -9685 -7072 -9676 -6368
rect -8972 -7072 -8963 -6368
rect -9685 -7081 -8963 -7072
rect -8692 -6392 -8676 -6328
rect -8612 -6392 -8596 -6328
rect -7280 -6328 -7184 -6292
rect -8692 -6408 -8596 -6392
rect -8692 -6472 -8676 -6408
rect -8612 -6472 -8596 -6408
rect -8692 -6488 -8596 -6472
rect -8692 -6552 -8676 -6488
rect -8612 -6552 -8596 -6488
rect -8692 -6568 -8596 -6552
rect -8692 -6632 -8676 -6568
rect -8612 -6632 -8596 -6568
rect -8692 -6648 -8596 -6632
rect -8692 -6712 -8676 -6648
rect -8612 -6712 -8596 -6648
rect -8692 -6728 -8596 -6712
rect -8692 -6792 -8676 -6728
rect -8612 -6792 -8596 -6728
rect -8692 -6808 -8596 -6792
rect -8692 -6872 -8676 -6808
rect -8612 -6872 -8596 -6808
rect -8692 -6888 -8596 -6872
rect -8692 -6952 -8676 -6888
rect -8612 -6952 -8596 -6888
rect -8692 -6968 -8596 -6952
rect -8692 -7032 -8676 -6968
rect -8612 -7032 -8596 -6968
rect -8692 -7048 -8596 -7032
rect -10104 -7148 -10008 -7112
rect -8692 -7112 -8676 -7048
rect -8612 -7112 -8596 -7048
rect -8273 -6368 -7551 -6359
rect -8273 -7072 -8264 -6368
rect -7560 -7072 -7551 -6368
rect -8273 -7081 -7551 -7072
rect -7280 -6392 -7264 -6328
rect -7200 -6392 -7184 -6328
rect -5868 -6328 -5772 -6292
rect -7280 -6408 -7184 -6392
rect -7280 -6472 -7264 -6408
rect -7200 -6472 -7184 -6408
rect -7280 -6488 -7184 -6472
rect -7280 -6552 -7264 -6488
rect -7200 -6552 -7184 -6488
rect -7280 -6568 -7184 -6552
rect -7280 -6632 -7264 -6568
rect -7200 -6632 -7184 -6568
rect -7280 -6648 -7184 -6632
rect -7280 -6712 -7264 -6648
rect -7200 -6712 -7184 -6648
rect -7280 -6728 -7184 -6712
rect -7280 -6792 -7264 -6728
rect -7200 -6792 -7184 -6728
rect -7280 -6808 -7184 -6792
rect -7280 -6872 -7264 -6808
rect -7200 -6872 -7184 -6808
rect -7280 -6888 -7184 -6872
rect -7280 -6952 -7264 -6888
rect -7200 -6952 -7184 -6888
rect -7280 -6968 -7184 -6952
rect -7280 -7032 -7264 -6968
rect -7200 -7032 -7184 -6968
rect -7280 -7048 -7184 -7032
rect -8692 -7148 -8596 -7112
rect -7280 -7112 -7264 -7048
rect -7200 -7112 -7184 -7048
rect -6861 -6368 -6139 -6359
rect -6861 -7072 -6852 -6368
rect -6148 -7072 -6139 -6368
rect -6861 -7081 -6139 -7072
rect -5868 -6392 -5852 -6328
rect -5788 -6392 -5772 -6328
rect -4456 -6328 -4360 -6292
rect -5868 -6408 -5772 -6392
rect -5868 -6472 -5852 -6408
rect -5788 -6472 -5772 -6408
rect -5868 -6488 -5772 -6472
rect -5868 -6552 -5852 -6488
rect -5788 -6552 -5772 -6488
rect -5868 -6568 -5772 -6552
rect -5868 -6632 -5852 -6568
rect -5788 -6632 -5772 -6568
rect -5868 -6648 -5772 -6632
rect -5868 -6712 -5852 -6648
rect -5788 -6712 -5772 -6648
rect -5868 -6728 -5772 -6712
rect -5868 -6792 -5852 -6728
rect -5788 -6792 -5772 -6728
rect -5868 -6808 -5772 -6792
rect -5868 -6872 -5852 -6808
rect -5788 -6872 -5772 -6808
rect -5868 -6888 -5772 -6872
rect -5868 -6952 -5852 -6888
rect -5788 -6952 -5772 -6888
rect -5868 -6968 -5772 -6952
rect -5868 -7032 -5852 -6968
rect -5788 -7032 -5772 -6968
rect -5868 -7048 -5772 -7032
rect -7280 -7148 -7184 -7112
rect -5868 -7112 -5852 -7048
rect -5788 -7112 -5772 -7048
rect -5449 -6368 -4727 -6359
rect -5449 -7072 -5440 -6368
rect -4736 -7072 -4727 -6368
rect -5449 -7081 -4727 -7072
rect -4456 -6392 -4440 -6328
rect -4376 -6392 -4360 -6328
rect -3044 -6328 -2948 -6292
rect -4456 -6408 -4360 -6392
rect -4456 -6472 -4440 -6408
rect -4376 -6472 -4360 -6408
rect -4456 -6488 -4360 -6472
rect -4456 -6552 -4440 -6488
rect -4376 -6552 -4360 -6488
rect -4456 -6568 -4360 -6552
rect -4456 -6632 -4440 -6568
rect -4376 -6632 -4360 -6568
rect -4456 -6648 -4360 -6632
rect -4456 -6712 -4440 -6648
rect -4376 -6712 -4360 -6648
rect -4456 -6728 -4360 -6712
rect -4456 -6792 -4440 -6728
rect -4376 -6792 -4360 -6728
rect -4456 -6808 -4360 -6792
rect -4456 -6872 -4440 -6808
rect -4376 -6872 -4360 -6808
rect -4456 -6888 -4360 -6872
rect -4456 -6952 -4440 -6888
rect -4376 -6952 -4360 -6888
rect -4456 -6968 -4360 -6952
rect -4456 -7032 -4440 -6968
rect -4376 -7032 -4360 -6968
rect -4456 -7048 -4360 -7032
rect -5868 -7148 -5772 -7112
rect -4456 -7112 -4440 -7048
rect -4376 -7112 -4360 -7048
rect -4037 -6368 -3315 -6359
rect -4037 -7072 -4028 -6368
rect -3324 -7072 -3315 -6368
rect -4037 -7081 -3315 -7072
rect -3044 -6392 -3028 -6328
rect -2964 -6392 -2948 -6328
rect -1632 -6328 -1536 -6292
rect -3044 -6408 -2948 -6392
rect -3044 -6472 -3028 -6408
rect -2964 -6472 -2948 -6408
rect -3044 -6488 -2948 -6472
rect -3044 -6552 -3028 -6488
rect -2964 -6552 -2948 -6488
rect -3044 -6568 -2948 -6552
rect -3044 -6632 -3028 -6568
rect -2964 -6632 -2948 -6568
rect -3044 -6648 -2948 -6632
rect -3044 -6712 -3028 -6648
rect -2964 -6712 -2948 -6648
rect -3044 -6728 -2948 -6712
rect -3044 -6792 -3028 -6728
rect -2964 -6792 -2948 -6728
rect -3044 -6808 -2948 -6792
rect -3044 -6872 -3028 -6808
rect -2964 -6872 -2948 -6808
rect -3044 -6888 -2948 -6872
rect -3044 -6952 -3028 -6888
rect -2964 -6952 -2948 -6888
rect -3044 -6968 -2948 -6952
rect -3044 -7032 -3028 -6968
rect -2964 -7032 -2948 -6968
rect -3044 -7048 -2948 -7032
rect -4456 -7148 -4360 -7112
rect -3044 -7112 -3028 -7048
rect -2964 -7112 -2948 -7048
rect -2625 -6368 -1903 -6359
rect -2625 -7072 -2616 -6368
rect -1912 -7072 -1903 -6368
rect -2625 -7081 -1903 -7072
rect -1632 -6392 -1616 -6328
rect -1552 -6392 -1536 -6328
rect -220 -6328 -124 -6292
rect -1632 -6408 -1536 -6392
rect -1632 -6472 -1616 -6408
rect -1552 -6472 -1536 -6408
rect -1632 -6488 -1536 -6472
rect -1632 -6552 -1616 -6488
rect -1552 -6552 -1536 -6488
rect -1632 -6568 -1536 -6552
rect -1632 -6632 -1616 -6568
rect -1552 -6632 -1536 -6568
rect -1632 -6648 -1536 -6632
rect -1632 -6712 -1616 -6648
rect -1552 -6712 -1536 -6648
rect -1632 -6728 -1536 -6712
rect -1632 -6792 -1616 -6728
rect -1552 -6792 -1536 -6728
rect -1632 -6808 -1536 -6792
rect -1632 -6872 -1616 -6808
rect -1552 -6872 -1536 -6808
rect -1632 -6888 -1536 -6872
rect -1632 -6952 -1616 -6888
rect -1552 -6952 -1536 -6888
rect -1632 -6968 -1536 -6952
rect -1632 -7032 -1616 -6968
rect -1552 -7032 -1536 -6968
rect -1632 -7048 -1536 -7032
rect -3044 -7148 -2948 -7112
rect -1632 -7112 -1616 -7048
rect -1552 -7112 -1536 -7048
rect -1213 -6368 -491 -6359
rect -1213 -7072 -1204 -6368
rect -500 -7072 -491 -6368
rect -1213 -7081 -491 -7072
rect -220 -6392 -204 -6328
rect -140 -6392 -124 -6328
rect 1192 -6328 1288 -6292
rect -220 -6408 -124 -6392
rect -220 -6472 -204 -6408
rect -140 -6472 -124 -6408
rect -220 -6488 -124 -6472
rect -220 -6552 -204 -6488
rect -140 -6552 -124 -6488
rect -220 -6568 -124 -6552
rect -220 -6632 -204 -6568
rect -140 -6632 -124 -6568
rect -220 -6648 -124 -6632
rect -220 -6712 -204 -6648
rect -140 -6712 -124 -6648
rect -220 -6728 -124 -6712
rect -220 -6792 -204 -6728
rect -140 -6792 -124 -6728
rect -220 -6808 -124 -6792
rect -220 -6872 -204 -6808
rect -140 -6872 -124 -6808
rect -220 -6888 -124 -6872
rect -220 -6952 -204 -6888
rect -140 -6952 -124 -6888
rect -220 -6968 -124 -6952
rect -220 -7032 -204 -6968
rect -140 -7032 -124 -6968
rect -220 -7048 -124 -7032
rect -1632 -7148 -1536 -7112
rect -220 -7112 -204 -7048
rect -140 -7112 -124 -7048
rect 199 -6368 921 -6359
rect 199 -7072 208 -6368
rect 912 -7072 921 -6368
rect 199 -7081 921 -7072
rect 1192 -6392 1208 -6328
rect 1272 -6392 1288 -6328
rect 2604 -6328 2700 -6292
rect 1192 -6408 1288 -6392
rect 1192 -6472 1208 -6408
rect 1272 -6472 1288 -6408
rect 1192 -6488 1288 -6472
rect 1192 -6552 1208 -6488
rect 1272 -6552 1288 -6488
rect 1192 -6568 1288 -6552
rect 1192 -6632 1208 -6568
rect 1272 -6632 1288 -6568
rect 1192 -6648 1288 -6632
rect 1192 -6712 1208 -6648
rect 1272 -6712 1288 -6648
rect 1192 -6728 1288 -6712
rect 1192 -6792 1208 -6728
rect 1272 -6792 1288 -6728
rect 1192 -6808 1288 -6792
rect 1192 -6872 1208 -6808
rect 1272 -6872 1288 -6808
rect 1192 -6888 1288 -6872
rect 1192 -6952 1208 -6888
rect 1272 -6952 1288 -6888
rect 1192 -6968 1288 -6952
rect 1192 -7032 1208 -6968
rect 1272 -7032 1288 -6968
rect 1192 -7048 1288 -7032
rect -220 -7148 -124 -7112
rect 1192 -7112 1208 -7048
rect 1272 -7112 1288 -7048
rect 1611 -6368 2333 -6359
rect 1611 -7072 1620 -6368
rect 2324 -7072 2333 -6368
rect 1611 -7081 2333 -7072
rect 2604 -6392 2620 -6328
rect 2684 -6392 2700 -6328
rect 4016 -6328 4112 -6292
rect 2604 -6408 2700 -6392
rect 2604 -6472 2620 -6408
rect 2684 -6472 2700 -6408
rect 2604 -6488 2700 -6472
rect 2604 -6552 2620 -6488
rect 2684 -6552 2700 -6488
rect 2604 -6568 2700 -6552
rect 2604 -6632 2620 -6568
rect 2684 -6632 2700 -6568
rect 2604 -6648 2700 -6632
rect 2604 -6712 2620 -6648
rect 2684 -6712 2700 -6648
rect 2604 -6728 2700 -6712
rect 2604 -6792 2620 -6728
rect 2684 -6792 2700 -6728
rect 2604 -6808 2700 -6792
rect 2604 -6872 2620 -6808
rect 2684 -6872 2700 -6808
rect 2604 -6888 2700 -6872
rect 2604 -6952 2620 -6888
rect 2684 -6952 2700 -6888
rect 2604 -6968 2700 -6952
rect 2604 -7032 2620 -6968
rect 2684 -7032 2700 -6968
rect 2604 -7048 2700 -7032
rect 1192 -7148 1288 -7112
rect 2604 -7112 2620 -7048
rect 2684 -7112 2700 -7048
rect 3023 -6368 3745 -6359
rect 3023 -7072 3032 -6368
rect 3736 -7072 3745 -6368
rect 3023 -7081 3745 -7072
rect 4016 -6392 4032 -6328
rect 4096 -6392 4112 -6328
rect 5428 -6328 5524 -6292
rect 4016 -6408 4112 -6392
rect 4016 -6472 4032 -6408
rect 4096 -6472 4112 -6408
rect 4016 -6488 4112 -6472
rect 4016 -6552 4032 -6488
rect 4096 -6552 4112 -6488
rect 4016 -6568 4112 -6552
rect 4016 -6632 4032 -6568
rect 4096 -6632 4112 -6568
rect 4016 -6648 4112 -6632
rect 4016 -6712 4032 -6648
rect 4096 -6712 4112 -6648
rect 4016 -6728 4112 -6712
rect 4016 -6792 4032 -6728
rect 4096 -6792 4112 -6728
rect 4016 -6808 4112 -6792
rect 4016 -6872 4032 -6808
rect 4096 -6872 4112 -6808
rect 4016 -6888 4112 -6872
rect 4016 -6952 4032 -6888
rect 4096 -6952 4112 -6888
rect 4016 -6968 4112 -6952
rect 4016 -7032 4032 -6968
rect 4096 -7032 4112 -6968
rect 4016 -7048 4112 -7032
rect 2604 -7148 2700 -7112
rect 4016 -7112 4032 -7048
rect 4096 -7112 4112 -7048
rect 4435 -6368 5157 -6359
rect 4435 -7072 4444 -6368
rect 5148 -7072 5157 -6368
rect 4435 -7081 5157 -7072
rect 5428 -6392 5444 -6328
rect 5508 -6392 5524 -6328
rect 6840 -6328 6936 -6292
rect 5428 -6408 5524 -6392
rect 5428 -6472 5444 -6408
rect 5508 -6472 5524 -6408
rect 5428 -6488 5524 -6472
rect 5428 -6552 5444 -6488
rect 5508 -6552 5524 -6488
rect 5428 -6568 5524 -6552
rect 5428 -6632 5444 -6568
rect 5508 -6632 5524 -6568
rect 5428 -6648 5524 -6632
rect 5428 -6712 5444 -6648
rect 5508 -6712 5524 -6648
rect 5428 -6728 5524 -6712
rect 5428 -6792 5444 -6728
rect 5508 -6792 5524 -6728
rect 5428 -6808 5524 -6792
rect 5428 -6872 5444 -6808
rect 5508 -6872 5524 -6808
rect 5428 -6888 5524 -6872
rect 5428 -6952 5444 -6888
rect 5508 -6952 5524 -6888
rect 5428 -6968 5524 -6952
rect 5428 -7032 5444 -6968
rect 5508 -7032 5524 -6968
rect 5428 -7048 5524 -7032
rect 4016 -7148 4112 -7112
rect 5428 -7112 5444 -7048
rect 5508 -7112 5524 -7048
rect 5847 -6368 6569 -6359
rect 5847 -7072 5856 -6368
rect 6560 -7072 6569 -6368
rect 5847 -7081 6569 -7072
rect 6840 -6392 6856 -6328
rect 6920 -6392 6936 -6328
rect 8252 -6328 8348 -6292
rect 6840 -6408 6936 -6392
rect 6840 -6472 6856 -6408
rect 6920 -6472 6936 -6408
rect 6840 -6488 6936 -6472
rect 6840 -6552 6856 -6488
rect 6920 -6552 6936 -6488
rect 6840 -6568 6936 -6552
rect 6840 -6632 6856 -6568
rect 6920 -6632 6936 -6568
rect 6840 -6648 6936 -6632
rect 6840 -6712 6856 -6648
rect 6920 -6712 6936 -6648
rect 6840 -6728 6936 -6712
rect 6840 -6792 6856 -6728
rect 6920 -6792 6936 -6728
rect 6840 -6808 6936 -6792
rect 6840 -6872 6856 -6808
rect 6920 -6872 6936 -6808
rect 6840 -6888 6936 -6872
rect 6840 -6952 6856 -6888
rect 6920 -6952 6936 -6888
rect 6840 -6968 6936 -6952
rect 6840 -7032 6856 -6968
rect 6920 -7032 6936 -6968
rect 6840 -7048 6936 -7032
rect 5428 -7148 5524 -7112
rect 6840 -7112 6856 -7048
rect 6920 -7112 6936 -7048
rect 7259 -6368 7981 -6359
rect 7259 -7072 7268 -6368
rect 7972 -7072 7981 -6368
rect 7259 -7081 7981 -7072
rect 8252 -6392 8268 -6328
rect 8332 -6392 8348 -6328
rect 9664 -6328 9760 -6292
rect 8252 -6408 8348 -6392
rect 8252 -6472 8268 -6408
rect 8332 -6472 8348 -6408
rect 8252 -6488 8348 -6472
rect 8252 -6552 8268 -6488
rect 8332 -6552 8348 -6488
rect 8252 -6568 8348 -6552
rect 8252 -6632 8268 -6568
rect 8332 -6632 8348 -6568
rect 8252 -6648 8348 -6632
rect 8252 -6712 8268 -6648
rect 8332 -6712 8348 -6648
rect 8252 -6728 8348 -6712
rect 8252 -6792 8268 -6728
rect 8332 -6792 8348 -6728
rect 8252 -6808 8348 -6792
rect 8252 -6872 8268 -6808
rect 8332 -6872 8348 -6808
rect 8252 -6888 8348 -6872
rect 8252 -6952 8268 -6888
rect 8332 -6952 8348 -6888
rect 8252 -6968 8348 -6952
rect 8252 -7032 8268 -6968
rect 8332 -7032 8348 -6968
rect 8252 -7048 8348 -7032
rect 6840 -7148 6936 -7112
rect 8252 -7112 8268 -7048
rect 8332 -7112 8348 -7048
rect 8671 -6368 9393 -6359
rect 8671 -7072 8680 -6368
rect 9384 -7072 9393 -6368
rect 8671 -7081 9393 -7072
rect 9664 -6392 9680 -6328
rect 9744 -6392 9760 -6328
rect 11076 -6328 11172 -6292
rect 9664 -6408 9760 -6392
rect 9664 -6472 9680 -6408
rect 9744 -6472 9760 -6408
rect 9664 -6488 9760 -6472
rect 9664 -6552 9680 -6488
rect 9744 -6552 9760 -6488
rect 9664 -6568 9760 -6552
rect 9664 -6632 9680 -6568
rect 9744 -6632 9760 -6568
rect 9664 -6648 9760 -6632
rect 9664 -6712 9680 -6648
rect 9744 -6712 9760 -6648
rect 9664 -6728 9760 -6712
rect 9664 -6792 9680 -6728
rect 9744 -6792 9760 -6728
rect 9664 -6808 9760 -6792
rect 9664 -6872 9680 -6808
rect 9744 -6872 9760 -6808
rect 9664 -6888 9760 -6872
rect 9664 -6952 9680 -6888
rect 9744 -6952 9760 -6888
rect 9664 -6968 9760 -6952
rect 9664 -7032 9680 -6968
rect 9744 -7032 9760 -6968
rect 9664 -7048 9760 -7032
rect 8252 -7148 8348 -7112
rect 9664 -7112 9680 -7048
rect 9744 -7112 9760 -7048
rect 10083 -6368 10805 -6359
rect 10083 -7072 10092 -6368
rect 10796 -7072 10805 -6368
rect 10083 -7081 10805 -7072
rect 11076 -6392 11092 -6328
rect 11156 -6392 11172 -6328
rect 12488 -6328 12584 -6292
rect 11076 -6408 11172 -6392
rect 11076 -6472 11092 -6408
rect 11156 -6472 11172 -6408
rect 11076 -6488 11172 -6472
rect 11076 -6552 11092 -6488
rect 11156 -6552 11172 -6488
rect 11076 -6568 11172 -6552
rect 11076 -6632 11092 -6568
rect 11156 -6632 11172 -6568
rect 11076 -6648 11172 -6632
rect 11076 -6712 11092 -6648
rect 11156 -6712 11172 -6648
rect 11076 -6728 11172 -6712
rect 11076 -6792 11092 -6728
rect 11156 -6792 11172 -6728
rect 11076 -6808 11172 -6792
rect 11076 -6872 11092 -6808
rect 11156 -6872 11172 -6808
rect 11076 -6888 11172 -6872
rect 11076 -6952 11092 -6888
rect 11156 -6952 11172 -6888
rect 11076 -6968 11172 -6952
rect 11076 -7032 11092 -6968
rect 11156 -7032 11172 -6968
rect 11076 -7048 11172 -7032
rect 9664 -7148 9760 -7112
rect 11076 -7112 11092 -7048
rect 11156 -7112 11172 -7048
rect 11495 -6368 12217 -6359
rect 11495 -7072 11504 -6368
rect 12208 -7072 12217 -6368
rect 11495 -7081 12217 -7072
rect 12488 -6392 12504 -6328
rect 12568 -6392 12584 -6328
rect 13900 -6328 13996 -6292
rect 12488 -6408 12584 -6392
rect 12488 -6472 12504 -6408
rect 12568 -6472 12584 -6408
rect 12488 -6488 12584 -6472
rect 12488 -6552 12504 -6488
rect 12568 -6552 12584 -6488
rect 12488 -6568 12584 -6552
rect 12488 -6632 12504 -6568
rect 12568 -6632 12584 -6568
rect 12488 -6648 12584 -6632
rect 12488 -6712 12504 -6648
rect 12568 -6712 12584 -6648
rect 12488 -6728 12584 -6712
rect 12488 -6792 12504 -6728
rect 12568 -6792 12584 -6728
rect 12488 -6808 12584 -6792
rect 12488 -6872 12504 -6808
rect 12568 -6872 12584 -6808
rect 12488 -6888 12584 -6872
rect 12488 -6952 12504 -6888
rect 12568 -6952 12584 -6888
rect 12488 -6968 12584 -6952
rect 12488 -7032 12504 -6968
rect 12568 -7032 12584 -6968
rect 12488 -7048 12584 -7032
rect 11076 -7148 11172 -7112
rect 12488 -7112 12504 -7048
rect 12568 -7112 12584 -7048
rect 12907 -6368 13629 -6359
rect 12907 -7072 12916 -6368
rect 13620 -7072 13629 -6368
rect 12907 -7081 13629 -7072
rect 13900 -6392 13916 -6328
rect 13980 -6392 13996 -6328
rect 15312 -6328 15408 -6292
rect 13900 -6408 13996 -6392
rect 13900 -6472 13916 -6408
rect 13980 -6472 13996 -6408
rect 13900 -6488 13996 -6472
rect 13900 -6552 13916 -6488
rect 13980 -6552 13996 -6488
rect 13900 -6568 13996 -6552
rect 13900 -6632 13916 -6568
rect 13980 -6632 13996 -6568
rect 13900 -6648 13996 -6632
rect 13900 -6712 13916 -6648
rect 13980 -6712 13996 -6648
rect 13900 -6728 13996 -6712
rect 13900 -6792 13916 -6728
rect 13980 -6792 13996 -6728
rect 13900 -6808 13996 -6792
rect 13900 -6872 13916 -6808
rect 13980 -6872 13996 -6808
rect 13900 -6888 13996 -6872
rect 13900 -6952 13916 -6888
rect 13980 -6952 13996 -6888
rect 13900 -6968 13996 -6952
rect 13900 -7032 13916 -6968
rect 13980 -7032 13996 -6968
rect 13900 -7048 13996 -7032
rect 12488 -7148 12584 -7112
rect 13900 -7112 13916 -7048
rect 13980 -7112 13996 -7048
rect 14319 -6368 15041 -6359
rect 14319 -7072 14328 -6368
rect 15032 -7072 15041 -6368
rect 14319 -7081 15041 -7072
rect 15312 -6392 15328 -6328
rect 15392 -6392 15408 -6328
rect 16724 -6328 16820 -6292
rect 15312 -6408 15408 -6392
rect 15312 -6472 15328 -6408
rect 15392 -6472 15408 -6408
rect 15312 -6488 15408 -6472
rect 15312 -6552 15328 -6488
rect 15392 -6552 15408 -6488
rect 15312 -6568 15408 -6552
rect 15312 -6632 15328 -6568
rect 15392 -6632 15408 -6568
rect 15312 -6648 15408 -6632
rect 15312 -6712 15328 -6648
rect 15392 -6712 15408 -6648
rect 15312 -6728 15408 -6712
rect 15312 -6792 15328 -6728
rect 15392 -6792 15408 -6728
rect 15312 -6808 15408 -6792
rect 15312 -6872 15328 -6808
rect 15392 -6872 15408 -6808
rect 15312 -6888 15408 -6872
rect 15312 -6952 15328 -6888
rect 15392 -6952 15408 -6888
rect 15312 -6968 15408 -6952
rect 15312 -7032 15328 -6968
rect 15392 -7032 15408 -6968
rect 15312 -7048 15408 -7032
rect 13900 -7148 13996 -7112
rect 15312 -7112 15328 -7048
rect 15392 -7112 15408 -7048
rect 15731 -6368 16453 -6359
rect 15731 -7072 15740 -6368
rect 16444 -7072 16453 -6368
rect 15731 -7081 16453 -7072
rect 16724 -6392 16740 -6328
rect 16804 -6392 16820 -6328
rect 18136 -6328 18232 -6292
rect 16724 -6408 16820 -6392
rect 16724 -6472 16740 -6408
rect 16804 -6472 16820 -6408
rect 16724 -6488 16820 -6472
rect 16724 -6552 16740 -6488
rect 16804 -6552 16820 -6488
rect 16724 -6568 16820 -6552
rect 16724 -6632 16740 -6568
rect 16804 -6632 16820 -6568
rect 16724 -6648 16820 -6632
rect 16724 -6712 16740 -6648
rect 16804 -6712 16820 -6648
rect 16724 -6728 16820 -6712
rect 16724 -6792 16740 -6728
rect 16804 -6792 16820 -6728
rect 16724 -6808 16820 -6792
rect 16724 -6872 16740 -6808
rect 16804 -6872 16820 -6808
rect 16724 -6888 16820 -6872
rect 16724 -6952 16740 -6888
rect 16804 -6952 16820 -6888
rect 16724 -6968 16820 -6952
rect 16724 -7032 16740 -6968
rect 16804 -7032 16820 -6968
rect 16724 -7048 16820 -7032
rect 15312 -7148 15408 -7112
rect 16724 -7112 16740 -7048
rect 16804 -7112 16820 -7048
rect 17143 -6368 17865 -6359
rect 17143 -7072 17152 -6368
rect 17856 -7072 17865 -6368
rect 17143 -7081 17865 -7072
rect 18136 -6392 18152 -6328
rect 18216 -6392 18232 -6328
rect 19548 -6328 19644 -6292
rect 18136 -6408 18232 -6392
rect 18136 -6472 18152 -6408
rect 18216 -6472 18232 -6408
rect 18136 -6488 18232 -6472
rect 18136 -6552 18152 -6488
rect 18216 -6552 18232 -6488
rect 18136 -6568 18232 -6552
rect 18136 -6632 18152 -6568
rect 18216 -6632 18232 -6568
rect 18136 -6648 18232 -6632
rect 18136 -6712 18152 -6648
rect 18216 -6712 18232 -6648
rect 18136 -6728 18232 -6712
rect 18136 -6792 18152 -6728
rect 18216 -6792 18232 -6728
rect 18136 -6808 18232 -6792
rect 18136 -6872 18152 -6808
rect 18216 -6872 18232 -6808
rect 18136 -6888 18232 -6872
rect 18136 -6952 18152 -6888
rect 18216 -6952 18232 -6888
rect 18136 -6968 18232 -6952
rect 18136 -7032 18152 -6968
rect 18216 -7032 18232 -6968
rect 18136 -7048 18232 -7032
rect 16724 -7148 16820 -7112
rect 18136 -7112 18152 -7048
rect 18216 -7112 18232 -7048
rect 18555 -6368 19277 -6359
rect 18555 -7072 18564 -6368
rect 19268 -7072 19277 -6368
rect 18555 -7081 19277 -7072
rect 19548 -6392 19564 -6328
rect 19628 -6392 19644 -6328
rect 20960 -6328 21056 -6292
rect 19548 -6408 19644 -6392
rect 19548 -6472 19564 -6408
rect 19628 -6472 19644 -6408
rect 19548 -6488 19644 -6472
rect 19548 -6552 19564 -6488
rect 19628 -6552 19644 -6488
rect 19548 -6568 19644 -6552
rect 19548 -6632 19564 -6568
rect 19628 -6632 19644 -6568
rect 19548 -6648 19644 -6632
rect 19548 -6712 19564 -6648
rect 19628 -6712 19644 -6648
rect 19548 -6728 19644 -6712
rect 19548 -6792 19564 -6728
rect 19628 -6792 19644 -6728
rect 19548 -6808 19644 -6792
rect 19548 -6872 19564 -6808
rect 19628 -6872 19644 -6808
rect 19548 -6888 19644 -6872
rect 19548 -6952 19564 -6888
rect 19628 -6952 19644 -6888
rect 19548 -6968 19644 -6952
rect 19548 -7032 19564 -6968
rect 19628 -7032 19644 -6968
rect 19548 -7048 19644 -7032
rect 18136 -7148 18232 -7112
rect 19548 -7112 19564 -7048
rect 19628 -7112 19644 -7048
rect 19967 -6368 20689 -6359
rect 19967 -7072 19976 -6368
rect 20680 -7072 20689 -6368
rect 19967 -7081 20689 -7072
rect 20960 -6392 20976 -6328
rect 21040 -6392 21056 -6328
rect 22372 -6328 22468 -6292
rect 20960 -6408 21056 -6392
rect 20960 -6472 20976 -6408
rect 21040 -6472 21056 -6408
rect 20960 -6488 21056 -6472
rect 20960 -6552 20976 -6488
rect 21040 -6552 21056 -6488
rect 20960 -6568 21056 -6552
rect 20960 -6632 20976 -6568
rect 21040 -6632 21056 -6568
rect 20960 -6648 21056 -6632
rect 20960 -6712 20976 -6648
rect 21040 -6712 21056 -6648
rect 20960 -6728 21056 -6712
rect 20960 -6792 20976 -6728
rect 21040 -6792 21056 -6728
rect 20960 -6808 21056 -6792
rect 20960 -6872 20976 -6808
rect 21040 -6872 21056 -6808
rect 20960 -6888 21056 -6872
rect 20960 -6952 20976 -6888
rect 21040 -6952 21056 -6888
rect 20960 -6968 21056 -6952
rect 20960 -7032 20976 -6968
rect 21040 -7032 21056 -6968
rect 20960 -7048 21056 -7032
rect 19548 -7148 19644 -7112
rect 20960 -7112 20976 -7048
rect 21040 -7112 21056 -7048
rect 21379 -6368 22101 -6359
rect 21379 -7072 21388 -6368
rect 22092 -7072 22101 -6368
rect 21379 -7081 22101 -7072
rect 22372 -6392 22388 -6328
rect 22452 -6392 22468 -6328
rect 23784 -6328 23880 -6292
rect 22372 -6408 22468 -6392
rect 22372 -6472 22388 -6408
rect 22452 -6472 22468 -6408
rect 22372 -6488 22468 -6472
rect 22372 -6552 22388 -6488
rect 22452 -6552 22468 -6488
rect 22372 -6568 22468 -6552
rect 22372 -6632 22388 -6568
rect 22452 -6632 22468 -6568
rect 22372 -6648 22468 -6632
rect 22372 -6712 22388 -6648
rect 22452 -6712 22468 -6648
rect 22372 -6728 22468 -6712
rect 22372 -6792 22388 -6728
rect 22452 -6792 22468 -6728
rect 22372 -6808 22468 -6792
rect 22372 -6872 22388 -6808
rect 22452 -6872 22468 -6808
rect 22372 -6888 22468 -6872
rect 22372 -6952 22388 -6888
rect 22452 -6952 22468 -6888
rect 22372 -6968 22468 -6952
rect 22372 -7032 22388 -6968
rect 22452 -7032 22468 -6968
rect 22372 -7048 22468 -7032
rect 20960 -7148 21056 -7112
rect 22372 -7112 22388 -7048
rect 22452 -7112 22468 -7048
rect 22791 -6368 23513 -6359
rect 22791 -7072 22800 -6368
rect 23504 -7072 23513 -6368
rect 22791 -7081 23513 -7072
rect 23784 -6392 23800 -6328
rect 23864 -6392 23880 -6328
rect 23784 -6408 23880 -6392
rect 23784 -6472 23800 -6408
rect 23864 -6472 23880 -6408
rect 23784 -6488 23880 -6472
rect 23784 -6552 23800 -6488
rect 23864 -6552 23880 -6488
rect 23784 -6568 23880 -6552
rect 23784 -6632 23800 -6568
rect 23864 -6632 23880 -6568
rect 23784 -6648 23880 -6632
rect 23784 -6712 23800 -6648
rect 23864 -6712 23880 -6648
rect 23784 -6728 23880 -6712
rect 23784 -6792 23800 -6728
rect 23864 -6792 23880 -6728
rect 23784 -6808 23880 -6792
rect 23784 -6872 23800 -6808
rect 23864 -6872 23880 -6808
rect 23784 -6888 23880 -6872
rect 23784 -6952 23800 -6888
rect 23864 -6952 23880 -6888
rect 23784 -6968 23880 -6952
rect 23784 -7032 23800 -6968
rect 23864 -7032 23880 -6968
rect 23784 -7048 23880 -7032
rect 22372 -7148 22468 -7112
rect 23784 -7112 23800 -7048
rect 23864 -7112 23880 -7048
rect 23784 -7148 23880 -7112
rect -22812 -7448 -22716 -7412
rect -23805 -7488 -23083 -7479
rect -23805 -8192 -23796 -7488
rect -23092 -8192 -23083 -7488
rect -23805 -8201 -23083 -8192
rect -22812 -7512 -22796 -7448
rect -22732 -7512 -22716 -7448
rect -21400 -7448 -21304 -7412
rect -22812 -7528 -22716 -7512
rect -22812 -7592 -22796 -7528
rect -22732 -7592 -22716 -7528
rect -22812 -7608 -22716 -7592
rect -22812 -7672 -22796 -7608
rect -22732 -7672 -22716 -7608
rect -22812 -7688 -22716 -7672
rect -22812 -7752 -22796 -7688
rect -22732 -7752 -22716 -7688
rect -22812 -7768 -22716 -7752
rect -22812 -7832 -22796 -7768
rect -22732 -7832 -22716 -7768
rect -22812 -7848 -22716 -7832
rect -22812 -7912 -22796 -7848
rect -22732 -7912 -22716 -7848
rect -22812 -7928 -22716 -7912
rect -22812 -7992 -22796 -7928
rect -22732 -7992 -22716 -7928
rect -22812 -8008 -22716 -7992
rect -22812 -8072 -22796 -8008
rect -22732 -8072 -22716 -8008
rect -22812 -8088 -22716 -8072
rect -22812 -8152 -22796 -8088
rect -22732 -8152 -22716 -8088
rect -22812 -8168 -22716 -8152
rect -22812 -8232 -22796 -8168
rect -22732 -8232 -22716 -8168
rect -22393 -7488 -21671 -7479
rect -22393 -8192 -22384 -7488
rect -21680 -8192 -21671 -7488
rect -22393 -8201 -21671 -8192
rect -21400 -7512 -21384 -7448
rect -21320 -7512 -21304 -7448
rect -19988 -7448 -19892 -7412
rect -21400 -7528 -21304 -7512
rect -21400 -7592 -21384 -7528
rect -21320 -7592 -21304 -7528
rect -21400 -7608 -21304 -7592
rect -21400 -7672 -21384 -7608
rect -21320 -7672 -21304 -7608
rect -21400 -7688 -21304 -7672
rect -21400 -7752 -21384 -7688
rect -21320 -7752 -21304 -7688
rect -21400 -7768 -21304 -7752
rect -21400 -7832 -21384 -7768
rect -21320 -7832 -21304 -7768
rect -21400 -7848 -21304 -7832
rect -21400 -7912 -21384 -7848
rect -21320 -7912 -21304 -7848
rect -21400 -7928 -21304 -7912
rect -21400 -7992 -21384 -7928
rect -21320 -7992 -21304 -7928
rect -21400 -8008 -21304 -7992
rect -21400 -8072 -21384 -8008
rect -21320 -8072 -21304 -8008
rect -21400 -8088 -21304 -8072
rect -21400 -8152 -21384 -8088
rect -21320 -8152 -21304 -8088
rect -21400 -8168 -21304 -8152
rect -22812 -8268 -22716 -8232
rect -21400 -8232 -21384 -8168
rect -21320 -8232 -21304 -8168
rect -20981 -7488 -20259 -7479
rect -20981 -8192 -20972 -7488
rect -20268 -8192 -20259 -7488
rect -20981 -8201 -20259 -8192
rect -19988 -7512 -19972 -7448
rect -19908 -7512 -19892 -7448
rect -18576 -7448 -18480 -7412
rect -19988 -7528 -19892 -7512
rect -19988 -7592 -19972 -7528
rect -19908 -7592 -19892 -7528
rect -19988 -7608 -19892 -7592
rect -19988 -7672 -19972 -7608
rect -19908 -7672 -19892 -7608
rect -19988 -7688 -19892 -7672
rect -19988 -7752 -19972 -7688
rect -19908 -7752 -19892 -7688
rect -19988 -7768 -19892 -7752
rect -19988 -7832 -19972 -7768
rect -19908 -7832 -19892 -7768
rect -19988 -7848 -19892 -7832
rect -19988 -7912 -19972 -7848
rect -19908 -7912 -19892 -7848
rect -19988 -7928 -19892 -7912
rect -19988 -7992 -19972 -7928
rect -19908 -7992 -19892 -7928
rect -19988 -8008 -19892 -7992
rect -19988 -8072 -19972 -8008
rect -19908 -8072 -19892 -8008
rect -19988 -8088 -19892 -8072
rect -19988 -8152 -19972 -8088
rect -19908 -8152 -19892 -8088
rect -19988 -8168 -19892 -8152
rect -21400 -8268 -21304 -8232
rect -19988 -8232 -19972 -8168
rect -19908 -8232 -19892 -8168
rect -19569 -7488 -18847 -7479
rect -19569 -8192 -19560 -7488
rect -18856 -8192 -18847 -7488
rect -19569 -8201 -18847 -8192
rect -18576 -7512 -18560 -7448
rect -18496 -7512 -18480 -7448
rect -17164 -7448 -17068 -7412
rect -18576 -7528 -18480 -7512
rect -18576 -7592 -18560 -7528
rect -18496 -7592 -18480 -7528
rect -18576 -7608 -18480 -7592
rect -18576 -7672 -18560 -7608
rect -18496 -7672 -18480 -7608
rect -18576 -7688 -18480 -7672
rect -18576 -7752 -18560 -7688
rect -18496 -7752 -18480 -7688
rect -18576 -7768 -18480 -7752
rect -18576 -7832 -18560 -7768
rect -18496 -7832 -18480 -7768
rect -18576 -7848 -18480 -7832
rect -18576 -7912 -18560 -7848
rect -18496 -7912 -18480 -7848
rect -18576 -7928 -18480 -7912
rect -18576 -7992 -18560 -7928
rect -18496 -7992 -18480 -7928
rect -18576 -8008 -18480 -7992
rect -18576 -8072 -18560 -8008
rect -18496 -8072 -18480 -8008
rect -18576 -8088 -18480 -8072
rect -18576 -8152 -18560 -8088
rect -18496 -8152 -18480 -8088
rect -18576 -8168 -18480 -8152
rect -19988 -8268 -19892 -8232
rect -18576 -8232 -18560 -8168
rect -18496 -8232 -18480 -8168
rect -18157 -7488 -17435 -7479
rect -18157 -8192 -18148 -7488
rect -17444 -8192 -17435 -7488
rect -18157 -8201 -17435 -8192
rect -17164 -7512 -17148 -7448
rect -17084 -7512 -17068 -7448
rect -15752 -7448 -15656 -7412
rect -17164 -7528 -17068 -7512
rect -17164 -7592 -17148 -7528
rect -17084 -7592 -17068 -7528
rect -17164 -7608 -17068 -7592
rect -17164 -7672 -17148 -7608
rect -17084 -7672 -17068 -7608
rect -17164 -7688 -17068 -7672
rect -17164 -7752 -17148 -7688
rect -17084 -7752 -17068 -7688
rect -17164 -7768 -17068 -7752
rect -17164 -7832 -17148 -7768
rect -17084 -7832 -17068 -7768
rect -17164 -7848 -17068 -7832
rect -17164 -7912 -17148 -7848
rect -17084 -7912 -17068 -7848
rect -17164 -7928 -17068 -7912
rect -17164 -7992 -17148 -7928
rect -17084 -7992 -17068 -7928
rect -17164 -8008 -17068 -7992
rect -17164 -8072 -17148 -8008
rect -17084 -8072 -17068 -8008
rect -17164 -8088 -17068 -8072
rect -17164 -8152 -17148 -8088
rect -17084 -8152 -17068 -8088
rect -17164 -8168 -17068 -8152
rect -18576 -8268 -18480 -8232
rect -17164 -8232 -17148 -8168
rect -17084 -8232 -17068 -8168
rect -16745 -7488 -16023 -7479
rect -16745 -8192 -16736 -7488
rect -16032 -8192 -16023 -7488
rect -16745 -8201 -16023 -8192
rect -15752 -7512 -15736 -7448
rect -15672 -7512 -15656 -7448
rect -14340 -7448 -14244 -7412
rect -15752 -7528 -15656 -7512
rect -15752 -7592 -15736 -7528
rect -15672 -7592 -15656 -7528
rect -15752 -7608 -15656 -7592
rect -15752 -7672 -15736 -7608
rect -15672 -7672 -15656 -7608
rect -15752 -7688 -15656 -7672
rect -15752 -7752 -15736 -7688
rect -15672 -7752 -15656 -7688
rect -15752 -7768 -15656 -7752
rect -15752 -7832 -15736 -7768
rect -15672 -7832 -15656 -7768
rect -15752 -7848 -15656 -7832
rect -15752 -7912 -15736 -7848
rect -15672 -7912 -15656 -7848
rect -15752 -7928 -15656 -7912
rect -15752 -7992 -15736 -7928
rect -15672 -7992 -15656 -7928
rect -15752 -8008 -15656 -7992
rect -15752 -8072 -15736 -8008
rect -15672 -8072 -15656 -8008
rect -15752 -8088 -15656 -8072
rect -15752 -8152 -15736 -8088
rect -15672 -8152 -15656 -8088
rect -15752 -8168 -15656 -8152
rect -17164 -8268 -17068 -8232
rect -15752 -8232 -15736 -8168
rect -15672 -8232 -15656 -8168
rect -15333 -7488 -14611 -7479
rect -15333 -8192 -15324 -7488
rect -14620 -8192 -14611 -7488
rect -15333 -8201 -14611 -8192
rect -14340 -7512 -14324 -7448
rect -14260 -7512 -14244 -7448
rect -12928 -7448 -12832 -7412
rect -14340 -7528 -14244 -7512
rect -14340 -7592 -14324 -7528
rect -14260 -7592 -14244 -7528
rect -14340 -7608 -14244 -7592
rect -14340 -7672 -14324 -7608
rect -14260 -7672 -14244 -7608
rect -14340 -7688 -14244 -7672
rect -14340 -7752 -14324 -7688
rect -14260 -7752 -14244 -7688
rect -14340 -7768 -14244 -7752
rect -14340 -7832 -14324 -7768
rect -14260 -7832 -14244 -7768
rect -14340 -7848 -14244 -7832
rect -14340 -7912 -14324 -7848
rect -14260 -7912 -14244 -7848
rect -14340 -7928 -14244 -7912
rect -14340 -7992 -14324 -7928
rect -14260 -7992 -14244 -7928
rect -14340 -8008 -14244 -7992
rect -14340 -8072 -14324 -8008
rect -14260 -8072 -14244 -8008
rect -14340 -8088 -14244 -8072
rect -14340 -8152 -14324 -8088
rect -14260 -8152 -14244 -8088
rect -14340 -8168 -14244 -8152
rect -15752 -8268 -15656 -8232
rect -14340 -8232 -14324 -8168
rect -14260 -8232 -14244 -8168
rect -13921 -7488 -13199 -7479
rect -13921 -8192 -13912 -7488
rect -13208 -8192 -13199 -7488
rect -13921 -8201 -13199 -8192
rect -12928 -7512 -12912 -7448
rect -12848 -7512 -12832 -7448
rect -11516 -7448 -11420 -7412
rect -12928 -7528 -12832 -7512
rect -12928 -7592 -12912 -7528
rect -12848 -7592 -12832 -7528
rect -12928 -7608 -12832 -7592
rect -12928 -7672 -12912 -7608
rect -12848 -7672 -12832 -7608
rect -12928 -7688 -12832 -7672
rect -12928 -7752 -12912 -7688
rect -12848 -7752 -12832 -7688
rect -12928 -7768 -12832 -7752
rect -12928 -7832 -12912 -7768
rect -12848 -7832 -12832 -7768
rect -12928 -7848 -12832 -7832
rect -12928 -7912 -12912 -7848
rect -12848 -7912 -12832 -7848
rect -12928 -7928 -12832 -7912
rect -12928 -7992 -12912 -7928
rect -12848 -7992 -12832 -7928
rect -12928 -8008 -12832 -7992
rect -12928 -8072 -12912 -8008
rect -12848 -8072 -12832 -8008
rect -12928 -8088 -12832 -8072
rect -12928 -8152 -12912 -8088
rect -12848 -8152 -12832 -8088
rect -12928 -8168 -12832 -8152
rect -14340 -8268 -14244 -8232
rect -12928 -8232 -12912 -8168
rect -12848 -8232 -12832 -8168
rect -12509 -7488 -11787 -7479
rect -12509 -8192 -12500 -7488
rect -11796 -8192 -11787 -7488
rect -12509 -8201 -11787 -8192
rect -11516 -7512 -11500 -7448
rect -11436 -7512 -11420 -7448
rect -10104 -7448 -10008 -7412
rect -11516 -7528 -11420 -7512
rect -11516 -7592 -11500 -7528
rect -11436 -7592 -11420 -7528
rect -11516 -7608 -11420 -7592
rect -11516 -7672 -11500 -7608
rect -11436 -7672 -11420 -7608
rect -11516 -7688 -11420 -7672
rect -11516 -7752 -11500 -7688
rect -11436 -7752 -11420 -7688
rect -11516 -7768 -11420 -7752
rect -11516 -7832 -11500 -7768
rect -11436 -7832 -11420 -7768
rect -11516 -7848 -11420 -7832
rect -11516 -7912 -11500 -7848
rect -11436 -7912 -11420 -7848
rect -11516 -7928 -11420 -7912
rect -11516 -7992 -11500 -7928
rect -11436 -7992 -11420 -7928
rect -11516 -8008 -11420 -7992
rect -11516 -8072 -11500 -8008
rect -11436 -8072 -11420 -8008
rect -11516 -8088 -11420 -8072
rect -11516 -8152 -11500 -8088
rect -11436 -8152 -11420 -8088
rect -11516 -8168 -11420 -8152
rect -12928 -8268 -12832 -8232
rect -11516 -8232 -11500 -8168
rect -11436 -8232 -11420 -8168
rect -11097 -7488 -10375 -7479
rect -11097 -8192 -11088 -7488
rect -10384 -8192 -10375 -7488
rect -11097 -8201 -10375 -8192
rect -10104 -7512 -10088 -7448
rect -10024 -7512 -10008 -7448
rect -8692 -7448 -8596 -7412
rect -10104 -7528 -10008 -7512
rect -10104 -7592 -10088 -7528
rect -10024 -7592 -10008 -7528
rect -10104 -7608 -10008 -7592
rect -10104 -7672 -10088 -7608
rect -10024 -7672 -10008 -7608
rect -10104 -7688 -10008 -7672
rect -10104 -7752 -10088 -7688
rect -10024 -7752 -10008 -7688
rect -10104 -7768 -10008 -7752
rect -10104 -7832 -10088 -7768
rect -10024 -7832 -10008 -7768
rect -10104 -7848 -10008 -7832
rect -10104 -7912 -10088 -7848
rect -10024 -7912 -10008 -7848
rect -10104 -7928 -10008 -7912
rect -10104 -7992 -10088 -7928
rect -10024 -7992 -10008 -7928
rect -10104 -8008 -10008 -7992
rect -10104 -8072 -10088 -8008
rect -10024 -8072 -10008 -8008
rect -10104 -8088 -10008 -8072
rect -10104 -8152 -10088 -8088
rect -10024 -8152 -10008 -8088
rect -10104 -8168 -10008 -8152
rect -11516 -8268 -11420 -8232
rect -10104 -8232 -10088 -8168
rect -10024 -8232 -10008 -8168
rect -9685 -7488 -8963 -7479
rect -9685 -8192 -9676 -7488
rect -8972 -8192 -8963 -7488
rect -9685 -8201 -8963 -8192
rect -8692 -7512 -8676 -7448
rect -8612 -7512 -8596 -7448
rect -7280 -7448 -7184 -7412
rect -8692 -7528 -8596 -7512
rect -8692 -7592 -8676 -7528
rect -8612 -7592 -8596 -7528
rect -8692 -7608 -8596 -7592
rect -8692 -7672 -8676 -7608
rect -8612 -7672 -8596 -7608
rect -8692 -7688 -8596 -7672
rect -8692 -7752 -8676 -7688
rect -8612 -7752 -8596 -7688
rect -8692 -7768 -8596 -7752
rect -8692 -7832 -8676 -7768
rect -8612 -7832 -8596 -7768
rect -8692 -7848 -8596 -7832
rect -8692 -7912 -8676 -7848
rect -8612 -7912 -8596 -7848
rect -8692 -7928 -8596 -7912
rect -8692 -7992 -8676 -7928
rect -8612 -7992 -8596 -7928
rect -8692 -8008 -8596 -7992
rect -8692 -8072 -8676 -8008
rect -8612 -8072 -8596 -8008
rect -8692 -8088 -8596 -8072
rect -8692 -8152 -8676 -8088
rect -8612 -8152 -8596 -8088
rect -8692 -8168 -8596 -8152
rect -10104 -8268 -10008 -8232
rect -8692 -8232 -8676 -8168
rect -8612 -8232 -8596 -8168
rect -8273 -7488 -7551 -7479
rect -8273 -8192 -8264 -7488
rect -7560 -8192 -7551 -7488
rect -8273 -8201 -7551 -8192
rect -7280 -7512 -7264 -7448
rect -7200 -7512 -7184 -7448
rect -5868 -7448 -5772 -7412
rect -7280 -7528 -7184 -7512
rect -7280 -7592 -7264 -7528
rect -7200 -7592 -7184 -7528
rect -7280 -7608 -7184 -7592
rect -7280 -7672 -7264 -7608
rect -7200 -7672 -7184 -7608
rect -7280 -7688 -7184 -7672
rect -7280 -7752 -7264 -7688
rect -7200 -7752 -7184 -7688
rect -7280 -7768 -7184 -7752
rect -7280 -7832 -7264 -7768
rect -7200 -7832 -7184 -7768
rect -7280 -7848 -7184 -7832
rect -7280 -7912 -7264 -7848
rect -7200 -7912 -7184 -7848
rect -7280 -7928 -7184 -7912
rect -7280 -7992 -7264 -7928
rect -7200 -7992 -7184 -7928
rect -7280 -8008 -7184 -7992
rect -7280 -8072 -7264 -8008
rect -7200 -8072 -7184 -8008
rect -7280 -8088 -7184 -8072
rect -7280 -8152 -7264 -8088
rect -7200 -8152 -7184 -8088
rect -7280 -8168 -7184 -8152
rect -8692 -8268 -8596 -8232
rect -7280 -8232 -7264 -8168
rect -7200 -8232 -7184 -8168
rect -6861 -7488 -6139 -7479
rect -6861 -8192 -6852 -7488
rect -6148 -8192 -6139 -7488
rect -6861 -8201 -6139 -8192
rect -5868 -7512 -5852 -7448
rect -5788 -7512 -5772 -7448
rect -4456 -7448 -4360 -7412
rect -5868 -7528 -5772 -7512
rect -5868 -7592 -5852 -7528
rect -5788 -7592 -5772 -7528
rect -5868 -7608 -5772 -7592
rect -5868 -7672 -5852 -7608
rect -5788 -7672 -5772 -7608
rect -5868 -7688 -5772 -7672
rect -5868 -7752 -5852 -7688
rect -5788 -7752 -5772 -7688
rect -5868 -7768 -5772 -7752
rect -5868 -7832 -5852 -7768
rect -5788 -7832 -5772 -7768
rect -5868 -7848 -5772 -7832
rect -5868 -7912 -5852 -7848
rect -5788 -7912 -5772 -7848
rect -5868 -7928 -5772 -7912
rect -5868 -7992 -5852 -7928
rect -5788 -7992 -5772 -7928
rect -5868 -8008 -5772 -7992
rect -5868 -8072 -5852 -8008
rect -5788 -8072 -5772 -8008
rect -5868 -8088 -5772 -8072
rect -5868 -8152 -5852 -8088
rect -5788 -8152 -5772 -8088
rect -5868 -8168 -5772 -8152
rect -7280 -8268 -7184 -8232
rect -5868 -8232 -5852 -8168
rect -5788 -8232 -5772 -8168
rect -5449 -7488 -4727 -7479
rect -5449 -8192 -5440 -7488
rect -4736 -8192 -4727 -7488
rect -5449 -8201 -4727 -8192
rect -4456 -7512 -4440 -7448
rect -4376 -7512 -4360 -7448
rect -3044 -7448 -2948 -7412
rect -4456 -7528 -4360 -7512
rect -4456 -7592 -4440 -7528
rect -4376 -7592 -4360 -7528
rect -4456 -7608 -4360 -7592
rect -4456 -7672 -4440 -7608
rect -4376 -7672 -4360 -7608
rect -4456 -7688 -4360 -7672
rect -4456 -7752 -4440 -7688
rect -4376 -7752 -4360 -7688
rect -4456 -7768 -4360 -7752
rect -4456 -7832 -4440 -7768
rect -4376 -7832 -4360 -7768
rect -4456 -7848 -4360 -7832
rect -4456 -7912 -4440 -7848
rect -4376 -7912 -4360 -7848
rect -4456 -7928 -4360 -7912
rect -4456 -7992 -4440 -7928
rect -4376 -7992 -4360 -7928
rect -4456 -8008 -4360 -7992
rect -4456 -8072 -4440 -8008
rect -4376 -8072 -4360 -8008
rect -4456 -8088 -4360 -8072
rect -4456 -8152 -4440 -8088
rect -4376 -8152 -4360 -8088
rect -4456 -8168 -4360 -8152
rect -5868 -8268 -5772 -8232
rect -4456 -8232 -4440 -8168
rect -4376 -8232 -4360 -8168
rect -4037 -7488 -3315 -7479
rect -4037 -8192 -4028 -7488
rect -3324 -8192 -3315 -7488
rect -4037 -8201 -3315 -8192
rect -3044 -7512 -3028 -7448
rect -2964 -7512 -2948 -7448
rect -1632 -7448 -1536 -7412
rect -3044 -7528 -2948 -7512
rect -3044 -7592 -3028 -7528
rect -2964 -7592 -2948 -7528
rect -3044 -7608 -2948 -7592
rect -3044 -7672 -3028 -7608
rect -2964 -7672 -2948 -7608
rect -3044 -7688 -2948 -7672
rect -3044 -7752 -3028 -7688
rect -2964 -7752 -2948 -7688
rect -3044 -7768 -2948 -7752
rect -3044 -7832 -3028 -7768
rect -2964 -7832 -2948 -7768
rect -3044 -7848 -2948 -7832
rect -3044 -7912 -3028 -7848
rect -2964 -7912 -2948 -7848
rect -3044 -7928 -2948 -7912
rect -3044 -7992 -3028 -7928
rect -2964 -7992 -2948 -7928
rect -3044 -8008 -2948 -7992
rect -3044 -8072 -3028 -8008
rect -2964 -8072 -2948 -8008
rect -3044 -8088 -2948 -8072
rect -3044 -8152 -3028 -8088
rect -2964 -8152 -2948 -8088
rect -3044 -8168 -2948 -8152
rect -4456 -8268 -4360 -8232
rect -3044 -8232 -3028 -8168
rect -2964 -8232 -2948 -8168
rect -2625 -7488 -1903 -7479
rect -2625 -8192 -2616 -7488
rect -1912 -8192 -1903 -7488
rect -2625 -8201 -1903 -8192
rect -1632 -7512 -1616 -7448
rect -1552 -7512 -1536 -7448
rect -220 -7448 -124 -7412
rect -1632 -7528 -1536 -7512
rect -1632 -7592 -1616 -7528
rect -1552 -7592 -1536 -7528
rect -1632 -7608 -1536 -7592
rect -1632 -7672 -1616 -7608
rect -1552 -7672 -1536 -7608
rect -1632 -7688 -1536 -7672
rect -1632 -7752 -1616 -7688
rect -1552 -7752 -1536 -7688
rect -1632 -7768 -1536 -7752
rect -1632 -7832 -1616 -7768
rect -1552 -7832 -1536 -7768
rect -1632 -7848 -1536 -7832
rect -1632 -7912 -1616 -7848
rect -1552 -7912 -1536 -7848
rect -1632 -7928 -1536 -7912
rect -1632 -7992 -1616 -7928
rect -1552 -7992 -1536 -7928
rect -1632 -8008 -1536 -7992
rect -1632 -8072 -1616 -8008
rect -1552 -8072 -1536 -8008
rect -1632 -8088 -1536 -8072
rect -1632 -8152 -1616 -8088
rect -1552 -8152 -1536 -8088
rect -1632 -8168 -1536 -8152
rect -3044 -8268 -2948 -8232
rect -1632 -8232 -1616 -8168
rect -1552 -8232 -1536 -8168
rect -1213 -7488 -491 -7479
rect -1213 -8192 -1204 -7488
rect -500 -8192 -491 -7488
rect -1213 -8201 -491 -8192
rect -220 -7512 -204 -7448
rect -140 -7512 -124 -7448
rect 1192 -7448 1288 -7412
rect -220 -7528 -124 -7512
rect -220 -7592 -204 -7528
rect -140 -7592 -124 -7528
rect -220 -7608 -124 -7592
rect -220 -7672 -204 -7608
rect -140 -7672 -124 -7608
rect -220 -7688 -124 -7672
rect -220 -7752 -204 -7688
rect -140 -7752 -124 -7688
rect -220 -7768 -124 -7752
rect -220 -7832 -204 -7768
rect -140 -7832 -124 -7768
rect -220 -7848 -124 -7832
rect -220 -7912 -204 -7848
rect -140 -7912 -124 -7848
rect -220 -7928 -124 -7912
rect -220 -7992 -204 -7928
rect -140 -7992 -124 -7928
rect -220 -8008 -124 -7992
rect -220 -8072 -204 -8008
rect -140 -8072 -124 -8008
rect -220 -8088 -124 -8072
rect -220 -8152 -204 -8088
rect -140 -8152 -124 -8088
rect -220 -8168 -124 -8152
rect -1632 -8268 -1536 -8232
rect -220 -8232 -204 -8168
rect -140 -8232 -124 -8168
rect 199 -7488 921 -7479
rect 199 -8192 208 -7488
rect 912 -8192 921 -7488
rect 199 -8201 921 -8192
rect 1192 -7512 1208 -7448
rect 1272 -7512 1288 -7448
rect 2604 -7448 2700 -7412
rect 1192 -7528 1288 -7512
rect 1192 -7592 1208 -7528
rect 1272 -7592 1288 -7528
rect 1192 -7608 1288 -7592
rect 1192 -7672 1208 -7608
rect 1272 -7672 1288 -7608
rect 1192 -7688 1288 -7672
rect 1192 -7752 1208 -7688
rect 1272 -7752 1288 -7688
rect 1192 -7768 1288 -7752
rect 1192 -7832 1208 -7768
rect 1272 -7832 1288 -7768
rect 1192 -7848 1288 -7832
rect 1192 -7912 1208 -7848
rect 1272 -7912 1288 -7848
rect 1192 -7928 1288 -7912
rect 1192 -7992 1208 -7928
rect 1272 -7992 1288 -7928
rect 1192 -8008 1288 -7992
rect 1192 -8072 1208 -8008
rect 1272 -8072 1288 -8008
rect 1192 -8088 1288 -8072
rect 1192 -8152 1208 -8088
rect 1272 -8152 1288 -8088
rect 1192 -8168 1288 -8152
rect -220 -8268 -124 -8232
rect 1192 -8232 1208 -8168
rect 1272 -8232 1288 -8168
rect 1611 -7488 2333 -7479
rect 1611 -8192 1620 -7488
rect 2324 -8192 2333 -7488
rect 1611 -8201 2333 -8192
rect 2604 -7512 2620 -7448
rect 2684 -7512 2700 -7448
rect 4016 -7448 4112 -7412
rect 2604 -7528 2700 -7512
rect 2604 -7592 2620 -7528
rect 2684 -7592 2700 -7528
rect 2604 -7608 2700 -7592
rect 2604 -7672 2620 -7608
rect 2684 -7672 2700 -7608
rect 2604 -7688 2700 -7672
rect 2604 -7752 2620 -7688
rect 2684 -7752 2700 -7688
rect 2604 -7768 2700 -7752
rect 2604 -7832 2620 -7768
rect 2684 -7832 2700 -7768
rect 2604 -7848 2700 -7832
rect 2604 -7912 2620 -7848
rect 2684 -7912 2700 -7848
rect 2604 -7928 2700 -7912
rect 2604 -7992 2620 -7928
rect 2684 -7992 2700 -7928
rect 2604 -8008 2700 -7992
rect 2604 -8072 2620 -8008
rect 2684 -8072 2700 -8008
rect 2604 -8088 2700 -8072
rect 2604 -8152 2620 -8088
rect 2684 -8152 2700 -8088
rect 2604 -8168 2700 -8152
rect 1192 -8268 1288 -8232
rect 2604 -8232 2620 -8168
rect 2684 -8232 2700 -8168
rect 3023 -7488 3745 -7479
rect 3023 -8192 3032 -7488
rect 3736 -8192 3745 -7488
rect 3023 -8201 3745 -8192
rect 4016 -7512 4032 -7448
rect 4096 -7512 4112 -7448
rect 5428 -7448 5524 -7412
rect 4016 -7528 4112 -7512
rect 4016 -7592 4032 -7528
rect 4096 -7592 4112 -7528
rect 4016 -7608 4112 -7592
rect 4016 -7672 4032 -7608
rect 4096 -7672 4112 -7608
rect 4016 -7688 4112 -7672
rect 4016 -7752 4032 -7688
rect 4096 -7752 4112 -7688
rect 4016 -7768 4112 -7752
rect 4016 -7832 4032 -7768
rect 4096 -7832 4112 -7768
rect 4016 -7848 4112 -7832
rect 4016 -7912 4032 -7848
rect 4096 -7912 4112 -7848
rect 4016 -7928 4112 -7912
rect 4016 -7992 4032 -7928
rect 4096 -7992 4112 -7928
rect 4016 -8008 4112 -7992
rect 4016 -8072 4032 -8008
rect 4096 -8072 4112 -8008
rect 4016 -8088 4112 -8072
rect 4016 -8152 4032 -8088
rect 4096 -8152 4112 -8088
rect 4016 -8168 4112 -8152
rect 2604 -8268 2700 -8232
rect 4016 -8232 4032 -8168
rect 4096 -8232 4112 -8168
rect 4435 -7488 5157 -7479
rect 4435 -8192 4444 -7488
rect 5148 -8192 5157 -7488
rect 4435 -8201 5157 -8192
rect 5428 -7512 5444 -7448
rect 5508 -7512 5524 -7448
rect 6840 -7448 6936 -7412
rect 5428 -7528 5524 -7512
rect 5428 -7592 5444 -7528
rect 5508 -7592 5524 -7528
rect 5428 -7608 5524 -7592
rect 5428 -7672 5444 -7608
rect 5508 -7672 5524 -7608
rect 5428 -7688 5524 -7672
rect 5428 -7752 5444 -7688
rect 5508 -7752 5524 -7688
rect 5428 -7768 5524 -7752
rect 5428 -7832 5444 -7768
rect 5508 -7832 5524 -7768
rect 5428 -7848 5524 -7832
rect 5428 -7912 5444 -7848
rect 5508 -7912 5524 -7848
rect 5428 -7928 5524 -7912
rect 5428 -7992 5444 -7928
rect 5508 -7992 5524 -7928
rect 5428 -8008 5524 -7992
rect 5428 -8072 5444 -8008
rect 5508 -8072 5524 -8008
rect 5428 -8088 5524 -8072
rect 5428 -8152 5444 -8088
rect 5508 -8152 5524 -8088
rect 5428 -8168 5524 -8152
rect 4016 -8268 4112 -8232
rect 5428 -8232 5444 -8168
rect 5508 -8232 5524 -8168
rect 5847 -7488 6569 -7479
rect 5847 -8192 5856 -7488
rect 6560 -8192 6569 -7488
rect 5847 -8201 6569 -8192
rect 6840 -7512 6856 -7448
rect 6920 -7512 6936 -7448
rect 8252 -7448 8348 -7412
rect 6840 -7528 6936 -7512
rect 6840 -7592 6856 -7528
rect 6920 -7592 6936 -7528
rect 6840 -7608 6936 -7592
rect 6840 -7672 6856 -7608
rect 6920 -7672 6936 -7608
rect 6840 -7688 6936 -7672
rect 6840 -7752 6856 -7688
rect 6920 -7752 6936 -7688
rect 6840 -7768 6936 -7752
rect 6840 -7832 6856 -7768
rect 6920 -7832 6936 -7768
rect 6840 -7848 6936 -7832
rect 6840 -7912 6856 -7848
rect 6920 -7912 6936 -7848
rect 6840 -7928 6936 -7912
rect 6840 -7992 6856 -7928
rect 6920 -7992 6936 -7928
rect 6840 -8008 6936 -7992
rect 6840 -8072 6856 -8008
rect 6920 -8072 6936 -8008
rect 6840 -8088 6936 -8072
rect 6840 -8152 6856 -8088
rect 6920 -8152 6936 -8088
rect 6840 -8168 6936 -8152
rect 5428 -8268 5524 -8232
rect 6840 -8232 6856 -8168
rect 6920 -8232 6936 -8168
rect 7259 -7488 7981 -7479
rect 7259 -8192 7268 -7488
rect 7972 -8192 7981 -7488
rect 7259 -8201 7981 -8192
rect 8252 -7512 8268 -7448
rect 8332 -7512 8348 -7448
rect 9664 -7448 9760 -7412
rect 8252 -7528 8348 -7512
rect 8252 -7592 8268 -7528
rect 8332 -7592 8348 -7528
rect 8252 -7608 8348 -7592
rect 8252 -7672 8268 -7608
rect 8332 -7672 8348 -7608
rect 8252 -7688 8348 -7672
rect 8252 -7752 8268 -7688
rect 8332 -7752 8348 -7688
rect 8252 -7768 8348 -7752
rect 8252 -7832 8268 -7768
rect 8332 -7832 8348 -7768
rect 8252 -7848 8348 -7832
rect 8252 -7912 8268 -7848
rect 8332 -7912 8348 -7848
rect 8252 -7928 8348 -7912
rect 8252 -7992 8268 -7928
rect 8332 -7992 8348 -7928
rect 8252 -8008 8348 -7992
rect 8252 -8072 8268 -8008
rect 8332 -8072 8348 -8008
rect 8252 -8088 8348 -8072
rect 8252 -8152 8268 -8088
rect 8332 -8152 8348 -8088
rect 8252 -8168 8348 -8152
rect 6840 -8268 6936 -8232
rect 8252 -8232 8268 -8168
rect 8332 -8232 8348 -8168
rect 8671 -7488 9393 -7479
rect 8671 -8192 8680 -7488
rect 9384 -8192 9393 -7488
rect 8671 -8201 9393 -8192
rect 9664 -7512 9680 -7448
rect 9744 -7512 9760 -7448
rect 11076 -7448 11172 -7412
rect 9664 -7528 9760 -7512
rect 9664 -7592 9680 -7528
rect 9744 -7592 9760 -7528
rect 9664 -7608 9760 -7592
rect 9664 -7672 9680 -7608
rect 9744 -7672 9760 -7608
rect 9664 -7688 9760 -7672
rect 9664 -7752 9680 -7688
rect 9744 -7752 9760 -7688
rect 9664 -7768 9760 -7752
rect 9664 -7832 9680 -7768
rect 9744 -7832 9760 -7768
rect 9664 -7848 9760 -7832
rect 9664 -7912 9680 -7848
rect 9744 -7912 9760 -7848
rect 9664 -7928 9760 -7912
rect 9664 -7992 9680 -7928
rect 9744 -7992 9760 -7928
rect 9664 -8008 9760 -7992
rect 9664 -8072 9680 -8008
rect 9744 -8072 9760 -8008
rect 9664 -8088 9760 -8072
rect 9664 -8152 9680 -8088
rect 9744 -8152 9760 -8088
rect 9664 -8168 9760 -8152
rect 8252 -8268 8348 -8232
rect 9664 -8232 9680 -8168
rect 9744 -8232 9760 -8168
rect 10083 -7488 10805 -7479
rect 10083 -8192 10092 -7488
rect 10796 -8192 10805 -7488
rect 10083 -8201 10805 -8192
rect 11076 -7512 11092 -7448
rect 11156 -7512 11172 -7448
rect 12488 -7448 12584 -7412
rect 11076 -7528 11172 -7512
rect 11076 -7592 11092 -7528
rect 11156 -7592 11172 -7528
rect 11076 -7608 11172 -7592
rect 11076 -7672 11092 -7608
rect 11156 -7672 11172 -7608
rect 11076 -7688 11172 -7672
rect 11076 -7752 11092 -7688
rect 11156 -7752 11172 -7688
rect 11076 -7768 11172 -7752
rect 11076 -7832 11092 -7768
rect 11156 -7832 11172 -7768
rect 11076 -7848 11172 -7832
rect 11076 -7912 11092 -7848
rect 11156 -7912 11172 -7848
rect 11076 -7928 11172 -7912
rect 11076 -7992 11092 -7928
rect 11156 -7992 11172 -7928
rect 11076 -8008 11172 -7992
rect 11076 -8072 11092 -8008
rect 11156 -8072 11172 -8008
rect 11076 -8088 11172 -8072
rect 11076 -8152 11092 -8088
rect 11156 -8152 11172 -8088
rect 11076 -8168 11172 -8152
rect 9664 -8268 9760 -8232
rect 11076 -8232 11092 -8168
rect 11156 -8232 11172 -8168
rect 11495 -7488 12217 -7479
rect 11495 -8192 11504 -7488
rect 12208 -8192 12217 -7488
rect 11495 -8201 12217 -8192
rect 12488 -7512 12504 -7448
rect 12568 -7512 12584 -7448
rect 13900 -7448 13996 -7412
rect 12488 -7528 12584 -7512
rect 12488 -7592 12504 -7528
rect 12568 -7592 12584 -7528
rect 12488 -7608 12584 -7592
rect 12488 -7672 12504 -7608
rect 12568 -7672 12584 -7608
rect 12488 -7688 12584 -7672
rect 12488 -7752 12504 -7688
rect 12568 -7752 12584 -7688
rect 12488 -7768 12584 -7752
rect 12488 -7832 12504 -7768
rect 12568 -7832 12584 -7768
rect 12488 -7848 12584 -7832
rect 12488 -7912 12504 -7848
rect 12568 -7912 12584 -7848
rect 12488 -7928 12584 -7912
rect 12488 -7992 12504 -7928
rect 12568 -7992 12584 -7928
rect 12488 -8008 12584 -7992
rect 12488 -8072 12504 -8008
rect 12568 -8072 12584 -8008
rect 12488 -8088 12584 -8072
rect 12488 -8152 12504 -8088
rect 12568 -8152 12584 -8088
rect 12488 -8168 12584 -8152
rect 11076 -8268 11172 -8232
rect 12488 -8232 12504 -8168
rect 12568 -8232 12584 -8168
rect 12907 -7488 13629 -7479
rect 12907 -8192 12916 -7488
rect 13620 -8192 13629 -7488
rect 12907 -8201 13629 -8192
rect 13900 -7512 13916 -7448
rect 13980 -7512 13996 -7448
rect 15312 -7448 15408 -7412
rect 13900 -7528 13996 -7512
rect 13900 -7592 13916 -7528
rect 13980 -7592 13996 -7528
rect 13900 -7608 13996 -7592
rect 13900 -7672 13916 -7608
rect 13980 -7672 13996 -7608
rect 13900 -7688 13996 -7672
rect 13900 -7752 13916 -7688
rect 13980 -7752 13996 -7688
rect 13900 -7768 13996 -7752
rect 13900 -7832 13916 -7768
rect 13980 -7832 13996 -7768
rect 13900 -7848 13996 -7832
rect 13900 -7912 13916 -7848
rect 13980 -7912 13996 -7848
rect 13900 -7928 13996 -7912
rect 13900 -7992 13916 -7928
rect 13980 -7992 13996 -7928
rect 13900 -8008 13996 -7992
rect 13900 -8072 13916 -8008
rect 13980 -8072 13996 -8008
rect 13900 -8088 13996 -8072
rect 13900 -8152 13916 -8088
rect 13980 -8152 13996 -8088
rect 13900 -8168 13996 -8152
rect 12488 -8268 12584 -8232
rect 13900 -8232 13916 -8168
rect 13980 -8232 13996 -8168
rect 14319 -7488 15041 -7479
rect 14319 -8192 14328 -7488
rect 15032 -8192 15041 -7488
rect 14319 -8201 15041 -8192
rect 15312 -7512 15328 -7448
rect 15392 -7512 15408 -7448
rect 16724 -7448 16820 -7412
rect 15312 -7528 15408 -7512
rect 15312 -7592 15328 -7528
rect 15392 -7592 15408 -7528
rect 15312 -7608 15408 -7592
rect 15312 -7672 15328 -7608
rect 15392 -7672 15408 -7608
rect 15312 -7688 15408 -7672
rect 15312 -7752 15328 -7688
rect 15392 -7752 15408 -7688
rect 15312 -7768 15408 -7752
rect 15312 -7832 15328 -7768
rect 15392 -7832 15408 -7768
rect 15312 -7848 15408 -7832
rect 15312 -7912 15328 -7848
rect 15392 -7912 15408 -7848
rect 15312 -7928 15408 -7912
rect 15312 -7992 15328 -7928
rect 15392 -7992 15408 -7928
rect 15312 -8008 15408 -7992
rect 15312 -8072 15328 -8008
rect 15392 -8072 15408 -8008
rect 15312 -8088 15408 -8072
rect 15312 -8152 15328 -8088
rect 15392 -8152 15408 -8088
rect 15312 -8168 15408 -8152
rect 13900 -8268 13996 -8232
rect 15312 -8232 15328 -8168
rect 15392 -8232 15408 -8168
rect 15731 -7488 16453 -7479
rect 15731 -8192 15740 -7488
rect 16444 -8192 16453 -7488
rect 15731 -8201 16453 -8192
rect 16724 -7512 16740 -7448
rect 16804 -7512 16820 -7448
rect 18136 -7448 18232 -7412
rect 16724 -7528 16820 -7512
rect 16724 -7592 16740 -7528
rect 16804 -7592 16820 -7528
rect 16724 -7608 16820 -7592
rect 16724 -7672 16740 -7608
rect 16804 -7672 16820 -7608
rect 16724 -7688 16820 -7672
rect 16724 -7752 16740 -7688
rect 16804 -7752 16820 -7688
rect 16724 -7768 16820 -7752
rect 16724 -7832 16740 -7768
rect 16804 -7832 16820 -7768
rect 16724 -7848 16820 -7832
rect 16724 -7912 16740 -7848
rect 16804 -7912 16820 -7848
rect 16724 -7928 16820 -7912
rect 16724 -7992 16740 -7928
rect 16804 -7992 16820 -7928
rect 16724 -8008 16820 -7992
rect 16724 -8072 16740 -8008
rect 16804 -8072 16820 -8008
rect 16724 -8088 16820 -8072
rect 16724 -8152 16740 -8088
rect 16804 -8152 16820 -8088
rect 16724 -8168 16820 -8152
rect 15312 -8268 15408 -8232
rect 16724 -8232 16740 -8168
rect 16804 -8232 16820 -8168
rect 17143 -7488 17865 -7479
rect 17143 -8192 17152 -7488
rect 17856 -8192 17865 -7488
rect 17143 -8201 17865 -8192
rect 18136 -7512 18152 -7448
rect 18216 -7512 18232 -7448
rect 19548 -7448 19644 -7412
rect 18136 -7528 18232 -7512
rect 18136 -7592 18152 -7528
rect 18216 -7592 18232 -7528
rect 18136 -7608 18232 -7592
rect 18136 -7672 18152 -7608
rect 18216 -7672 18232 -7608
rect 18136 -7688 18232 -7672
rect 18136 -7752 18152 -7688
rect 18216 -7752 18232 -7688
rect 18136 -7768 18232 -7752
rect 18136 -7832 18152 -7768
rect 18216 -7832 18232 -7768
rect 18136 -7848 18232 -7832
rect 18136 -7912 18152 -7848
rect 18216 -7912 18232 -7848
rect 18136 -7928 18232 -7912
rect 18136 -7992 18152 -7928
rect 18216 -7992 18232 -7928
rect 18136 -8008 18232 -7992
rect 18136 -8072 18152 -8008
rect 18216 -8072 18232 -8008
rect 18136 -8088 18232 -8072
rect 18136 -8152 18152 -8088
rect 18216 -8152 18232 -8088
rect 18136 -8168 18232 -8152
rect 16724 -8268 16820 -8232
rect 18136 -8232 18152 -8168
rect 18216 -8232 18232 -8168
rect 18555 -7488 19277 -7479
rect 18555 -8192 18564 -7488
rect 19268 -8192 19277 -7488
rect 18555 -8201 19277 -8192
rect 19548 -7512 19564 -7448
rect 19628 -7512 19644 -7448
rect 20960 -7448 21056 -7412
rect 19548 -7528 19644 -7512
rect 19548 -7592 19564 -7528
rect 19628 -7592 19644 -7528
rect 19548 -7608 19644 -7592
rect 19548 -7672 19564 -7608
rect 19628 -7672 19644 -7608
rect 19548 -7688 19644 -7672
rect 19548 -7752 19564 -7688
rect 19628 -7752 19644 -7688
rect 19548 -7768 19644 -7752
rect 19548 -7832 19564 -7768
rect 19628 -7832 19644 -7768
rect 19548 -7848 19644 -7832
rect 19548 -7912 19564 -7848
rect 19628 -7912 19644 -7848
rect 19548 -7928 19644 -7912
rect 19548 -7992 19564 -7928
rect 19628 -7992 19644 -7928
rect 19548 -8008 19644 -7992
rect 19548 -8072 19564 -8008
rect 19628 -8072 19644 -8008
rect 19548 -8088 19644 -8072
rect 19548 -8152 19564 -8088
rect 19628 -8152 19644 -8088
rect 19548 -8168 19644 -8152
rect 18136 -8268 18232 -8232
rect 19548 -8232 19564 -8168
rect 19628 -8232 19644 -8168
rect 19967 -7488 20689 -7479
rect 19967 -8192 19976 -7488
rect 20680 -8192 20689 -7488
rect 19967 -8201 20689 -8192
rect 20960 -7512 20976 -7448
rect 21040 -7512 21056 -7448
rect 22372 -7448 22468 -7412
rect 20960 -7528 21056 -7512
rect 20960 -7592 20976 -7528
rect 21040 -7592 21056 -7528
rect 20960 -7608 21056 -7592
rect 20960 -7672 20976 -7608
rect 21040 -7672 21056 -7608
rect 20960 -7688 21056 -7672
rect 20960 -7752 20976 -7688
rect 21040 -7752 21056 -7688
rect 20960 -7768 21056 -7752
rect 20960 -7832 20976 -7768
rect 21040 -7832 21056 -7768
rect 20960 -7848 21056 -7832
rect 20960 -7912 20976 -7848
rect 21040 -7912 21056 -7848
rect 20960 -7928 21056 -7912
rect 20960 -7992 20976 -7928
rect 21040 -7992 21056 -7928
rect 20960 -8008 21056 -7992
rect 20960 -8072 20976 -8008
rect 21040 -8072 21056 -8008
rect 20960 -8088 21056 -8072
rect 20960 -8152 20976 -8088
rect 21040 -8152 21056 -8088
rect 20960 -8168 21056 -8152
rect 19548 -8268 19644 -8232
rect 20960 -8232 20976 -8168
rect 21040 -8232 21056 -8168
rect 21379 -7488 22101 -7479
rect 21379 -8192 21388 -7488
rect 22092 -8192 22101 -7488
rect 21379 -8201 22101 -8192
rect 22372 -7512 22388 -7448
rect 22452 -7512 22468 -7448
rect 23784 -7448 23880 -7412
rect 22372 -7528 22468 -7512
rect 22372 -7592 22388 -7528
rect 22452 -7592 22468 -7528
rect 22372 -7608 22468 -7592
rect 22372 -7672 22388 -7608
rect 22452 -7672 22468 -7608
rect 22372 -7688 22468 -7672
rect 22372 -7752 22388 -7688
rect 22452 -7752 22468 -7688
rect 22372 -7768 22468 -7752
rect 22372 -7832 22388 -7768
rect 22452 -7832 22468 -7768
rect 22372 -7848 22468 -7832
rect 22372 -7912 22388 -7848
rect 22452 -7912 22468 -7848
rect 22372 -7928 22468 -7912
rect 22372 -7992 22388 -7928
rect 22452 -7992 22468 -7928
rect 22372 -8008 22468 -7992
rect 22372 -8072 22388 -8008
rect 22452 -8072 22468 -8008
rect 22372 -8088 22468 -8072
rect 22372 -8152 22388 -8088
rect 22452 -8152 22468 -8088
rect 22372 -8168 22468 -8152
rect 20960 -8268 21056 -8232
rect 22372 -8232 22388 -8168
rect 22452 -8232 22468 -8168
rect 22791 -7488 23513 -7479
rect 22791 -8192 22800 -7488
rect 23504 -8192 23513 -7488
rect 22791 -8201 23513 -8192
rect 23784 -7512 23800 -7448
rect 23864 -7512 23880 -7448
rect 23784 -7528 23880 -7512
rect 23784 -7592 23800 -7528
rect 23864 -7592 23880 -7528
rect 23784 -7608 23880 -7592
rect 23784 -7672 23800 -7608
rect 23864 -7672 23880 -7608
rect 23784 -7688 23880 -7672
rect 23784 -7752 23800 -7688
rect 23864 -7752 23880 -7688
rect 23784 -7768 23880 -7752
rect 23784 -7832 23800 -7768
rect 23864 -7832 23880 -7768
rect 23784 -7848 23880 -7832
rect 23784 -7912 23800 -7848
rect 23864 -7912 23880 -7848
rect 23784 -7928 23880 -7912
rect 23784 -7992 23800 -7928
rect 23864 -7992 23880 -7928
rect 23784 -8008 23880 -7992
rect 23784 -8072 23800 -8008
rect 23864 -8072 23880 -8008
rect 23784 -8088 23880 -8072
rect 23784 -8152 23800 -8088
rect 23864 -8152 23880 -8088
rect 23784 -8168 23880 -8152
rect 22372 -8268 22468 -8232
rect 23784 -8232 23800 -8168
rect 23864 -8232 23880 -8168
rect 23784 -8268 23880 -8232
rect -22812 -8568 -22716 -8532
rect -23805 -8608 -23083 -8599
rect -23805 -9312 -23796 -8608
rect -23092 -9312 -23083 -8608
rect -23805 -9321 -23083 -9312
rect -22812 -8632 -22796 -8568
rect -22732 -8632 -22716 -8568
rect -21400 -8568 -21304 -8532
rect -22812 -8648 -22716 -8632
rect -22812 -8712 -22796 -8648
rect -22732 -8712 -22716 -8648
rect -22812 -8728 -22716 -8712
rect -22812 -8792 -22796 -8728
rect -22732 -8792 -22716 -8728
rect -22812 -8808 -22716 -8792
rect -22812 -8872 -22796 -8808
rect -22732 -8872 -22716 -8808
rect -22812 -8888 -22716 -8872
rect -22812 -8952 -22796 -8888
rect -22732 -8952 -22716 -8888
rect -22812 -8968 -22716 -8952
rect -22812 -9032 -22796 -8968
rect -22732 -9032 -22716 -8968
rect -22812 -9048 -22716 -9032
rect -22812 -9112 -22796 -9048
rect -22732 -9112 -22716 -9048
rect -22812 -9128 -22716 -9112
rect -22812 -9192 -22796 -9128
rect -22732 -9192 -22716 -9128
rect -22812 -9208 -22716 -9192
rect -22812 -9272 -22796 -9208
rect -22732 -9272 -22716 -9208
rect -22812 -9288 -22716 -9272
rect -22812 -9352 -22796 -9288
rect -22732 -9352 -22716 -9288
rect -22393 -8608 -21671 -8599
rect -22393 -9312 -22384 -8608
rect -21680 -9312 -21671 -8608
rect -22393 -9321 -21671 -9312
rect -21400 -8632 -21384 -8568
rect -21320 -8632 -21304 -8568
rect -19988 -8568 -19892 -8532
rect -21400 -8648 -21304 -8632
rect -21400 -8712 -21384 -8648
rect -21320 -8712 -21304 -8648
rect -21400 -8728 -21304 -8712
rect -21400 -8792 -21384 -8728
rect -21320 -8792 -21304 -8728
rect -21400 -8808 -21304 -8792
rect -21400 -8872 -21384 -8808
rect -21320 -8872 -21304 -8808
rect -21400 -8888 -21304 -8872
rect -21400 -8952 -21384 -8888
rect -21320 -8952 -21304 -8888
rect -21400 -8968 -21304 -8952
rect -21400 -9032 -21384 -8968
rect -21320 -9032 -21304 -8968
rect -21400 -9048 -21304 -9032
rect -21400 -9112 -21384 -9048
rect -21320 -9112 -21304 -9048
rect -21400 -9128 -21304 -9112
rect -21400 -9192 -21384 -9128
rect -21320 -9192 -21304 -9128
rect -21400 -9208 -21304 -9192
rect -21400 -9272 -21384 -9208
rect -21320 -9272 -21304 -9208
rect -21400 -9288 -21304 -9272
rect -22812 -9388 -22716 -9352
rect -21400 -9352 -21384 -9288
rect -21320 -9352 -21304 -9288
rect -20981 -8608 -20259 -8599
rect -20981 -9312 -20972 -8608
rect -20268 -9312 -20259 -8608
rect -20981 -9321 -20259 -9312
rect -19988 -8632 -19972 -8568
rect -19908 -8632 -19892 -8568
rect -18576 -8568 -18480 -8532
rect -19988 -8648 -19892 -8632
rect -19988 -8712 -19972 -8648
rect -19908 -8712 -19892 -8648
rect -19988 -8728 -19892 -8712
rect -19988 -8792 -19972 -8728
rect -19908 -8792 -19892 -8728
rect -19988 -8808 -19892 -8792
rect -19988 -8872 -19972 -8808
rect -19908 -8872 -19892 -8808
rect -19988 -8888 -19892 -8872
rect -19988 -8952 -19972 -8888
rect -19908 -8952 -19892 -8888
rect -19988 -8968 -19892 -8952
rect -19988 -9032 -19972 -8968
rect -19908 -9032 -19892 -8968
rect -19988 -9048 -19892 -9032
rect -19988 -9112 -19972 -9048
rect -19908 -9112 -19892 -9048
rect -19988 -9128 -19892 -9112
rect -19988 -9192 -19972 -9128
rect -19908 -9192 -19892 -9128
rect -19988 -9208 -19892 -9192
rect -19988 -9272 -19972 -9208
rect -19908 -9272 -19892 -9208
rect -19988 -9288 -19892 -9272
rect -21400 -9388 -21304 -9352
rect -19988 -9352 -19972 -9288
rect -19908 -9352 -19892 -9288
rect -19569 -8608 -18847 -8599
rect -19569 -9312 -19560 -8608
rect -18856 -9312 -18847 -8608
rect -19569 -9321 -18847 -9312
rect -18576 -8632 -18560 -8568
rect -18496 -8632 -18480 -8568
rect -17164 -8568 -17068 -8532
rect -18576 -8648 -18480 -8632
rect -18576 -8712 -18560 -8648
rect -18496 -8712 -18480 -8648
rect -18576 -8728 -18480 -8712
rect -18576 -8792 -18560 -8728
rect -18496 -8792 -18480 -8728
rect -18576 -8808 -18480 -8792
rect -18576 -8872 -18560 -8808
rect -18496 -8872 -18480 -8808
rect -18576 -8888 -18480 -8872
rect -18576 -8952 -18560 -8888
rect -18496 -8952 -18480 -8888
rect -18576 -8968 -18480 -8952
rect -18576 -9032 -18560 -8968
rect -18496 -9032 -18480 -8968
rect -18576 -9048 -18480 -9032
rect -18576 -9112 -18560 -9048
rect -18496 -9112 -18480 -9048
rect -18576 -9128 -18480 -9112
rect -18576 -9192 -18560 -9128
rect -18496 -9192 -18480 -9128
rect -18576 -9208 -18480 -9192
rect -18576 -9272 -18560 -9208
rect -18496 -9272 -18480 -9208
rect -18576 -9288 -18480 -9272
rect -19988 -9388 -19892 -9352
rect -18576 -9352 -18560 -9288
rect -18496 -9352 -18480 -9288
rect -18157 -8608 -17435 -8599
rect -18157 -9312 -18148 -8608
rect -17444 -9312 -17435 -8608
rect -18157 -9321 -17435 -9312
rect -17164 -8632 -17148 -8568
rect -17084 -8632 -17068 -8568
rect -15752 -8568 -15656 -8532
rect -17164 -8648 -17068 -8632
rect -17164 -8712 -17148 -8648
rect -17084 -8712 -17068 -8648
rect -17164 -8728 -17068 -8712
rect -17164 -8792 -17148 -8728
rect -17084 -8792 -17068 -8728
rect -17164 -8808 -17068 -8792
rect -17164 -8872 -17148 -8808
rect -17084 -8872 -17068 -8808
rect -17164 -8888 -17068 -8872
rect -17164 -8952 -17148 -8888
rect -17084 -8952 -17068 -8888
rect -17164 -8968 -17068 -8952
rect -17164 -9032 -17148 -8968
rect -17084 -9032 -17068 -8968
rect -17164 -9048 -17068 -9032
rect -17164 -9112 -17148 -9048
rect -17084 -9112 -17068 -9048
rect -17164 -9128 -17068 -9112
rect -17164 -9192 -17148 -9128
rect -17084 -9192 -17068 -9128
rect -17164 -9208 -17068 -9192
rect -17164 -9272 -17148 -9208
rect -17084 -9272 -17068 -9208
rect -17164 -9288 -17068 -9272
rect -18576 -9388 -18480 -9352
rect -17164 -9352 -17148 -9288
rect -17084 -9352 -17068 -9288
rect -16745 -8608 -16023 -8599
rect -16745 -9312 -16736 -8608
rect -16032 -9312 -16023 -8608
rect -16745 -9321 -16023 -9312
rect -15752 -8632 -15736 -8568
rect -15672 -8632 -15656 -8568
rect -14340 -8568 -14244 -8532
rect -15752 -8648 -15656 -8632
rect -15752 -8712 -15736 -8648
rect -15672 -8712 -15656 -8648
rect -15752 -8728 -15656 -8712
rect -15752 -8792 -15736 -8728
rect -15672 -8792 -15656 -8728
rect -15752 -8808 -15656 -8792
rect -15752 -8872 -15736 -8808
rect -15672 -8872 -15656 -8808
rect -15752 -8888 -15656 -8872
rect -15752 -8952 -15736 -8888
rect -15672 -8952 -15656 -8888
rect -15752 -8968 -15656 -8952
rect -15752 -9032 -15736 -8968
rect -15672 -9032 -15656 -8968
rect -15752 -9048 -15656 -9032
rect -15752 -9112 -15736 -9048
rect -15672 -9112 -15656 -9048
rect -15752 -9128 -15656 -9112
rect -15752 -9192 -15736 -9128
rect -15672 -9192 -15656 -9128
rect -15752 -9208 -15656 -9192
rect -15752 -9272 -15736 -9208
rect -15672 -9272 -15656 -9208
rect -15752 -9288 -15656 -9272
rect -17164 -9388 -17068 -9352
rect -15752 -9352 -15736 -9288
rect -15672 -9352 -15656 -9288
rect -15333 -8608 -14611 -8599
rect -15333 -9312 -15324 -8608
rect -14620 -9312 -14611 -8608
rect -15333 -9321 -14611 -9312
rect -14340 -8632 -14324 -8568
rect -14260 -8632 -14244 -8568
rect -12928 -8568 -12832 -8532
rect -14340 -8648 -14244 -8632
rect -14340 -8712 -14324 -8648
rect -14260 -8712 -14244 -8648
rect -14340 -8728 -14244 -8712
rect -14340 -8792 -14324 -8728
rect -14260 -8792 -14244 -8728
rect -14340 -8808 -14244 -8792
rect -14340 -8872 -14324 -8808
rect -14260 -8872 -14244 -8808
rect -14340 -8888 -14244 -8872
rect -14340 -8952 -14324 -8888
rect -14260 -8952 -14244 -8888
rect -14340 -8968 -14244 -8952
rect -14340 -9032 -14324 -8968
rect -14260 -9032 -14244 -8968
rect -14340 -9048 -14244 -9032
rect -14340 -9112 -14324 -9048
rect -14260 -9112 -14244 -9048
rect -14340 -9128 -14244 -9112
rect -14340 -9192 -14324 -9128
rect -14260 -9192 -14244 -9128
rect -14340 -9208 -14244 -9192
rect -14340 -9272 -14324 -9208
rect -14260 -9272 -14244 -9208
rect -14340 -9288 -14244 -9272
rect -15752 -9388 -15656 -9352
rect -14340 -9352 -14324 -9288
rect -14260 -9352 -14244 -9288
rect -13921 -8608 -13199 -8599
rect -13921 -9312 -13912 -8608
rect -13208 -9312 -13199 -8608
rect -13921 -9321 -13199 -9312
rect -12928 -8632 -12912 -8568
rect -12848 -8632 -12832 -8568
rect -11516 -8568 -11420 -8532
rect -12928 -8648 -12832 -8632
rect -12928 -8712 -12912 -8648
rect -12848 -8712 -12832 -8648
rect -12928 -8728 -12832 -8712
rect -12928 -8792 -12912 -8728
rect -12848 -8792 -12832 -8728
rect -12928 -8808 -12832 -8792
rect -12928 -8872 -12912 -8808
rect -12848 -8872 -12832 -8808
rect -12928 -8888 -12832 -8872
rect -12928 -8952 -12912 -8888
rect -12848 -8952 -12832 -8888
rect -12928 -8968 -12832 -8952
rect -12928 -9032 -12912 -8968
rect -12848 -9032 -12832 -8968
rect -12928 -9048 -12832 -9032
rect -12928 -9112 -12912 -9048
rect -12848 -9112 -12832 -9048
rect -12928 -9128 -12832 -9112
rect -12928 -9192 -12912 -9128
rect -12848 -9192 -12832 -9128
rect -12928 -9208 -12832 -9192
rect -12928 -9272 -12912 -9208
rect -12848 -9272 -12832 -9208
rect -12928 -9288 -12832 -9272
rect -14340 -9388 -14244 -9352
rect -12928 -9352 -12912 -9288
rect -12848 -9352 -12832 -9288
rect -12509 -8608 -11787 -8599
rect -12509 -9312 -12500 -8608
rect -11796 -9312 -11787 -8608
rect -12509 -9321 -11787 -9312
rect -11516 -8632 -11500 -8568
rect -11436 -8632 -11420 -8568
rect -10104 -8568 -10008 -8532
rect -11516 -8648 -11420 -8632
rect -11516 -8712 -11500 -8648
rect -11436 -8712 -11420 -8648
rect -11516 -8728 -11420 -8712
rect -11516 -8792 -11500 -8728
rect -11436 -8792 -11420 -8728
rect -11516 -8808 -11420 -8792
rect -11516 -8872 -11500 -8808
rect -11436 -8872 -11420 -8808
rect -11516 -8888 -11420 -8872
rect -11516 -8952 -11500 -8888
rect -11436 -8952 -11420 -8888
rect -11516 -8968 -11420 -8952
rect -11516 -9032 -11500 -8968
rect -11436 -9032 -11420 -8968
rect -11516 -9048 -11420 -9032
rect -11516 -9112 -11500 -9048
rect -11436 -9112 -11420 -9048
rect -11516 -9128 -11420 -9112
rect -11516 -9192 -11500 -9128
rect -11436 -9192 -11420 -9128
rect -11516 -9208 -11420 -9192
rect -11516 -9272 -11500 -9208
rect -11436 -9272 -11420 -9208
rect -11516 -9288 -11420 -9272
rect -12928 -9388 -12832 -9352
rect -11516 -9352 -11500 -9288
rect -11436 -9352 -11420 -9288
rect -11097 -8608 -10375 -8599
rect -11097 -9312 -11088 -8608
rect -10384 -9312 -10375 -8608
rect -11097 -9321 -10375 -9312
rect -10104 -8632 -10088 -8568
rect -10024 -8632 -10008 -8568
rect -8692 -8568 -8596 -8532
rect -10104 -8648 -10008 -8632
rect -10104 -8712 -10088 -8648
rect -10024 -8712 -10008 -8648
rect -10104 -8728 -10008 -8712
rect -10104 -8792 -10088 -8728
rect -10024 -8792 -10008 -8728
rect -10104 -8808 -10008 -8792
rect -10104 -8872 -10088 -8808
rect -10024 -8872 -10008 -8808
rect -10104 -8888 -10008 -8872
rect -10104 -8952 -10088 -8888
rect -10024 -8952 -10008 -8888
rect -10104 -8968 -10008 -8952
rect -10104 -9032 -10088 -8968
rect -10024 -9032 -10008 -8968
rect -10104 -9048 -10008 -9032
rect -10104 -9112 -10088 -9048
rect -10024 -9112 -10008 -9048
rect -10104 -9128 -10008 -9112
rect -10104 -9192 -10088 -9128
rect -10024 -9192 -10008 -9128
rect -10104 -9208 -10008 -9192
rect -10104 -9272 -10088 -9208
rect -10024 -9272 -10008 -9208
rect -10104 -9288 -10008 -9272
rect -11516 -9388 -11420 -9352
rect -10104 -9352 -10088 -9288
rect -10024 -9352 -10008 -9288
rect -9685 -8608 -8963 -8599
rect -9685 -9312 -9676 -8608
rect -8972 -9312 -8963 -8608
rect -9685 -9321 -8963 -9312
rect -8692 -8632 -8676 -8568
rect -8612 -8632 -8596 -8568
rect -7280 -8568 -7184 -8532
rect -8692 -8648 -8596 -8632
rect -8692 -8712 -8676 -8648
rect -8612 -8712 -8596 -8648
rect -8692 -8728 -8596 -8712
rect -8692 -8792 -8676 -8728
rect -8612 -8792 -8596 -8728
rect -8692 -8808 -8596 -8792
rect -8692 -8872 -8676 -8808
rect -8612 -8872 -8596 -8808
rect -8692 -8888 -8596 -8872
rect -8692 -8952 -8676 -8888
rect -8612 -8952 -8596 -8888
rect -8692 -8968 -8596 -8952
rect -8692 -9032 -8676 -8968
rect -8612 -9032 -8596 -8968
rect -8692 -9048 -8596 -9032
rect -8692 -9112 -8676 -9048
rect -8612 -9112 -8596 -9048
rect -8692 -9128 -8596 -9112
rect -8692 -9192 -8676 -9128
rect -8612 -9192 -8596 -9128
rect -8692 -9208 -8596 -9192
rect -8692 -9272 -8676 -9208
rect -8612 -9272 -8596 -9208
rect -8692 -9288 -8596 -9272
rect -10104 -9388 -10008 -9352
rect -8692 -9352 -8676 -9288
rect -8612 -9352 -8596 -9288
rect -8273 -8608 -7551 -8599
rect -8273 -9312 -8264 -8608
rect -7560 -9312 -7551 -8608
rect -8273 -9321 -7551 -9312
rect -7280 -8632 -7264 -8568
rect -7200 -8632 -7184 -8568
rect -5868 -8568 -5772 -8532
rect -7280 -8648 -7184 -8632
rect -7280 -8712 -7264 -8648
rect -7200 -8712 -7184 -8648
rect -7280 -8728 -7184 -8712
rect -7280 -8792 -7264 -8728
rect -7200 -8792 -7184 -8728
rect -7280 -8808 -7184 -8792
rect -7280 -8872 -7264 -8808
rect -7200 -8872 -7184 -8808
rect -7280 -8888 -7184 -8872
rect -7280 -8952 -7264 -8888
rect -7200 -8952 -7184 -8888
rect -7280 -8968 -7184 -8952
rect -7280 -9032 -7264 -8968
rect -7200 -9032 -7184 -8968
rect -7280 -9048 -7184 -9032
rect -7280 -9112 -7264 -9048
rect -7200 -9112 -7184 -9048
rect -7280 -9128 -7184 -9112
rect -7280 -9192 -7264 -9128
rect -7200 -9192 -7184 -9128
rect -7280 -9208 -7184 -9192
rect -7280 -9272 -7264 -9208
rect -7200 -9272 -7184 -9208
rect -7280 -9288 -7184 -9272
rect -8692 -9388 -8596 -9352
rect -7280 -9352 -7264 -9288
rect -7200 -9352 -7184 -9288
rect -6861 -8608 -6139 -8599
rect -6861 -9312 -6852 -8608
rect -6148 -9312 -6139 -8608
rect -6861 -9321 -6139 -9312
rect -5868 -8632 -5852 -8568
rect -5788 -8632 -5772 -8568
rect -4456 -8568 -4360 -8532
rect -5868 -8648 -5772 -8632
rect -5868 -8712 -5852 -8648
rect -5788 -8712 -5772 -8648
rect -5868 -8728 -5772 -8712
rect -5868 -8792 -5852 -8728
rect -5788 -8792 -5772 -8728
rect -5868 -8808 -5772 -8792
rect -5868 -8872 -5852 -8808
rect -5788 -8872 -5772 -8808
rect -5868 -8888 -5772 -8872
rect -5868 -8952 -5852 -8888
rect -5788 -8952 -5772 -8888
rect -5868 -8968 -5772 -8952
rect -5868 -9032 -5852 -8968
rect -5788 -9032 -5772 -8968
rect -5868 -9048 -5772 -9032
rect -5868 -9112 -5852 -9048
rect -5788 -9112 -5772 -9048
rect -5868 -9128 -5772 -9112
rect -5868 -9192 -5852 -9128
rect -5788 -9192 -5772 -9128
rect -5868 -9208 -5772 -9192
rect -5868 -9272 -5852 -9208
rect -5788 -9272 -5772 -9208
rect -5868 -9288 -5772 -9272
rect -7280 -9388 -7184 -9352
rect -5868 -9352 -5852 -9288
rect -5788 -9352 -5772 -9288
rect -5449 -8608 -4727 -8599
rect -5449 -9312 -5440 -8608
rect -4736 -9312 -4727 -8608
rect -5449 -9321 -4727 -9312
rect -4456 -8632 -4440 -8568
rect -4376 -8632 -4360 -8568
rect -3044 -8568 -2948 -8532
rect -4456 -8648 -4360 -8632
rect -4456 -8712 -4440 -8648
rect -4376 -8712 -4360 -8648
rect -4456 -8728 -4360 -8712
rect -4456 -8792 -4440 -8728
rect -4376 -8792 -4360 -8728
rect -4456 -8808 -4360 -8792
rect -4456 -8872 -4440 -8808
rect -4376 -8872 -4360 -8808
rect -4456 -8888 -4360 -8872
rect -4456 -8952 -4440 -8888
rect -4376 -8952 -4360 -8888
rect -4456 -8968 -4360 -8952
rect -4456 -9032 -4440 -8968
rect -4376 -9032 -4360 -8968
rect -4456 -9048 -4360 -9032
rect -4456 -9112 -4440 -9048
rect -4376 -9112 -4360 -9048
rect -4456 -9128 -4360 -9112
rect -4456 -9192 -4440 -9128
rect -4376 -9192 -4360 -9128
rect -4456 -9208 -4360 -9192
rect -4456 -9272 -4440 -9208
rect -4376 -9272 -4360 -9208
rect -4456 -9288 -4360 -9272
rect -5868 -9388 -5772 -9352
rect -4456 -9352 -4440 -9288
rect -4376 -9352 -4360 -9288
rect -4037 -8608 -3315 -8599
rect -4037 -9312 -4028 -8608
rect -3324 -9312 -3315 -8608
rect -4037 -9321 -3315 -9312
rect -3044 -8632 -3028 -8568
rect -2964 -8632 -2948 -8568
rect -1632 -8568 -1536 -8532
rect -3044 -8648 -2948 -8632
rect -3044 -8712 -3028 -8648
rect -2964 -8712 -2948 -8648
rect -3044 -8728 -2948 -8712
rect -3044 -8792 -3028 -8728
rect -2964 -8792 -2948 -8728
rect -3044 -8808 -2948 -8792
rect -3044 -8872 -3028 -8808
rect -2964 -8872 -2948 -8808
rect -3044 -8888 -2948 -8872
rect -3044 -8952 -3028 -8888
rect -2964 -8952 -2948 -8888
rect -3044 -8968 -2948 -8952
rect -3044 -9032 -3028 -8968
rect -2964 -9032 -2948 -8968
rect -3044 -9048 -2948 -9032
rect -3044 -9112 -3028 -9048
rect -2964 -9112 -2948 -9048
rect -3044 -9128 -2948 -9112
rect -3044 -9192 -3028 -9128
rect -2964 -9192 -2948 -9128
rect -3044 -9208 -2948 -9192
rect -3044 -9272 -3028 -9208
rect -2964 -9272 -2948 -9208
rect -3044 -9288 -2948 -9272
rect -4456 -9388 -4360 -9352
rect -3044 -9352 -3028 -9288
rect -2964 -9352 -2948 -9288
rect -2625 -8608 -1903 -8599
rect -2625 -9312 -2616 -8608
rect -1912 -9312 -1903 -8608
rect -2625 -9321 -1903 -9312
rect -1632 -8632 -1616 -8568
rect -1552 -8632 -1536 -8568
rect -220 -8568 -124 -8532
rect -1632 -8648 -1536 -8632
rect -1632 -8712 -1616 -8648
rect -1552 -8712 -1536 -8648
rect -1632 -8728 -1536 -8712
rect -1632 -8792 -1616 -8728
rect -1552 -8792 -1536 -8728
rect -1632 -8808 -1536 -8792
rect -1632 -8872 -1616 -8808
rect -1552 -8872 -1536 -8808
rect -1632 -8888 -1536 -8872
rect -1632 -8952 -1616 -8888
rect -1552 -8952 -1536 -8888
rect -1632 -8968 -1536 -8952
rect -1632 -9032 -1616 -8968
rect -1552 -9032 -1536 -8968
rect -1632 -9048 -1536 -9032
rect -1632 -9112 -1616 -9048
rect -1552 -9112 -1536 -9048
rect -1632 -9128 -1536 -9112
rect -1632 -9192 -1616 -9128
rect -1552 -9192 -1536 -9128
rect -1632 -9208 -1536 -9192
rect -1632 -9272 -1616 -9208
rect -1552 -9272 -1536 -9208
rect -1632 -9288 -1536 -9272
rect -3044 -9388 -2948 -9352
rect -1632 -9352 -1616 -9288
rect -1552 -9352 -1536 -9288
rect -1213 -8608 -491 -8599
rect -1213 -9312 -1204 -8608
rect -500 -9312 -491 -8608
rect -1213 -9321 -491 -9312
rect -220 -8632 -204 -8568
rect -140 -8632 -124 -8568
rect 1192 -8568 1288 -8532
rect -220 -8648 -124 -8632
rect -220 -8712 -204 -8648
rect -140 -8712 -124 -8648
rect -220 -8728 -124 -8712
rect -220 -8792 -204 -8728
rect -140 -8792 -124 -8728
rect -220 -8808 -124 -8792
rect -220 -8872 -204 -8808
rect -140 -8872 -124 -8808
rect -220 -8888 -124 -8872
rect -220 -8952 -204 -8888
rect -140 -8952 -124 -8888
rect -220 -8968 -124 -8952
rect -220 -9032 -204 -8968
rect -140 -9032 -124 -8968
rect -220 -9048 -124 -9032
rect -220 -9112 -204 -9048
rect -140 -9112 -124 -9048
rect -220 -9128 -124 -9112
rect -220 -9192 -204 -9128
rect -140 -9192 -124 -9128
rect -220 -9208 -124 -9192
rect -220 -9272 -204 -9208
rect -140 -9272 -124 -9208
rect -220 -9288 -124 -9272
rect -1632 -9388 -1536 -9352
rect -220 -9352 -204 -9288
rect -140 -9352 -124 -9288
rect 199 -8608 921 -8599
rect 199 -9312 208 -8608
rect 912 -9312 921 -8608
rect 199 -9321 921 -9312
rect 1192 -8632 1208 -8568
rect 1272 -8632 1288 -8568
rect 2604 -8568 2700 -8532
rect 1192 -8648 1288 -8632
rect 1192 -8712 1208 -8648
rect 1272 -8712 1288 -8648
rect 1192 -8728 1288 -8712
rect 1192 -8792 1208 -8728
rect 1272 -8792 1288 -8728
rect 1192 -8808 1288 -8792
rect 1192 -8872 1208 -8808
rect 1272 -8872 1288 -8808
rect 1192 -8888 1288 -8872
rect 1192 -8952 1208 -8888
rect 1272 -8952 1288 -8888
rect 1192 -8968 1288 -8952
rect 1192 -9032 1208 -8968
rect 1272 -9032 1288 -8968
rect 1192 -9048 1288 -9032
rect 1192 -9112 1208 -9048
rect 1272 -9112 1288 -9048
rect 1192 -9128 1288 -9112
rect 1192 -9192 1208 -9128
rect 1272 -9192 1288 -9128
rect 1192 -9208 1288 -9192
rect 1192 -9272 1208 -9208
rect 1272 -9272 1288 -9208
rect 1192 -9288 1288 -9272
rect -220 -9388 -124 -9352
rect 1192 -9352 1208 -9288
rect 1272 -9352 1288 -9288
rect 1611 -8608 2333 -8599
rect 1611 -9312 1620 -8608
rect 2324 -9312 2333 -8608
rect 1611 -9321 2333 -9312
rect 2604 -8632 2620 -8568
rect 2684 -8632 2700 -8568
rect 4016 -8568 4112 -8532
rect 2604 -8648 2700 -8632
rect 2604 -8712 2620 -8648
rect 2684 -8712 2700 -8648
rect 2604 -8728 2700 -8712
rect 2604 -8792 2620 -8728
rect 2684 -8792 2700 -8728
rect 2604 -8808 2700 -8792
rect 2604 -8872 2620 -8808
rect 2684 -8872 2700 -8808
rect 2604 -8888 2700 -8872
rect 2604 -8952 2620 -8888
rect 2684 -8952 2700 -8888
rect 2604 -8968 2700 -8952
rect 2604 -9032 2620 -8968
rect 2684 -9032 2700 -8968
rect 2604 -9048 2700 -9032
rect 2604 -9112 2620 -9048
rect 2684 -9112 2700 -9048
rect 2604 -9128 2700 -9112
rect 2604 -9192 2620 -9128
rect 2684 -9192 2700 -9128
rect 2604 -9208 2700 -9192
rect 2604 -9272 2620 -9208
rect 2684 -9272 2700 -9208
rect 2604 -9288 2700 -9272
rect 1192 -9388 1288 -9352
rect 2604 -9352 2620 -9288
rect 2684 -9352 2700 -9288
rect 3023 -8608 3745 -8599
rect 3023 -9312 3032 -8608
rect 3736 -9312 3745 -8608
rect 3023 -9321 3745 -9312
rect 4016 -8632 4032 -8568
rect 4096 -8632 4112 -8568
rect 5428 -8568 5524 -8532
rect 4016 -8648 4112 -8632
rect 4016 -8712 4032 -8648
rect 4096 -8712 4112 -8648
rect 4016 -8728 4112 -8712
rect 4016 -8792 4032 -8728
rect 4096 -8792 4112 -8728
rect 4016 -8808 4112 -8792
rect 4016 -8872 4032 -8808
rect 4096 -8872 4112 -8808
rect 4016 -8888 4112 -8872
rect 4016 -8952 4032 -8888
rect 4096 -8952 4112 -8888
rect 4016 -8968 4112 -8952
rect 4016 -9032 4032 -8968
rect 4096 -9032 4112 -8968
rect 4016 -9048 4112 -9032
rect 4016 -9112 4032 -9048
rect 4096 -9112 4112 -9048
rect 4016 -9128 4112 -9112
rect 4016 -9192 4032 -9128
rect 4096 -9192 4112 -9128
rect 4016 -9208 4112 -9192
rect 4016 -9272 4032 -9208
rect 4096 -9272 4112 -9208
rect 4016 -9288 4112 -9272
rect 2604 -9388 2700 -9352
rect 4016 -9352 4032 -9288
rect 4096 -9352 4112 -9288
rect 4435 -8608 5157 -8599
rect 4435 -9312 4444 -8608
rect 5148 -9312 5157 -8608
rect 4435 -9321 5157 -9312
rect 5428 -8632 5444 -8568
rect 5508 -8632 5524 -8568
rect 6840 -8568 6936 -8532
rect 5428 -8648 5524 -8632
rect 5428 -8712 5444 -8648
rect 5508 -8712 5524 -8648
rect 5428 -8728 5524 -8712
rect 5428 -8792 5444 -8728
rect 5508 -8792 5524 -8728
rect 5428 -8808 5524 -8792
rect 5428 -8872 5444 -8808
rect 5508 -8872 5524 -8808
rect 5428 -8888 5524 -8872
rect 5428 -8952 5444 -8888
rect 5508 -8952 5524 -8888
rect 5428 -8968 5524 -8952
rect 5428 -9032 5444 -8968
rect 5508 -9032 5524 -8968
rect 5428 -9048 5524 -9032
rect 5428 -9112 5444 -9048
rect 5508 -9112 5524 -9048
rect 5428 -9128 5524 -9112
rect 5428 -9192 5444 -9128
rect 5508 -9192 5524 -9128
rect 5428 -9208 5524 -9192
rect 5428 -9272 5444 -9208
rect 5508 -9272 5524 -9208
rect 5428 -9288 5524 -9272
rect 4016 -9388 4112 -9352
rect 5428 -9352 5444 -9288
rect 5508 -9352 5524 -9288
rect 5847 -8608 6569 -8599
rect 5847 -9312 5856 -8608
rect 6560 -9312 6569 -8608
rect 5847 -9321 6569 -9312
rect 6840 -8632 6856 -8568
rect 6920 -8632 6936 -8568
rect 8252 -8568 8348 -8532
rect 6840 -8648 6936 -8632
rect 6840 -8712 6856 -8648
rect 6920 -8712 6936 -8648
rect 6840 -8728 6936 -8712
rect 6840 -8792 6856 -8728
rect 6920 -8792 6936 -8728
rect 6840 -8808 6936 -8792
rect 6840 -8872 6856 -8808
rect 6920 -8872 6936 -8808
rect 6840 -8888 6936 -8872
rect 6840 -8952 6856 -8888
rect 6920 -8952 6936 -8888
rect 6840 -8968 6936 -8952
rect 6840 -9032 6856 -8968
rect 6920 -9032 6936 -8968
rect 6840 -9048 6936 -9032
rect 6840 -9112 6856 -9048
rect 6920 -9112 6936 -9048
rect 6840 -9128 6936 -9112
rect 6840 -9192 6856 -9128
rect 6920 -9192 6936 -9128
rect 6840 -9208 6936 -9192
rect 6840 -9272 6856 -9208
rect 6920 -9272 6936 -9208
rect 6840 -9288 6936 -9272
rect 5428 -9388 5524 -9352
rect 6840 -9352 6856 -9288
rect 6920 -9352 6936 -9288
rect 7259 -8608 7981 -8599
rect 7259 -9312 7268 -8608
rect 7972 -9312 7981 -8608
rect 7259 -9321 7981 -9312
rect 8252 -8632 8268 -8568
rect 8332 -8632 8348 -8568
rect 9664 -8568 9760 -8532
rect 8252 -8648 8348 -8632
rect 8252 -8712 8268 -8648
rect 8332 -8712 8348 -8648
rect 8252 -8728 8348 -8712
rect 8252 -8792 8268 -8728
rect 8332 -8792 8348 -8728
rect 8252 -8808 8348 -8792
rect 8252 -8872 8268 -8808
rect 8332 -8872 8348 -8808
rect 8252 -8888 8348 -8872
rect 8252 -8952 8268 -8888
rect 8332 -8952 8348 -8888
rect 8252 -8968 8348 -8952
rect 8252 -9032 8268 -8968
rect 8332 -9032 8348 -8968
rect 8252 -9048 8348 -9032
rect 8252 -9112 8268 -9048
rect 8332 -9112 8348 -9048
rect 8252 -9128 8348 -9112
rect 8252 -9192 8268 -9128
rect 8332 -9192 8348 -9128
rect 8252 -9208 8348 -9192
rect 8252 -9272 8268 -9208
rect 8332 -9272 8348 -9208
rect 8252 -9288 8348 -9272
rect 6840 -9388 6936 -9352
rect 8252 -9352 8268 -9288
rect 8332 -9352 8348 -9288
rect 8671 -8608 9393 -8599
rect 8671 -9312 8680 -8608
rect 9384 -9312 9393 -8608
rect 8671 -9321 9393 -9312
rect 9664 -8632 9680 -8568
rect 9744 -8632 9760 -8568
rect 11076 -8568 11172 -8532
rect 9664 -8648 9760 -8632
rect 9664 -8712 9680 -8648
rect 9744 -8712 9760 -8648
rect 9664 -8728 9760 -8712
rect 9664 -8792 9680 -8728
rect 9744 -8792 9760 -8728
rect 9664 -8808 9760 -8792
rect 9664 -8872 9680 -8808
rect 9744 -8872 9760 -8808
rect 9664 -8888 9760 -8872
rect 9664 -8952 9680 -8888
rect 9744 -8952 9760 -8888
rect 9664 -8968 9760 -8952
rect 9664 -9032 9680 -8968
rect 9744 -9032 9760 -8968
rect 9664 -9048 9760 -9032
rect 9664 -9112 9680 -9048
rect 9744 -9112 9760 -9048
rect 9664 -9128 9760 -9112
rect 9664 -9192 9680 -9128
rect 9744 -9192 9760 -9128
rect 9664 -9208 9760 -9192
rect 9664 -9272 9680 -9208
rect 9744 -9272 9760 -9208
rect 9664 -9288 9760 -9272
rect 8252 -9388 8348 -9352
rect 9664 -9352 9680 -9288
rect 9744 -9352 9760 -9288
rect 10083 -8608 10805 -8599
rect 10083 -9312 10092 -8608
rect 10796 -9312 10805 -8608
rect 10083 -9321 10805 -9312
rect 11076 -8632 11092 -8568
rect 11156 -8632 11172 -8568
rect 12488 -8568 12584 -8532
rect 11076 -8648 11172 -8632
rect 11076 -8712 11092 -8648
rect 11156 -8712 11172 -8648
rect 11076 -8728 11172 -8712
rect 11076 -8792 11092 -8728
rect 11156 -8792 11172 -8728
rect 11076 -8808 11172 -8792
rect 11076 -8872 11092 -8808
rect 11156 -8872 11172 -8808
rect 11076 -8888 11172 -8872
rect 11076 -8952 11092 -8888
rect 11156 -8952 11172 -8888
rect 11076 -8968 11172 -8952
rect 11076 -9032 11092 -8968
rect 11156 -9032 11172 -8968
rect 11076 -9048 11172 -9032
rect 11076 -9112 11092 -9048
rect 11156 -9112 11172 -9048
rect 11076 -9128 11172 -9112
rect 11076 -9192 11092 -9128
rect 11156 -9192 11172 -9128
rect 11076 -9208 11172 -9192
rect 11076 -9272 11092 -9208
rect 11156 -9272 11172 -9208
rect 11076 -9288 11172 -9272
rect 9664 -9388 9760 -9352
rect 11076 -9352 11092 -9288
rect 11156 -9352 11172 -9288
rect 11495 -8608 12217 -8599
rect 11495 -9312 11504 -8608
rect 12208 -9312 12217 -8608
rect 11495 -9321 12217 -9312
rect 12488 -8632 12504 -8568
rect 12568 -8632 12584 -8568
rect 13900 -8568 13996 -8532
rect 12488 -8648 12584 -8632
rect 12488 -8712 12504 -8648
rect 12568 -8712 12584 -8648
rect 12488 -8728 12584 -8712
rect 12488 -8792 12504 -8728
rect 12568 -8792 12584 -8728
rect 12488 -8808 12584 -8792
rect 12488 -8872 12504 -8808
rect 12568 -8872 12584 -8808
rect 12488 -8888 12584 -8872
rect 12488 -8952 12504 -8888
rect 12568 -8952 12584 -8888
rect 12488 -8968 12584 -8952
rect 12488 -9032 12504 -8968
rect 12568 -9032 12584 -8968
rect 12488 -9048 12584 -9032
rect 12488 -9112 12504 -9048
rect 12568 -9112 12584 -9048
rect 12488 -9128 12584 -9112
rect 12488 -9192 12504 -9128
rect 12568 -9192 12584 -9128
rect 12488 -9208 12584 -9192
rect 12488 -9272 12504 -9208
rect 12568 -9272 12584 -9208
rect 12488 -9288 12584 -9272
rect 11076 -9388 11172 -9352
rect 12488 -9352 12504 -9288
rect 12568 -9352 12584 -9288
rect 12907 -8608 13629 -8599
rect 12907 -9312 12916 -8608
rect 13620 -9312 13629 -8608
rect 12907 -9321 13629 -9312
rect 13900 -8632 13916 -8568
rect 13980 -8632 13996 -8568
rect 15312 -8568 15408 -8532
rect 13900 -8648 13996 -8632
rect 13900 -8712 13916 -8648
rect 13980 -8712 13996 -8648
rect 13900 -8728 13996 -8712
rect 13900 -8792 13916 -8728
rect 13980 -8792 13996 -8728
rect 13900 -8808 13996 -8792
rect 13900 -8872 13916 -8808
rect 13980 -8872 13996 -8808
rect 13900 -8888 13996 -8872
rect 13900 -8952 13916 -8888
rect 13980 -8952 13996 -8888
rect 13900 -8968 13996 -8952
rect 13900 -9032 13916 -8968
rect 13980 -9032 13996 -8968
rect 13900 -9048 13996 -9032
rect 13900 -9112 13916 -9048
rect 13980 -9112 13996 -9048
rect 13900 -9128 13996 -9112
rect 13900 -9192 13916 -9128
rect 13980 -9192 13996 -9128
rect 13900 -9208 13996 -9192
rect 13900 -9272 13916 -9208
rect 13980 -9272 13996 -9208
rect 13900 -9288 13996 -9272
rect 12488 -9388 12584 -9352
rect 13900 -9352 13916 -9288
rect 13980 -9352 13996 -9288
rect 14319 -8608 15041 -8599
rect 14319 -9312 14328 -8608
rect 15032 -9312 15041 -8608
rect 14319 -9321 15041 -9312
rect 15312 -8632 15328 -8568
rect 15392 -8632 15408 -8568
rect 16724 -8568 16820 -8532
rect 15312 -8648 15408 -8632
rect 15312 -8712 15328 -8648
rect 15392 -8712 15408 -8648
rect 15312 -8728 15408 -8712
rect 15312 -8792 15328 -8728
rect 15392 -8792 15408 -8728
rect 15312 -8808 15408 -8792
rect 15312 -8872 15328 -8808
rect 15392 -8872 15408 -8808
rect 15312 -8888 15408 -8872
rect 15312 -8952 15328 -8888
rect 15392 -8952 15408 -8888
rect 15312 -8968 15408 -8952
rect 15312 -9032 15328 -8968
rect 15392 -9032 15408 -8968
rect 15312 -9048 15408 -9032
rect 15312 -9112 15328 -9048
rect 15392 -9112 15408 -9048
rect 15312 -9128 15408 -9112
rect 15312 -9192 15328 -9128
rect 15392 -9192 15408 -9128
rect 15312 -9208 15408 -9192
rect 15312 -9272 15328 -9208
rect 15392 -9272 15408 -9208
rect 15312 -9288 15408 -9272
rect 13900 -9388 13996 -9352
rect 15312 -9352 15328 -9288
rect 15392 -9352 15408 -9288
rect 15731 -8608 16453 -8599
rect 15731 -9312 15740 -8608
rect 16444 -9312 16453 -8608
rect 15731 -9321 16453 -9312
rect 16724 -8632 16740 -8568
rect 16804 -8632 16820 -8568
rect 18136 -8568 18232 -8532
rect 16724 -8648 16820 -8632
rect 16724 -8712 16740 -8648
rect 16804 -8712 16820 -8648
rect 16724 -8728 16820 -8712
rect 16724 -8792 16740 -8728
rect 16804 -8792 16820 -8728
rect 16724 -8808 16820 -8792
rect 16724 -8872 16740 -8808
rect 16804 -8872 16820 -8808
rect 16724 -8888 16820 -8872
rect 16724 -8952 16740 -8888
rect 16804 -8952 16820 -8888
rect 16724 -8968 16820 -8952
rect 16724 -9032 16740 -8968
rect 16804 -9032 16820 -8968
rect 16724 -9048 16820 -9032
rect 16724 -9112 16740 -9048
rect 16804 -9112 16820 -9048
rect 16724 -9128 16820 -9112
rect 16724 -9192 16740 -9128
rect 16804 -9192 16820 -9128
rect 16724 -9208 16820 -9192
rect 16724 -9272 16740 -9208
rect 16804 -9272 16820 -9208
rect 16724 -9288 16820 -9272
rect 15312 -9388 15408 -9352
rect 16724 -9352 16740 -9288
rect 16804 -9352 16820 -9288
rect 17143 -8608 17865 -8599
rect 17143 -9312 17152 -8608
rect 17856 -9312 17865 -8608
rect 17143 -9321 17865 -9312
rect 18136 -8632 18152 -8568
rect 18216 -8632 18232 -8568
rect 19548 -8568 19644 -8532
rect 18136 -8648 18232 -8632
rect 18136 -8712 18152 -8648
rect 18216 -8712 18232 -8648
rect 18136 -8728 18232 -8712
rect 18136 -8792 18152 -8728
rect 18216 -8792 18232 -8728
rect 18136 -8808 18232 -8792
rect 18136 -8872 18152 -8808
rect 18216 -8872 18232 -8808
rect 18136 -8888 18232 -8872
rect 18136 -8952 18152 -8888
rect 18216 -8952 18232 -8888
rect 18136 -8968 18232 -8952
rect 18136 -9032 18152 -8968
rect 18216 -9032 18232 -8968
rect 18136 -9048 18232 -9032
rect 18136 -9112 18152 -9048
rect 18216 -9112 18232 -9048
rect 18136 -9128 18232 -9112
rect 18136 -9192 18152 -9128
rect 18216 -9192 18232 -9128
rect 18136 -9208 18232 -9192
rect 18136 -9272 18152 -9208
rect 18216 -9272 18232 -9208
rect 18136 -9288 18232 -9272
rect 16724 -9388 16820 -9352
rect 18136 -9352 18152 -9288
rect 18216 -9352 18232 -9288
rect 18555 -8608 19277 -8599
rect 18555 -9312 18564 -8608
rect 19268 -9312 19277 -8608
rect 18555 -9321 19277 -9312
rect 19548 -8632 19564 -8568
rect 19628 -8632 19644 -8568
rect 20960 -8568 21056 -8532
rect 19548 -8648 19644 -8632
rect 19548 -8712 19564 -8648
rect 19628 -8712 19644 -8648
rect 19548 -8728 19644 -8712
rect 19548 -8792 19564 -8728
rect 19628 -8792 19644 -8728
rect 19548 -8808 19644 -8792
rect 19548 -8872 19564 -8808
rect 19628 -8872 19644 -8808
rect 19548 -8888 19644 -8872
rect 19548 -8952 19564 -8888
rect 19628 -8952 19644 -8888
rect 19548 -8968 19644 -8952
rect 19548 -9032 19564 -8968
rect 19628 -9032 19644 -8968
rect 19548 -9048 19644 -9032
rect 19548 -9112 19564 -9048
rect 19628 -9112 19644 -9048
rect 19548 -9128 19644 -9112
rect 19548 -9192 19564 -9128
rect 19628 -9192 19644 -9128
rect 19548 -9208 19644 -9192
rect 19548 -9272 19564 -9208
rect 19628 -9272 19644 -9208
rect 19548 -9288 19644 -9272
rect 18136 -9388 18232 -9352
rect 19548 -9352 19564 -9288
rect 19628 -9352 19644 -9288
rect 19967 -8608 20689 -8599
rect 19967 -9312 19976 -8608
rect 20680 -9312 20689 -8608
rect 19967 -9321 20689 -9312
rect 20960 -8632 20976 -8568
rect 21040 -8632 21056 -8568
rect 22372 -8568 22468 -8532
rect 20960 -8648 21056 -8632
rect 20960 -8712 20976 -8648
rect 21040 -8712 21056 -8648
rect 20960 -8728 21056 -8712
rect 20960 -8792 20976 -8728
rect 21040 -8792 21056 -8728
rect 20960 -8808 21056 -8792
rect 20960 -8872 20976 -8808
rect 21040 -8872 21056 -8808
rect 20960 -8888 21056 -8872
rect 20960 -8952 20976 -8888
rect 21040 -8952 21056 -8888
rect 20960 -8968 21056 -8952
rect 20960 -9032 20976 -8968
rect 21040 -9032 21056 -8968
rect 20960 -9048 21056 -9032
rect 20960 -9112 20976 -9048
rect 21040 -9112 21056 -9048
rect 20960 -9128 21056 -9112
rect 20960 -9192 20976 -9128
rect 21040 -9192 21056 -9128
rect 20960 -9208 21056 -9192
rect 20960 -9272 20976 -9208
rect 21040 -9272 21056 -9208
rect 20960 -9288 21056 -9272
rect 19548 -9388 19644 -9352
rect 20960 -9352 20976 -9288
rect 21040 -9352 21056 -9288
rect 21379 -8608 22101 -8599
rect 21379 -9312 21388 -8608
rect 22092 -9312 22101 -8608
rect 21379 -9321 22101 -9312
rect 22372 -8632 22388 -8568
rect 22452 -8632 22468 -8568
rect 23784 -8568 23880 -8532
rect 22372 -8648 22468 -8632
rect 22372 -8712 22388 -8648
rect 22452 -8712 22468 -8648
rect 22372 -8728 22468 -8712
rect 22372 -8792 22388 -8728
rect 22452 -8792 22468 -8728
rect 22372 -8808 22468 -8792
rect 22372 -8872 22388 -8808
rect 22452 -8872 22468 -8808
rect 22372 -8888 22468 -8872
rect 22372 -8952 22388 -8888
rect 22452 -8952 22468 -8888
rect 22372 -8968 22468 -8952
rect 22372 -9032 22388 -8968
rect 22452 -9032 22468 -8968
rect 22372 -9048 22468 -9032
rect 22372 -9112 22388 -9048
rect 22452 -9112 22468 -9048
rect 22372 -9128 22468 -9112
rect 22372 -9192 22388 -9128
rect 22452 -9192 22468 -9128
rect 22372 -9208 22468 -9192
rect 22372 -9272 22388 -9208
rect 22452 -9272 22468 -9208
rect 22372 -9288 22468 -9272
rect 20960 -9388 21056 -9352
rect 22372 -9352 22388 -9288
rect 22452 -9352 22468 -9288
rect 22791 -8608 23513 -8599
rect 22791 -9312 22800 -8608
rect 23504 -9312 23513 -8608
rect 22791 -9321 23513 -9312
rect 23784 -8632 23800 -8568
rect 23864 -8632 23880 -8568
rect 23784 -8648 23880 -8632
rect 23784 -8712 23800 -8648
rect 23864 -8712 23880 -8648
rect 23784 -8728 23880 -8712
rect 23784 -8792 23800 -8728
rect 23864 -8792 23880 -8728
rect 23784 -8808 23880 -8792
rect 23784 -8872 23800 -8808
rect 23864 -8872 23880 -8808
rect 23784 -8888 23880 -8872
rect 23784 -8952 23800 -8888
rect 23864 -8952 23880 -8888
rect 23784 -8968 23880 -8952
rect 23784 -9032 23800 -8968
rect 23864 -9032 23880 -8968
rect 23784 -9048 23880 -9032
rect 23784 -9112 23800 -9048
rect 23864 -9112 23880 -9048
rect 23784 -9128 23880 -9112
rect 23784 -9192 23800 -9128
rect 23864 -9192 23880 -9128
rect 23784 -9208 23880 -9192
rect 23784 -9272 23800 -9208
rect 23864 -9272 23880 -9208
rect 23784 -9288 23880 -9272
rect 22372 -9388 22468 -9352
rect 23784 -9352 23800 -9288
rect 23864 -9352 23880 -9288
rect 23784 -9388 23880 -9352
rect -22812 -9688 -22716 -9652
rect -23805 -9728 -23083 -9719
rect -23805 -10432 -23796 -9728
rect -23092 -10432 -23083 -9728
rect -23805 -10441 -23083 -10432
rect -22812 -9752 -22796 -9688
rect -22732 -9752 -22716 -9688
rect -21400 -9688 -21304 -9652
rect -22812 -9768 -22716 -9752
rect -22812 -9832 -22796 -9768
rect -22732 -9832 -22716 -9768
rect -22812 -9848 -22716 -9832
rect -22812 -9912 -22796 -9848
rect -22732 -9912 -22716 -9848
rect -22812 -9928 -22716 -9912
rect -22812 -9992 -22796 -9928
rect -22732 -9992 -22716 -9928
rect -22812 -10008 -22716 -9992
rect -22812 -10072 -22796 -10008
rect -22732 -10072 -22716 -10008
rect -22812 -10088 -22716 -10072
rect -22812 -10152 -22796 -10088
rect -22732 -10152 -22716 -10088
rect -22812 -10168 -22716 -10152
rect -22812 -10232 -22796 -10168
rect -22732 -10232 -22716 -10168
rect -22812 -10248 -22716 -10232
rect -22812 -10312 -22796 -10248
rect -22732 -10312 -22716 -10248
rect -22812 -10328 -22716 -10312
rect -22812 -10392 -22796 -10328
rect -22732 -10392 -22716 -10328
rect -22812 -10408 -22716 -10392
rect -22812 -10472 -22796 -10408
rect -22732 -10472 -22716 -10408
rect -22393 -9728 -21671 -9719
rect -22393 -10432 -22384 -9728
rect -21680 -10432 -21671 -9728
rect -22393 -10441 -21671 -10432
rect -21400 -9752 -21384 -9688
rect -21320 -9752 -21304 -9688
rect -19988 -9688 -19892 -9652
rect -21400 -9768 -21304 -9752
rect -21400 -9832 -21384 -9768
rect -21320 -9832 -21304 -9768
rect -21400 -9848 -21304 -9832
rect -21400 -9912 -21384 -9848
rect -21320 -9912 -21304 -9848
rect -21400 -9928 -21304 -9912
rect -21400 -9992 -21384 -9928
rect -21320 -9992 -21304 -9928
rect -21400 -10008 -21304 -9992
rect -21400 -10072 -21384 -10008
rect -21320 -10072 -21304 -10008
rect -21400 -10088 -21304 -10072
rect -21400 -10152 -21384 -10088
rect -21320 -10152 -21304 -10088
rect -21400 -10168 -21304 -10152
rect -21400 -10232 -21384 -10168
rect -21320 -10232 -21304 -10168
rect -21400 -10248 -21304 -10232
rect -21400 -10312 -21384 -10248
rect -21320 -10312 -21304 -10248
rect -21400 -10328 -21304 -10312
rect -21400 -10392 -21384 -10328
rect -21320 -10392 -21304 -10328
rect -21400 -10408 -21304 -10392
rect -22812 -10508 -22716 -10472
rect -21400 -10472 -21384 -10408
rect -21320 -10472 -21304 -10408
rect -20981 -9728 -20259 -9719
rect -20981 -10432 -20972 -9728
rect -20268 -10432 -20259 -9728
rect -20981 -10441 -20259 -10432
rect -19988 -9752 -19972 -9688
rect -19908 -9752 -19892 -9688
rect -18576 -9688 -18480 -9652
rect -19988 -9768 -19892 -9752
rect -19988 -9832 -19972 -9768
rect -19908 -9832 -19892 -9768
rect -19988 -9848 -19892 -9832
rect -19988 -9912 -19972 -9848
rect -19908 -9912 -19892 -9848
rect -19988 -9928 -19892 -9912
rect -19988 -9992 -19972 -9928
rect -19908 -9992 -19892 -9928
rect -19988 -10008 -19892 -9992
rect -19988 -10072 -19972 -10008
rect -19908 -10072 -19892 -10008
rect -19988 -10088 -19892 -10072
rect -19988 -10152 -19972 -10088
rect -19908 -10152 -19892 -10088
rect -19988 -10168 -19892 -10152
rect -19988 -10232 -19972 -10168
rect -19908 -10232 -19892 -10168
rect -19988 -10248 -19892 -10232
rect -19988 -10312 -19972 -10248
rect -19908 -10312 -19892 -10248
rect -19988 -10328 -19892 -10312
rect -19988 -10392 -19972 -10328
rect -19908 -10392 -19892 -10328
rect -19988 -10408 -19892 -10392
rect -21400 -10508 -21304 -10472
rect -19988 -10472 -19972 -10408
rect -19908 -10472 -19892 -10408
rect -19569 -9728 -18847 -9719
rect -19569 -10432 -19560 -9728
rect -18856 -10432 -18847 -9728
rect -19569 -10441 -18847 -10432
rect -18576 -9752 -18560 -9688
rect -18496 -9752 -18480 -9688
rect -17164 -9688 -17068 -9652
rect -18576 -9768 -18480 -9752
rect -18576 -9832 -18560 -9768
rect -18496 -9832 -18480 -9768
rect -18576 -9848 -18480 -9832
rect -18576 -9912 -18560 -9848
rect -18496 -9912 -18480 -9848
rect -18576 -9928 -18480 -9912
rect -18576 -9992 -18560 -9928
rect -18496 -9992 -18480 -9928
rect -18576 -10008 -18480 -9992
rect -18576 -10072 -18560 -10008
rect -18496 -10072 -18480 -10008
rect -18576 -10088 -18480 -10072
rect -18576 -10152 -18560 -10088
rect -18496 -10152 -18480 -10088
rect -18576 -10168 -18480 -10152
rect -18576 -10232 -18560 -10168
rect -18496 -10232 -18480 -10168
rect -18576 -10248 -18480 -10232
rect -18576 -10312 -18560 -10248
rect -18496 -10312 -18480 -10248
rect -18576 -10328 -18480 -10312
rect -18576 -10392 -18560 -10328
rect -18496 -10392 -18480 -10328
rect -18576 -10408 -18480 -10392
rect -19988 -10508 -19892 -10472
rect -18576 -10472 -18560 -10408
rect -18496 -10472 -18480 -10408
rect -18157 -9728 -17435 -9719
rect -18157 -10432 -18148 -9728
rect -17444 -10432 -17435 -9728
rect -18157 -10441 -17435 -10432
rect -17164 -9752 -17148 -9688
rect -17084 -9752 -17068 -9688
rect -15752 -9688 -15656 -9652
rect -17164 -9768 -17068 -9752
rect -17164 -9832 -17148 -9768
rect -17084 -9832 -17068 -9768
rect -17164 -9848 -17068 -9832
rect -17164 -9912 -17148 -9848
rect -17084 -9912 -17068 -9848
rect -17164 -9928 -17068 -9912
rect -17164 -9992 -17148 -9928
rect -17084 -9992 -17068 -9928
rect -17164 -10008 -17068 -9992
rect -17164 -10072 -17148 -10008
rect -17084 -10072 -17068 -10008
rect -17164 -10088 -17068 -10072
rect -17164 -10152 -17148 -10088
rect -17084 -10152 -17068 -10088
rect -17164 -10168 -17068 -10152
rect -17164 -10232 -17148 -10168
rect -17084 -10232 -17068 -10168
rect -17164 -10248 -17068 -10232
rect -17164 -10312 -17148 -10248
rect -17084 -10312 -17068 -10248
rect -17164 -10328 -17068 -10312
rect -17164 -10392 -17148 -10328
rect -17084 -10392 -17068 -10328
rect -17164 -10408 -17068 -10392
rect -18576 -10508 -18480 -10472
rect -17164 -10472 -17148 -10408
rect -17084 -10472 -17068 -10408
rect -16745 -9728 -16023 -9719
rect -16745 -10432 -16736 -9728
rect -16032 -10432 -16023 -9728
rect -16745 -10441 -16023 -10432
rect -15752 -9752 -15736 -9688
rect -15672 -9752 -15656 -9688
rect -14340 -9688 -14244 -9652
rect -15752 -9768 -15656 -9752
rect -15752 -9832 -15736 -9768
rect -15672 -9832 -15656 -9768
rect -15752 -9848 -15656 -9832
rect -15752 -9912 -15736 -9848
rect -15672 -9912 -15656 -9848
rect -15752 -9928 -15656 -9912
rect -15752 -9992 -15736 -9928
rect -15672 -9992 -15656 -9928
rect -15752 -10008 -15656 -9992
rect -15752 -10072 -15736 -10008
rect -15672 -10072 -15656 -10008
rect -15752 -10088 -15656 -10072
rect -15752 -10152 -15736 -10088
rect -15672 -10152 -15656 -10088
rect -15752 -10168 -15656 -10152
rect -15752 -10232 -15736 -10168
rect -15672 -10232 -15656 -10168
rect -15752 -10248 -15656 -10232
rect -15752 -10312 -15736 -10248
rect -15672 -10312 -15656 -10248
rect -15752 -10328 -15656 -10312
rect -15752 -10392 -15736 -10328
rect -15672 -10392 -15656 -10328
rect -15752 -10408 -15656 -10392
rect -17164 -10508 -17068 -10472
rect -15752 -10472 -15736 -10408
rect -15672 -10472 -15656 -10408
rect -15333 -9728 -14611 -9719
rect -15333 -10432 -15324 -9728
rect -14620 -10432 -14611 -9728
rect -15333 -10441 -14611 -10432
rect -14340 -9752 -14324 -9688
rect -14260 -9752 -14244 -9688
rect -12928 -9688 -12832 -9652
rect -14340 -9768 -14244 -9752
rect -14340 -9832 -14324 -9768
rect -14260 -9832 -14244 -9768
rect -14340 -9848 -14244 -9832
rect -14340 -9912 -14324 -9848
rect -14260 -9912 -14244 -9848
rect -14340 -9928 -14244 -9912
rect -14340 -9992 -14324 -9928
rect -14260 -9992 -14244 -9928
rect -14340 -10008 -14244 -9992
rect -14340 -10072 -14324 -10008
rect -14260 -10072 -14244 -10008
rect -14340 -10088 -14244 -10072
rect -14340 -10152 -14324 -10088
rect -14260 -10152 -14244 -10088
rect -14340 -10168 -14244 -10152
rect -14340 -10232 -14324 -10168
rect -14260 -10232 -14244 -10168
rect -14340 -10248 -14244 -10232
rect -14340 -10312 -14324 -10248
rect -14260 -10312 -14244 -10248
rect -14340 -10328 -14244 -10312
rect -14340 -10392 -14324 -10328
rect -14260 -10392 -14244 -10328
rect -14340 -10408 -14244 -10392
rect -15752 -10508 -15656 -10472
rect -14340 -10472 -14324 -10408
rect -14260 -10472 -14244 -10408
rect -13921 -9728 -13199 -9719
rect -13921 -10432 -13912 -9728
rect -13208 -10432 -13199 -9728
rect -13921 -10441 -13199 -10432
rect -12928 -9752 -12912 -9688
rect -12848 -9752 -12832 -9688
rect -11516 -9688 -11420 -9652
rect -12928 -9768 -12832 -9752
rect -12928 -9832 -12912 -9768
rect -12848 -9832 -12832 -9768
rect -12928 -9848 -12832 -9832
rect -12928 -9912 -12912 -9848
rect -12848 -9912 -12832 -9848
rect -12928 -9928 -12832 -9912
rect -12928 -9992 -12912 -9928
rect -12848 -9992 -12832 -9928
rect -12928 -10008 -12832 -9992
rect -12928 -10072 -12912 -10008
rect -12848 -10072 -12832 -10008
rect -12928 -10088 -12832 -10072
rect -12928 -10152 -12912 -10088
rect -12848 -10152 -12832 -10088
rect -12928 -10168 -12832 -10152
rect -12928 -10232 -12912 -10168
rect -12848 -10232 -12832 -10168
rect -12928 -10248 -12832 -10232
rect -12928 -10312 -12912 -10248
rect -12848 -10312 -12832 -10248
rect -12928 -10328 -12832 -10312
rect -12928 -10392 -12912 -10328
rect -12848 -10392 -12832 -10328
rect -12928 -10408 -12832 -10392
rect -14340 -10508 -14244 -10472
rect -12928 -10472 -12912 -10408
rect -12848 -10472 -12832 -10408
rect -12509 -9728 -11787 -9719
rect -12509 -10432 -12500 -9728
rect -11796 -10432 -11787 -9728
rect -12509 -10441 -11787 -10432
rect -11516 -9752 -11500 -9688
rect -11436 -9752 -11420 -9688
rect -10104 -9688 -10008 -9652
rect -11516 -9768 -11420 -9752
rect -11516 -9832 -11500 -9768
rect -11436 -9832 -11420 -9768
rect -11516 -9848 -11420 -9832
rect -11516 -9912 -11500 -9848
rect -11436 -9912 -11420 -9848
rect -11516 -9928 -11420 -9912
rect -11516 -9992 -11500 -9928
rect -11436 -9992 -11420 -9928
rect -11516 -10008 -11420 -9992
rect -11516 -10072 -11500 -10008
rect -11436 -10072 -11420 -10008
rect -11516 -10088 -11420 -10072
rect -11516 -10152 -11500 -10088
rect -11436 -10152 -11420 -10088
rect -11516 -10168 -11420 -10152
rect -11516 -10232 -11500 -10168
rect -11436 -10232 -11420 -10168
rect -11516 -10248 -11420 -10232
rect -11516 -10312 -11500 -10248
rect -11436 -10312 -11420 -10248
rect -11516 -10328 -11420 -10312
rect -11516 -10392 -11500 -10328
rect -11436 -10392 -11420 -10328
rect -11516 -10408 -11420 -10392
rect -12928 -10508 -12832 -10472
rect -11516 -10472 -11500 -10408
rect -11436 -10472 -11420 -10408
rect -11097 -9728 -10375 -9719
rect -11097 -10432 -11088 -9728
rect -10384 -10432 -10375 -9728
rect -11097 -10441 -10375 -10432
rect -10104 -9752 -10088 -9688
rect -10024 -9752 -10008 -9688
rect -8692 -9688 -8596 -9652
rect -10104 -9768 -10008 -9752
rect -10104 -9832 -10088 -9768
rect -10024 -9832 -10008 -9768
rect -10104 -9848 -10008 -9832
rect -10104 -9912 -10088 -9848
rect -10024 -9912 -10008 -9848
rect -10104 -9928 -10008 -9912
rect -10104 -9992 -10088 -9928
rect -10024 -9992 -10008 -9928
rect -10104 -10008 -10008 -9992
rect -10104 -10072 -10088 -10008
rect -10024 -10072 -10008 -10008
rect -10104 -10088 -10008 -10072
rect -10104 -10152 -10088 -10088
rect -10024 -10152 -10008 -10088
rect -10104 -10168 -10008 -10152
rect -10104 -10232 -10088 -10168
rect -10024 -10232 -10008 -10168
rect -10104 -10248 -10008 -10232
rect -10104 -10312 -10088 -10248
rect -10024 -10312 -10008 -10248
rect -10104 -10328 -10008 -10312
rect -10104 -10392 -10088 -10328
rect -10024 -10392 -10008 -10328
rect -10104 -10408 -10008 -10392
rect -11516 -10508 -11420 -10472
rect -10104 -10472 -10088 -10408
rect -10024 -10472 -10008 -10408
rect -9685 -9728 -8963 -9719
rect -9685 -10432 -9676 -9728
rect -8972 -10432 -8963 -9728
rect -9685 -10441 -8963 -10432
rect -8692 -9752 -8676 -9688
rect -8612 -9752 -8596 -9688
rect -7280 -9688 -7184 -9652
rect -8692 -9768 -8596 -9752
rect -8692 -9832 -8676 -9768
rect -8612 -9832 -8596 -9768
rect -8692 -9848 -8596 -9832
rect -8692 -9912 -8676 -9848
rect -8612 -9912 -8596 -9848
rect -8692 -9928 -8596 -9912
rect -8692 -9992 -8676 -9928
rect -8612 -9992 -8596 -9928
rect -8692 -10008 -8596 -9992
rect -8692 -10072 -8676 -10008
rect -8612 -10072 -8596 -10008
rect -8692 -10088 -8596 -10072
rect -8692 -10152 -8676 -10088
rect -8612 -10152 -8596 -10088
rect -8692 -10168 -8596 -10152
rect -8692 -10232 -8676 -10168
rect -8612 -10232 -8596 -10168
rect -8692 -10248 -8596 -10232
rect -8692 -10312 -8676 -10248
rect -8612 -10312 -8596 -10248
rect -8692 -10328 -8596 -10312
rect -8692 -10392 -8676 -10328
rect -8612 -10392 -8596 -10328
rect -8692 -10408 -8596 -10392
rect -10104 -10508 -10008 -10472
rect -8692 -10472 -8676 -10408
rect -8612 -10472 -8596 -10408
rect -8273 -9728 -7551 -9719
rect -8273 -10432 -8264 -9728
rect -7560 -10432 -7551 -9728
rect -8273 -10441 -7551 -10432
rect -7280 -9752 -7264 -9688
rect -7200 -9752 -7184 -9688
rect -5868 -9688 -5772 -9652
rect -7280 -9768 -7184 -9752
rect -7280 -9832 -7264 -9768
rect -7200 -9832 -7184 -9768
rect -7280 -9848 -7184 -9832
rect -7280 -9912 -7264 -9848
rect -7200 -9912 -7184 -9848
rect -7280 -9928 -7184 -9912
rect -7280 -9992 -7264 -9928
rect -7200 -9992 -7184 -9928
rect -7280 -10008 -7184 -9992
rect -7280 -10072 -7264 -10008
rect -7200 -10072 -7184 -10008
rect -7280 -10088 -7184 -10072
rect -7280 -10152 -7264 -10088
rect -7200 -10152 -7184 -10088
rect -7280 -10168 -7184 -10152
rect -7280 -10232 -7264 -10168
rect -7200 -10232 -7184 -10168
rect -7280 -10248 -7184 -10232
rect -7280 -10312 -7264 -10248
rect -7200 -10312 -7184 -10248
rect -7280 -10328 -7184 -10312
rect -7280 -10392 -7264 -10328
rect -7200 -10392 -7184 -10328
rect -7280 -10408 -7184 -10392
rect -8692 -10508 -8596 -10472
rect -7280 -10472 -7264 -10408
rect -7200 -10472 -7184 -10408
rect -6861 -9728 -6139 -9719
rect -6861 -10432 -6852 -9728
rect -6148 -10432 -6139 -9728
rect -6861 -10441 -6139 -10432
rect -5868 -9752 -5852 -9688
rect -5788 -9752 -5772 -9688
rect -4456 -9688 -4360 -9652
rect -5868 -9768 -5772 -9752
rect -5868 -9832 -5852 -9768
rect -5788 -9832 -5772 -9768
rect -5868 -9848 -5772 -9832
rect -5868 -9912 -5852 -9848
rect -5788 -9912 -5772 -9848
rect -5868 -9928 -5772 -9912
rect -5868 -9992 -5852 -9928
rect -5788 -9992 -5772 -9928
rect -5868 -10008 -5772 -9992
rect -5868 -10072 -5852 -10008
rect -5788 -10072 -5772 -10008
rect -5868 -10088 -5772 -10072
rect -5868 -10152 -5852 -10088
rect -5788 -10152 -5772 -10088
rect -5868 -10168 -5772 -10152
rect -5868 -10232 -5852 -10168
rect -5788 -10232 -5772 -10168
rect -5868 -10248 -5772 -10232
rect -5868 -10312 -5852 -10248
rect -5788 -10312 -5772 -10248
rect -5868 -10328 -5772 -10312
rect -5868 -10392 -5852 -10328
rect -5788 -10392 -5772 -10328
rect -5868 -10408 -5772 -10392
rect -7280 -10508 -7184 -10472
rect -5868 -10472 -5852 -10408
rect -5788 -10472 -5772 -10408
rect -5449 -9728 -4727 -9719
rect -5449 -10432 -5440 -9728
rect -4736 -10432 -4727 -9728
rect -5449 -10441 -4727 -10432
rect -4456 -9752 -4440 -9688
rect -4376 -9752 -4360 -9688
rect -3044 -9688 -2948 -9652
rect -4456 -9768 -4360 -9752
rect -4456 -9832 -4440 -9768
rect -4376 -9832 -4360 -9768
rect -4456 -9848 -4360 -9832
rect -4456 -9912 -4440 -9848
rect -4376 -9912 -4360 -9848
rect -4456 -9928 -4360 -9912
rect -4456 -9992 -4440 -9928
rect -4376 -9992 -4360 -9928
rect -4456 -10008 -4360 -9992
rect -4456 -10072 -4440 -10008
rect -4376 -10072 -4360 -10008
rect -4456 -10088 -4360 -10072
rect -4456 -10152 -4440 -10088
rect -4376 -10152 -4360 -10088
rect -4456 -10168 -4360 -10152
rect -4456 -10232 -4440 -10168
rect -4376 -10232 -4360 -10168
rect -4456 -10248 -4360 -10232
rect -4456 -10312 -4440 -10248
rect -4376 -10312 -4360 -10248
rect -4456 -10328 -4360 -10312
rect -4456 -10392 -4440 -10328
rect -4376 -10392 -4360 -10328
rect -4456 -10408 -4360 -10392
rect -5868 -10508 -5772 -10472
rect -4456 -10472 -4440 -10408
rect -4376 -10472 -4360 -10408
rect -4037 -9728 -3315 -9719
rect -4037 -10432 -4028 -9728
rect -3324 -10432 -3315 -9728
rect -4037 -10441 -3315 -10432
rect -3044 -9752 -3028 -9688
rect -2964 -9752 -2948 -9688
rect -1632 -9688 -1536 -9652
rect -3044 -9768 -2948 -9752
rect -3044 -9832 -3028 -9768
rect -2964 -9832 -2948 -9768
rect -3044 -9848 -2948 -9832
rect -3044 -9912 -3028 -9848
rect -2964 -9912 -2948 -9848
rect -3044 -9928 -2948 -9912
rect -3044 -9992 -3028 -9928
rect -2964 -9992 -2948 -9928
rect -3044 -10008 -2948 -9992
rect -3044 -10072 -3028 -10008
rect -2964 -10072 -2948 -10008
rect -3044 -10088 -2948 -10072
rect -3044 -10152 -3028 -10088
rect -2964 -10152 -2948 -10088
rect -3044 -10168 -2948 -10152
rect -3044 -10232 -3028 -10168
rect -2964 -10232 -2948 -10168
rect -3044 -10248 -2948 -10232
rect -3044 -10312 -3028 -10248
rect -2964 -10312 -2948 -10248
rect -3044 -10328 -2948 -10312
rect -3044 -10392 -3028 -10328
rect -2964 -10392 -2948 -10328
rect -3044 -10408 -2948 -10392
rect -4456 -10508 -4360 -10472
rect -3044 -10472 -3028 -10408
rect -2964 -10472 -2948 -10408
rect -2625 -9728 -1903 -9719
rect -2625 -10432 -2616 -9728
rect -1912 -10432 -1903 -9728
rect -2625 -10441 -1903 -10432
rect -1632 -9752 -1616 -9688
rect -1552 -9752 -1536 -9688
rect -220 -9688 -124 -9652
rect -1632 -9768 -1536 -9752
rect -1632 -9832 -1616 -9768
rect -1552 -9832 -1536 -9768
rect -1632 -9848 -1536 -9832
rect -1632 -9912 -1616 -9848
rect -1552 -9912 -1536 -9848
rect -1632 -9928 -1536 -9912
rect -1632 -9992 -1616 -9928
rect -1552 -9992 -1536 -9928
rect -1632 -10008 -1536 -9992
rect -1632 -10072 -1616 -10008
rect -1552 -10072 -1536 -10008
rect -1632 -10088 -1536 -10072
rect -1632 -10152 -1616 -10088
rect -1552 -10152 -1536 -10088
rect -1632 -10168 -1536 -10152
rect -1632 -10232 -1616 -10168
rect -1552 -10232 -1536 -10168
rect -1632 -10248 -1536 -10232
rect -1632 -10312 -1616 -10248
rect -1552 -10312 -1536 -10248
rect -1632 -10328 -1536 -10312
rect -1632 -10392 -1616 -10328
rect -1552 -10392 -1536 -10328
rect -1632 -10408 -1536 -10392
rect -3044 -10508 -2948 -10472
rect -1632 -10472 -1616 -10408
rect -1552 -10472 -1536 -10408
rect -1213 -9728 -491 -9719
rect -1213 -10432 -1204 -9728
rect -500 -10432 -491 -9728
rect -1213 -10441 -491 -10432
rect -220 -9752 -204 -9688
rect -140 -9752 -124 -9688
rect 1192 -9688 1288 -9652
rect -220 -9768 -124 -9752
rect -220 -9832 -204 -9768
rect -140 -9832 -124 -9768
rect -220 -9848 -124 -9832
rect -220 -9912 -204 -9848
rect -140 -9912 -124 -9848
rect -220 -9928 -124 -9912
rect -220 -9992 -204 -9928
rect -140 -9992 -124 -9928
rect -220 -10008 -124 -9992
rect -220 -10072 -204 -10008
rect -140 -10072 -124 -10008
rect -220 -10088 -124 -10072
rect -220 -10152 -204 -10088
rect -140 -10152 -124 -10088
rect -220 -10168 -124 -10152
rect -220 -10232 -204 -10168
rect -140 -10232 -124 -10168
rect -220 -10248 -124 -10232
rect -220 -10312 -204 -10248
rect -140 -10312 -124 -10248
rect -220 -10328 -124 -10312
rect -220 -10392 -204 -10328
rect -140 -10392 -124 -10328
rect -220 -10408 -124 -10392
rect -1632 -10508 -1536 -10472
rect -220 -10472 -204 -10408
rect -140 -10472 -124 -10408
rect 199 -9728 921 -9719
rect 199 -10432 208 -9728
rect 912 -10432 921 -9728
rect 199 -10441 921 -10432
rect 1192 -9752 1208 -9688
rect 1272 -9752 1288 -9688
rect 2604 -9688 2700 -9652
rect 1192 -9768 1288 -9752
rect 1192 -9832 1208 -9768
rect 1272 -9832 1288 -9768
rect 1192 -9848 1288 -9832
rect 1192 -9912 1208 -9848
rect 1272 -9912 1288 -9848
rect 1192 -9928 1288 -9912
rect 1192 -9992 1208 -9928
rect 1272 -9992 1288 -9928
rect 1192 -10008 1288 -9992
rect 1192 -10072 1208 -10008
rect 1272 -10072 1288 -10008
rect 1192 -10088 1288 -10072
rect 1192 -10152 1208 -10088
rect 1272 -10152 1288 -10088
rect 1192 -10168 1288 -10152
rect 1192 -10232 1208 -10168
rect 1272 -10232 1288 -10168
rect 1192 -10248 1288 -10232
rect 1192 -10312 1208 -10248
rect 1272 -10312 1288 -10248
rect 1192 -10328 1288 -10312
rect 1192 -10392 1208 -10328
rect 1272 -10392 1288 -10328
rect 1192 -10408 1288 -10392
rect -220 -10508 -124 -10472
rect 1192 -10472 1208 -10408
rect 1272 -10472 1288 -10408
rect 1611 -9728 2333 -9719
rect 1611 -10432 1620 -9728
rect 2324 -10432 2333 -9728
rect 1611 -10441 2333 -10432
rect 2604 -9752 2620 -9688
rect 2684 -9752 2700 -9688
rect 4016 -9688 4112 -9652
rect 2604 -9768 2700 -9752
rect 2604 -9832 2620 -9768
rect 2684 -9832 2700 -9768
rect 2604 -9848 2700 -9832
rect 2604 -9912 2620 -9848
rect 2684 -9912 2700 -9848
rect 2604 -9928 2700 -9912
rect 2604 -9992 2620 -9928
rect 2684 -9992 2700 -9928
rect 2604 -10008 2700 -9992
rect 2604 -10072 2620 -10008
rect 2684 -10072 2700 -10008
rect 2604 -10088 2700 -10072
rect 2604 -10152 2620 -10088
rect 2684 -10152 2700 -10088
rect 2604 -10168 2700 -10152
rect 2604 -10232 2620 -10168
rect 2684 -10232 2700 -10168
rect 2604 -10248 2700 -10232
rect 2604 -10312 2620 -10248
rect 2684 -10312 2700 -10248
rect 2604 -10328 2700 -10312
rect 2604 -10392 2620 -10328
rect 2684 -10392 2700 -10328
rect 2604 -10408 2700 -10392
rect 1192 -10508 1288 -10472
rect 2604 -10472 2620 -10408
rect 2684 -10472 2700 -10408
rect 3023 -9728 3745 -9719
rect 3023 -10432 3032 -9728
rect 3736 -10432 3745 -9728
rect 3023 -10441 3745 -10432
rect 4016 -9752 4032 -9688
rect 4096 -9752 4112 -9688
rect 5428 -9688 5524 -9652
rect 4016 -9768 4112 -9752
rect 4016 -9832 4032 -9768
rect 4096 -9832 4112 -9768
rect 4016 -9848 4112 -9832
rect 4016 -9912 4032 -9848
rect 4096 -9912 4112 -9848
rect 4016 -9928 4112 -9912
rect 4016 -9992 4032 -9928
rect 4096 -9992 4112 -9928
rect 4016 -10008 4112 -9992
rect 4016 -10072 4032 -10008
rect 4096 -10072 4112 -10008
rect 4016 -10088 4112 -10072
rect 4016 -10152 4032 -10088
rect 4096 -10152 4112 -10088
rect 4016 -10168 4112 -10152
rect 4016 -10232 4032 -10168
rect 4096 -10232 4112 -10168
rect 4016 -10248 4112 -10232
rect 4016 -10312 4032 -10248
rect 4096 -10312 4112 -10248
rect 4016 -10328 4112 -10312
rect 4016 -10392 4032 -10328
rect 4096 -10392 4112 -10328
rect 4016 -10408 4112 -10392
rect 2604 -10508 2700 -10472
rect 4016 -10472 4032 -10408
rect 4096 -10472 4112 -10408
rect 4435 -9728 5157 -9719
rect 4435 -10432 4444 -9728
rect 5148 -10432 5157 -9728
rect 4435 -10441 5157 -10432
rect 5428 -9752 5444 -9688
rect 5508 -9752 5524 -9688
rect 6840 -9688 6936 -9652
rect 5428 -9768 5524 -9752
rect 5428 -9832 5444 -9768
rect 5508 -9832 5524 -9768
rect 5428 -9848 5524 -9832
rect 5428 -9912 5444 -9848
rect 5508 -9912 5524 -9848
rect 5428 -9928 5524 -9912
rect 5428 -9992 5444 -9928
rect 5508 -9992 5524 -9928
rect 5428 -10008 5524 -9992
rect 5428 -10072 5444 -10008
rect 5508 -10072 5524 -10008
rect 5428 -10088 5524 -10072
rect 5428 -10152 5444 -10088
rect 5508 -10152 5524 -10088
rect 5428 -10168 5524 -10152
rect 5428 -10232 5444 -10168
rect 5508 -10232 5524 -10168
rect 5428 -10248 5524 -10232
rect 5428 -10312 5444 -10248
rect 5508 -10312 5524 -10248
rect 5428 -10328 5524 -10312
rect 5428 -10392 5444 -10328
rect 5508 -10392 5524 -10328
rect 5428 -10408 5524 -10392
rect 4016 -10508 4112 -10472
rect 5428 -10472 5444 -10408
rect 5508 -10472 5524 -10408
rect 5847 -9728 6569 -9719
rect 5847 -10432 5856 -9728
rect 6560 -10432 6569 -9728
rect 5847 -10441 6569 -10432
rect 6840 -9752 6856 -9688
rect 6920 -9752 6936 -9688
rect 8252 -9688 8348 -9652
rect 6840 -9768 6936 -9752
rect 6840 -9832 6856 -9768
rect 6920 -9832 6936 -9768
rect 6840 -9848 6936 -9832
rect 6840 -9912 6856 -9848
rect 6920 -9912 6936 -9848
rect 6840 -9928 6936 -9912
rect 6840 -9992 6856 -9928
rect 6920 -9992 6936 -9928
rect 6840 -10008 6936 -9992
rect 6840 -10072 6856 -10008
rect 6920 -10072 6936 -10008
rect 6840 -10088 6936 -10072
rect 6840 -10152 6856 -10088
rect 6920 -10152 6936 -10088
rect 6840 -10168 6936 -10152
rect 6840 -10232 6856 -10168
rect 6920 -10232 6936 -10168
rect 6840 -10248 6936 -10232
rect 6840 -10312 6856 -10248
rect 6920 -10312 6936 -10248
rect 6840 -10328 6936 -10312
rect 6840 -10392 6856 -10328
rect 6920 -10392 6936 -10328
rect 6840 -10408 6936 -10392
rect 5428 -10508 5524 -10472
rect 6840 -10472 6856 -10408
rect 6920 -10472 6936 -10408
rect 7259 -9728 7981 -9719
rect 7259 -10432 7268 -9728
rect 7972 -10432 7981 -9728
rect 7259 -10441 7981 -10432
rect 8252 -9752 8268 -9688
rect 8332 -9752 8348 -9688
rect 9664 -9688 9760 -9652
rect 8252 -9768 8348 -9752
rect 8252 -9832 8268 -9768
rect 8332 -9832 8348 -9768
rect 8252 -9848 8348 -9832
rect 8252 -9912 8268 -9848
rect 8332 -9912 8348 -9848
rect 8252 -9928 8348 -9912
rect 8252 -9992 8268 -9928
rect 8332 -9992 8348 -9928
rect 8252 -10008 8348 -9992
rect 8252 -10072 8268 -10008
rect 8332 -10072 8348 -10008
rect 8252 -10088 8348 -10072
rect 8252 -10152 8268 -10088
rect 8332 -10152 8348 -10088
rect 8252 -10168 8348 -10152
rect 8252 -10232 8268 -10168
rect 8332 -10232 8348 -10168
rect 8252 -10248 8348 -10232
rect 8252 -10312 8268 -10248
rect 8332 -10312 8348 -10248
rect 8252 -10328 8348 -10312
rect 8252 -10392 8268 -10328
rect 8332 -10392 8348 -10328
rect 8252 -10408 8348 -10392
rect 6840 -10508 6936 -10472
rect 8252 -10472 8268 -10408
rect 8332 -10472 8348 -10408
rect 8671 -9728 9393 -9719
rect 8671 -10432 8680 -9728
rect 9384 -10432 9393 -9728
rect 8671 -10441 9393 -10432
rect 9664 -9752 9680 -9688
rect 9744 -9752 9760 -9688
rect 11076 -9688 11172 -9652
rect 9664 -9768 9760 -9752
rect 9664 -9832 9680 -9768
rect 9744 -9832 9760 -9768
rect 9664 -9848 9760 -9832
rect 9664 -9912 9680 -9848
rect 9744 -9912 9760 -9848
rect 9664 -9928 9760 -9912
rect 9664 -9992 9680 -9928
rect 9744 -9992 9760 -9928
rect 9664 -10008 9760 -9992
rect 9664 -10072 9680 -10008
rect 9744 -10072 9760 -10008
rect 9664 -10088 9760 -10072
rect 9664 -10152 9680 -10088
rect 9744 -10152 9760 -10088
rect 9664 -10168 9760 -10152
rect 9664 -10232 9680 -10168
rect 9744 -10232 9760 -10168
rect 9664 -10248 9760 -10232
rect 9664 -10312 9680 -10248
rect 9744 -10312 9760 -10248
rect 9664 -10328 9760 -10312
rect 9664 -10392 9680 -10328
rect 9744 -10392 9760 -10328
rect 9664 -10408 9760 -10392
rect 8252 -10508 8348 -10472
rect 9664 -10472 9680 -10408
rect 9744 -10472 9760 -10408
rect 10083 -9728 10805 -9719
rect 10083 -10432 10092 -9728
rect 10796 -10432 10805 -9728
rect 10083 -10441 10805 -10432
rect 11076 -9752 11092 -9688
rect 11156 -9752 11172 -9688
rect 12488 -9688 12584 -9652
rect 11076 -9768 11172 -9752
rect 11076 -9832 11092 -9768
rect 11156 -9832 11172 -9768
rect 11076 -9848 11172 -9832
rect 11076 -9912 11092 -9848
rect 11156 -9912 11172 -9848
rect 11076 -9928 11172 -9912
rect 11076 -9992 11092 -9928
rect 11156 -9992 11172 -9928
rect 11076 -10008 11172 -9992
rect 11076 -10072 11092 -10008
rect 11156 -10072 11172 -10008
rect 11076 -10088 11172 -10072
rect 11076 -10152 11092 -10088
rect 11156 -10152 11172 -10088
rect 11076 -10168 11172 -10152
rect 11076 -10232 11092 -10168
rect 11156 -10232 11172 -10168
rect 11076 -10248 11172 -10232
rect 11076 -10312 11092 -10248
rect 11156 -10312 11172 -10248
rect 11076 -10328 11172 -10312
rect 11076 -10392 11092 -10328
rect 11156 -10392 11172 -10328
rect 11076 -10408 11172 -10392
rect 9664 -10508 9760 -10472
rect 11076 -10472 11092 -10408
rect 11156 -10472 11172 -10408
rect 11495 -9728 12217 -9719
rect 11495 -10432 11504 -9728
rect 12208 -10432 12217 -9728
rect 11495 -10441 12217 -10432
rect 12488 -9752 12504 -9688
rect 12568 -9752 12584 -9688
rect 13900 -9688 13996 -9652
rect 12488 -9768 12584 -9752
rect 12488 -9832 12504 -9768
rect 12568 -9832 12584 -9768
rect 12488 -9848 12584 -9832
rect 12488 -9912 12504 -9848
rect 12568 -9912 12584 -9848
rect 12488 -9928 12584 -9912
rect 12488 -9992 12504 -9928
rect 12568 -9992 12584 -9928
rect 12488 -10008 12584 -9992
rect 12488 -10072 12504 -10008
rect 12568 -10072 12584 -10008
rect 12488 -10088 12584 -10072
rect 12488 -10152 12504 -10088
rect 12568 -10152 12584 -10088
rect 12488 -10168 12584 -10152
rect 12488 -10232 12504 -10168
rect 12568 -10232 12584 -10168
rect 12488 -10248 12584 -10232
rect 12488 -10312 12504 -10248
rect 12568 -10312 12584 -10248
rect 12488 -10328 12584 -10312
rect 12488 -10392 12504 -10328
rect 12568 -10392 12584 -10328
rect 12488 -10408 12584 -10392
rect 11076 -10508 11172 -10472
rect 12488 -10472 12504 -10408
rect 12568 -10472 12584 -10408
rect 12907 -9728 13629 -9719
rect 12907 -10432 12916 -9728
rect 13620 -10432 13629 -9728
rect 12907 -10441 13629 -10432
rect 13900 -9752 13916 -9688
rect 13980 -9752 13996 -9688
rect 15312 -9688 15408 -9652
rect 13900 -9768 13996 -9752
rect 13900 -9832 13916 -9768
rect 13980 -9832 13996 -9768
rect 13900 -9848 13996 -9832
rect 13900 -9912 13916 -9848
rect 13980 -9912 13996 -9848
rect 13900 -9928 13996 -9912
rect 13900 -9992 13916 -9928
rect 13980 -9992 13996 -9928
rect 13900 -10008 13996 -9992
rect 13900 -10072 13916 -10008
rect 13980 -10072 13996 -10008
rect 13900 -10088 13996 -10072
rect 13900 -10152 13916 -10088
rect 13980 -10152 13996 -10088
rect 13900 -10168 13996 -10152
rect 13900 -10232 13916 -10168
rect 13980 -10232 13996 -10168
rect 13900 -10248 13996 -10232
rect 13900 -10312 13916 -10248
rect 13980 -10312 13996 -10248
rect 13900 -10328 13996 -10312
rect 13900 -10392 13916 -10328
rect 13980 -10392 13996 -10328
rect 13900 -10408 13996 -10392
rect 12488 -10508 12584 -10472
rect 13900 -10472 13916 -10408
rect 13980 -10472 13996 -10408
rect 14319 -9728 15041 -9719
rect 14319 -10432 14328 -9728
rect 15032 -10432 15041 -9728
rect 14319 -10441 15041 -10432
rect 15312 -9752 15328 -9688
rect 15392 -9752 15408 -9688
rect 16724 -9688 16820 -9652
rect 15312 -9768 15408 -9752
rect 15312 -9832 15328 -9768
rect 15392 -9832 15408 -9768
rect 15312 -9848 15408 -9832
rect 15312 -9912 15328 -9848
rect 15392 -9912 15408 -9848
rect 15312 -9928 15408 -9912
rect 15312 -9992 15328 -9928
rect 15392 -9992 15408 -9928
rect 15312 -10008 15408 -9992
rect 15312 -10072 15328 -10008
rect 15392 -10072 15408 -10008
rect 15312 -10088 15408 -10072
rect 15312 -10152 15328 -10088
rect 15392 -10152 15408 -10088
rect 15312 -10168 15408 -10152
rect 15312 -10232 15328 -10168
rect 15392 -10232 15408 -10168
rect 15312 -10248 15408 -10232
rect 15312 -10312 15328 -10248
rect 15392 -10312 15408 -10248
rect 15312 -10328 15408 -10312
rect 15312 -10392 15328 -10328
rect 15392 -10392 15408 -10328
rect 15312 -10408 15408 -10392
rect 13900 -10508 13996 -10472
rect 15312 -10472 15328 -10408
rect 15392 -10472 15408 -10408
rect 15731 -9728 16453 -9719
rect 15731 -10432 15740 -9728
rect 16444 -10432 16453 -9728
rect 15731 -10441 16453 -10432
rect 16724 -9752 16740 -9688
rect 16804 -9752 16820 -9688
rect 18136 -9688 18232 -9652
rect 16724 -9768 16820 -9752
rect 16724 -9832 16740 -9768
rect 16804 -9832 16820 -9768
rect 16724 -9848 16820 -9832
rect 16724 -9912 16740 -9848
rect 16804 -9912 16820 -9848
rect 16724 -9928 16820 -9912
rect 16724 -9992 16740 -9928
rect 16804 -9992 16820 -9928
rect 16724 -10008 16820 -9992
rect 16724 -10072 16740 -10008
rect 16804 -10072 16820 -10008
rect 16724 -10088 16820 -10072
rect 16724 -10152 16740 -10088
rect 16804 -10152 16820 -10088
rect 16724 -10168 16820 -10152
rect 16724 -10232 16740 -10168
rect 16804 -10232 16820 -10168
rect 16724 -10248 16820 -10232
rect 16724 -10312 16740 -10248
rect 16804 -10312 16820 -10248
rect 16724 -10328 16820 -10312
rect 16724 -10392 16740 -10328
rect 16804 -10392 16820 -10328
rect 16724 -10408 16820 -10392
rect 15312 -10508 15408 -10472
rect 16724 -10472 16740 -10408
rect 16804 -10472 16820 -10408
rect 17143 -9728 17865 -9719
rect 17143 -10432 17152 -9728
rect 17856 -10432 17865 -9728
rect 17143 -10441 17865 -10432
rect 18136 -9752 18152 -9688
rect 18216 -9752 18232 -9688
rect 19548 -9688 19644 -9652
rect 18136 -9768 18232 -9752
rect 18136 -9832 18152 -9768
rect 18216 -9832 18232 -9768
rect 18136 -9848 18232 -9832
rect 18136 -9912 18152 -9848
rect 18216 -9912 18232 -9848
rect 18136 -9928 18232 -9912
rect 18136 -9992 18152 -9928
rect 18216 -9992 18232 -9928
rect 18136 -10008 18232 -9992
rect 18136 -10072 18152 -10008
rect 18216 -10072 18232 -10008
rect 18136 -10088 18232 -10072
rect 18136 -10152 18152 -10088
rect 18216 -10152 18232 -10088
rect 18136 -10168 18232 -10152
rect 18136 -10232 18152 -10168
rect 18216 -10232 18232 -10168
rect 18136 -10248 18232 -10232
rect 18136 -10312 18152 -10248
rect 18216 -10312 18232 -10248
rect 18136 -10328 18232 -10312
rect 18136 -10392 18152 -10328
rect 18216 -10392 18232 -10328
rect 18136 -10408 18232 -10392
rect 16724 -10508 16820 -10472
rect 18136 -10472 18152 -10408
rect 18216 -10472 18232 -10408
rect 18555 -9728 19277 -9719
rect 18555 -10432 18564 -9728
rect 19268 -10432 19277 -9728
rect 18555 -10441 19277 -10432
rect 19548 -9752 19564 -9688
rect 19628 -9752 19644 -9688
rect 20960 -9688 21056 -9652
rect 19548 -9768 19644 -9752
rect 19548 -9832 19564 -9768
rect 19628 -9832 19644 -9768
rect 19548 -9848 19644 -9832
rect 19548 -9912 19564 -9848
rect 19628 -9912 19644 -9848
rect 19548 -9928 19644 -9912
rect 19548 -9992 19564 -9928
rect 19628 -9992 19644 -9928
rect 19548 -10008 19644 -9992
rect 19548 -10072 19564 -10008
rect 19628 -10072 19644 -10008
rect 19548 -10088 19644 -10072
rect 19548 -10152 19564 -10088
rect 19628 -10152 19644 -10088
rect 19548 -10168 19644 -10152
rect 19548 -10232 19564 -10168
rect 19628 -10232 19644 -10168
rect 19548 -10248 19644 -10232
rect 19548 -10312 19564 -10248
rect 19628 -10312 19644 -10248
rect 19548 -10328 19644 -10312
rect 19548 -10392 19564 -10328
rect 19628 -10392 19644 -10328
rect 19548 -10408 19644 -10392
rect 18136 -10508 18232 -10472
rect 19548 -10472 19564 -10408
rect 19628 -10472 19644 -10408
rect 19967 -9728 20689 -9719
rect 19967 -10432 19976 -9728
rect 20680 -10432 20689 -9728
rect 19967 -10441 20689 -10432
rect 20960 -9752 20976 -9688
rect 21040 -9752 21056 -9688
rect 22372 -9688 22468 -9652
rect 20960 -9768 21056 -9752
rect 20960 -9832 20976 -9768
rect 21040 -9832 21056 -9768
rect 20960 -9848 21056 -9832
rect 20960 -9912 20976 -9848
rect 21040 -9912 21056 -9848
rect 20960 -9928 21056 -9912
rect 20960 -9992 20976 -9928
rect 21040 -9992 21056 -9928
rect 20960 -10008 21056 -9992
rect 20960 -10072 20976 -10008
rect 21040 -10072 21056 -10008
rect 20960 -10088 21056 -10072
rect 20960 -10152 20976 -10088
rect 21040 -10152 21056 -10088
rect 20960 -10168 21056 -10152
rect 20960 -10232 20976 -10168
rect 21040 -10232 21056 -10168
rect 20960 -10248 21056 -10232
rect 20960 -10312 20976 -10248
rect 21040 -10312 21056 -10248
rect 20960 -10328 21056 -10312
rect 20960 -10392 20976 -10328
rect 21040 -10392 21056 -10328
rect 20960 -10408 21056 -10392
rect 19548 -10508 19644 -10472
rect 20960 -10472 20976 -10408
rect 21040 -10472 21056 -10408
rect 21379 -9728 22101 -9719
rect 21379 -10432 21388 -9728
rect 22092 -10432 22101 -9728
rect 21379 -10441 22101 -10432
rect 22372 -9752 22388 -9688
rect 22452 -9752 22468 -9688
rect 23784 -9688 23880 -9652
rect 22372 -9768 22468 -9752
rect 22372 -9832 22388 -9768
rect 22452 -9832 22468 -9768
rect 22372 -9848 22468 -9832
rect 22372 -9912 22388 -9848
rect 22452 -9912 22468 -9848
rect 22372 -9928 22468 -9912
rect 22372 -9992 22388 -9928
rect 22452 -9992 22468 -9928
rect 22372 -10008 22468 -9992
rect 22372 -10072 22388 -10008
rect 22452 -10072 22468 -10008
rect 22372 -10088 22468 -10072
rect 22372 -10152 22388 -10088
rect 22452 -10152 22468 -10088
rect 22372 -10168 22468 -10152
rect 22372 -10232 22388 -10168
rect 22452 -10232 22468 -10168
rect 22372 -10248 22468 -10232
rect 22372 -10312 22388 -10248
rect 22452 -10312 22468 -10248
rect 22372 -10328 22468 -10312
rect 22372 -10392 22388 -10328
rect 22452 -10392 22468 -10328
rect 22372 -10408 22468 -10392
rect 20960 -10508 21056 -10472
rect 22372 -10472 22388 -10408
rect 22452 -10472 22468 -10408
rect 22791 -9728 23513 -9719
rect 22791 -10432 22800 -9728
rect 23504 -10432 23513 -9728
rect 22791 -10441 23513 -10432
rect 23784 -9752 23800 -9688
rect 23864 -9752 23880 -9688
rect 23784 -9768 23880 -9752
rect 23784 -9832 23800 -9768
rect 23864 -9832 23880 -9768
rect 23784 -9848 23880 -9832
rect 23784 -9912 23800 -9848
rect 23864 -9912 23880 -9848
rect 23784 -9928 23880 -9912
rect 23784 -9992 23800 -9928
rect 23864 -9992 23880 -9928
rect 23784 -10008 23880 -9992
rect 23784 -10072 23800 -10008
rect 23864 -10072 23880 -10008
rect 23784 -10088 23880 -10072
rect 23784 -10152 23800 -10088
rect 23864 -10152 23880 -10088
rect 23784 -10168 23880 -10152
rect 23784 -10232 23800 -10168
rect 23864 -10232 23880 -10168
rect 23784 -10248 23880 -10232
rect 23784 -10312 23800 -10248
rect 23864 -10312 23880 -10248
rect 23784 -10328 23880 -10312
rect 23784 -10392 23800 -10328
rect 23864 -10392 23880 -10328
rect 23784 -10408 23880 -10392
rect 22372 -10508 22468 -10472
rect 23784 -10472 23800 -10408
rect 23864 -10472 23880 -10408
rect 23784 -10508 23880 -10472
rect -22812 -10808 -22716 -10772
rect -23805 -10848 -23083 -10839
rect -23805 -11552 -23796 -10848
rect -23092 -11552 -23083 -10848
rect -23805 -11561 -23083 -11552
rect -22812 -10872 -22796 -10808
rect -22732 -10872 -22716 -10808
rect -21400 -10808 -21304 -10772
rect -22812 -10888 -22716 -10872
rect -22812 -10952 -22796 -10888
rect -22732 -10952 -22716 -10888
rect -22812 -10968 -22716 -10952
rect -22812 -11032 -22796 -10968
rect -22732 -11032 -22716 -10968
rect -22812 -11048 -22716 -11032
rect -22812 -11112 -22796 -11048
rect -22732 -11112 -22716 -11048
rect -22812 -11128 -22716 -11112
rect -22812 -11192 -22796 -11128
rect -22732 -11192 -22716 -11128
rect -22812 -11208 -22716 -11192
rect -22812 -11272 -22796 -11208
rect -22732 -11272 -22716 -11208
rect -22812 -11288 -22716 -11272
rect -22812 -11352 -22796 -11288
rect -22732 -11352 -22716 -11288
rect -22812 -11368 -22716 -11352
rect -22812 -11432 -22796 -11368
rect -22732 -11432 -22716 -11368
rect -22812 -11448 -22716 -11432
rect -22812 -11512 -22796 -11448
rect -22732 -11512 -22716 -11448
rect -22812 -11528 -22716 -11512
rect -22812 -11592 -22796 -11528
rect -22732 -11592 -22716 -11528
rect -22393 -10848 -21671 -10839
rect -22393 -11552 -22384 -10848
rect -21680 -11552 -21671 -10848
rect -22393 -11561 -21671 -11552
rect -21400 -10872 -21384 -10808
rect -21320 -10872 -21304 -10808
rect -19988 -10808 -19892 -10772
rect -21400 -10888 -21304 -10872
rect -21400 -10952 -21384 -10888
rect -21320 -10952 -21304 -10888
rect -21400 -10968 -21304 -10952
rect -21400 -11032 -21384 -10968
rect -21320 -11032 -21304 -10968
rect -21400 -11048 -21304 -11032
rect -21400 -11112 -21384 -11048
rect -21320 -11112 -21304 -11048
rect -21400 -11128 -21304 -11112
rect -21400 -11192 -21384 -11128
rect -21320 -11192 -21304 -11128
rect -21400 -11208 -21304 -11192
rect -21400 -11272 -21384 -11208
rect -21320 -11272 -21304 -11208
rect -21400 -11288 -21304 -11272
rect -21400 -11352 -21384 -11288
rect -21320 -11352 -21304 -11288
rect -21400 -11368 -21304 -11352
rect -21400 -11432 -21384 -11368
rect -21320 -11432 -21304 -11368
rect -21400 -11448 -21304 -11432
rect -21400 -11512 -21384 -11448
rect -21320 -11512 -21304 -11448
rect -21400 -11528 -21304 -11512
rect -22812 -11628 -22716 -11592
rect -21400 -11592 -21384 -11528
rect -21320 -11592 -21304 -11528
rect -20981 -10848 -20259 -10839
rect -20981 -11552 -20972 -10848
rect -20268 -11552 -20259 -10848
rect -20981 -11561 -20259 -11552
rect -19988 -10872 -19972 -10808
rect -19908 -10872 -19892 -10808
rect -18576 -10808 -18480 -10772
rect -19988 -10888 -19892 -10872
rect -19988 -10952 -19972 -10888
rect -19908 -10952 -19892 -10888
rect -19988 -10968 -19892 -10952
rect -19988 -11032 -19972 -10968
rect -19908 -11032 -19892 -10968
rect -19988 -11048 -19892 -11032
rect -19988 -11112 -19972 -11048
rect -19908 -11112 -19892 -11048
rect -19988 -11128 -19892 -11112
rect -19988 -11192 -19972 -11128
rect -19908 -11192 -19892 -11128
rect -19988 -11208 -19892 -11192
rect -19988 -11272 -19972 -11208
rect -19908 -11272 -19892 -11208
rect -19988 -11288 -19892 -11272
rect -19988 -11352 -19972 -11288
rect -19908 -11352 -19892 -11288
rect -19988 -11368 -19892 -11352
rect -19988 -11432 -19972 -11368
rect -19908 -11432 -19892 -11368
rect -19988 -11448 -19892 -11432
rect -19988 -11512 -19972 -11448
rect -19908 -11512 -19892 -11448
rect -19988 -11528 -19892 -11512
rect -21400 -11628 -21304 -11592
rect -19988 -11592 -19972 -11528
rect -19908 -11592 -19892 -11528
rect -19569 -10848 -18847 -10839
rect -19569 -11552 -19560 -10848
rect -18856 -11552 -18847 -10848
rect -19569 -11561 -18847 -11552
rect -18576 -10872 -18560 -10808
rect -18496 -10872 -18480 -10808
rect -17164 -10808 -17068 -10772
rect -18576 -10888 -18480 -10872
rect -18576 -10952 -18560 -10888
rect -18496 -10952 -18480 -10888
rect -18576 -10968 -18480 -10952
rect -18576 -11032 -18560 -10968
rect -18496 -11032 -18480 -10968
rect -18576 -11048 -18480 -11032
rect -18576 -11112 -18560 -11048
rect -18496 -11112 -18480 -11048
rect -18576 -11128 -18480 -11112
rect -18576 -11192 -18560 -11128
rect -18496 -11192 -18480 -11128
rect -18576 -11208 -18480 -11192
rect -18576 -11272 -18560 -11208
rect -18496 -11272 -18480 -11208
rect -18576 -11288 -18480 -11272
rect -18576 -11352 -18560 -11288
rect -18496 -11352 -18480 -11288
rect -18576 -11368 -18480 -11352
rect -18576 -11432 -18560 -11368
rect -18496 -11432 -18480 -11368
rect -18576 -11448 -18480 -11432
rect -18576 -11512 -18560 -11448
rect -18496 -11512 -18480 -11448
rect -18576 -11528 -18480 -11512
rect -19988 -11628 -19892 -11592
rect -18576 -11592 -18560 -11528
rect -18496 -11592 -18480 -11528
rect -18157 -10848 -17435 -10839
rect -18157 -11552 -18148 -10848
rect -17444 -11552 -17435 -10848
rect -18157 -11561 -17435 -11552
rect -17164 -10872 -17148 -10808
rect -17084 -10872 -17068 -10808
rect -15752 -10808 -15656 -10772
rect -17164 -10888 -17068 -10872
rect -17164 -10952 -17148 -10888
rect -17084 -10952 -17068 -10888
rect -17164 -10968 -17068 -10952
rect -17164 -11032 -17148 -10968
rect -17084 -11032 -17068 -10968
rect -17164 -11048 -17068 -11032
rect -17164 -11112 -17148 -11048
rect -17084 -11112 -17068 -11048
rect -17164 -11128 -17068 -11112
rect -17164 -11192 -17148 -11128
rect -17084 -11192 -17068 -11128
rect -17164 -11208 -17068 -11192
rect -17164 -11272 -17148 -11208
rect -17084 -11272 -17068 -11208
rect -17164 -11288 -17068 -11272
rect -17164 -11352 -17148 -11288
rect -17084 -11352 -17068 -11288
rect -17164 -11368 -17068 -11352
rect -17164 -11432 -17148 -11368
rect -17084 -11432 -17068 -11368
rect -17164 -11448 -17068 -11432
rect -17164 -11512 -17148 -11448
rect -17084 -11512 -17068 -11448
rect -17164 -11528 -17068 -11512
rect -18576 -11628 -18480 -11592
rect -17164 -11592 -17148 -11528
rect -17084 -11592 -17068 -11528
rect -16745 -10848 -16023 -10839
rect -16745 -11552 -16736 -10848
rect -16032 -11552 -16023 -10848
rect -16745 -11561 -16023 -11552
rect -15752 -10872 -15736 -10808
rect -15672 -10872 -15656 -10808
rect -14340 -10808 -14244 -10772
rect -15752 -10888 -15656 -10872
rect -15752 -10952 -15736 -10888
rect -15672 -10952 -15656 -10888
rect -15752 -10968 -15656 -10952
rect -15752 -11032 -15736 -10968
rect -15672 -11032 -15656 -10968
rect -15752 -11048 -15656 -11032
rect -15752 -11112 -15736 -11048
rect -15672 -11112 -15656 -11048
rect -15752 -11128 -15656 -11112
rect -15752 -11192 -15736 -11128
rect -15672 -11192 -15656 -11128
rect -15752 -11208 -15656 -11192
rect -15752 -11272 -15736 -11208
rect -15672 -11272 -15656 -11208
rect -15752 -11288 -15656 -11272
rect -15752 -11352 -15736 -11288
rect -15672 -11352 -15656 -11288
rect -15752 -11368 -15656 -11352
rect -15752 -11432 -15736 -11368
rect -15672 -11432 -15656 -11368
rect -15752 -11448 -15656 -11432
rect -15752 -11512 -15736 -11448
rect -15672 -11512 -15656 -11448
rect -15752 -11528 -15656 -11512
rect -17164 -11628 -17068 -11592
rect -15752 -11592 -15736 -11528
rect -15672 -11592 -15656 -11528
rect -15333 -10848 -14611 -10839
rect -15333 -11552 -15324 -10848
rect -14620 -11552 -14611 -10848
rect -15333 -11561 -14611 -11552
rect -14340 -10872 -14324 -10808
rect -14260 -10872 -14244 -10808
rect -12928 -10808 -12832 -10772
rect -14340 -10888 -14244 -10872
rect -14340 -10952 -14324 -10888
rect -14260 -10952 -14244 -10888
rect -14340 -10968 -14244 -10952
rect -14340 -11032 -14324 -10968
rect -14260 -11032 -14244 -10968
rect -14340 -11048 -14244 -11032
rect -14340 -11112 -14324 -11048
rect -14260 -11112 -14244 -11048
rect -14340 -11128 -14244 -11112
rect -14340 -11192 -14324 -11128
rect -14260 -11192 -14244 -11128
rect -14340 -11208 -14244 -11192
rect -14340 -11272 -14324 -11208
rect -14260 -11272 -14244 -11208
rect -14340 -11288 -14244 -11272
rect -14340 -11352 -14324 -11288
rect -14260 -11352 -14244 -11288
rect -14340 -11368 -14244 -11352
rect -14340 -11432 -14324 -11368
rect -14260 -11432 -14244 -11368
rect -14340 -11448 -14244 -11432
rect -14340 -11512 -14324 -11448
rect -14260 -11512 -14244 -11448
rect -14340 -11528 -14244 -11512
rect -15752 -11628 -15656 -11592
rect -14340 -11592 -14324 -11528
rect -14260 -11592 -14244 -11528
rect -13921 -10848 -13199 -10839
rect -13921 -11552 -13912 -10848
rect -13208 -11552 -13199 -10848
rect -13921 -11561 -13199 -11552
rect -12928 -10872 -12912 -10808
rect -12848 -10872 -12832 -10808
rect -11516 -10808 -11420 -10772
rect -12928 -10888 -12832 -10872
rect -12928 -10952 -12912 -10888
rect -12848 -10952 -12832 -10888
rect -12928 -10968 -12832 -10952
rect -12928 -11032 -12912 -10968
rect -12848 -11032 -12832 -10968
rect -12928 -11048 -12832 -11032
rect -12928 -11112 -12912 -11048
rect -12848 -11112 -12832 -11048
rect -12928 -11128 -12832 -11112
rect -12928 -11192 -12912 -11128
rect -12848 -11192 -12832 -11128
rect -12928 -11208 -12832 -11192
rect -12928 -11272 -12912 -11208
rect -12848 -11272 -12832 -11208
rect -12928 -11288 -12832 -11272
rect -12928 -11352 -12912 -11288
rect -12848 -11352 -12832 -11288
rect -12928 -11368 -12832 -11352
rect -12928 -11432 -12912 -11368
rect -12848 -11432 -12832 -11368
rect -12928 -11448 -12832 -11432
rect -12928 -11512 -12912 -11448
rect -12848 -11512 -12832 -11448
rect -12928 -11528 -12832 -11512
rect -14340 -11628 -14244 -11592
rect -12928 -11592 -12912 -11528
rect -12848 -11592 -12832 -11528
rect -12509 -10848 -11787 -10839
rect -12509 -11552 -12500 -10848
rect -11796 -11552 -11787 -10848
rect -12509 -11561 -11787 -11552
rect -11516 -10872 -11500 -10808
rect -11436 -10872 -11420 -10808
rect -10104 -10808 -10008 -10772
rect -11516 -10888 -11420 -10872
rect -11516 -10952 -11500 -10888
rect -11436 -10952 -11420 -10888
rect -11516 -10968 -11420 -10952
rect -11516 -11032 -11500 -10968
rect -11436 -11032 -11420 -10968
rect -11516 -11048 -11420 -11032
rect -11516 -11112 -11500 -11048
rect -11436 -11112 -11420 -11048
rect -11516 -11128 -11420 -11112
rect -11516 -11192 -11500 -11128
rect -11436 -11192 -11420 -11128
rect -11516 -11208 -11420 -11192
rect -11516 -11272 -11500 -11208
rect -11436 -11272 -11420 -11208
rect -11516 -11288 -11420 -11272
rect -11516 -11352 -11500 -11288
rect -11436 -11352 -11420 -11288
rect -11516 -11368 -11420 -11352
rect -11516 -11432 -11500 -11368
rect -11436 -11432 -11420 -11368
rect -11516 -11448 -11420 -11432
rect -11516 -11512 -11500 -11448
rect -11436 -11512 -11420 -11448
rect -11516 -11528 -11420 -11512
rect -12928 -11628 -12832 -11592
rect -11516 -11592 -11500 -11528
rect -11436 -11592 -11420 -11528
rect -11097 -10848 -10375 -10839
rect -11097 -11552 -11088 -10848
rect -10384 -11552 -10375 -10848
rect -11097 -11561 -10375 -11552
rect -10104 -10872 -10088 -10808
rect -10024 -10872 -10008 -10808
rect -8692 -10808 -8596 -10772
rect -10104 -10888 -10008 -10872
rect -10104 -10952 -10088 -10888
rect -10024 -10952 -10008 -10888
rect -10104 -10968 -10008 -10952
rect -10104 -11032 -10088 -10968
rect -10024 -11032 -10008 -10968
rect -10104 -11048 -10008 -11032
rect -10104 -11112 -10088 -11048
rect -10024 -11112 -10008 -11048
rect -10104 -11128 -10008 -11112
rect -10104 -11192 -10088 -11128
rect -10024 -11192 -10008 -11128
rect -10104 -11208 -10008 -11192
rect -10104 -11272 -10088 -11208
rect -10024 -11272 -10008 -11208
rect -10104 -11288 -10008 -11272
rect -10104 -11352 -10088 -11288
rect -10024 -11352 -10008 -11288
rect -10104 -11368 -10008 -11352
rect -10104 -11432 -10088 -11368
rect -10024 -11432 -10008 -11368
rect -10104 -11448 -10008 -11432
rect -10104 -11512 -10088 -11448
rect -10024 -11512 -10008 -11448
rect -10104 -11528 -10008 -11512
rect -11516 -11628 -11420 -11592
rect -10104 -11592 -10088 -11528
rect -10024 -11592 -10008 -11528
rect -9685 -10848 -8963 -10839
rect -9685 -11552 -9676 -10848
rect -8972 -11552 -8963 -10848
rect -9685 -11561 -8963 -11552
rect -8692 -10872 -8676 -10808
rect -8612 -10872 -8596 -10808
rect -7280 -10808 -7184 -10772
rect -8692 -10888 -8596 -10872
rect -8692 -10952 -8676 -10888
rect -8612 -10952 -8596 -10888
rect -8692 -10968 -8596 -10952
rect -8692 -11032 -8676 -10968
rect -8612 -11032 -8596 -10968
rect -8692 -11048 -8596 -11032
rect -8692 -11112 -8676 -11048
rect -8612 -11112 -8596 -11048
rect -8692 -11128 -8596 -11112
rect -8692 -11192 -8676 -11128
rect -8612 -11192 -8596 -11128
rect -8692 -11208 -8596 -11192
rect -8692 -11272 -8676 -11208
rect -8612 -11272 -8596 -11208
rect -8692 -11288 -8596 -11272
rect -8692 -11352 -8676 -11288
rect -8612 -11352 -8596 -11288
rect -8692 -11368 -8596 -11352
rect -8692 -11432 -8676 -11368
rect -8612 -11432 -8596 -11368
rect -8692 -11448 -8596 -11432
rect -8692 -11512 -8676 -11448
rect -8612 -11512 -8596 -11448
rect -8692 -11528 -8596 -11512
rect -10104 -11628 -10008 -11592
rect -8692 -11592 -8676 -11528
rect -8612 -11592 -8596 -11528
rect -8273 -10848 -7551 -10839
rect -8273 -11552 -8264 -10848
rect -7560 -11552 -7551 -10848
rect -8273 -11561 -7551 -11552
rect -7280 -10872 -7264 -10808
rect -7200 -10872 -7184 -10808
rect -5868 -10808 -5772 -10772
rect -7280 -10888 -7184 -10872
rect -7280 -10952 -7264 -10888
rect -7200 -10952 -7184 -10888
rect -7280 -10968 -7184 -10952
rect -7280 -11032 -7264 -10968
rect -7200 -11032 -7184 -10968
rect -7280 -11048 -7184 -11032
rect -7280 -11112 -7264 -11048
rect -7200 -11112 -7184 -11048
rect -7280 -11128 -7184 -11112
rect -7280 -11192 -7264 -11128
rect -7200 -11192 -7184 -11128
rect -7280 -11208 -7184 -11192
rect -7280 -11272 -7264 -11208
rect -7200 -11272 -7184 -11208
rect -7280 -11288 -7184 -11272
rect -7280 -11352 -7264 -11288
rect -7200 -11352 -7184 -11288
rect -7280 -11368 -7184 -11352
rect -7280 -11432 -7264 -11368
rect -7200 -11432 -7184 -11368
rect -7280 -11448 -7184 -11432
rect -7280 -11512 -7264 -11448
rect -7200 -11512 -7184 -11448
rect -7280 -11528 -7184 -11512
rect -8692 -11628 -8596 -11592
rect -7280 -11592 -7264 -11528
rect -7200 -11592 -7184 -11528
rect -6861 -10848 -6139 -10839
rect -6861 -11552 -6852 -10848
rect -6148 -11552 -6139 -10848
rect -6861 -11561 -6139 -11552
rect -5868 -10872 -5852 -10808
rect -5788 -10872 -5772 -10808
rect -4456 -10808 -4360 -10772
rect -5868 -10888 -5772 -10872
rect -5868 -10952 -5852 -10888
rect -5788 -10952 -5772 -10888
rect -5868 -10968 -5772 -10952
rect -5868 -11032 -5852 -10968
rect -5788 -11032 -5772 -10968
rect -5868 -11048 -5772 -11032
rect -5868 -11112 -5852 -11048
rect -5788 -11112 -5772 -11048
rect -5868 -11128 -5772 -11112
rect -5868 -11192 -5852 -11128
rect -5788 -11192 -5772 -11128
rect -5868 -11208 -5772 -11192
rect -5868 -11272 -5852 -11208
rect -5788 -11272 -5772 -11208
rect -5868 -11288 -5772 -11272
rect -5868 -11352 -5852 -11288
rect -5788 -11352 -5772 -11288
rect -5868 -11368 -5772 -11352
rect -5868 -11432 -5852 -11368
rect -5788 -11432 -5772 -11368
rect -5868 -11448 -5772 -11432
rect -5868 -11512 -5852 -11448
rect -5788 -11512 -5772 -11448
rect -5868 -11528 -5772 -11512
rect -7280 -11628 -7184 -11592
rect -5868 -11592 -5852 -11528
rect -5788 -11592 -5772 -11528
rect -5449 -10848 -4727 -10839
rect -5449 -11552 -5440 -10848
rect -4736 -11552 -4727 -10848
rect -5449 -11561 -4727 -11552
rect -4456 -10872 -4440 -10808
rect -4376 -10872 -4360 -10808
rect -3044 -10808 -2948 -10772
rect -4456 -10888 -4360 -10872
rect -4456 -10952 -4440 -10888
rect -4376 -10952 -4360 -10888
rect -4456 -10968 -4360 -10952
rect -4456 -11032 -4440 -10968
rect -4376 -11032 -4360 -10968
rect -4456 -11048 -4360 -11032
rect -4456 -11112 -4440 -11048
rect -4376 -11112 -4360 -11048
rect -4456 -11128 -4360 -11112
rect -4456 -11192 -4440 -11128
rect -4376 -11192 -4360 -11128
rect -4456 -11208 -4360 -11192
rect -4456 -11272 -4440 -11208
rect -4376 -11272 -4360 -11208
rect -4456 -11288 -4360 -11272
rect -4456 -11352 -4440 -11288
rect -4376 -11352 -4360 -11288
rect -4456 -11368 -4360 -11352
rect -4456 -11432 -4440 -11368
rect -4376 -11432 -4360 -11368
rect -4456 -11448 -4360 -11432
rect -4456 -11512 -4440 -11448
rect -4376 -11512 -4360 -11448
rect -4456 -11528 -4360 -11512
rect -5868 -11628 -5772 -11592
rect -4456 -11592 -4440 -11528
rect -4376 -11592 -4360 -11528
rect -4037 -10848 -3315 -10839
rect -4037 -11552 -4028 -10848
rect -3324 -11552 -3315 -10848
rect -4037 -11561 -3315 -11552
rect -3044 -10872 -3028 -10808
rect -2964 -10872 -2948 -10808
rect -1632 -10808 -1536 -10772
rect -3044 -10888 -2948 -10872
rect -3044 -10952 -3028 -10888
rect -2964 -10952 -2948 -10888
rect -3044 -10968 -2948 -10952
rect -3044 -11032 -3028 -10968
rect -2964 -11032 -2948 -10968
rect -3044 -11048 -2948 -11032
rect -3044 -11112 -3028 -11048
rect -2964 -11112 -2948 -11048
rect -3044 -11128 -2948 -11112
rect -3044 -11192 -3028 -11128
rect -2964 -11192 -2948 -11128
rect -3044 -11208 -2948 -11192
rect -3044 -11272 -3028 -11208
rect -2964 -11272 -2948 -11208
rect -3044 -11288 -2948 -11272
rect -3044 -11352 -3028 -11288
rect -2964 -11352 -2948 -11288
rect -3044 -11368 -2948 -11352
rect -3044 -11432 -3028 -11368
rect -2964 -11432 -2948 -11368
rect -3044 -11448 -2948 -11432
rect -3044 -11512 -3028 -11448
rect -2964 -11512 -2948 -11448
rect -3044 -11528 -2948 -11512
rect -4456 -11628 -4360 -11592
rect -3044 -11592 -3028 -11528
rect -2964 -11592 -2948 -11528
rect -2625 -10848 -1903 -10839
rect -2625 -11552 -2616 -10848
rect -1912 -11552 -1903 -10848
rect -2625 -11561 -1903 -11552
rect -1632 -10872 -1616 -10808
rect -1552 -10872 -1536 -10808
rect -220 -10808 -124 -10772
rect -1632 -10888 -1536 -10872
rect -1632 -10952 -1616 -10888
rect -1552 -10952 -1536 -10888
rect -1632 -10968 -1536 -10952
rect -1632 -11032 -1616 -10968
rect -1552 -11032 -1536 -10968
rect -1632 -11048 -1536 -11032
rect -1632 -11112 -1616 -11048
rect -1552 -11112 -1536 -11048
rect -1632 -11128 -1536 -11112
rect -1632 -11192 -1616 -11128
rect -1552 -11192 -1536 -11128
rect -1632 -11208 -1536 -11192
rect -1632 -11272 -1616 -11208
rect -1552 -11272 -1536 -11208
rect -1632 -11288 -1536 -11272
rect -1632 -11352 -1616 -11288
rect -1552 -11352 -1536 -11288
rect -1632 -11368 -1536 -11352
rect -1632 -11432 -1616 -11368
rect -1552 -11432 -1536 -11368
rect -1632 -11448 -1536 -11432
rect -1632 -11512 -1616 -11448
rect -1552 -11512 -1536 -11448
rect -1632 -11528 -1536 -11512
rect -3044 -11628 -2948 -11592
rect -1632 -11592 -1616 -11528
rect -1552 -11592 -1536 -11528
rect -1213 -10848 -491 -10839
rect -1213 -11552 -1204 -10848
rect -500 -11552 -491 -10848
rect -1213 -11561 -491 -11552
rect -220 -10872 -204 -10808
rect -140 -10872 -124 -10808
rect 1192 -10808 1288 -10772
rect -220 -10888 -124 -10872
rect -220 -10952 -204 -10888
rect -140 -10952 -124 -10888
rect -220 -10968 -124 -10952
rect -220 -11032 -204 -10968
rect -140 -11032 -124 -10968
rect -220 -11048 -124 -11032
rect -220 -11112 -204 -11048
rect -140 -11112 -124 -11048
rect -220 -11128 -124 -11112
rect -220 -11192 -204 -11128
rect -140 -11192 -124 -11128
rect -220 -11208 -124 -11192
rect -220 -11272 -204 -11208
rect -140 -11272 -124 -11208
rect -220 -11288 -124 -11272
rect -220 -11352 -204 -11288
rect -140 -11352 -124 -11288
rect -220 -11368 -124 -11352
rect -220 -11432 -204 -11368
rect -140 -11432 -124 -11368
rect -220 -11448 -124 -11432
rect -220 -11512 -204 -11448
rect -140 -11512 -124 -11448
rect -220 -11528 -124 -11512
rect -1632 -11628 -1536 -11592
rect -220 -11592 -204 -11528
rect -140 -11592 -124 -11528
rect 199 -10848 921 -10839
rect 199 -11552 208 -10848
rect 912 -11552 921 -10848
rect 199 -11561 921 -11552
rect 1192 -10872 1208 -10808
rect 1272 -10872 1288 -10808
rect 2604 -10808 2700 -10772
rect 1192 -10888 1288 -10872
rect 1192 -10952 1208 -10888
rect 1272 -10952 1288 -10888
rect 1192 -10968 1288 -10952
rect 1192 -11032 1208 -10968
rect 1272 -11032 1288 -10968
rect 1192 -11048 1288 -11032
rect 1192 -11112 1208 -11048
rect 1272 -11112 1288 -11048
rect 1192 -11128 1288 -11112
rect 1192 -11192 1208 -11128
rect 1272 -11192 1288 -11128
rect 1192 -11208 1288 -11192
rect 1192 -11272 1208 -11208
rect 1272 -11272 1288 -11208
rect 1192 -11288 1288 -11272
rect 1192 -11352 1208 -11288
rect 1272 -11352 1288 -11288
rect 1192 -11368 1288 -11352
rect 1192 -11432 1208 -11368
rect 1272 -11432 1288 -11368
rect 1192 -11448 1288 -11432
rect 1192 -11512 1208 -11448
rect 1272 -11512 1288 -11448
rect 1192 -11528 1288 -11512
rect -220 -11628 -124 -11592
rect 1192 -11592 1208 -11528
rect 1272 -11592 1288 -11528
rect 1611 -10848 2333 -10839
rect 1611 -11552 1620 -10848
rect 2324 -11552 2333 -10848
rect 1611 -11561 2333 -11552
rect 2604 -10872 2620 -10808
rect 2684 -10872 2700 -10808
rect 4016 -10808 4112 -10772
rect 2604 -10888 2700 -10872
rect 2604 -10952 2620 -10888
rect 2684 -10952 2700 -10888
rect 2604 -10968 2700 -10952
rect 2604 -11032 2620 -10968
rect 2684 -11032 2700 -10968
rect 2604 -11048 2700 -11032
rect 2604 -11112 2620 -11048
rect 2684 -11112 2700 -11048
rect 2604 -11128 2700 -11112
rect 2604 -11192 2620 -11128
rect 2684 -11192 2700 -11128
rect 2604 -11208 2700 -11192
rect 2604 -11272 2620 -11208
rect 2684 -11272 2700 -11208
rect 2604 -11288 2700 -11272
rect 2604 -11352 2620 -11288
rect 2684 -11352 2700 -11288
rect 2604 -11368 2700 -11352
rect 2604 -11432 2620 -11368
rect 2684 -11432 2700 -11368
rect 2604 -11448 2700 -11432
rect 2604 -11512 2620 -11448
rect 2684 -11512 2700 -11448
rect 2604 -11528 2700 -11512
rect 1192 -11628 1288 -11592
rect 2604 -11592 2620 -11528
rect 2684 -11592 2700 -11528
rect 3023 -10848 3745 -10839
rect 3023 -11552 3032 -10848
rect 3736 -11552 3745 -10848
rect 3023 -11561 3745 -11552
rect 4016 -10872 4032 -10808
rect 4096 -10872 4112 -10808
rect 5428 -10808 5524 -10772
rect 4016 -10888 4112 -10872
rect 4016 -10952 4032 -10888
rect 4096 -10952 4112 -10888
rect 4016 -10968 4112 -10952
rect 4016 -11032 4032 -10968
rect 4096 -11032 4112 -10968
rect 4016 -11048 4112 -11032
rect 4016 -11112 4032 -11048
rect 4096 -11112 4112 -11048
rect 4016 -11128 4112 -11112
rect 4016 -11192 4032 -11128
rect 4096 -11192 4112 -11128
rect 4016 -11208 4112 -11192
rect 4016 -11272 4032 -11208
rect 4096 -11272 4112 -11208
rect 4016 -11288 4112 -11272
rect 4016 -11352 4032 -11288
rect 4096 -11352 4112 -11288
rect 4016 -11368 4112 -11352
rect 4016 -11432 4032 -11368
rect 4096 -11432 4112 -11368
rect 4016 -11448 4112 -11432
rect 4016 -11512 4032 -11448
rect 4096 -11512 4112 -11448
rect 4016 -11528 4112 -11512
rect 2604 -11628 2700 -11592
rect 4016 -11592 4032 -11528
rect 4096 -11592 4112 -11528
rect 4435 -10848 5157 -10839
rect 4435 -11552 4444 -10848
rect 5148 -11552 5157 -10848
rect 4435 -11561 5157 -11552
rect 5428 -10872 5444 -10808
rect 5508 -10872 5524 -10808
rect 6840 -10808 6936 -10772
rect 5428 -10888 5524 -10872
rect 5428 -10952 5444 -10888
rect 5508 -10952 5524 -10888
rect 5428 -10968 5524 -10952
rect 5428 -11032 5444 -10968
rect 5508 -11032 5524 -10968
rect 5428 -11048 5524 -11032
rect 5428 -11112 5444 -11048
rect 5508 -11112 5524 -11048
rect 5428 -11128 5524 -11112
rect 5428 -11192 5444 -11128
rect 5508 -11192 5524 -11128
rect 5428 -11208 5524 -11192
rect 5428 -11272 5444 -11208
rect 5508 -11272 5524 -11208
rect 5428 -11288 5524 -11272
rect 5428 -11352 5444 -11288
rect 5508 -11352 5524 -11288
rect 5428 -11368 5524 -11352
rect 5428 -11432 5444 -11368
rect 5508 -11432 5524 -11368
rect 5428 -11448 5524 -11432
rect 5428 -11512 5444 -11448
rect 5508 -11512 5524 -11448
rect 5428 -11528 5524 -11512
rect 4016 -11628 4112 -11592
rect 5428 -11592 5444 -11528
rect 5508 -11592 5524 -11528
rect 5847 -10848 6569 -10839
rect 5847 -11552 5856 -10848
rect 6560 -11552 6569 -10848
rect 5847 -11561 6569 -11552
rect 6840 -10872 6856 -10808
rect 6920 -10872 6936 -10808
rect 8252 -10808 8348 -10772
rect 6840 -10888 6936 -10872
rect 6840 -10952 6856 -10888
rect 6920 -10952 6936 -10888
rect 6840 -10968 6936 -10952
rect 6840 -11032 6856 -10968
rect 6920 -11032 6936 -10968
rect 6840 -11048 6936 -11032
rect 6840 -11112 6856 -11048
rect 6920 -11112 6936 -11048
rect 6840 -11128 6936 -11112
rect 6840 -11192 6856 -11128
rect 6920 -11192 6936 -11128
rect 6840 -11208 6936 -11192
rect 6840 -11272 6856 -11208
rect 6920 -11272 6936 -11208
rect 6840 -11288 6936 -11272
rect 6840 -11352 6856 -11288
rect 6920 -11352 6936 -11288
rect 6840 -11368 6936 -11352
rect 6840 -11432 6856 -11368
rect 6920 -11432 6936 -11368
rect 6840 -11448 6936 -11432
rect 6840 -11512 6856 -11448
rect 6920 -11512 6936 -11448
rect 6840 -11528 6936 -11512
rect 5428 -11628 5524 -11592
rect 6840 -11592 6856 -11528
rect 6920 -11592 6936 -11528
rect 7259 -10848 7981 -10839
rect 7259 -11552 7268 -10848
rect 7972 -11552 7981 -10848
rect 7259 -11561 7981 -11552
rect 8252 -10872 8268 -10808
rect 8332 -10872 8348 -10808
rect 9664 -10808 9760 -10772
rect 8252 -10888 8348 -10872
rect 8252 -10952 8268 -10888
rect 8332 -10952 8348 -10888
rect 8252 -10968 8348 -10952
rect 8252 -11032 8268 -10968
rect 8332 -11032 8348 -10968
rect 8252 -11048 8348 -11032
rect 8252 -11112 8268 -11048
rect 8332 -11112 8348 -11048
rect 8252 -11128 8348 -11112
rect 8252 -11192 8268 -11128
rect 8332 -11192 8348 -11128
rect 8252 -11208 8348 -11192
rect 8252 -11272 8268 -11208
rect 8332 -11272 8348 -11208
rect 8252 -11288 8348 -11272
rect 8252 -11352 8268 -11288
rect 8332 -11352 8348 -11288
rect 8252 -11368 8348 -11352
rect 8252 -11432 8268 -11368
rect 8332 -11432 8348 -11368
rect 8252 -11448 8348 -11432
rect 8252 -11512 8268 -11448
rect 8332 -11512 8348 -11448
rect 8252 -11528 8348 -11512
rect 6840 -11628 6936 -11592
rect 8252 -11592 8268 -11528
rect 8332 -11592 8348 -11528
rect 8671 -10848 9393 -10839
rect 8671 -11552 8680 -10848
rect 9384 -11552 9393 -10848
rect 8671 -11561 9393 -11552
rect 9664 -10872 9680 -10808
rect 9744 -10872 9760 -10808
rect 11076 -10808 11172 -10772
rect 9664 -10888 9760 -10872
rect 9664 -10952 9680 -10888
rect 9744 -10952 9760 -10888
rect 9664 -10968 9760 -10952
rect 9664 -11032 9680 -10968
rect 9744 -11032 9760 -10968
rect 9664 -11048 9760 -11032
rect 9664 -11112 9680 -11048
rect 9744 -11112 9760 -11048
rect 9664 -11128 9760 -11112
rect 9664 -11192 9680 -11128
rect 9744 -11192 9760 -11128
rect 9664 -11208 9760 -11192
rect 9664 -11272 9680 -11208
rect 9744 -11272 9760 -11208
rect 9664 -11288 9760 -11272
rect 9664 -11352 9680 -11288
rect 9744 -11352 9760 -11288
rect 9664 -11368 9760 -11352
rect 9664 -11432 9680 -11368
rect 9744 -11432 9760 -11368
rect 9664 -11448 9760 -11432
rect 9664 -11512 9680 -11448
rect 9744 -11512 9760 -11448
rect 9664 -11528 9760 -11512
rect 8252 -11628 8348 -11592
rect 9664 -11592 9680 -11528
rect 9744 -11592 9760 -11528
rect 10083 -10848 10805 -10839
rect 10083 -11552 10092 -10848
rect 10796 -11552 10805 -10848
rect 10083 -11561 10805 -11552
rect 11076 -10872 11092 -10808
rect 11156 -10872 11172 -10808
rect 12488 -10808 12584 -10772
rect 11076 -10888 11172 -10872
rect 11076 -10952 11092 -10888
rect 11156 -10952 11172 -10888
rect 11076 -10968 11172 -10952
rect 11076 -11032 11092 -10968
rect 11156 -11032 11172 -10968
rect 11076 -11048 11172 -11032
rect 11076 -11112 11092 -11048
rect 11156 -11112 11172 -11048
rect 11076 -11128 11172 -11112
rect 11076 -11192 11092 -11128
rect 11156 -11192 11172 -11128
rect 11076 -11208 11172 -11192
rect 11076 -11272 11092 -11208
rect 11156 -11272 11172 -11208
rect 11076 -11288 11172 -11272
rect 11076 -11352 11092 -11288
rect 11156 -11352 11172 -11288
rect 11076 -11368 11172 -11352
rect 11076 -11432 11092 -11368
rect 11156 -11432 11172 -11368
rect 11076 -11448 11172 -11432
rect 11076 -11512 11092 -11448
rect 11156 -11512 11172 -11448
rect 11076 -11528 11172 -11512
rect 9664 -11628 9760 -11592
rect 11076 -11592 11092 -11528
rect 11156 -11592 11172 -11528
rect 11495 -10848 12217 -10839
rect 11495 -11552 11504 -10848
rect 12208 -11552 12217 -10848
rect 11495 -11561 12217 -11552
rect 12488 -10872 12504 -10808
rect 12568 -10872 12584 -10808
rect 13900 -10808 13996 -10772
rect 12488 -10888 12584 -10872
rect 12488 -10952 12504 -10888
rect 12568 -10952 12584 -10888
rect 12488 -10968 12584 -10952
rect 12488 -11032 12504 -10968
rect 12568 -11032 12584 -10968
rect 12488 -11048 12584 -11032
rect 12488 -11112 12504 -11048
rect 12568 -11112 12584 -11048
rect 12488 -11128 12584 -11112
rect 12488 -11192 12504 -11128
rect 12568 -11192 12584 -11128
rect 12488 -11208 12584 -11192
rect 12488 -11272 12504 -11208
rect 12568 -11272 12584 -11208
rect 12488 -11288 12584 -11272
rect 12488 -11352 12504 -11288
rect 12568 -11352 12584 -11288
rect 12488 -11368 12584 -11352
rect 12488 -11432 12504 -11368
rect 12568 -11432 12584 -11368
rect 12488 -11448 12584 -11432
rect 12488 -11512 12504 -11448
rect 12568 -11512 12584 -11448
rect 12488 -11528 12584 -11512
rect 11076 -11628 11172 -11592
rect 12488 -11592 12504 -11528
rect 12568 -11592 12584 -11528
rect 12907 -10848 13629 -10839
rect 12907 -11552 12916 -10848
rect 13620 -11552 13629 -10848
rect 12907 -11561 13629 -11552
rect 13900 -10872 13916 -10808
rect 13980 -10872 13996 -10808
rect 15312 -10808 15408 -10772
rect 13900 -10888 13996 -10872
rect 13900 -10952 13916 -10888
rect 13980 -10952 13996 -10888
rect 13900 -10968 13996 -10952
rect 13900 -11032 13916 -10968
rect 13980 -11032 13996 -10968
rect 13900 -11048 13996 -11032
rect 13900 -11112 13916 -11048
rect 13980 -11112 13996 -11048
rect 13900 -11128 13996 -11112
rect 13900 -11192 13916 -11128
rect 13980 -11192 13996 -11128
rect 13900 -11208 13996 -11192
rect 13900 -11272 13916 -11208
rect 13980 -11272 13996 -11208
rect 13900 -11288 13996 -11272
rect 13900 -11352 13916 -11288
rect 13980 -11352 13996 -11288
rect 13900 -11368 13996 -11352
rect 13900 -11432 13916 -11368
rect 13980 -11432 13996 -11368
rect 13900 -11448 13996 -11432
rect 13900 -11512 13916 -11448
rect 13980 -11512 13996 -11448
rect 13900 -11528 13996 -11512
rect 12488 -11628 12584 -11592
rect 13900 -11592 13916 -11528
rect 13980 -11592 13996 -11528
rect 14319 -10848 15041 -10839
rect 14319 -11552 14328 -10848
rect 15032 -11552 15041 -10848
rect 14319 -11561 15041 -11552
rect 15312 -10872 15328 -10808
rect 15392 -10872 15408 -10808
rect 16724 -10808 16820 -10772
rect 15312 -10888 15408 -10872
rect 15312 -10952 15328 -10888
rect 15392 -10952 15408 -10888
rect 15312 -10968 15408 -10952
rect 15312 -11032 15328 -10968
rect 15392 -11032 15408 -10968
rect 15312 -11048 15408 -11032
rect 15312 -11112 15328 -11048
rect 15392 -11112 15408 -11048
rect 15312 -11128 15408 -11112
rect 15312 -11192 15328 -11128
rect 15392 -11192 15408 -11128
rect 15312 -11208 15408 -11192
rect 15312 -11272 15328 -11208
rect 15392 -11272 15408 -11208
rect 15312 -11288 15408 -11272
rect 15312 -11352 15328 -11288
rect 15392 -11352 15408 -11288
rect 15312 -11368 15408 -11352
rect 15312 -11432 15328 -11368
rect 15392 -11432 15408 -11368
rect 15312 -11448 15408 -11432
rect 15312 -11512 15328 -11448
rect 15392 -11512 15408 -11448
rect 15312 -11528 15408 -11512
rect 13900 -11628 13996 -11592
rect 15312 -11592 15328 -11528
rect 15392 -11592 15408 -11528
rect 15731 -10848 16453 -10839
rect 15731 -11552 15740 -10848
rect 16444 -11552 16453 -10848
rect 15731 -11561 16453 -11552
rect 16724 -10872 16740 -10808
rect 16804 -10872 16820 -10808
rect 18136 -10808 18232 -10772
rect 16724 -10888 16820 -10872
rect 16724 -10952 16740 -10888
rect 16804 -10952 16820 -10888
rect 16724 -10968 16820 -10952
rect 16724 -11032 16740 -10968
rect 16804 -11032 16820 -10968
rect 16724 -11048 16820 -11032
rect 16724 -11112 16740 -11048
rect 16804 -11112 16820 -11048
rect 16724 -11128 16820 -11112
rect 16724 -11192 16740 -11128
rect 16804 -11192 16820 -11128
rect 16724 -11208 16820 -11192
rect 16724 -11272 16740 -11208
rect 16804 -11272 16820 -11208
rect 16724 -11288 16820 -11272
rect 16724 -11352 16740 -11288
rect 16804 -11352 16820 -11288
rect 16724 -11368 16820 -11352
rect 16724 -11432 16740 -11368
rect 16804 -11432 16820 -11368
rect 16724 -11448 16820 -11432
rect 16724 -11512 16740 -11448
rect 16804 -11512 16820 -11448
rect 16724 -11528 16820 -11512
rect 15312 -11628 15408 -11592
rect 16724 -11592 16740 -11528
rect 16804 -11592 16820 -11528
rect 17143 -10848 17865 -10839
rect 17143 -11552 17152 -10848
rect 17856 -11552 17865 -10848
rect 17143 -11561 17865 -11552
rect 18136 -10872 18152 -10808
rect 18216 -10872 18232 -10808
rect 19548 -10808 19644 -10772
rect 18136 -10888 18232 -10872
rect 18136 -10952 18152 -10888
rect 18216 -10952 18232 -10888
rect 18136 -10968 18232 -10952
rect 18136 -11032 18152 -10968
rect 18216 -11032 18232 -10968
rect 18136 -11048 18232 -11032
rect 18136 -11112 18152 -11048
rect 18216 -11112 18232 -11048
rect 18136 -11128 18232 -11112
rect 18136 -11192 18152 -11128
rect 18216 -11192 18232 -11128
rect 18136 -11208 18232 -11192
rect 18136 -11272 18152 -11208
rect 18216 -11272 18232 -11208
rect 18136 -11288 18232 -11272
rect 18136 -11352 18152 -11288
rect 18216 -11352 18232 -11288
rect 18136 -11368 18232 -11352
rect 18136 -11432 18152 -11368
rect 18216 -11432 18232 -11368
rect 18136 -11448 18232 -11432
rect 18136 -11512 18152 -11448
rect 18216 -11512 18232 -11448
rect 18136 -11528 18232 -11512
rect 16724 -11628 16820 -11592
rect 18136 -11592 18152 -11528
rect 18216 -11592 18232 -11528
rect 18555 -10848 19277 -10839
rect 18555 -11552 18564 -10848
rect 19268 -11552 19277 -10848
rect 18555 -11561 19277 -11552
rect 19548 -10872 19564 -10808
rect 19628 -10872 19644 -10808
rect 20960 -10808 21056 -10772
rect 19548 -10888 19644 -10872
rect 19548 -10952 19564 -10888
rect 19628 -10952 19644 -10888
rect 19548 -10968 19644 -10952
rect 19548 -11032 19564 -10968
rect 19628 -11032 19644 -10968
rect 19548 -11048 19644 -11032
rect 19548 -11112 19564 -11048
rect 19628 -11112 19644 -11048
rect 19548 -11128 19644 -11112
rect 19548 -11192 19564 -11128
rect 19628 -11192 19644 -11128
rect 19548 -11208 19644 -11192
rect 19548 -11272 19564 -11208
rect 19628 -11272 19644 -11208
rect 19548 -11288 19644 -11272
rect 19548 -11352 19564 -11288
rect 19628 -11352 19644 -11288
rect 19548 -11368 19644 -11352
rect 19548 -11432 19564 -11368
rect 19628 -11432 19644 -11368
rect 19548 -11448 19644 -11432
rect 19548 -11512 19564 -11448
rect 19628 -11512 19644 -11448
rect 19548 -11528 19644 -11512
rect 18136 -11628 18232 -11592
rect 19548 -11592 19564 -11528
rect 19628 -11592 19644 -11528
rect 19967 -10848 20689 -10839
rect 19967 -11552 19976 -10848
rect 20680 -11552 20689 -10848
rect 19967 -11561 20689 -11552
rect 20960 -10872 20976 -10808
rect 21040 -10872 21056 -10808
rect 22372 -10808 22468 -10772
rect 20960 -10888 21056 -10872
rect 20960 -10952 20976 -10888
rect 21040 -10952 21056 -10888
rect 20960 -10968 21056 -10952
rect 20960 -11032 20976 -10968
rect 21040 -11032 21056 -10968
rect 20960 -11048 21056 -11032
rect 20960 -11112 20976 -11048
rect 21040 -11112 21056 -11048
rect 20960 -11128 21056 -11112
rect 20960 -11192 20976 -11128
rect 21040 -11192 21056 -11128
rect 20960 -11208 21056 -11192
rect 20960 -11272 20976 -11208
rect 21040 -11272 21056 -11208
rect 20960 -11288 21056 -11272
rect 20960 -11352 20976 -11288
rect 21040 -11352 21056 -11288
rect 20960 -11368 21056 -11352
rect 20960 -11432 20976 -11368
rect 21040 -11432 21056 -11368
rect 20960 -11448 21056 -11432
rect 20960 -11512 20976 -11448
rect 21040 -11512 21056 -11448
rect 20960 -11528 21056 -11512
rect 19548 -11628 19644 -11592
rect 20960 -11592 20976 -11528
rect 21040 -11592 21056 -11528
rect 21379 -10848 22101 -10839
rect 21379 -11552 21388 -10848
rect 22092 -11552 22101 -10848
rect 21379 -11561 22101 -11552
rect 22372 -10872 22388 -10808
rect 22452 -10872 22468 -10808
rect 23784 -10808 23880 -10772
rect 22372 -10888 22468 -10872
rect 22372 -10952 22388 -10888
rect 22452 -10952 22468 -10888
rect 22372 -10968 22468 -10952
rect 22372 -11032 22388 -10968
rect 22452 -11032 22468 -10968
rect 22372 -11048 22468 -11032
rect 22372 -11112 22388 -11048
rect 22452 -11112 22468 -11048
rect 22372 -11128 22468 -11112
rect 22372 -11192 22388 -11128
rect 22452 -11192 22468 -11128
rect 22372 -11208 22468 -11192
rect 22372 -11272 22388 -11208
rect 22452 -11272 22468 -11208
rect 22372 -11288 22468 -11272
rect 22372 -11352 22388 -11288
rect 22452 -11352 22468 -11288
rect 22372 -11368 22468 -11352
rect 22372 -11432 22388 -11368
rect 22452 -11432 22468 -11368
rect 22372 -11448 22468 -11432
rect 22372 -11512 22388 -11448
rect 22452 -11512 22468 -11448
rect 22372 -11528 22468 -11512
rect 20960 -11628 21056 -11592
rect 22372 -11592 22388 -11528
rect 22452 -11592 22468 -11528
rect 22791 -10848 23513 -10839
rect 22791 -11552 22800 -10848
rect 23504 -11552 23513 -10848
rect 22791 -11561 23513 -11552
rect 23784 -10872 23800 -10808
rect 23864 -10872 23880 -10808
rect 23784 -10888 23880 -10872
rect 23784 -10952 23800 -10888
rect 23864 -10952 23880 -10888
rect 23784 -10968 23880 -10952
rect 23784 -11032 23800 -10968
rect 23864 -11032 23880 -10968
rect 23784 -11048 23880 -11032
rect 23784 -11112 23800 -11048
rect 23864 -11112 23880 -11048
rect 23784 -11128 23880 -11112
rect 23784 -11192 23800 -11128
rect 23864 -11192 23880 -11128
rect 23784 -11208 23880 -11192
rect 23784 -11272 23800 -11208
rect 23864 -11272 23880 -11208
rect 23784 -11288 23880 -11272
rect 23784 -11352 23800 -11288
rect 23864 -11352 23880 -11288
rect 23784 -11368 23880 -11352
rect 23784 -11432 23800 -11368
rect 23864 -11432 23880 -11368
rect 23784 -11448 23880 -11432
rect 23784 -11512 23800 -11448
rect 23864 -11512 23880 -11448
rect 23784 -11528 23880 -11512
rect 22372 -11628 22468 -11592
rect 23784 -11592 23800 -11528
rect 23864 -11592 23880 -11528
rect 23784 -11628 23880 -11592
rect -22812 -11928 -22716 -11892
rect -23805 -11968 -23083 -11959
rect -23805 -12672 -23796 -11968
rect -23092 -12672 -23083 -11968
rect -23805 -12681 -23083 -12672
rect -22812 -11992 -22796 -11928
rect -22732 -11992 -22716 -11928
rect -21400 -11928 -21304 -11892
rect -22812 -12008 -22716 -11992
rect -22812 -12072 -22796 -12008
rect -22732 -12072 -22716 -12008
rect -22812 -12088 -22716 -12072
rect -22812 -12152 -22796 -12088
rect -22732 -12152 -22716 -12088
rect -22812 -12168 -22716 -12152
rect -22812 -12232 -22796 -12168
rect -22732 -12232 -22716 -12168
rect -22812 -12248 -22716 -12232
rect -22812 -12312 -22796 -12248
rect -22732 -12312 -22716 -12248
rect -22812 -12328 -22716 -12312
rect -22812 -12392 -22796 -12328
rect -22732 -12392 -22716 -12328
rect -22812 -12408 -22716 -12392
rect -22812 -12472 -22796 -12408
rect -22732 -12472 -22716 -12408
rect -22812 -12488 -22716 -12472
rect -22812 -12552 -22796 -12488
rect -22732 -12552 -22716 -12488
rect -22812 -12568 -22716 -12552
rect -22812 -12632 -22796 -12568
rect -22732 -12632 -22716 -12568
rect -22812 -12648 -22716 -12632
rect -22812 -12712 -22796 -12648
rect -22732 -12712 -22716 -12648
rect -22393 -11968 -21671 -11959
rect -22393 -12672 -22384 -11968
rect -21680 -12672 -21671 -11968
rect -22393 -12681 -21671 -12672
rect -21400 -11992 -21384 -11928
rect -21320 -11992 -21304 -11928
rect -19988 -11928 -19892 -11892
rect -21400 -12008 -21304 -11992
rect -21400 -12072 -21384 -12008
rect -21320 -12072 -21304 -12008
rect -21400 -12088 -21304 -12072
rect -21400 -12152 -21384 -12088
rect -21320 -12152 -21304 -12088
rect -21400 -12168 -21304 -12152
rect -21400 -12232 -21384 -12168
rect -21320 -12232 -21304 -12168
rect -21400 -12248 -21304 -12232
rect -21400 -12312 -21384 -12248
rect -21320 -12312 -21304 -12248
rect -21400 -12328 -21304 -12312
rect -21400 -12392 -21384 -12328
rect -21320 -12392 -21304 -12328
rect -21400 -12408 -21304 -12392
rect -21400 -12472 -21384 -12408
rect -21320 -12472 -21304 -12408
rect -21400 -12488 -21304 -12472
rect -21400 -12552 -21384 -12488
rect -21320 -12552 -21304 -12488
rect -21400 -12568 -21304 -12552
rect -21400 -12632 -21384 -12568
rect -21320 -12632 -21304 -12568
rect -21400 -12648 -21304 -12632
rect -22812 -12748 -22716 -12712
rect -21400 -12712 -21384 -12648
rect -21320 -12712 -21304 -12648
rect -20981 -11968 -20259 -11959
rect -20981 -12672 -20972 -11968
rect -20268 -12672 -20259 -11968
rect -20981 -12681 -20259 -12672
rect -19988 -11992 -19972 -11928
rect -19908 -11992 -19892 -11928
rect -18576 -11928 -18480 -11892
rect -19988 -12008 -19892 -11992
rect -19988 -12072 -19972 -12008
rect -19908 -12072 -19892 -12008
rect -19988 -12088 -19892 -12072
rect -19988 -12152 -19972 -12088
rect -19908 -12152 -19892 -12088
rect -19988 -12168 -19892 -12152
rect -19988 -12232 -19972 -12168
rect -19908 -12232 -19892 -12168
rect -19988 -12248 -19892 -12232
rect -19988 -12312 -19972 -12248
rect -19908 -12312 -19892 -12248
rect -19988 -12328 -19892 -12312
rect -19988 -12392 -19972 -12328
rect -19908 -12392 -19892 -12328
rect -19988 -12408 -19892 -12392
rect -19988 -12472 -19972 -12408
rect -19908 -12472 -19892 -12408
rect -19988 -12488 -19892 -12472
rect -19988 -12552 -19972 -12488
rect -19908 -12552 -19892 -12488
rect -19988 -12568 -19892 -12552
rect -19988 -12632 -19972 -12568
rect -19908 -12632 -19892 -12568
rect -19988 -12648 -19892 -12632
rect -21400 -12748 -21304 -12712
rect -19988 -12712 -19972 -12648
rect -19908 -12712 -19892 -12648
rect -19569 -11968 -18847 -11959
rect -19569 -12672 -19560 -11968
rect -18856 -12672 -18847 -11968
rect -19569 -12681 -18847 -12672
rect -18576 -11992 -18560 -11928
rect -18496 -11992 -18480 -11928
rect -17164 -11928 -17068 -11892
rect -18576 -12008 -18480 -11992
rect -18576 -12072 -18560 -12008
rect -18496 -12072 -18480 -12008
rect -18576 -12088 -18480 -12072
rect -18576 -12152 -18560 -12088
rect -18496 -12152 -18480 -12088
rect -18576 -12168 -18480 -12152
rect -18576 -12232 -18560 -12168
rect -18496 -12232 -18480 -12168
rect -18576 -12248 -18480 -12232
rect -18576 -12312 -18560 -12248
rect -18496 -12312 -18480 -12248
rect -18576 -12328 -18480 -12312
rect -18576 -12392 -18560 -12328
rect -18496 -12392 -18480 -12328
rect -18576 -12408 -18480 -12392
rect -18576 -12472 -18560 -12408
rect -18496 -12472 -18480 -12408
rect -18576 -12488 -18480 -12472
rect -18576 -12552 -18560 -12488
rect -18496 -12552 -18480 -12488
rect -18576 -12568 -18480 -12552
rect -18576 -12632 -18560 -12568
rect -18496 -12632 -18480 -12568
rect -18576 -12648 -18480 -12632
rect -19988 -12748 -19892 -12712
rect -18576 -12712 -18560 -12648
rect -18496 -12712 -18480 -12648
rect -18157 -11968 -17435 -11959
rect -18157 -12672 -18148 -11968
rect -17444 -12672 -17435 -11968
rect -18157 -12681 -17435 -12672
rect -17164 -11992 -17148 -11928
rect -17084 -11992 -17068 -11928
rect -15752 -11928 -15656 -11892
rect -17164 -12008 -17068 -11992
rect -17164 -12072 -17148 -12008
rect -17084 -12072 -17068 -12008
rect -17164 -12088 -17068 -12072
rect -17164 -12152 -17148 -12088
rect -17084 -12152 -17068 -12088
rect -17164 -12168 -17068 -12152
rect -17164 -12232 -17148 -12168
rect -17084 -12232 -17068 -12168
rect -17164 -12248 -17068 -12232
rect -17164 -12312 -17148 -12248
rect -17084 -12312 -17068 -12248
rect -17164 -12328 -17068 -12312
rect -17164 -12392 -17148 -12328
rect -17084 -12392 -17068 -12328
rect -17164 -12408 -17068 -12392
rect -17164 -12472 -17148 -12408
rect -17084 -12472 -17068 -12408
rect -17164 -12488 -17068 -12472
rect -17164 -12552 -17148 -12488
rect -17084 -12552 -17068 -12488
rect -17164 -12568 -17068 -12552
rect -17164 -12632 -17148 -12568
rect -17084 -12632 -17068 -12568
rect -17164 -12648 -17068 -12632
rect -18576 -12748 -18480 -12712
rect -17164 -12712 -17148 -12648
rect -17084 -12712 -17068 -12648
rect -16745 -11968 -16023 -11959
rect -16745 -12672 -16736 -11968
rect -16032 -12672 -16023 -11968
rect -16745 -12681 -16023 -12672
rect -15752 -11992 -15736 -11928
rect -15672 -11992 -15656 -11928
rect -14340 -11928 -14244 -11892
rect -15752 -12008 -15656 -11992
rect -15752 -12072 -15736 -12008
rect -15672 -12072 -15656 -12008
rect -15752 -12088 -15656 -12072
rect -15752 -12152 -15736 -12088
rect -15672 -12152 -15656 -12088
rect -15752 -12168 -15656 -12152
rect -15752 -12232 -15736 -12168
rect -15672 -12232 -15656 -12168
rect -15752 -12248 -15656 -12232
rect -15752 -12312 -15736 -12248
rect -15672 -12312 -15656 -12248
rect -15752 -12328 -15656 -12312
rect -15752 -12392 -15736 -12328
rect -15672 -12392 -15656 -12328
rect -15752 -12408 -15656 -12392
rect -15752 -12472 -15736 -12408
rect -15672 -12472 -15656 -12408
rect -15752 -12488 -15656 -12472
rect -15752 -12552 -15736 -12488
rect -15672 -12552 -15656 -12488
rect -15752 -12568 -15656 -12552
rect -15752 -12632 -15736 -12568
rect -15672 -12632 -15656 -12568
rect -15752 -12648 -15656 -12632
rect -17164 -12748 -17068 -12712
rect -15752 -12712 -15736 -12648
rect -15672 -12712 -15656 -12648
rect -15333 -11968 -14611 -11959
rect -15333 -12672 -15324 -11968
rect -14620 -12672 -14611 -11968
rect -15333 -12681 -14611 -12672
rect -14340 -11992 -14324 -11928
rect -14260 -11992 -14244 -11928
rect -12928 -11928 -12832 -11892
rect -14340 -12008 -14244 -11992
rect -14340 -12072 -14324 -12008
rect -14260 -12072 -14244 -12008
rect -14340 -12088 -14244 -12072
rect -14340 -12152 -14324 -12088
rect -14260 -12152 -14244 -12088
rect -14340 -12168 -14244 -12152
rect -14340 -12232 -14324 -12168
rect -14260 -12232 -14244 -12168
rect -14340 -12248 -14244 -12232
rect -14340 -12312 -14324 -12248
rect -14260 -12312 -14244 -12248
rect -14340 -12328 -14244 -12312
rect -14340 -12392 -14324 -12328
rect -14260 -12392 -14244 -12328
rect -14340 -12408 -14244 -12392
rect -14340 -12472 -14324 -12408
rect -14260 -12472 -14244 -12408
rect -14340 -12488 -14244 -12472
rect -14340 -12552 -14324 -12488
rect -14260 -12552 -14244 -12488
rect -14340 -12568 -14244 -12552
rect -14340 -12632 -14324 -12568
rect -14260 -12632 -14244 -12568
rect -14340 -12648 -14244 -12632
rect -15752 -12748 -15656 -12712
rect -14340 -12712 -14324 -12648
rect -14260 -12712 -14244 -12648
rect -13921 -11968 -13199 -11959
rect -13921 -12672 -13912 -11968
rect -13208 -12672 -13199 -11968
rect -13921 -12681 -13199 -12672
rect -12928 -11992 -12912 -11928
rect -12848 -11992 -12832 -11928
rect -11516 -11928 -11420 -11892
rect -12928 -12008 -12832 -11992
rect -12928 -12072 -12912 -12008
rect -12848 -12072 -12832 -12008
rect -12928 -12088 -12832 -12072
rect -12928 -12152 -12912 -12088
rect -12848 -12152 -12832 -12088
rect -12928 -12168 -12832 -12152
rect -12928 -12232 -12912 -12168
rect -12848 -12232 -12832 -12168
rect -12928 -12248 -12832 -12232
rect -12928 -12312 -12912 -12248
rect -12848 -12312 -12832 -12248
rect -12928 -12328 -12832 -12312
rect -12928 -12392 -12912 -12328
rect -12848 -12392 -12832 -12328
rect -12928 -12408 -12832 -12392
rect -12928 -12472 -12912 -12408
rect -12848 -12472 -12832 -12408
rect -12928 -12488 -12832 -12472
rect -12928 -12552 -12912 -12488
rect -12848 -12552 -12832 -12488
rect -12928 -12568 -12832 -12552
rect -12928 -12632 -12912 -12568
rect -12848 -12632 -12832 -12568
rect -12928 -12648 -12832 -12632
rect -14340 -12748 -14244 -12712
rect -12928 -12712 -12912 -12648
rect -12848 -12712 -12832 -12648
rect -12509 -11968 -11787 -11959
rect -12509 -12672 -12500 -11968
rect -11796 -12672 -11787 -11968
rect -12509 -12681 -11787 -12672
rect -11516 -11992 -11500 -11928
rect -11436 -11992 -11420 -11928
rect -10104 -11928 -10008 -11892
rect -11516 -12008 -11420 -11992
rect -11516 -12072 -11500 -12008
rect -11436 -12072 -11420 -12008
rect -11516 -12088 -11420 -12072
rect -11516 -12152 -11500 -12088
rect -11436 -12152 -11420 -12088
rect -11516 -12168 -11420 -12152
rect -11516 -12232 -11500 -12168
rect -11436 -12232 -11420 -12168
rect -11516 -12248 -11420 -12232
rect -11516 -12312 -11500 -12248
rect -11436 -12312 -11420 -12248
rect -11516 -12328 -11420 -12312
rect -11516 -12392 -11500 -12328
rect -11436 -12392 -11420 -12328
rect -11516 -12408 -11420 -12392
rect -11516 -12472 -11500 -12408
rect -11436 -12472 -11420 -12408
rect -11516 -12488 -11420 -12472
rect -11516 -12552 -11500 -12488
rect -11436 -12552 -11420 -12488
rect -11516 -12568 -11420 -12552
rect -11516 -12632 -11500 -12568
rect -11436 -12632 -11420 -12568
rect -11516 -12648 -11420 -12632
rect -12928 -12748 -12832 -12712
rect -11516 -12712 -11500 -12648
rect -11436 -12712 -11420 -12648
rect -11097 -11968 -10375 -11959
rect -11097 -12672 -11088 -11968
rect -10384 -12672 -10375 -11968
rect -11097 -12681 -10375 -12672
rect -10104 -11992 -10088 -11928
rect -10024 -11992 -10008 -11928
rect -8692 -11928 -8596 -11892
rect -10104 -12008 -10008 -11992
rect -10104 -12072 -10088 -12008
rect -10024 -12072 -10008 -12008
rect -10104 -12088 -10008 -12072
rect -10104 -12152 -10088 -12088
rect -10024 -12152 -10008 -12088
rect -10104 -12168 -10008 -12152
rect -10104 -12232 -10088 -12168
rect -10024 -12232 -10008 -12168
rect -10104 -12248 -10008 -12232
rect -10104 -12312 -10088 -12248
rect -10024 -12312 -10008 -12248
rect -10104 -12328 -10008 -12312
rect -10104 -12392 -10088 -12328
rect -10024 -12392 -10008 -12328
rect -10104 -12408 -10008 -12392
rect -10104 -12472 -10088 -12408
rect -10024 -12472 -10008 -12408
rect -10104 -12488 -10008 -12472
rect -10104 -12552 -10088 -12488
rect -10024 -12552 -10008 -12488
rect -10104 -12568 -10008 -12552
rect -10104 -12632 -10088 -12568
rect -10024 -12632 -10008 -12568
rect -10104 -12648 -10008 -12632
rect -11516 -12748 -11420 -12712
rect -10104 -12712 -10088 -12648
rect -10024 -12712 -10008 -12648
rect -9685 -11968 -8963 -11959
rect -9685 -12672 -9676 -11968
rect -8972 -12672 -8963 -11968
rect -9685 -12681 -8963 -12672
rect -8692 -11992 -8676 -11928
rect -8612 -11992 -8596 -11928
rect -7280 -11928 -7184 -11892
rect -8692 -12008 -8596 -11992
rect -8692 -12072 -8676 -12008
rect -8612 -12072 -8596 -12008
rect -8692 -12088 -8596 -12072
rect -8692 -12152 -8676 -12088
rect -8612 -12152 -8596 -12088
rect -8692 -12168 -8596 -12152
rect -8692 -12232 -8676 -12168
rect -8612 -12232 -8596 -12168
rect -8692 -12248 -8596 -12232
rect -8692 -12312 -8676 -12248
rect -8612 -12312 -8596 -12248
rect -8692 -12328 -8596 -12312
rect -8692 -12392 -8676 -12328
rect -8612 -12392 -8596 -12328
rect -8692 -12408 -8596 -12392
rect -8692 -12472 -8676 -12408
rect -8612 -12472 -8596 -12408
rect -8692 -12488 -8596 -12472
rect -8692 -12552 -8676 -12488
rect -8612 -12552 -8596 -12488
rect -8692 -12568 -8596 -12552
rect -8692 -12632 -8676 -12568
rect -8612 -12632 -8596 -12568
rect -8692 -12648 -8596 -12632
rect -10104 -12748 -10008 -12712
rect -8692 -12712 -8676 -12648
rect -8612 -12712 -8596 -12648
rect -8273 -11968 -7551 -11959
rect -8273 -12672 -8264 -11968
rect -7560 -12672 -7551 -11968
rect -8273 -12681 -7551 -12672
rect -7280 -11992 -7264 -11928
rect -7200 -11992 -7184 -11928
rect -5868 -11928 -5772 -11892
rect -7280 -12008 -7184 -11992
rect -7280 -12072 -7264 -12008
rect -7200 -12072 -7184 -12008
rect -7280 -12088 -7184 -12072
rect -7280 -12152 -7264 -12088
rect -7200 -12152 -7184 -12088
rect -7280 -12168 -7184 -12152
rect -7280 -12232 -7264 -12168
rect -7200 -12232 -7184 -12168
rect -7280 -12248 -7184 -12232
rect -7280 -12312 -7264 -12248
rect -7200 -12312 -7184 -12248
rect -7280 -12328 -7184 -12312
rect -7280 -12392 -7264 -12328
rect -7200 -12392 -7184 -12328
rect -7280 -12408 -7184 -12392
rect -7280 -12472 -7264 -12408
rect -7200 -12472 -7184 -12408
rect -7280 -12488 -7184 -12472
rect -7280 -12552 -7264 -12488
rect -7200 -12552 -7184 -12488
rect -7280 -12568 -7184 -12552
rect -7280 -12632 -7264 -12568
rect -7200 -12632 -7184 -12568
rect -7280 -12648 -7184 -12632
rect -8692 -12748 -8596 -12712
rect -7280 -12712 -7264 -12648
rect -7200 -12712 -7184 -12648
rect -6861 -11968 -6139 -11959
rect -6861 -12672 -6852 -11968
rect -6148 -12672 -6139 -11968
rect -6861 -12681 -6139 -12672
rect -5868 -11992 -5852 -11928
rect -5788 -11992 -5772 -11928
rect -4456 -11928 -4360 -11892
rect -5868 -12008 -5772 -11992
rect -5868 -12072 -5852 -12008
rect -5788 -12072 -5772 -12008
rect -5868 -12088 -5772 -12072
rect -5868 -12152 -5852 -12088
rect -5788 -12152 -5772 -12088
rect -5868 -12168 -5772 -12152
rect -5868 -12232 -5852 -12168
rect -5788 -12232 -5772 -12168
rect -5868 -12248 -5772 -12232
rect -5868 -12312 -5852 -12248
rect -5788 -12312 -5772 -12248
rect -5868 -12328 -5772 -12312
rect -5868 -12392 -5852 -12328
rect -5788 -12392 -5772 -12328
rect -5868 -12408 -5772 -12392
rect -5868 -12472 -5852 -12408
rect -5788 -12472 -5772 -12408
rect -5868 -12488 -5772 -12472
rect -5868 -12552 -5852 -12488
rect -5788 -12552 -5772 -12488
rect -5868 -12568 -5772 -12552
rect -5868 -12632 -5852 -12568
rect -5788 -12632 -5772 -12568
rect -5868 -12648 -5772 -12632
rect -7280 -12748 -7184 -12712
rect -5868 -12712 -5852 -12648
rect -5788 -12712 -5772 -12648
rect -5449 -11968 -4727 -11959
rect -5449 -12672 -5440 -11968
rect -4736 -12672 -4727 -11968
rect -5449 -12681 -4727 -12672
rect -4456 -11992 -4440 -11928
rect -4376 -11992 -4360 -11928
rect -3044 -11928 -2948 -11892
rect -4456 -12008 -4360 -11992
rect -4456 -12072 -4440 -12008
rect -4376 -12072 -4360 -12008
rect -4456 -12088 -4360 -12072
rect -4456 -12152 -4440 -12088
rect -4376 -12152 -4360 -12088
rect -4456 -12168 -4360 -12152
rect -4456 -12232 -4440 -12168
rect -4376 -12232 -4360 -12168
rect -4456 -12248 -4360 -12232
rect -4456 -12312 -4440 -12248
rect -4376 -12312 -4360 -12248
rect -4456 -12328 -4360 -12312
rect -4456 -12392 -4440 -12328
rect -4376 -12392 -4360 -12328
rect -4456 -12408 -4360 -12392
rect -4456 -12472 -4440 -12408
rect -4376 -12472 -4360 -12408
rect -4456 -12488 -4360 -12472
rect -4456 -12552 -4440 -12488
rect -4376 -12552 -4360 -12488
rect -4456 -12568 -4360 -12552
rect -4456 -12632 -4440 -12568
rect -4376 -12632 -4360 -12568
rect -4456 -12648 -4360 -12632
rect -5868 -12748 -5772 -12712
rect -4456 -12712 -4440 -12648
rect -4376 -12712 -4360 -12648
rect -4037 -11968 -3315 -11959
rect -4037 -12672 -4028 -11968
rect -3324 -12672 -3315 -11968
rect -4037 -12681 -3315 -12672
rect -3044 -11992 -3028 -11928
rect -2964 -11992 -2948 -11928
rect -1632 -11928 -1536 -11892
rect -3044 -12008 -2948 -11992
rect -3044 -12072 -3028 -12008
rect -2964 -12072 -2948 -12008
rect -3044 -12088 -2948 -12072
rect -3044 -12152 -3028 -12088
rect -2964 -12152 -2948 -12088
rect -3044 -12168 -2948 -12152
rect -3044 -12232 -3028 -12168
rect -2964 -12232 -2948 -12168
rect -3044 -12248 -2948 -12232
rect -3044 -12312 -3028 -12248
rect -2964 -12312 -2948 -12248
rect -3044 -12328 -2948 -12312
rect -3044 -12392 -3028 -12328
rect -2964 -12392 -2948 -12328
rect -3044 -12408 -2948 -12392
rect -3044 -12472 -3028 -12408
rect -2964 -12472 -2948 -12408
rect -3044 -12488 -2948 -12472
rect -3044 -12552 -3028 -12488
rect -2964 -12552 -2948 -12488
rect -3044 -12568 -2948 -12552
rect -3044 -12632 -3028 -12568
rect -2964 -12632 -2948 -12568
rect -3044 -12648 -2948 -12632
rect -4456 -12748 -4360 -12712
rect -3044 -12712 -3028 -12648
rect -2964 -12712 -2948 -12648
rect -2625 -11968 -1903 -11959
rect -2625 -12672 -2616 -11968
rect -1912 -12672 -1903 -11968
rect -2625 -12681 -1903 -12672
rect -1632 -11992 -1616 -11928
rect -1552 -11992 -1536 -11928
rect -220 -11928 -124 -11892
rect -1632 -12008 -1536 -11992
rect -1632 -12072 -1616 -12008
rect -1552 -12072 -1536 -12008
rect -1632 -12088 -1536 -12072
rect -1632 -12152 -1616 -12088
rect -1552 -12152 -1536 -12088
rect -1632 -12168 -1536 -12152
rect -1632 -12232 -1616 -12168
rect -1552 -12232 -1536 -12168
rect -1632 -12248 -1536 -12232
rect -1632 -12312 -1616 -12248
rect -1552 -12312 -1536 -12248
rect -1632 -12328 -1536 -12312
rect -1632 -12392 -1616 -12328
rect -1552 -12392 -1536 -12328
rect -1632 -12408 -1536 -12392
rect -1632 -12472 -1616 -12408
rect -1552 -12472 -1536 -12408
rect -1632 -12488 -1536 -12472
rect -1632 -12552 -1616 -12488
rect -1552 -12552 -1536 -12488
rect -1632 -12568 -1536 -12552
rect -1632 -12632 -1616 -12568
rect -1552 -12632 -1536 -12568
rect -1632 -12648 -1536 -12632
rect -3044 -12748 -2948 -12712
rect -1632 -12712 -1616 -12648
rect -1552 -12712 -1536 -12648
rect -1213 -11968 -491 -11959
rect -1213 -12672 -1204 -11968
rect -500 -12672 -491 -11968
rect -1213 -12681 -491 -12672
rect -220 -11992 -204 -11928
rect -140 -11992 -124 -11928
rect 1192 -11928 1288 -11892
rect -220 -12008 -124 -11992
rect -220 -12072 -204 -12008
rect -140 -12072 -124 -12008
rect -220 -12088 -124 -12072
rect -220 -12152 -204 -12088
rect -140 -12152 -124 -12088
rect -220 -12168 -124 -12152
rect -220 -12232 -204 -12168
rect -140 -12232 -124 -12168
rect -220 -12248 -124 -12232
rect -220 -12312 -204 -12248
rect -140 -12312 -124 -12248
rect -220 -12328 -124 -12312
rect -220 -12392 -204 -12328
rect -140 -12392 -124 -12328
rect -220 -12408 -124 -12392
rect -220 -12472 -204 -12408
rect -140 -12472 -124 -12408
rect -220 -12488 -124 -12472
rect -220 -12552 -204 -12488
rect -140 -12552 -124 -12488
rect -220 -12568 -124 -12552
rect -220 -12632 -204 -12568
rect -140 -12632 -124 -12568
rect -220 -12648 -124 -12632
rect -1632 -12748 -1536 -12712
rect -220 -12712 -204 -12648
rect -140 -12712 -124 -12648
rect 199 -11968 921 -11959
rect 199 -12672 208 -11968
rect 912 -12672 921 -11968
rect 199 -12681 921 -12672
rect 1192 -11992 1208 -11928
rect 1272 -11992 1288 -11928
rect 2604 -11928 2700 -11892
rect 1192 -12008 1288 -11992
rect 1192 -12072 1208 -12008
rect 1272 -12072 1288 -12008
rect 1192 -12088 1288 -12072
rect 1192 -12152 1208 -12088
rect 1272 -12152 1288 -12088
rect 1192 -12168 1288 -12152
rect 1192 -12232 1208 -12168
rect 1272 -12232 1288 -12168
rect 1192 -12248 1288 -12232
rect 1192 -12312 1208 -12248
rect 1272 -12312 1288 -12248
rect 1192 -12328 1288 -12312
rect 1192 -12392 1208 -12328
rect 1272 -12392 1288 -12328
rect 1192 -12408 1288 -12392
rect 1192 -12472 1208 -12408
rect 1272 -12472 1288 -12408
rect 1192 -12488 1288 -12472
rect 1192 -12552 1208 -12488
rect 1272 -12552 1288 -12488
rect 1192 -12568 1288 -12552
rect 1192 -12632 1208 -12568
rect 1272 -12632 1288 -12568
rect 1192 -12648 1288 -12632
rect -220 -12748 -124 -12712
rect 1192 -12712 1208 -12648
rect 1272 -12712 1288 -12648
rect 1611 -11968 2333 -11959
rect 1611 -12672 1620 -11968
rect 2324 -12672 2333 -11968
rect 1611 -12681 2333 -12672
rect 2604 -11992 2620 -11928
rect 2684 -11992 2700 -11928
rect 4016 -11928 4112 -11892
rect 2604 -12008 2700 -11992
rect 2604 -12072 2620 -12008
rect 2684 -12072 2700 -12008
rect 2604 -12088 2700 -12072
rect 2604 -12152 2620 -12088
rect 2684 -12152 2700 -12088
rect 2604 -12168 2700 -12152
rect 2604 -12232 2620 -12168
rect 2684 -12232 2700 -12168
rect 2604 -12248 2700 -12232
rect 2604 -12312 2620 -12248
rect 2684 -12312 2700 -12248
rect 2604 -12328 2700 -12312
rect 2604 -12392 2620 -12328
rect 2684 -12392 2700 -12328
rect 2604 -12408 2700 -12392
rect 2604 -12472 2620 -12408
rect 2684 -12472 2700 -12408
rect 2604 -12488 2700 -12472
rect 2604 -12552 2620 -12488
rect 2684 -12552 2700 -12488
rect 2604 -12568 2700 -12552
rect 2604 -12632 2620 -12568
rect 2684 -12632 2700 -12568
rect 2604 -12648 2700 -12632
rect 1192 -12748 1288 -12712
rect 2604 -12712 2620 -12648
rect 2684 -12712 2700 -12648
rect 3023 -11968 3745 -11959
rect 3023 -12672 3032 -11968
rect 3736 -12672 3745 -11968
rect 3023 -12681 3745 -12672
rect 4016 -11992 4032 -11928
rect 4096 -11992 4112 -11928
rect 5428 -11928 5524 -11892
rect 4016 -12008 4112 -11992
rect 4016 -12072 4032 -12008
rect 4096 -12072 4112 -12008
rect 4016 -12088 4112 -12072
rect 4016 -12152 4032 -12088
rect 4096 -12152 4112 -12088
rect 4016 -12168 4112 -12152
rect 4016 -12232 4032 -12168
rect 4096 -12232 4112 -12168
rect 4016 -12248 4112 -12232
rect 4016 -12312 4032 -12248
rect 4096 -12312 4112 -12248
rect 4016 -12328 4112 -12312
rect 4016 -12392 4032 -12328
rect 4096 -12392 4112 -12328
rect 4016 -12408 4112 -12392
rect 4016 -12472 4032 -12408
rect 4096 -12472 4112 -12408
rect 4016 -12488 4112 -12472
rect 4016 -12552 4032 -12488
rect 4096 -12552 4112 -12488
rect 4016 -12568 4112 -12552
rect 4016 -12632 4032 -12568
rect 4096 -12632 4112 -12568
rect 4016 -12648 4112 -12632
rect 2604 -12748 2700 -12712
rect 4016 -12712 4032 -12648
rect 4096 -12712 4112 -12648
rect 4435 -11968 5157 -11959
rect 4435 -12672 4444 -11968
rect 5148 -12672 5157 -11968
rect 4435 -12681 5157 -12672
rect 5428 -11992 5444 -11928
rect 5508 -11992 5524 -11928
rect 6840 -11928 6936 -11892
rect 5428 -12008 5524 -11992
rect 5428 -12072 5444 -12008
rect 5508 -12072 5524 -12008
rect 5428 -12088 5524 -12072
rect 5428 -12152 5444 -12088
rect 5508 -12152 5524 -12088
rect 5428 -12168 5524 -12152
rect 5428 -12232 5444 -12168
rect 5508 -12232 5524 -12168
rect 5428 -12248 5524 -12232
rect 5428 -12312 5444 -12248
rect 5508 -12312 5524 -12248
rect 5428 -12328 5524 -12312
rect 5428 -12392 5444 -12328
rect 5508 -12392 5524 -12328
rect 5428 -12408 5524 -12392
rect 5428 -12472 5444 -12408
rect 5508 -12472 5524 -12408
rect 5428 -12488 5524 -12472
rect 5428 -12552 5444 -12488
rect 5508 -12552 5524 -12488
rect 5428 -12568 5524 -12552
rect 5428 -12632 5444 -12568
rect 5508 -12632 5524 -12568
rect 5428 -12648 5524 -12632
rect 4016 -12748 4112 -12712
rect 5428 -12712 5444 -12648
rect 5508 -12712 5524 -12648
rect 5847 -11968 6569 -11959
rect 5847 -12672 5856 -11968
rect 6560 -12672 6569 -11968
rect 5847 -12681 6569 -12672
rect 6840 -11992 6856 -11928
rect 6920 -11992 6936 -11928
rect 8252 -11928 8348 -11892
rect 6840 -12008 6936 -11992
rect 6840 -12072 6856 -12008
rect 6920 -12072 6936 -12008
rect 6840 -12088 6936 -12072
rect 6840 -12152 6856 -12088
rect 6920 -12152 6936 -12088
rect 6840 -12168 6936 -12152
rect 6840 -12232 6856 -12168
rect 6920 -12232 6936 -12168
rect 6840 -12248 6936 -12232
rect 6840 -12312 6856 -12248
rect 6920 -12312 6936 -12248
rect 6840 -12328 6936 -12312
rect 6840 -12392 6856 -12328
rect 6920 -12392 6936 -12328
rect 6840 -12408 6936 -12392
rect 6840 -12472 6856 -12408
rect 6920 -12472 6936 -12408
rect 6840 -12488 6936 -12472
rect 6840 -12552 6856 -12488
rect 6920 -12552 6936 -12488
rect 6840 -12568 6936 -12552
rect 6840 -12632 6856 -12568
rect 6920 -12632 6936 -12568
rect 6840 -12648 6936 -12632
rect 5428 -12748 5524 -12712
rect 6840 -12712 6856 -12648
rect 6920 -12712 6936 -12648
rect 7259 -11968 7981 -11959
rect 7259 -12672 7268 -11968
rect 7972 -12672 7981 -11968
rect 7259 -12681 7981 -12672
rect 8252 -11992 8268 -11928
rect 8332 -11992 8348 -11928
rect 9664 -11928 9760 -11892
rect 8252 -12008 8348 -11992
rect 8252 -12072 8268 -12008
rect 8332 -12072 8348 -12008
rect 8252 -12088 8348 -12072
rect 8252 -12152 8268 -12088
rect 8332 -12152 8348 -12088
rect 8252 -12168 8348 -12152
rect 8252 -12232 8268 -12168
rect 8332 -12232 8348 -12168
rect 8252 -12248 8348 -12232
rect 8252 -12312 8268 -12248
rect 8332 -12312 8348 -12248
rect 8252 -12328 8348 -12312
rect 8252 -12392 8268 -12328
rect 8332 -12392 8348 -12328
rect 8252 -12408 8348 -12392
rect 8252 -12472 8268 -12408
rect 8332 -12472 8348 -12408
rect 8252 -12488 8348 -12472
rect 8252 -12552 8268 -12488
rect 8332 -12552 8348 -12488
rect 8252 -12568 8348 -12552
rect 8252 -12632 8268 -12568
rect 8332 -12632 8348 -12568
rect 8252 -12648 8348 -12632
rect 6840 -12748 6936 -12712
rect 8252 -12712 8268 -12648
rect 8332 -12712 8348 -12648
rect 8671 -11968 9393 -11959
rect 8671 -12672 8680 -11968
rect 9384 -12672 9393 -11968
rect 8671 -12681 9393 -12672
rect 9664 -11992 9680 -11928
rect 9744 -11992 9760 -11928
rect 11076 -11928 11172 -11892
rect 9664 -12008 9760 -11992
rect 9664 -12072 9680 -12008
rect 9744 -12072 9760 -12008
rect 9664 -12088 9760 -12072
rect 9664 -12152 9680 -12088
rect 9744 -12152 9760 -12088
rect 9664 -12168 9760 -12152
rect 9664 -12232 9680 -12168
rect 9744 -12232 9760 -12168
rect 9664 -12248 9760 -12232
rect 9664 -12312 9680 -12248
rect 9744 -12312 9760 -12248
rect 9664 -12328 9760 -12312
rect 9664 -12392 9680 -12328
rect 9744 -12392 9760 -12328
rect 9664 -12408 9760 -12392
rect 9664 -12472 9680 -12408
rect 9744 -12472 9760 -12408
rect 9664 -12488 9760 -12472
rect 9664 -12552 9680 -12488
rect 9744 -12552 9760 -12488
rect 9664 -12568 9760 -12552
rect 9664 -12632 9680 -12568
rect 9744 -12632 9760 -12568
rect 9664 -12648 9760 -12632
rect 8252 -12748 8348 -12712
rect 9664 -12712 9680 -12648
rect 9744 -12712 9760 -12648
rect 10083 -11968 10805 -11959
rect 10083 -12672 10092 -11968
rect 10796 -12672 10805 -11968
rect 10083 -12681 10805 -12672
rect 11076 -11992 11092 -11928
rect 11156 -11992 11172 -11928
rect 12488 -11928 12584 -11892
rect 11076 -12008 11172 -11992
rect 11076 -12072 11092 -12008
rect 11156 -12072 11172 -12008
rect 11076 -12088 11172 -12072
rect 11076 -12152 11092 -12088
rect 11156 -12152 11172 -12088
rect 11076 -12168 11172 -12152
rect 11076 -12232 11092 -12168
rect 11156 -12232 11172 -12168
rect 11076 -12248 11172 -12232
rect 11076 -12312 11092 -12248
rect 11156 -12312 11172 -12248
rect 11076 -12328 11172 -12312
rect 11076 -12392 11092 -12328
rect 11156 -12392 11172 -12328
rect 11076 -12408 11172 -12392
rect 11076 -12472 11092 -12408
rect 11156 -12472 11172 -12408
rect 11076 -12488 11172 -12472
rect 11076 -12552 11092 -12488
rect 11156 -12552 11172 -12488
rect 11076 -12568 11172 -12552
rect 11076 -12632 11092 -12568
rect 11156 -12632 11172 -12568
rect 11076 -12648 11172 -12632
rect 9664 -12748 9760 -12712
rect 11076 -12712 11092 -12648
rect 11156 -12712 11172 -12648
rect 11495 -11968 12217 -11959
rect 11495 -12672 11504 -11968
rect 12208 -12672 12217 -11968
rect 11495 -12681 12217 -12672
rect 12488 -11992 12504 -11928
rect 12568 -11992 12584 -11928
rect 13900 -11928 13996 -11892
rect 12488 -12008 12584 -11992
rect 12488 -12072 12504 -12008
rect 12568 -12072 12584 -12008
rect 12488 -12088 12584 -12072
rect 12488 -12152 12504 -12088
rect 12568 -12152 12584 -12088
rect 12488 -12168 12584 -12152
rect 12488 -12232 12504 -12168
rect 12568 -12232 12584 -12168
rect 12488 -12248 12584 -12232
rect 12488 -12312 12504 -12248
rect 12568 -12312 12584 -12248
rect 12488 -12328 12584 -12312
rect 12488 -12392 12504 -12328
rect 12568 -12392 12584 -12328
rect 12488 -12408 12584 -12392
rect 12488 -12472 12504 -12408
rect 12568 -12472 12584 -12408
rect 12488 -12488 12584 -12472
rect 12488 -12552 12504 -12488
rect 12568 -12552 12584 -12488
rect 12488 -12568 12584 -12552
rect 12488 -12632 12504 -12568
rect 12568 -12632 12584 -12568
rect 12488 -12648 12584 -12632
rect 11076 -12748 11172 -12712
rect 12488 -12712 12504 -12648
rect 12568 -12712 12584 -12648
rect 12907 -11968 13629 -11959
rect 12907 -12672 12916 -11968
rect 13620 -12672 13629 -11968
rect 12907 -12681 13629 -12672
rect 13900 -11992 13916 -11928
rect 13980 -11992 13996 -11928
rect 15312 -11928 15408 -11892
rect 13900 -12008 13996 -11992
rect 13900 -12072 13916 -12008
rect 13980 -12072 13996 -12008
rect 13900 -12088 13996 -12072
rect 13900 -12152 13916 -12088
rect 13980 -12152 13996 -12088
rect 13900 -12168 13996 -12152
rect 13900 -12232 13916 -12168
rect 13980 -12232 13996 -12168
rect 13900 -12248 13996 -12232
rect 13900 -12312 13916 -12248
rect 13980 -12312 13996 -12248
rect 13900 -12328 13996 -12312
rect 13900 -12392 13916 -12328
rect 13980 -12392 13996 -12328
rect 13900 -12408 13996 -12392
rect 13900 -12472 13916 -12408
rect 13980 -12472 13996 -12408
rect 13900 -12488 13996 -12472
rect 13900 -12552 13916 -12488
rect 13980 -12552 13996 -12488
rect 13900 -12568 13996 -12552
rect 13900 -12632 13916 -12568
rect 13980 -12632 13996 -12568
rect 13900 -12648 13996 -12632
rect 12488 -12748 12584 -12712
rect 13900 -12712 13916 -12648
rect 13980 -12712 13996 -12648
rect 14319 -11968 15041 -11959
rect 14319 -12672 14328 -11968
rect 15032 -12672 15041 -11968
rect 14319 -12681 15041 -12672
rect 15312 -11992 15328 -11928
rect 15392 -11992 15408 -11928
rect 16724 -11928 16820 -11892
rect 15312 -12008 15408 -11992
rect 15312 -12072 15328 -12008
rect 15392 -12072 15408 -12008
rect 15312 -12088 15408 -12072
rect 15312 -12152 15328 -12088
rect 15392 -12152 15408 -12088
rect 15312 -12168 15408 -12152
rect 15312 -12232 15328 -12168
rect 15392 -12232 15408 -12168
rect 15312 -12248 15408 -12232
rect 15312 -12312 15328 -12248
rect 15392 -12312 15408 -12248
rect 15312 -12328 15408 -12312
rect 15312 -12392 15328 -12328
rect 15392 -12392 15408 -12328
rect 15312 -12408 15408 -12392
rect 15312 -12472 15328 -12408
rect 15392 -12472 15408 -12408
rect 15312 -12488 15408 -12472
rect 15312 -12552 15328 -12488
rect 15392 -12552 15408 -12488
rect 15312 -12568 15408 -12552
rect 15312 -12632 15328 -12568
rect 15392 -12632 15408 -12568
rect 15312 -12648 15408 -12632
rect 13900 -12748 13996 -12712
rect 15312 -12712 15328 -12648
rect 15392 -12712 15408 -12648
rect 15731 -11968 16453 -11959
rect 15731 -12672 15740 -11968
rect 16444 -12672 16453 -11968
rect 15731 -12681 16453 -12672
rect 16724 -11992 16740 -11928
rect 16804 -11992 16820 -11928
rect 18136 -11928 18232 -11892
rect 16724 -12008 16820 -11992
rect 16724 -12072 16740 -12008
rect 16804 -12072 16820 -12008
rect 16724 -12088 16820 -12072
rect 16724 -12152 16740 -12088
rect 16804 -12152 16820 -12088
rect 16724 -12168 16820 -12152
rect 16724 -12232 16740 -12168
rect 16804 -12232 16820 -12168
rect 16724 -12248 16820 -12232
rect 16724 -12312 16740 -12248
rect 16804 -12312 16820 -12248
rect 16724 -12328 16820 -12312
rect 16724 -12392 16740 -12328
rect 16804 -12392 16820 -12328
rect 16724 -12408 16820 -12392
rect 16724 -12472 16740 -12408
rect 16804 -12472 16820 -12408
rect 16724 -12488 16820 -12472
rect 16724 -12552 16740 -12488
rect 16804 -12552 16820 -12488
rect 16724 -12568 16820 -12552
rect 16724 -12632 16740 -12568
rect 16804 -12632 16820 -12568
rect 16724 -12648 16820 -12632
rect 15312 -12748 15408 -12712
rect 16724 -12712 16740 -12648
rect 16804 -12712 16820 -12648
rect 17143 -11968 17865 -11959
rect 17143 -12672 17152 -11968
rect 17856 -12672 17865 -11968
rect 17143 -12681 17865 -12672
rect 18136 -11992 18152 -11928
rect 18216 -11992 18232 -11928
rect 19548 -11928 19644 -11892
rect 18136 -12008 18232 -11992
rect 18136 -12072 18152 -12008
rect 18216 -12072 18232 -12008
rect 18136 -12088 18232 -12072
rect 18136 -12152 18152 -12088
rect 18216 -12152 18232 -12088
rect 18136 -12168 18232 -12152
rect 18136 -12232 18152 -12168
rect 18216 -12232 18232 -12168
rect 18136 -12248 18232 -12232
rect 18136 -12312 18152 -12248
rect 18216 -12312 18232 -12248
rect 18136 -12328 18232 -12312
rect 18136 -12392 18152 -12328
rect 18216 -12392 18232 -12328
rect 18136 -12408 18232 -12392
rect 18136 -12472 18152 -12408
rect 18216 -12472 18232 -12408
rect 18136 -12488 18232 -12472
rect 18136 -12552 18152 -12488
rect 18216 -12552 18232 -12488
rect 18136 -12568 18232 -12552
rect 18136 -12632 18152 -12568
rect 18216 -12632 18232 -12568
rect 18136 -12648 18232 -12632
rect 16724 -12748 16820 -12712
rect 18136 -12712 18152 -12648
rect 18216 -12712 18232 -12648
rect 18555 -11968 19277 -11959
rect 18555 -12672 18564 -11968
rect 19268 -12672 19277 -11968
rect 18555 -12681 19277 -12672
rect 19548 -11992 19564 -11928
rect 19628 -11992 19644 -11928
rect 20960 -11928 21056 -11892
rect 19548 -12008 19644 -11992
rect 19548 -12072 19564 -12008
rect 19628 -12072 19644 -12008
rect 19548 -12088 19644 -12072
rect 19548 -12152 19564 -12088
rect 19628 -12152 19644 -12088
rect 19548 -12168 19644 -12152
rect 19548 -12232 19564 -12168
rect 19628 -12232 19644 -12168
rect 19548 -12248 19644 -12232
rect 19548 -12312 19564 -12248
rect 19628 -12312 19644 -12248
rect 19548 -12328 19644 -12312
rect 19548 -12392 19564 -12328
rect 19628 -12392 19644 -12328
rect 19548 -12408 19644 -12392
rect 19548 -12472 19564 -12408
rect 19628 -12472 19644 -12408
rect 19548 -12488 19644 -12472
rect 19548 -12552 19564 -12488
rect 19628 -12552 19644 -12488
rect 19548 -12568 19644 -12552
rect 19548 -12632 19564 -12568
rect 19628 -12632 19644 -12568
rect 19548 -12648 19644 -12632
rect 18136 -12748 18232 -12712
rect 19548 -12712 19564 -12648
rect 19628 -12712 19644 -12648
rect 19967 -11968 20689 -11959
rect 19967 -12672 19976 -11968
rect 20680 -12672 20689 -11968
rect 19967 -12681 20689 -12672
rect 20960 -11992 20976 -11928
rect 21040 -11992 21056 -11928
rect 22372 -11928 22468 -11892
rect 20960 -12008 21056 -11992
rect 20960 -12072 20976 -12008
rect 21040 -12072 21056 -12008
rect 20960 -12088 21056 -12072
rect 20960 -12152 20976 -12088
rect 21040 -12152 21056 -12088
rect 20960 -12168 21056 -12152
rect 20960 -12232 20976 -12168
rect 21040 -12232 21056 -12168
rect 20960 -12248 21056 -12232
rect 20960 -12312 20976 -12248
rect 21040 -12312 21056 -12248
rect 20960 -12328 21056 -12312
rect 20960 -12392 20976 -12328
rect 21040 -12392 21056 -12328
rect 20960 -12408 21056 -12392
rect 20960 -12472 20976 -12408
rect 21040 -12472 21056 -12408
rect 20960 -12488 21056 -12472
rect 20960 -12552 20976 -12488
rect 21040 -12552 21056 -12488
rect 20960 -12568 21056 -12552
rect 20960 -12632 20976 -12568
rect 21040 -12632 21056 -12568
rect 20960 -12648 21056 -12632
rect 19548 -12748 19644 -12712
rect 20960 -12712 20976 -12648
rect 21040 -12712 21056 -12648
rect 21379 -11968 22101 -11959
rect 21379 -12672 21388 -11968
rect 22092 -12672 22101 -11968
rect 21379 -12681 22101 -12672
rect 22372 -11992 22388 -11928
rect 22452 -11992 22468 -11928
rect 23784 -11928 23880 -11892
rect 22372 -12008 22468 -11992
rect 22372 -12072 22388 -12008
rect 22452 -12072 22468 -12008
rect 22372 -12088 22468 -12072
rect 22372 -12152 22388 -12088
rect 22452 -12152 22468 -12088
rect 22372 -12168 22468 -12152
rect 22372 -12232 22388 -12168
rect 22452 -12232 22468 -12168
rect 22372 -12248 22468 -12232
rect 22372 -12312 22388 -12248
rect 22452 -12312 22468 -12248
rect 22372 -12328 22468 -12312
rect 22372 -12392 22388 -12328
rect 22452 -12392 22468 -12328
rect 22372 -12408 22468 -12392
rect 22372 -12472 22388 -12408
rect 22452 -12472 22468 -12408
rect 22372 -12488 22468 -12472
rect 22372 -12552 22388 -12488
rect 22452 -12552 22468 -12488
rect 22372 -12568 22468 -12552
rect 22372 -12632 22388 -12568
rect 22452 -12632 22468 -12568
rect 22372 -12648 22468 -12632
rect 20960 -12748 21056 -12712
rect 22372 -12712 22388 -12648
rect 22452 -12712 22468 -12648
rect 22791 -11968 23513 -11959
rect 22791 -12672 22800 -11968
rect 23504 -12672 23513 -11968
rect 22791 -12681 23513 -12672
rect 23784 -11992 23800 -11928
rect 23864 -11992 23880 -11928
rect 23784 -12008 23880 -11992
rect 23784 -12072 23800 -12008
rect 23864 -12072 23880 -12008
rect 23784 -12088 23880 -12072
rect 23784 -12152 23800 -12088
rect 23864 -12152 23880 -12088
rect 23784 -12168 23880 -12152
rect 23784 -12232 23800 -12168
rect 23864 -12232 23880 -12168
rect 23784 -12248 23880 -12232
rect 23784 -12312 23800 -12248
rect 23864 -12312 23880 -12248
rect 23784 -12328 23880 -12312
rect 23784 -12392 23800 -12328
rect 23864 -12392 23880 -12328
rect 23784 -12408 23880 -12392
rect 23784 -12472 23800 -12408
rect 23864 -12472 23880 -12408
rect 23784 -12488 23880 -12472
rect 23784 -12552 23800 -12488
rect 23864 -12552 23880 -12488
rect 23784 -12568 23880 -12552
rect 23784 -12632 23800 -12568
rect 23864 -12632 23880 -12568
rect 23784 -12648 23880 -12632
rect 22372 -12748 22468 -12712
rect 23784 -12712 23800 -12648
rect 23864 -12712 23880 -12648
rect 23784 -12748 23880 -12712
rect -22812 -13048 -22716 -13012
rect -23805 -13088 -23083 -13079
rect -23805 -13792 -23796 -13088
rect -23092 -13792 -23083 -13088
rect -23805 -13801 -23083 -13792
rect -22812 -13112 -22796 -13048
rect -22732 -13112 -22716 -13048
rect -21400 -13048 -21304 -13012
rect -22812 -13128 -22716 -13112
rect -22812 -13192 -22796 -13128
rect -22732 -13192 -22716 -13128
rect -22812 -13208 -22716 -13192
rect -22812 -13272 -22796 -13208
rect -22732 -13272 -22716 -13208
rect -22812 -13288 -22716 -13272
rect -22812 -13352 -22796 -13288
rect -22732 -13352 -22716 -13288
rect -22812 -13368 -22716 -13352
rect -22812 -13432 -22796 -13368
rect -22732 -13432 -22716 -13368
rect -22812 -13448 -22716 -13432
rect -22812 -13512 -22796 -13448
rect -22732 -13512 -22716 -13448
rect -22812 -13528 -22716 -13512
rect -22812 -13592 -22796 -13528
rect -22732 -13592 -22716 -13528
rect -22812 -13608 -22716 -13592
rect -22812 -13672 -22796 -13608
rect -22732 -13672 -22716 -13608
rect -22812 -13688 -22716 -13672
rect -22812 -13752 -22796 -13688
rect -22732 -13752 -22716 -13688
rect -22812 -13768 -22716 -13752
rect -22812 -13832 -22796 -13768
rect -22732 -13832 -22716 -13768
rect -22393 -13088 -21671 -13079
rect -22393 -13792 -22384 -13088
rect -21680 -13792 -21671 -13088
rect -22393 -13801 -21671 -13792
rect -21400 -13112 -21384 -13048
rect -21320 -13112 -21304 -13048
rect -19988 -13048 -19892 -13012
rect -21400 -13128 -21304 -13112
rect -21400 -13192 -21384 -13128
rect -21320 -13192 -21304 -13128
rect -21400 -13208 -21304 -13192
rect -21400 -13272 -21384 -13208
rect -21320 -13272 -21304 -13208
rect -21400 -13288 -21304 -13272
rect -21400 -13352 -21384 -13288
rect -21320 -13352 -21304 -13288
rect -21400 -13368 -21304 -13352
rect -21400 -13432 -21384 -13368
rect -21320 -13432 -21304 -13368
rect -21400 -13448 -21304 -13432
rect -21400 -13512 -21384 -13448
rect -21320 -13512 -21304 -13448
rect -21400 -13528 -21304 -13512
rect -21400 -13592 -21384 -13528
rect -21320 -13592 -21304 -13528
rect -21400 -13608 -21304 -13592
rect -21400 -13672 -21384 -13608
rect -21320 -13672 -21304 -13608
rect -21400 -13688 -21304 -13672
rect -21400 -13752 -21384 -13688
rect -21320 -13752 -21304 -13688
rect -21400 -13768 -21304 -13752
rect -22812 -13868 -22716 -13832
rect -21400 -13832 -21384 -13768
rect -21320 -13832 -21304 -13768
rect -20981 -13088 -20259 -13079
rect -20981 -13792 -20972 -13088
rect -20268 -13792 -20259 -13088
rect -20981 -13801 -20259 -13792
rect -19988 -13112 -19972 -13048
rect -19908 -13112 -19892 -13048
rect -18576 -13048 -18480 -13012
rect -19988 -13128 -19892 -13112
rect -19988 -13192 -19972 -13128
rect -19908 -13192 -19892 -13128
rect -19988 -13208 -19892 -13192
rect -19988 -13272 -19972 -13208
rect -19908 -13272 -19892 -13208
rect -19988 -13288 -19892 -13272
rect -19988 -13352 -19972 -13288
rect -19908 -13352 -19892 -13288
rect -19988 -13368 -19892 -13352
rect -19988 -13432 -19972 -13368
rect -19908 -13432 -19892 -13368
rect -19988 -13448 -19892 -13432
rect -19988 -13512 -19972 -13448
rect -19908 -13512 -19892 -13448
rect -19988 -13528 -19892 -13512
rect -19988 -13592 -19972 -13528
rect -19908 -13592 -19892 -13528
rect -19988 -13608 -19892 -13592
rect -19988 -13672 -19972 -13608
rect -19908 -13672 -19892 -13608
rect -19988 -13688 -19892 -13672
rect -19988 -13752 -19972 -13688
rect -19908 -13752 -19892 -13688
rect -19988 -13768 -19892 -13752
rect -21400 -13868 -21304 -13832
rect -19988 -13832 -19972 -13768
rect -19908 -13832 -19892 -13768
rect -19569 -13088 -18847 -13079
rect -19569 -13792 -19560 -13088
rect -18856 -13792 -18847 -13088
rect -19569 -13801 -18847 -13792
rect -18576 -13112 -18560 -13048
rect -18496 -13112 -18480 -13048
rect -17164 -13048 -17068 -13012
rect -18576 -13128 -18480 -13112
rect -18576 -13192 -18560 -13128
rect -18496 -13192 -18480 -13128
rect -18576 -13208 -18480 -13192
rect -18576 -13272 -18560 -13208
rect -18496 -13272 -18480 -13208
rect -18576 -13288 -18480 -13272
rect -18576 -13352 -18560 -13288
rect -18496 -13352 -18480 -13288
rect -18576 -13368 -18480 -13352
rect -18576 -13432 -18560 -13368
rect -18496 -13432 -18480 -13368
rect -18576 -13448 -18480 -13432
rect -18576 -13512 -18560 -13448
rect -18496 -13512 -18480 -13448
rect -18576 -13528 -18480 -13512
rect -18576 -13592 -18560 -13528
rect -18496 -13592 -18480 -13528
rect -18576 -13608 -18480 -13592
rect -18576 -13672 -18560 -13608
rect -18496 -13672 -18480 -13608
rect -18576 -13688 -18480 -13672
rect -18576 -13752 -18560 -13688
rect -18496 -13752 -18480 -13688
rect -18576 -13768 -18480 -13752
rect -19988 -13868 -19892 -13832
rect -18576 -13832 -18560 -13768
rect -18496 -13832 -18480 -13768
rect -18157 -13088 -17435 -13079
rect -18157 -13792 -18148 -13088
rect -17444 -13792 -17435 -13088
rect -18157 -13801 -17435 -13792
rect -17164 -13112 -17148 -13048
rect -17084 -13112 -17068 -13048
rect -15752 -13048 -15656 -13012
rect -17164 -13128 -17068 -13112
rect -17164 -13192 -17148 -13128
rect -17084 -13192 -17068 -13128
rect -17164 -13208 -17068 -13192
rect -17164 -13272 -17148 -13208
rect -17084 -13272 -17068 -13208
rect -17164 -13288 -17068 -13272
rect -17164 -13352 -17148 -13288
rect -17084 -13352 -17068 -13288
rect -17164 -13368 -17068 -13352
rect -17164 -13432 -17148 -13368
rect -17084 -13432 -17068 -13368
rect -17164 -13448 -17068 -13432
rect -17164 -13512 -17148 -13448
rect -17084 -13512 -17068 -13448
rect -17164 -13528 -17068 -13512
rect -17164 -13592 -17148 -13528
rect -17084 -13592 -17068 -13528
rect -17164 -13608 -17068 -13592
rect -17164 -13672 -17148 -13608
rect -17084 -13672 -17068 -13608
rect -17164 -13688 -17068 -13672
rect -17164 -13752 -17148 -13688
rect -17084 -13752 -17068 -13688
rect -17164 -13768 -17068 -13752
rect -18576 -13868 -18480 -13832
rect -17164 -13832 -17148 -13768
rect -17084 -13832 -17068 -13768
rect -16745 -13088 -16023 -13079
rect -16745 -13792 -16736 -13088
rect -16032 -13792 -16023 -13088
rect -16745 -13801 -16023 -13792
rect -15752 -13112 -15736 -13048
rect -15672 -13112 -15656 -13048
rect -14340 -13048 -14244 -13012
rect -15752 -13128 -15656 -13112
rect -15752 -13192 -15736 -13128
rect -15672 -13192 -15656 -13128
rect -15752 -13208 -15656 -13192
rect -15752 -13272 -15736 -13208
rect -15672 -13272 -15656 -13208
rect -15752 -13288 -15656 -13272
rect -15752 -13352 -15736 -13288
rect -15672 -13352 -15656 -13288
rect -15752 -13368 -15656 -13352
rect -15752 -13432 -15736 -13368
rect -15672 -13432 -15656 -13368
rect -15752 -13448 -15656 -13432
rect -15752 -13512 -15736 -13448
rect -15672 -13512 -15656 -13448
rect -15752 -13528 -15656 -13512
rect -15752 -13592 -15736 -13528
rect -15672 -13592 -15656 -13528
rect -15752 -13608 -15656 -13592
rect -15752 -13672 -15736 -13608
rect -15672 -13672 -15656 -13608
rect -15752 -13688 -15656 -13672
rect -15752 -13752 -15736 -13688
rect -15672 -13752 -15656 -13688
rect -15752 -13768 -15656 -13752
rect -17164 -13868 -17068 -13832
rect -15752 -13832 -15736 -13768
rect -15672 -13832 -15656 -13768
rect -15333 -13088 -14611 -13079
rect -15333 -13792 -15324 -13088
rect -14620 -13792 -14611 -13088
rect -15333 -13801 -14611 -13792
rect -14340 -13112 -14324 -13048
rect -14260 -13112 -14244 -13048
rect -12928 -13048 -12832 -13012
rect -14340 -13128 -14244 -13112
rect -14340 -13192 -14324 -13128
rect -14260 -13192 -14244 -13128
rect -14340 -13208 -14244 -13192
rect -14340 -13272 -14324 -13208
rect -14260 -13272 -14244 -13208
rect -14340 -13288 -14244 -13272
rect -14340 -13352 -14324 -13288
rect -14260 -13352 -14244 -13288
rect -14340 -13368 -14244 -13352
rect -14340 -13432 -14324 -13368
rect -14260 -13432 -14244 -13368
rect -14340 -13448 -14244 -13432
rect -14340 -13512 -14324 -13448
rect -14260 -13512 -14244 -13448
rect -14340 -13528 -14244 -13512
rect -14340 -13592 -14324 -13528
rect -14260 -13592 -14244 -13528
rect -14340 -13608 -14244 -13592
rect -14340 -13672 -14324 -13608
rect -14260 -13672 -14244 -13608
rect -14340 -13688 -14244 -13672
rect -14340 -13752 -14324 -13688
rect -14260 -13752 -14244 -13688
rect -14340 -13768 -14244 -13752
rect -15752 -13868 -15656 -13832
rect -14340 -13832 -14324 -13768
rect -14260 -13832 -14244 -13768
rect -13921 -13088 -13199 -13079
rect -13921 -13792 -13912 -13088
rect -13208 -13792 -13199 -13088
rect -13921 -13801 -13199 -13792
rect -12928 -13112 -12912 -13048
rect -12848 -13112 -12832 -13048
rect -11516 -13048 -11420 -13012
rect -12928 -13128 -12832 -13112
rect -12928 -13192 -12912 -13128
rect -12848 -13192 -12832 -13128
rect -12928 -13208 -12832 -13192
rect -12928 -13272 -12912 -13208
rect -12848 -13272 -12832 -13208
rect -12928 -13288 -12832 -13272
rect -12928 -13352 -12912 -13288
rect -12848 -13352 -12832 -13288
rect -12928 -13368 -12832 -13352
rect -12928 -13432 -12912 -13368
rect -12848 -13432 -12832 -13368
rect -12928 -13448 -12832 -13432
rect -12928 -13512 -12912 -13448
rect -12848 -13512 -12832 -13448
rect -12928 -13528 -12832 -13512
rect -12928 -13592 -12912 -13528
rect -12848 -13592 -12832 -13528
rect -12928 -13608 -12832 -13592
rect -12928 -13672 -12912 -13608
rect -12848 -13672 -12832 -13608
rect -12928 -13688 -12832 -13672
rect -12928 -13752 -12912 -13688
rect -12848 -13752 -12832 -13688
rect -12928 -13768 -12832 -13752
rect -14340 -13868 -14244 -13832
rect -12928 -13832 -12912 -13768
rect -12848 -13832 -12832 -13768
rect -12509 -13088 -11787 -13079
rect -12509 -13792 -12500 -13088
rect -11796 -13792 -11787 -13088
rect -12509 -13801 -11787 -13792
rect -11516 -13112 -11500 -13048
rect -11436 -13112 -11420 -13048
rect -10104 -13048 -10008 -13012
rect -11516 -13128 -11420 -13112
rect -11516 -13192 -11500 -13128
rect -11436 -13192 -11420 -13128
rect -11516 -13208 -11420 -13192
rect -11516 -13272 -11500 -13208
rect -11436 -13272 -11420 -13208
rect -11516 -13288 -11420 -13272
rect -11516 -13352 -11500 -13288
rect -11436 -13352 -11420 -13288
rect -11516 -13368 -11420 -13352
rect -11516 -13432 -11500 -13368
rect -11436 -13432 -11420 -13368
rect -11516 -13448 -11420 -13432
rect -11516 -13512 -11500 -13448
rect -11436 -13512 -11420 -13448
rect -11516 -13528 -11420 -13512
rect -11516 -13592 -11500 -13528
rect -11436 -13592 -11420 -13528
rect -11516 -13608 -11420 -13592
rect -11516 -13672 -11500 -13608
rect -11436 -13672 -11420 -13608
rect -11516 -13688 -11420 -13672
rect -11516 -13752 -11500 -13688
rect -11436 -13752 -11420 -13688
rect -11516 -13768 -11420 -13752
rect -12928 -13868 -12832 -13832
rect -11516 -13832 -11500 -13768
rect -11436 -13832 -11420 -13768
rect -11097 -13088 -10375 -13079
rect -11097 -13792 -11088 -13088
rect -10384 -13792 -10375 -13088
rect -11097 -13801 -10375 -13792
rect -10104 -13112 -10088 -13048
rect -10024 -13112 -10008 -13048
rect -8692 -13048 -8596 -13012
rect -10104 -13128 -10008 -13112
rect -10104 -13192 -10088 -13128
rect -10024 -13192 -10008 -13128
rect -10104 -13208 -10008 -13192
rect -10104 -13272 -10088 -13208
rect -10024 -13272 -10008 -13208
rect -10104 -13288 -10008 -13272
rect -10104 -13352 -10088 -13288
rect -10024 -13352 -10008 -13288
rect -10104 -13368 -10008 -13352
rect -10104 -13432 -10088 -13368
rect -10024 -13432 -10008 -13368
rect -10104 -13448 -10008 -13432
rect -10104 -13512 -10088 -13448
rect -10024 -13512 -10008 -13448
rect -10104 -13528 -10008 -13512
rect -10104 -13592 -10088 -13528
rect -10024 -13592 -10008 -13528
rect -10104 -13608 -10008 -13592
rect -10104 -13672 -10088 -13608
rect -10024 -13672 -10008 -13608
rect -10104 -13688 -10008 -13672
rect -10104 -13752 -10088 -13688
rect -10024 -13752 -10008 -13688
rect -10104 -13768 -10008 -13752
rect -11516 -13868 -11420 -13832
rect -10104 -13832 -10088 -13768
rect -10024 -13832 -10008 -13768
rect -9685 -13088 -8963 -13079
rect -9685 -13792 -9676 -13088
rect -8972 -13792 -8963 -13088
rect -9685 -13801 -8963 -13792
rect -8692 -13112 -8676 -13048
rect -8612 -13112 -8596 -13048
rect -7280 -13048 -7184 -13012
rect -8692 -13128 -8596 -13112
rect -8692 -13192 -8676 -13128
rect -8612 -13192 -8596 -13128
rect -8692 -13208 -8596 -13192
rect -8692 -13272 -8676 -13208
rect -8612 -13272 -8596 -13208
rect -8692 -13288 -8596 -13272
rect -8692 -13352 -8676 -13288
rect -8612 -13352 -8596 -13288
rect -8692 -13368 -8596 -13352
rect -8692 -13432 -8676 -13368
rect -8612 -13432 -8596 -13368
rect -8692 -13448 -8596 -13432
rect -8692 -13512 -8676 -13448
rect -8612 -13512 -8596 -13448
rect -8692 -13528 -8596 -13512
rect -8692 -13592 -8676 -13528
rect -8612 -13592 -8596 -13528
rect -8692 -13608 -8596 -13592
rect -8692 -13672 -8676 -13608
rect -8612 -13672 -8596 -13608
rect -8692 -13688 -8596 -13672
rect -8692 -13752 -8676 -13688
rect -8612 -13752 -8596 -13688
rect -8692 -13768 -8596 -13752
rect -10104 -13868 -10008 -13832
rect -8692 -13832 -8676 -13768
rect -8612 -13832 -8596 -13768
rect -8273 -13088 -7551 -13079
rect -8273 -13792 -8264 -13088
rect -7560 -13792 -7551 -13088
rect -8273 -13801 -7551 -13792
rect -7280 -13112 -7264 -13048
rect -7200 -13112 -7184 -13048
rect -5868 -13048 -5772 -13012
rect -7280 -13128 -7184 -13112
rect -7280 -13192 -7264 -13128
rect -7200 -13192 -7184 -13128
rect -7280 -13208 -7184 -13192
rect -7280 -13272 -7264 -13208
rect -7200 -13272 -7184 -13208
rect -7280 -13288 -7184 -13272
rect -7280 -13352 -7264 -13288
rect -7200 -13352 -7184 -13288
rect -7280 -13368 -7184 -13352
rect -7280 -13432 -7264 -13368
rect -7200 -13432 -7184 -13368
rect -7280 -13448 -7184 -13432
rect -7280 -13512 -7264 -13448
rect -7200 -13512 -7184 -13448
rect -7280 -13528 -7184 -13512
rect -7280 -13592 -7264 -13528
rect -7200 -13592 -7184 -13528
rect -7280 -13608 -7184 -13592
rect -7280 -13672 -7264 -13608
rect -7200 -13672 -7184 -13608
rect -7280 -13688 -7184 -13672
rect -7280 -13752 -7264 -13688
rect -7200 -13752 -7184 -13688
rect -7280 -13768 -7184 -13752
rect -8692 -13868 -8596 -13832
rect -7280 -13832 -7264 -13768
rect -7200 -13832 -7184 -13768
rect -6861 -13088 -6139 -13079
rect -6861 -13792 -6852 -13088
rect -6148 -13792 -6139 -13088
rect -6861 -13801 -6139 -13792
rect -5868 -13112 -5852 -13048
rect -5788 -13112 -5772 -13048
rect -4456 -13048 -4360 -13012
rect -5868 -13128 -5772 -13112
rect -5868 -13192 -5852 -13128
rect -5788 -13192 -5772 -13128
rect -5868 -13208 -5772 -13192
rect -5868 -13272 -5852 -13208
rect -5788 -13272 -5772 -13208
rect -5868 -13288 -5772 -13272
rect -5868 -13352 -5852 -13288
rect -5788 -13352 -5772 -13288
rect -5868 -13368 -5772 -13352
rect -5868 -13432 -5852 -13368
rect -5788 -13432 -5772 -13368
rect -5868 -13448 -5772 -13432
rect -5868 -13512 -5852 -13448
rect -5788 -13512 -5772 -13448
rect -5868 -13528 -5772 -13512
rect -5868 -13592 -5852 -13528
rect -5788 -13592 -5772 -13528
rect -5868 -13608 -5772 -13592
rect -5868 -13672 -5852 -13608
rect -5788 -13672 -5772 -13608
rect -5868 -13688 -5772 -13672
rect -5868 -13752 -5852 -13688
rect -5788 -13752 -5772 -13688
rect -5868 -13768 -5772 -13752
rect -7280 -13868 -7184 -13832
rect -5868 -13832 -5852 -13768
rect -5788 -13832 -5772 -13768
rect -5449 -13088 -4727 -13079
rect -5449 -13792 -5440 -13088
rect -4736 -13792 -4727 -13088
rect -5449 -13801 -4727 -13792
rect -4456 -13112 -4440 -13048
rect -4376 -13112 -4360 -13048
rect -3044 -13048 -2948 -13012
rect -4456 -13128 -4360 -13112
rect -4456 -13192 -4440 -13128
rect -4376 -13192 -4360 -13128
rect -4456 -13208 -4360 -13192
rect -4456 -13272 -4440 -13208
rect -4376 -13272 -4360 -13208
rect -4456 -13288 -4360 -13272
rect -4456 -13352 -4440 -13288
rect -4376 -13352 -4360 -13288
rect -4456 -13368 -4360 -13352
rect -4456 -13432 -4440 -13368
rect -4376 -13432 -4360 -13368
rect -4456 -13448 -4360 -13432
rect -4456 -13512 -4440 -13448
rect -4376 -13512 -4360 -13448
rect -4456 -13528 -4360 -13512
rect -4456 -13592 -4440 -13528
rect -4376 -13592 -4360 -13528
rect -4456 -13608 -4360 -13592
rect -4456 -13672 -4440 -13608
rect -4376 -13672 -4360 -13608
rect -4456 -13688 -4360 -13672
rect -4456 -13752 -4440 -13688
rect -4376 -13752 -4360 -13688
rect -4456 -13768 -4360 -13752
rect -5868 -13868 -5772 -13832
rect -4456 -13832 -4440 -13768
rect -4376 -13832 -4360 -13768
rect -4037 -13088 -3315 -13079
rect -4037 -13792 -4028 -13088
rect -3324 -13792 -3315 -13088
rect -4037 -13801 -3315 -13792
rect -3044 -13112 -3028 -13048
rect -2964 -13112 -2948 -13048
rect -1632 -13048 -1536 -13012
rect -3044 -13128 -2948 -13112
rect -3044 -13192 -3028 -13128
rect -2964 -13192 -2948 -13128
rect -3044 -13208 -2948 -13192
rect -3044 -13272 -3028 -13208
rect -2964 -13272 -2948 -13208
rect -3044 -13288 -2948 -13272
rect -3044 -13352 -3028 -13288
rect -2964 -13352 -2948 -13288
rect -3044 -13368 -2948 -13352
rect -3044 -13432 -3028 -13368
rect -2964 -13432 -2948 -13368
rect -3044 -13448 -2948 -13432
rect -3044 -13512 -3028 -13448
rect -2964 -13512 -2948 -13448
rect -3044 -13528 -2948 -13512
rect -3044 -13592 -3028 -13528
rect -2964 -13592 -2948 -13528
rect -3044 -13608 -2948 -13592
rect -3044 -13672 -3028 -13608
rect -2964 -13672 -2948 -13608
rect -3044 -13688 -2948 -13672
rect -3044 -13752 -3028 -13688
rect -2964 -13752 -2948 -13688
rect -3044 -13768 -2948 -13752
rect -4456 -13868 -4360 -13832
rect -3044 -13832 -3028 -13768
rect -2964 -13832 -2948 -13768
rect -2625 -13088 -1903 -13079
rect -2625 -13792 -2616 -13088
rect -1912 -13792 -1903 -13088
rect -2625 -13801 -1903 -13792
rect -1632 -13112 -1616 -13048
rect -1552 -13112 -1536 -13048
rect -220 -13048 -124 -13012
rect -1632 -13128 -1536 -13112
rect -1632 -13192 -1616 -13128
rect -1552 -13192 -1536 -13128
rect -1632 -13208 -1536 -13192
rect -1632 -13272 -1616 -13208
rect -1552 -13272 -1536 -13208
rect -1632 -13288 -1536 -13272
rect -1632 -13352 -1616 -13288
rect -1552 -13352 -1536 -13288
rect -1632 -13368 -1536 -13352
rect -1632 -13432 -1616 -13368
rect -1552 -13432 -1536 -13368
rect -1632 -13448 -1536 -13432
rect -1632 -13512 -1616 -13448
rect -1552 -13512 -1536 -13448
rect -1632 -13528 -1536 -13512
rect -1632 -13592 -1616 -13528
rect -1552 -13592 -1536 -13528
rect -1632 -13608 -1536 -13592
rect -1632 -13672 -1616 -13608
rect -1552 -13672 -1536 -13608
rect -1632 -13688 -1536 -13672
rect -1632 -13752 -1616 -13688
rect -1552 -13752 -1536 -13688
rect -1632 -13768 -1536 -13752
rect -3044 -13868 -2948 -13832
rect -1632 -13832 -1616 -13768
rect -1552 -13832 -1536 -13768
rect -1213 -13088 -491 -13079
rect -1213 -13792 -1204 -13088
rect -500 -13792 -491 -13088
rect -1213 -13801 -491 -13792
rect -220 -13112 -204 -13048
rect -140 -13112 -124 -13048
rect 1192 -13048 1288 -13012
rect -220 -13128 -124 -13112
rect -220 -13192 -204 -13128
rect -140 -13192 -124 -13128
rect -220 -13208 -124 -13192
rect -220 -13272 -204 -13208
rect -140 -13272 -124 -13208
rect -220 -13288 -124 -13272
rect -220 -13352 -204 -13288
rect -140 -13352 -124 -13288
rect -220 -13368 -124 -13352
rect -220 -13432 -204 -13368
rect -140 -13432 -124 -13368
rect -220 -13448 -124 -13432
rect -220 -13512 -204 -13448
rect -140 -13512 -124 -13448
rect -220 -13528 -124 -13512
rect -220 -13592 -204 -13528
rect -140 -13592 -124 -13528
rect -220 -13608 -124 -13592
rect -220 -13672 -204 -13608
rect -140 -13672 -124 -13608
rect -220 -13688 -124 -13672
rect -220 -13752 -204 -13688
rect -140 -13752 -124 -13688
rect -220 -13768 -124 -13752
rect -1632 -13868 -1536 -13832
rect -220 -13832 -204 -13768
rect -140 -13832 -124 -13768
rect 199 -13088 921 -13079
rect 199 -13792 208 -13088
rect 912 -13792 921 -13088
rect 199 -13801 921 -13792
rect 1192 -13112 1208 -13048
rect 1272 -13112 1288 -13048
rect 2604 -13048 2700 -13012
rect 1192 -13128 1288 -13112
rect 1192 -13192 1208 -13128
rect 1272 -13192 1288 -13128
rect 1192 -13208 1288 -13192
rect 1192 -13272 1208 -13208
rect 1272 -13272 1288 -13208
rect 1192 -13288 1288 -13272
rect 1192 -13352 1208 -13288
rect 1272 -13352 1288 -13288
rect 1192 -13368 1288 -13352
rect 1192 -13432 1208 -13368
rect 1272 -13432 1288 -13368
rect 1192 -13448 1288 -13432
rect 1192 -13512 1208 -13448
rect 1272 -13512 1288 -13448
rect 1192 -13528 1288 -13512
rect 1192 -13592 1208 -13528
rect 1272 -13592 1288 -13528
rect 1192 -13608 1288 -13592
rect 1192 -13672 1208 -13608
rect 1272 -13672 1288 -13608
rect 1192 -13688 1288 -13672
rect 1192 -13752 1208 -13688
rect 1272 -13752 1288 -13688
rect 1192 -13768 1288 -13752
rect -220 -13868 -124 -13832
rect 1192 -13832 1208 -13768
rect 1272 -13832 1288 -13768
rect 1611 -13088 2333 -13079
rect 1611 -13792 1620 -13088
rect 2324 -13792 2333 -13088
rect 1611 -13801 2333 -13792
rect 2604 -13112 2620 -13048
rect 2684 -13112 2700 -13048
rect 4016 -13048 4112 -13012
rect 2604 -13128 2700 -13112
rect 2604 -13192 2620 -13128
rect 2684 -13192 2700 -13128
rect 2604 -13208 2700 -13192
rect 2604 -13272 2620 -13208
rect 2684 -13272 2700 -13208
rect 2604 -13288 2700 -13272
rect 2604 -13352 2620 -13288
rect 2684 -13352 2700 -13288
rect 2604 -13368 2700 -13352
rect 2604 -13432 2620 -13368
rect 2684 -13432 2700 -13368
rect 2604 -13448 2700 -13432
rect 2604 -13512 2620 -13448
rect 2684 -13512 2700 -13448
rect 2604 -13528 2700 -13512
rect 2604 -13592 2620 -13528
rect 2684 -13592 2700 -13528
rect 2604 -13608 2700 -13592
rect 2604 -13672 2620 -13608
rect 2684 -13672 2700 -13608
rect 2604 -13688 2700 -13672
rect 2604 -13752 2620 -13688
rect 2684 -13752 2700 -13688
rect 2604 -13768 2700 -13752
rect 1192 -13868 1288 -13832
rect 2604 -13832 2620 -13768
rect 2684 -13832 2700 -13768
rect 3023 -13088 3745 -13079
rect 3023 -13792 3032 -13088
rect 3736 -13792 3745 -13088
rect 3023 -13801 3745 -13792
rect 4016 -13112 4032 -13048
rect 4096 -13112 4112 -13048
rect 5428 -13048 5524 -13012
rect 4016 -13128 4112 -13112
rect 4016 -13192 4032 -13128
rect 4096 -13192 4112 -13128
rect 4016 -13208 4112 -13192
rect 4016 -13272 4032 -13208
rect 4096 -13272 4112 -13208
rect 4016 -13288 4112 -13272
rect 4016 -13352 4032 -13288
rect 4096 -13352 4112 -13288
rect 4016 -13368 4112 -13352
rect 4016 -13432 4032 -13368
rect 4096 -13432 4112 -13368
rect 4016 -13448 4112 -13432
rect 4016 -13512 4032 -13448
rect 4096 -13512 4112 -13448
rect 4016 -13528 4112 -13512
rect 4016 -13592 4032 -13528
rect 4096 -13592 4112 -13528
rect 4016 -13608 4112 -13592
rect 4016 -13672 4032 -13608
rect 4096 -13672 4112 -13608
rect 4016 -13688 4112 -13672
rect 4016 -13752 4032 -13688
rect 4096 -13752 4112 -13688
rect 4016 -13768 4112 -13752
rect 2604 -13868 2700 -13832
rect 4016 -13832 4032 -13768
rect 4096 -13832 4112 -13768
rect 4435 -13088 5157 -13079
rect 4435 -13792 4444 -13088
rect 5148 -13792 5157 -13088
rect 4435 -13801 5157 -13792
rect 5428 -13112 5444 -13048
rect 5508 -13112 5524 -13048
rect 6840 -13048 6936 -13012
rect 5428 -13128 5524 -13112
rect 5428 -13192 5444 -13128
rect 5508 -13192 5524 -13128
rect 5428 -13208 5524 -13192
rect 5428 -13272 5444 -13208
rect 5508 -13272 5524 -13208
rect 5428 -13288 5524 -13272
rect 5428 -13352 5444 -13288
rect 5508 -13352 5524 -13288
rect 5428 -13368 5524 -13352
rect 5428 -13432 5444 -13368
rect 5508 -13432 5524 -13368
rect 5428 -13448 5524 -13432
rect 5428 -13512 5444 -13448
rect 5508 -13512 5524 -13448
rect 5428 -13528 5524 -13512
rect 5428 -13592 5444 -13528
rect 5508 -13592 5524 -13528
rect 5428 -13608 5524 -13592
rect 5428 -13672 5444 -13608
rect 5508 -13672 5524 -13608
rect 5428 -13688 5524 -13672
rect 5428 -13752 5444 -13688
rect 5508 -13752 5524 -13688
rect 5428 -13768 5524 -13752
rect 4016 -13868 4112 -13832
rect 5428 -13832 5444 -13768
rect 5508 -13832 5524 -13768
rect 5847 -13088 6569 -13079
rect 5847 -13792 5856 -13088
rect 6560 -13792 6569 -13088
rect 5847 -13801 6569 -13792
rect 6840 -13112 6856 -13048
rect 6920 -13112 6936 -13048
rect 8252 -13048 8348 -13012
rect 6840 -13128 6936 -13112
rect 6840 -13192 6856 -13128
rect 6920 -13192 6936 -13128
rect 6840 -13208 6936 -13192
rect 6840 -13272 6856 -13208
rect 6920 -13272 6936 -13208
rect 6840 -13288 6936 -13272
rect 6840 -13352 6856 -13288
rect 6920 -13352 6936 -13288
rect 6840 -13368 6936 -13352
rect 6840 -13432 6856 -13368
rect 6920 -13432 6936 -13368
rect 6840 -13448 6936 -13432
rect 6840 -13512 6856 -13448
rect 6920 -13512 6936 -13448
rect 6840 -13528 6936 -13512
rect 6840 -13592 6856 -13528
rect 6920 -13592 6936 -13528
rect 6840 -13608 6936 -13592
rect 6840 -13672 6856 -13608
rect 6920 -13672 6936 -13608
rect 6840 -13688 6936 -13672
rect 6840 -13752 6856 -13688
rect 6920 -13752 6936 -13688
rect 6840 -13768 6936 -13752
rect 5428 -13868 5524 -13832
rect 6840 -13832 6856 -13768
rect 6920 -13832 6936 -13768
rect 7259 -13088 7981 -13079
rect 7259 -13792 7268 -13088
rect 7972 -13792 7981 -13088
rect 7259 -13801 7981 -13792
rect 8252 -13112 8268 -13048
rect 8332 -13112 8348 -13048
rect 9664 -13048 9760 -13012
rect 8252 -13128 8348 -13112
rect 8252 -13192 8268 -13128
rect 8332 -13192 8348 -13128
rect 8252 -13208 8348 -13192
rect 8252 -13272 8268 -13208
rect 8332 -13272 8348 -13208
rect 8252 -13288 8348 -13272
rect 8252 -13352 8268 -13288
rect 8332 -13352 8348 -13288
rect 8252 -13368 8348 -13352
rect 8252 -13432 8268 -13368
rect 8332 -13432 8348 -13368
rect 8252 -13448 8348 -13432
rect 8252 -13512 8268 -13448
rect 8332 -13512 8348 -13448
rect 8252 -13528 8348 -13512
rect 8252 -13592 8268 -13528
rect 8332 -13592 8348 -13528
rect 8252 -13608 8348 -13592
rect 8252 -13672 8268 -13608
rect 8332 -13672 8348 -13608
rect 8252 -13688 8348 -13672
rect 8252 -13752 8268 -13688
rect 8332 -13752 8348 -13688
rect 8252 -13768 8348 -13752
rect 6840 -13868 6936 -13832
rect 8252 -13832 8268 -13768
rect 8332 -13832 8348 -13768
rect 8671 -13088 9393 -13079
rect 8671 -13792 8680 -13088
rect 9384 -13792 9393 -13088
rect 8671 -13801 9393 -13792
rect 9664 -13112 9680 -13048
rect 9744 -13112 9760 -13048
rect 11076 -13048 11172 -13012
rect 9664 -13128 9760 -13112
rect 9664 -13192 9680 -13128
rect 9744 -13192 9760 -13128
rect 9664 -13208 9760 -13192
rect 9664 -13272 9680 -13208
rect 9744 -13272 9760 -13208
rect 9664 -13288 9760 -13272
rect 9664 -13352 9680 -13288
rect 9744 -13352 9760 -13288
rect 9664 -13368 9760 -13352
rect 9664 -13432 9680 -13368
rect 9744 -13432 9760 -13368
rect 9664 -13448 9760 -13432
rect 9664 -13512 9680 -13448
rect 9744 -13512 9760 -13448
rect 9664 -13528 9760 -13512
rect 9664 -13592 9680 -13528
rect 9744 -13592 9760 -13528
rect 9664 -13608 9760 -13592
rect 9664 -13672 9680 -13608
rect 9744 -13672 9760 -13608
rect 9664 -13688 9760 -13672
rect 9664 -13752 9680 -13688
rect 9744 -13752 9760 -13688
rect 9664 -13768 9760 -13752
rect 8252 -13868 8348 -13832
rect 9664 -13832 9680 -13768
rect 9744 -13832 9760 -13768
rect 10083 -13088 10805 -13079
rect 10083 -13792 10092 -13088
rect 10796 -13792 10805 -13088
rect 10083 -13801 10805 -13792
rect 11076 -13112 11092 -13048
rect 11156 -13112 11172 -13048
rect 12488 -13048 12584 -13012
rect 11076 -13128 11172 -13112
rect 11076 -13192 11092 -13128
rect 11156 -13192 11172 -13128
rect 11076 -13208 11172 -13192
rect 11076 -13272 11092 -13208
rect 11156 -13272 11172 -13208
rect 11076 -13288 11172 -13272
rect 11076 -13352 11092 -13288
rect 11156 -13352 11172 -13288
rect 11076 -13368 11172 -13352
rect 11076 -13432 11092 -13368
rect 11156 -13432 11172 -13368
rect 11076 -13448 11172 -13432
rect 11076 -13512 11092 -13448
rect 11156 -13512 11172 -13448
rect 11076 -13528 11172 -13512
rect 11076 -13592 11092 -13528
rect 11156 -13592 11172 -13528
rect 11076 -13608 11172 -13592
rect 11076 -13672 11092 -13608
rect 11156 -13672 11172 -13608
rect 11076 -13688 11172 -13672
rect 11076 -13752 11092 -13688
rect 11156 -13752 11172 -13688
rect 11076 -13768 11172 -13752
rect 9664 -13868 9760 -13832
rect 11076 -13832 11092 -13768
rect 11156 -13832 11172 -13768
rect 11495 -13088 12217 -13079
rect 11495 -13792 11504 -13088
rect 12208 -13792 12217 -13088
rect 11495 -13801 12217 -13792
rect 12488 -13112 12504 -13048
rect 12568 -13112 12584 -13048
rect 13900 -13048 13996 -13012
rect 12488 -13128 12584 -13112
rect 12488 -13192 12504 -13128
rect 12568 -13192 12584 -13128
rect 12488 -13208 12584 -13192
rect 12488 -13272 12504 -13208
rect 12568 -13272 12584 -13208
rect 12488 -13288 12584 -13272
rect 12488 -13352 12504 -13288
rect 12568 -13352 12584 -13288
rect 12488 -13368 12584 -13352
rect 12488 -13432 12504 -13368
rect 12568 -13432 12584 -13368
rect 12488 -13448 12584 -13432
rect 12488 -13512 12504 -13448
rect 12568 -13512 12584 -13448
rect 12488 -13528 12584 -13512
rect 12488 -13592 12504 -13528
rect 12568 -13592 12584 -13528
rect 12488 -13608 12584 -13592
rect 12488 -13672 12504 -13608
rect 12568 -13672 12584 -13608
rect 12488 -13688 12584 -13672
rect 12488 -13752 12504 -13688
rect 12568 -13752 12584 -13688
rect 12488 -13768 12584 -13752
rect 11076 -13868 11172 -13832
rect 12488 -13832 12504 -13768
rect 12568 -13832 12584 -13768
rect 12907 -13088 13629 -13079
rect 12907 -13792 12916 -13088
rect 13620 -13792 13629 -13088
rect 12907 -13801 13629 -13792
rect 13900 -13112 13916 -13048
rect 13980 -13112 13996 -13048
rect 15312 -13048 15408 -13012
rect 13900 -13128 13996 -13112
rect 13900 -13192 13916 -13128
rect 13980 -13192 13996 -13128
rect 13900 -13208 13996 -13192
rect 13900 -13272 13916 -13208
rect 13980 -13272 13996 -13208
rect 13900 -13288 13996 -13272
rect 13900 -13352 13916 -13288
rect 13980 -13352 13996 -13288
rect 13900 -13368 13996 -13352
rect 13900 -13432 13916 -13368
rect 13980 -13432 13996 -13368
rect 13900 -13448 13996 -13432
rect 13900 -13512 13916 -13448
rect 13980 -13512 13996 -13448
rect 13900 -13528 13996 -13512
rect 13900 -13592 13916 -13528
rect 13980 -13592 13996 -13528
rect 13900 -13608 13996 -13592
rect 13900 -13672 13916 -13608
rect 13980 -13672 13996 -13608
rect 13900 -13688 13996 -13672
rect 13900 -13752 13916 -13688
rect 13980 -13752 13996 -13688
rect 13900 -13768 13996 -13752
rect 12488 -13868 12584 -13832
rect 13900 -13832 13916 -13768
rect 13980 -13832 13996 -13768
rect 14319 -13088 15041 -13079
rect 14319 -13792 14328 -13088
rect 15032 -13792 15041 -13088
rect 14319 -13801 15041 -13792
rect 15312 -13112 15328 -13048
rect 15392 -13112 15408 -13048
rect 16724 -13048 16820 -13012
rect 15312 -13128 15408 -13112
rect 15312 -13192 15328 -13128
rect 15392 -13192 15408 -13128
rect 15312 -13208 15408 -13192
rect 15312 -13272 15328 -13208
rect 15392 -13272 15408 -13208
rect 15312 -13288 15408 -13272
rect 15312 -13352 15328 -13288
rect 15392 -13352 15408 -13288
rect 15312 -13368 15408 -13352
rect 15312 -13432 15328 -13368
rect 15392 -13432 15408 -13368
rect 15312 -13448 15408 -13432
rect 15312 -13512 15328 -13448
rect 15392 -13512 15408 -13448
rect 15312 -13528 15408 -13512
rect 15312 -13592 15328 -13528
rect 15392 -13592 15408 -13528
rect 15312 -13608 15408 -13592
rect 15312 -13672 15328 -13608
rect 15392 -13672 15408 -13608
rect 15312 -13688 15408 -13672
rect 15312 -13752 15328 -13688
rect 15392 -13752 15408 -13688
rect 15312 -13768 15408 -13752
rect 13900 -13868 13996 -13832
rect 15312 -13832 15328 -13768
rect 15392 -13832 15408 -13768
rect 15731 -13088 16453 -13079
rect 15731 -13792 15740 -13088
rect 16444 -13792 16453 -13088
rect 15731 -13801 16453 -13792
rect 16724 -13112 16740 -13048
rect 16804 -13112 16820 -13048
rect 18136 -13048 18232 -13012
rect 16724 -13128 16820 -13112
rect 16724 -13192 16740 -13128
rect 16804 -13192 16820 -13128
rect 16724 -13208 16820 -13192
rect 16724 -13272 16740 -13208
rect 16804 -13272 16820 -13208
rect 16724 -13288 16820 -13272
rect 16724 -13352 16740 -13288
rect 16804 -13352 16820 -13288
rect 16724 -13368 16820 -13352
rect 16724 -13432 16740 -13368
rect 16804 -13432 16820 -13368
rect 16724 -13448 16820 -13432
rect 16724 -13512 16740 -13448
rect 16804 -13512 16820 -13448
rect 16724 -13528 16820 -13512
rect 16724 -13592 16740 -13528
rect 16804 -13592 16820 -13528
rect 16724 -13608 16820 -13592
rect 16724 -13672 16740 -13608
rect 16804 -13672 16820 -13608
rect 16724 -13688 16820 -13672
rect 16724 -13752 16740 -13688
rect 16804 -13752 16820 -13688
rect 16724 -13768 16820 -13752
rect 15312 -13868 15408 -13832
rect 16724 -13832 16740 -13768
rect 16804 -13832 16820 -13768
rect 17143 -13088 17865 -13079
rect 17143 -13792 17152 -13088
rect 17856 -13792 17865 -13088
rect 17143 -13801 17865 -13792
rect 18136 -13112 18152 -13048
rect 18216 -13112 18232 -13048
rect 19548 -13048 19644 -13012
rect 18136 -13128 18232 -13112
rect 18136 -13192 18152 -13128
rect 18216 -13192 18232 -13128
rect 18136 -13208 18232 -13192
rect 18136 -13272 18152 -13208
rect 18216 -13272 18232 -13208
rect 18136 -13288 18232 -13272
rect 18136 -13352 18152 -13288
rect 18216 -13352 18232 -13288
rect 18136 -13368 18232 -13352
rect 18136 -13432 18152 -13368
rect 18216 -13432 18232 -13368
rect 18136 -13448 18232 -13432
rect 18136 -13512 18152 -13448
rect 18216 -13512 18232 -13448
rect 18136 -13528 18232 -13512
rect 18136 -13592 18152 -13528
rect 18216 -13592 18232 -13528
rect 18136 -13608 18232 -13592
rect 18136 -13672 18152 -13608
rect 18216 -13672 18232 -13608
rect 18136 -13688 18232 -13672
rect 18136 -13752 18152 -13688
rect 18216 -13752 18232 -13688
rect 18136 -13768 18232 -13752
rect 16724 -13868 16820 -13832
rect 18136 -13832 18152 -13768
rect 18216 -13832 18232 -13768
rect 18555 -13088 19277 -13079
rect 18555 -13792 18564 -13088
rect 19268 -13792 19277 -13088
rect 18555 -13801 19277 -13792
rect 19548 -13112 19564 -13048
rect 19628 -13112 19644 -13048
rect 20960 -13048 21056 -13012
rect 19548 -13128 19644 -13112
rect 19548 -13192 19564 -13128
rect 19628 -13192 19644 -13128
rect 19548 -13208 19644 -13192
rect 19548 -13272 19564 -13208
rect 19628 -13272 19644 -13208
rect 19548 -13288 19644 -13272
rect 19548 -13352 19564 -13288
rect 19628 -13352 19644 -13288
rect 19548 -13368 19644 -13352
rect 19548 -13432 19564 -13368
rect 19628 -13432 19644 -13368
rect 19548 -13448 19644 -13432
rect 19548 -13512 19564 -13448
rect 19628 -13512 19644 -13448
rect 19548 -13528 19644 -13512
rect 19548 -13592 19564 -13528
rect 19628 -13592 19644 -13528
rect 19548 -13608 19644 -13592
rect 19548 -13672 19564 -13608
rect 19628 -13672 19644 -13608
rect 19548 -13688 19644 -13672
rect 19548 -13752 19564 -13688
rect 19628 -13752 19644 -13688
rect 19548 -13768 19644 -13752
rect 18136 -13868 18232 -13832
rect 19548 -13832 19564 -13768
rect 19628 -13832 19644 -13768
rect 19967 -13088 20689 -13079
rect 19967 -13792 19976 -13088
rect 20680 -13792 20689 -13088
rect 19967 -13801 20689 -13792
rect 20960 -13112 20976 -13048
rect 21040 -13112 21056 -13048
rect 22372 -13048 22468 -13012
rect 20960 -13128 21056 -13112
rect 20960 -13192 20976 -13128
rect 21040 -13192 21056 -13128
rect 20960 -13208 21056 -13192
rect 20960 -13272 20976 -13208
rect 21040 -13272 21056 -13208
rect 20960 -13288 21056 -13272
rect 20960 -13352 20976 -13288
rect 21040 -13352 21056 -13288
rect 20960 -13368 21056 -13352
rect 20960 -13432 20976 -13368
rect 21040 -13432 21056 -13368
rect 20960 -13448 21056 -13432
rect 20960 -13512 20976 -13448
rect 21040 -13512 21056 -13448
rect 20960 -13528 21056 -13512
rect 20960 -13592 20976 -13528
rect 21040 -13592 21056 -13528
rect 20960 -13608 21056 -13592
rect 20960 -13672 20976 -13608
rect 21040 -13672 21056 -13608
rect 20960 -13688 21056 -13672
rect 20960 -13752 20976 -13688
rect 21040 -13752 21056 -13688
rect 20960 -13768 21056 -13752
rect 19548 -13868 19644 -13832
rect 20960 -13832 20976 -13768
rect 21040 -13832 21056 -13768
rect 21379 -13088 22101 -13079
rect 21379 -13792 21388 -13088
rect 22092 -13792 22101 -13088
rect 21379 -13801 22101 -13792
rect 22372 -13112 22388 -13048
rect 22452 -13112 22468 -13048
rect 23784 -13048 23880 -13012
rect 22372 -13128 22468 -13112
rect 22372 -13192 22388 -13128
rect 22452 -13192 22468 -13128
rect 22372 -13208 22468 -13192
rect 22372 -13272 22388 -13208
rect 22452 -13272 22468 -13208
rect 22372 -13288 22468 -13272
rect 22372 -13352 22388 -13288
rect 22452 -13352 22468 -13288
rect 22372 -13368 22468 -13352
rect 22372 -13432 22388 -13368
rect 22452 -13432 22468 -13368
rect 22372 -13448 22468 -13432
rect 22372 -13512 22388 -13448
rect 22452 -13512 22468 -13448
rect 22372 -13528 22468 -13512
rect 22372 -13592 22388 -13528
rect 22452 -13592 22468 -13528
rect 22372 -13608 22468 -13592
rect 22372 -13672 22388 -13608
rect 22452 -13672 22468 -13608
rect 22372 -13688 22468 -13672
rect 22372 -13752 22388 -13688
rect 22452 -13752 22468 -13688
rect 22372 -13768 22468 -13752
rect 20960 -13868 21056 -13832
rect 22372 -13832 22388 -13768
rect 22452 -13832 22468 -13768
rect 22791 -13088 23513 -13079
rect 22791 -13792 22800 -13088
rect 23504 -13792 23513 -13088
rect 22791 -13801 23513 -13792
rect 23784 -13112 23800 -13048
rect 23864 -13112 23880 -13048
rect 23784 -13128 23880 -13112
rect 23784 -13192 23800 -13128
rect 23864 -13192 23880 -13128
rect 23784 -13208 23880 -13192
rect 23784 -13272 23800 -13208
rect 23864 -13272 23880 -13208
rect 23784 -13288 23880 -13272
rect 23784 -13352 23800 -13288
rect 23864 -13352 23880 -13288
rect 23784 -13368 23880 -13352
rect 23784 -13432 23800 -13368
rect 23864 -13432 23880 -13368
rect 23784 -13448 23880 -13432
rect 23784 -13512 23800 -13448
rect 23864 -13512 23880 -13448
rect 23784 -13528 23880 -13512
rect 23784 -13592 23800 -13528
rect 23864 -13592 23880 -13528
rect 23784 -13608 23880 -13592
rect 23784 -13672 23800 -13608
rect 23864 -13672 23880 -13608
rect 23784 -13688 23880 -13672
rect 23784 -13752 23800 -13688
rect 23864 -13752 23880 -13688
rect 23784 -13768 23880 -13752
rect 22372 -13868 22468 -13832
rect 23784 -13832 23800 -13768
rect 23864 -13832 23880 -13768
rect 23784 -13868 23880 -13832
rect -22812 -14168 -22716 -14132
rect -23805 -14208 -23083 -14199
rect -23805 -14912 -23796 -14208
rect -23092 -14912 -23083 -14208
rect -23805 -14921 -23083 -14912
rect -22812 -14232 -22796 -14168
rect -22732 -14232 -22716 -14168
rect -21400 -14168 -21304 -14132
rect -22812 -14248 -22716 -14232
rect -22812 -14312 -22796 -14248
rect -22732 -14312 -22716 -14248
rect -22812 -14328 -22716 -14312
rect -22812 -14392 -22796 -14328
rect -22732 -14392 -22716 -14328
rect -22812 -14408 -22716 -14392
rect -22812 -14472 -22796 -14408
rect -22732 -14472 -22716 -14408
rect -22812 -14488 -22716 -14472
rect -22812 -14552 -22796 -14488
rect -22732 -14552 -22716 -14488
rect -22812 -14568 -22716 -14552
rect -22812 -14632 -22796 -14568
rect -22732 -14632 -22716 -14568
rect -22812 -14648 -22716 -14632
rect -22812 -14712 -22796 -14648
rect -22732 -14712 -22716 -14648
rect -22812 -14728 -22716 -14712
rect -22812 -14792 -22796 -14728
rect -22732 -14792 -22716 -14728
rect -22812 -14808 -22716 -14792
rect -22812 -14872 -22796 -14808
rect -22732 -14872 -22716 -14808
rect -22812 -14888 -22716 -14872
rect -22812 -14952 -22796 -14888
rect -22732 -14952 -22716 -14888
rect -22393 -14208 -21671 -14199
rect -22393 -14912 -22384 -14208
rect -21680 -14912 -21671 -14208
rect -22393 -14921 -21671 -14912
rect -21400 -14232 -21384 -14168
rect -21320 -14232 -21304 -14168
rect -19988 -14168 -19892 -14132
rect -21400 -14248 -21304 -14232
rect -21400 -14312 -21384 -14248
rect -21320 -14312 -21304 -14248
rect -21400 -14328 -21304 -14312
rect -21400 -14392 -21384 -14328
rect -21320 -14392 -21304 -14328
rect -21400 -14408 -21304 -14392
rect -21400 -14472 -21384 -14408
rect -21320 -14472 -21304 -14408
rect -21400 -14488 -21304 -14472
rect -21400 -14552 -21384 -14488
rect -21320 -14552 -21304 -14488
rect -21400 -14568 -21304 -14552
rect -21400 -14632 -21384 -14568
rect -21320 -14632 -21304 -14568
rect -21400 -14648 -21304 -14632
rect -21400 -14712 -21384 -14648
rect -21320 -14712 -21304 -14648
rect -21400 -14728 -21304 -14712
rect -21400 -14792 -21384 -14728
rect -21320 -14792 -21304 -14728
rect -21400 -14808 -21304 -14792
rect -21400 -14872 -21384 -14808
rect -21320 -14872 -21304 -14808
rect -21400 -14888 -21304 -14872
rect -22812 -14988 -22716 -14952
rect -21400 -14952 -21384 -14888
rect -21320 -14952 -21304 -14888
rect -20981 -14208 -20259 -14199
rect -20981 -14912 -20972 -14208
rect -20268 -14912 -20259 -14208
rect -20981 -14921 -20259 -14912
rect -19988 -14232 -19972 -14168
rect -19908 -14232 -19892 -14168
rect -18576 -14168 -18480 -14132
rect -19988 -14248 -19892 -14232
rect -19988 -14312 -19972 -14248
rect -19908 -14312 -19892 -14248
rect -19988 -14328 -19892 -14312
rect -19988 -14392 -19972 -14328
rect -19908 -14392 -19892 -14328
rect -19988 -14408 -19892 -14392
rect -19988 -14472 -19972 -14408
rect -19908 -14472 -19892 -14408
rect -19988 -14488 -19892 -14472
rect -19988 -14552 -19972 -14488
rect -19908 -14552 -19892 -14488
rect -19988 -14568 -19892 -14552
rect -19988 -14632 -19972 -14568
rect -19908 -14632 -19892 -14568
rect -19988 -14648 -19892 -14632
rect -19988 -14712 -19972 -14648
rect -19908 -14712 -19892 -14648
rect -19988 -14728 -19892 -14712
rect -19988 -14792 -19972 -14728
rect -19908 -14792 -19892 -14728
rect -19988 -14808 -19892 -14792
rect -19988 -14872 -19972 -14808
rect -19908 -14872 -19892 -14808
rect -19988 -14888 -19892 -14872
rect -21400 -14988 -21304 -14952
rect -19988 -14952 -19972 -14888
rect -19908 -14952 -19892 -14888
rect -19569 -14208 -18847 -14199
rect -19569 -14912 -19560 -14208
rect -18856 -14912 -18847 -14208
rect -19569 -14921 -18847 -14912
rect -18576 -14232 -18560 -14168
rect -18496 -14232 -18480 -14168
rect -17164 -14168 -17068 -14132
rect -18576 -14248 -18480 -14232
rect -18576 -14312 -18560 -14248
rect -18496 -14312 -18480 -14248
rect -18576 -14328 -18480 -14312
rect -18576 -14392 -18560 -14328
rect -18496 -14392 -18480 -14328
rect -18576 -14408 -18480 -14392
rect -18576 -14472 -18560 -14408
rect -18496 -14472 -18480 -14408
rect -18576 -14488 -18480 -14472
rect -18576 -14552 -18560 -14488
rect -18496 -14552 -18480 -14488
rect -18576 -14568 -18480 -14552
rect -18576 -14632 -18560 -14568
rect -18496 -14632 -18480 -14568
rect -18576 -14648 -18480 -14632
rect -18576 -14712 -18560 -14648
rect -18496 -14712 -18480 -14648
rect -18576 -14728 -18480 -14712
rect -18576 -14792 -18560 -14728
rect -18496 -14792 -18480 -14728
rect -18576 -14808 -18480 -14792
rect -18576 -14872 -18560 -14808
rect -18496 -14872 -18480 -14808
rect -18576 -14888 -18480 -14872
rect -19988 -14988 -19892 -14952
rect -18576 -14952 -18560 -14888
rect -18496 -14952 -18480 -14888
rect -18157 -14208 -17435 -14199
rect -18157 -14912 -18148 -14208
rect -17444 -14912 -17435 -14208
rect -18157 -14921 -17435 -14912
rect -17164 -14232 -17148 -14168
rect -17084 -14232 -17068 -14168
rect -15752 -14168 -15656 -14132
rect -17164 -14248 -17068 -14232
rect -17164 -14312 -17148 -14248
rect -17084 -14312 -17068 -14248
rect -17164 -14328 -17068 -14312
rect -17164 -14392 -17148 -14328
rect -17084 -14392 -17068 -14328
rect -17164 -14408 -17068 -14392
rect -17164 -14472 -17148 -14408
rect -17084 -14472 -17068 -14408
rect -17164 -14488 -17068 -14472
rect -17164 -14552 -17148 -14488
rect -17084 -14552 -17068 -14488
rect -17164 -14568 -17068 -14552
rect -17164 -14632 -17148 -14568
rect -17084 -14632 -17068 -14568
rect -17164 -14648 -17068 -14632
rect -17164 -14712 -17148 -14648
rect -17084 -14712 -17068 -14648
rect -17164 -14728 -17068 -14712
rect -17164 -14792 -17148 -14728
rect -17084 -14792 -17068 -14728
rect -17164 -14808 -17068 -14792
rect -17164 -14872 -17148 -14808
rect -17084 -14872 -17068 -14808
rect -17164 -14888 -17068 -14872
rect -18576 -14988 -18480 -14952
rect -17164 -14952 -17148 -14888
rect -17084 -14952 -17068 -14888
rect -16745 -14208 -16023 -14199
rect -16745 -14912 -16736 -14208
rect -16032 -14912 -16023 -14208
rect -16745 -14921 -16023 -14912
rect -15752 -14232 -15736 -14168
rect -15672 -14232 -15656 -14168
rect -14340 -14168 -14244 -14132
rect -15752 -14248 -15656 -14232
rect -15752 -14312 -15736 -14248
rect -15672 -14312 -15656 -14248
rect -15752 -14328 -15656 -14312
rect -15752 -14392 -15736 -14328
rect -15672 -14392 -15656 -14328
rect -15752 -14408 -15656 -14392
rect -15752 -14472 -15736 -14408
rect -15672 -14472 -15656 -14408
rect -15752 -14488 -15656 -14472
rect -15752 -14552 -15736 -14488
rect -15672 -14552 -15656 -14488
rect -15752 -14568 -15656 -14552
rect -15752 -14632 -15736 -14568
rect -15672 -14632 -15656 -14568
rect -15752 -14648 -15656 -14632
rect -15752 -14712 -15736 -14648
rect -15672 -14712 -15656 -14648
rect -15752 -14728 -15656 -14712
rect -15752 -14792 -15736 -14728
rect -15672 -14792 -15656 -14728
rect -15752 -14808 -15656 -14792
rect -15752 -14872 -15736 -14808
rect -15672 -14872 -15656 -14808
rect -15752 -14888 -15656 -14872
rect -17164 -14988 -17068 -14952
rect -15752 -14952 -15736 -14888
rect -15672 -14952 -15656 -14888
rect -15333 -14208 -14611 -14199
rect -15333 -14912 -15324 -14208
rect -14620 -14912 -14611 -14208
rect -15333 -14921 -14611 -14912
rect -14340 -14232 -14324 -14168
rect -14260 -14232 -14244 -14168
rect -12928 -14168 -12832 -14132
rect -14340 -14248 -14244 -14232
rect -14340 -14312 -14324 -14248
rect -14260 -14312 -14244 -14248
rect -14340 -14328 -14244 -14312
rect -14340 -14392 -14324 -14328
rect -14260 -14392 -14244 -14328
rect -14340 -14408 -14244 -14392
rect -14340 -14472 -14324 -14408
rect -14260 -14472 -14244 -14408
rect -14340 -14488 -14244 -14472
rect -14340 -14552 -14324 -14488
rect -14260 -14552 -14244 -14488
rect -14340 -14568 -14244 -14552
rect -14340 -14632 -14324 -14568
rect -14260 -14632 -14244 -14568
rect -14340 -14648 -14244 -14632
rect -14340 -14712 -14324 -14648
rect -14260 -14712 -14244 -14648
rect -14340 -14728 -14244 -14712
rect -14340 -14792 -14324 -14728
rect -14260 -14792 -14244 -14728
rect -14340 -14808 -14244 -14792
rect -14340 -14872 -14324 -14808
rect -14260 -14872 -14244 -14808
rect -14340 -14888 -14244 -14872
rect -15752 -14988 -15656 -14952
rect -14340 -14952 -14324 -14888
rect -14260 -14952 -14244 -14888
rect -13921 -14208 -13199 -14199
rect -13921 -14912 -13912 -14208
rect -13208 -14912 -13199 -14208
rect -13921 -14921 -13199 -14912
rect -12928 -14232 -12912 -14168
rect -12848 -14232 -12832 -14168
rect -11516 -14168 -11420 -14132
rect -12928 -14248 -12832 -14232
rect -12928 -14312 -12912 -14248
rect -12848 -14312 -12832 -14248
rect -12928 -14328 -12832 -14312
rect -12928 -14392 -12912 -14328
rect -12848 -14392 -12832 -14328
rect -12928 -14408 -12832 -14392
rect -12928 -14472 -12912 -14408
rect -12848 -14472 -12832 -14408
rect -12928 -14488 -12832 -14472
rect -12928 -14552 -12912 -14488
rect -12848 -14552 -12832 -14488
rect -12928 -14568 -12832 -14552
rect -12928 -14632 -12912 -14568
rect -12848 -14632 -12832 -14568
rect -12928 -14648 -12832 -14632
rect -12928 -14712 -12912 -14648
rect -12848 -14712 -12832 -14648
rect -12928 -14728 -12832 -14712
rect -12928 -14792 -12912 -14728
rect -12848 -14792 -12832 -14728
rect -12928 -14808 -12832 -14792
rect -12928 -14872 -12912 -14808
rect -12848 -14872 -12832 -14808
rect -12928 -14888 -12832 -14872
rect -14340 -14988 -14244 -14952
rect -12928 -14952 -12912 -14888
rect -12848 -14952 -12832 -14888
rect -12509 -14208 -11787 -14199
rect -12509 -14912 -12500 -14208
rect -11796 -14912 -11787 -14208
rect -12509 -14921 -11787 -14912
rect -11516 -14232 -11500 -14168
rect -11436 -14232 -11420 -14168
rect -10104 -14168 -10008 -14132
rect -11516 -14248 -11420 -14232
rect -11516 -14312 -11500 -14248
rect -11436 -14312 -11420 -14248
rect -11516 -14328 -11420 -14312
rect -11516 -14392 -11500 -14328
rect -11436 -14392 -11420 -14328
rect -11516 -14408 -11420 -14392
rect -11516 -14472 -11500 -14408
rect -11436 -14472 -11420 -14408
rect -11516 -14488 -11420 -14472
rect -11516 -14552 -11500 -14488
rect -11436 -14552 -11420 -14488
rect -11516 -14568 -11420 -14552
rect -11516 -14632 -11500 -14568
rect -11436 -14632 -11420 -14568
rect -11516 -14648 -11420 -14632
rect -11516 -14712 -11500 -14648
rect -11436 -14712 -11420 -14648
rect -11516 -14728 -11420 -14712
rect -11516 -14792 -11500 -14728
rect -11436 -14792 -11420 -14728
rect -11516 -14808 -11420 -14792
rect -11516 -14872 -11500 -14808
rect -11436 -14872 -11420 -14808
rect -11516 -14888 -11420 -14872
rect -12928 -14988 -12832 -14952
rect -11516 -14952 -11500 -14888
rect -11436 -14952 -11420 -14888
rect -11097 -14208 -10375 -14199
rect -11097 -14912 -11088 -14208
rect -10384 -14912 -10375 -14208
rect -11097 -14921 -10375 -14912
rect -10104 -14232 -10088 -14168
rect -10024 -14232 -10008 -14168
rect -8692 -14168 -8596 -14132
rect -10104 -14248 -10008 -14232
rect -10104 -14312 -10088 -14248
rect -10024 -14312 -10008 -14248
rect -10104 -14328 -10008 -14312
rect -10104 -14392 -10088 -14328
rect -10024 -14392 -10008 -14328
rect -10104 -14408 -10008 -14392
rect -10104 -14472 -10088 -14408
rect -10024 -14472 -10008 -14408
rect -10104 -14488 -10008 -14472
rect -10104 -14552 -10088 -14488
rect -10024 -14552 -10008 -14488
rect -10104 -14568 -10008 -14552
rect -10104 -14632 -10088 -14568
rect -10024 -14632 -10008 -14568
rect -10104 -14648 -10008 -14632
rect -10104 -14712 -10088 -14648
rect -10024 -14712 -10008 -14648
rect -10104 -14728 -10008 -14712
rect -10104 -14792 -10088 -14728
rect -10024 -14792 -10008 -14728
rect -10104 -14808 -10008 -14792
rect -10104 -14872 -10088 -14808
rect -10024 -14872 -10008 -14808
rect -10104 -14888 -10008 -14872
rect -11516 -14988 -11420 -14952
rect -10104 -14952 -10088 -14888
rect -10024 -14952 -10008 -14888
rect -9685 -14208 -8963 -14199
rect -9685 -14912 -9676 -14208
rect -8972 -14912 -8963 -14208
rect -9685 -14921 -8963 -14912
rect -8692 -14232 -8676 -14168
rect -8612 -14232 -8596 -14168
rect -7280 -14168 -7184 -14132
rect -8692 -14248 -8596 -14232
rect -8692 -14312 -8676 -14248
rect -8612 -14312 -8596 -14248
rect -8692 -14328 -8596 -14312
rect -8692 -14392 -8676 -14328
rect -8612 -14392 -8596 -14328
rect -8692 -14408 -8596 -14392
rect -8692 -14472 -8676 -14408
rect -8612 -14472 -8596 -14408
rect -8692 -14488 -8596 -14472
rect -8692 -14552 -8676 -14488
rect -8612 -14552 -8596 -14488
rect -8692 -14568 -8596 -14552
rect -8692 -14632 -8676 -14568
rect -8612 -14632 -8596 -14568
rect -8692 -14648 -8596 -14632
rect -8692 -14712 -8676 -14648
rect -8612 -14712 -8596 -14648
rect -8692 -14728 -8596 -14712
rect -8692 -14792 -8676 -14728
rect -8612 -14792 -8596 -14728
rect -8692 -14808 -8596 -14792
rect -8692 -14872 -8676 -14808
rect -8612 -14872 -8596 -14808
rect -8692 -14888 -8596 -14872
rect -10104 -14988 -10008 -14952
rect -8692 -14952 -8676 -14888
rect -8612 -14952 -8596 -14888
rect -8273 -14208 -7551 -14199
rect -8273 -14912 -8264 -14208
rect -7560 -14912 -7551 -14208
rect -8273 -14921 -7551 -14912
rect -7280 -14232 -7264 -14168
rect -7200 -14232 -7184 -14168
rect -5868 -14168 -5772 -14132
rect -7280 -14248 -7184 -14232
rect -7280 -14312 -7264 -14248
rect -7200 -14312 -7184 -14248
rect -7280 -14328 -7184 -14312
rect -7280 -14392 -7264 -14328
rect -7200 -14392 -7184 -14328
rect -7280 -14408 -7184 -14392
rect -7280 -14472 -7264 -14408
rect -7200 -14472 -7184 -14408
rect -7280 -14488 -7184 -14472
rect -7280 -14552 -7264 -14488
rect -7200 -14552 -7184 -14488
rect -7280 -14568 -7184 -14552
rect -7280 -14632 -7264 -14568
rect -7200 -14632 -7184 -14568
rect -7280 -14648 -7184 -14632
rect -7280 -14712 -7264 -14648
rect -7200 -14712 -7184 -14648
rect -7280 -14728 -7184 -14712
rect -7280 -14792 -7264 -14728
rect -7200 -14792 -7184 -14728
rect -7280 -14808 -7184 -14792
rect -7280 -14872 -7264 -14808
rect -7200 -14872 -7184 -14808
rect -7280 -14888 -7184 -14872
rect -8692 -14988 -8596 -14952
rect -7280 -14952 -7264 -14888
rect -7200 -14952 -7184 -14888
rect -6861 -14208 -6139 -14199
rect -6861 -14912 -6852 -14208
rect -6148 -14912 -6139 -14208
rect -6861 -14921 -6139 -14912
rect -5868 -14232 -5852 -14168
rect -5788 -14232 -5772 -14168
rect -4456 -14168 -4360 -14132
rect -5868 -14248 -5772 -14232
rect -5868 -14312 -5852 -14248
rect -5788 -14312 -5772 -14248
rect -5868 -14328 -5772 -14312
rect -5868 -14392 -5852 -14328
rect -5788 -14392 -5772 -14328
rect -5868 -14408 -5772 -14392
rect -5868 -14472 -5852 -14408
rect -5788 -14472 -5772 -14408
rect -5868 -14488 -5772 -14472
rect -5868 -14552 -5852 -14488
rect -5788 -14552 -5772 -14488
rect -5868 -14568 -5772 -14552
rect -5868 -14632 -5852 -14568
rect -5788 -14632 -5772 -14568
rect -5868 -14648 -5772 -14632
rect -5868 -14712 -5852 -14648
rect -5788 -14712 -5772 -14648
rect -5868 -14728 -5772 -14712
rect -5868 -14792 -5852 -14728
rect -5788 -14792 -5772 -14728
rect -5868 -14808 -5772 -14792
rect -5868 -14872 -5852 -14808
rect -5788 -14872 -5772 -14808
rect -5868 -14888 -5772 -14872
rect -7280 -14988 -7184 -14952
rect -5868 -14952 -5852 -14888
rect -5788 -14952 -5772 -14888
rect -5449 -14208 -4727 -14199
rect -5449 -14912 -5440 -14208
rect -4736 -14912 -4727 -14208
rect -5449 -14921 -4727 -14912
rect -4456 -14232 -4440 -14168
rect -4376 -14232 -4360 -14168
rect -3044 -14168 -2948 -14132
rect -4456 -14248 -4360 -14232
rect -4456 -14312 -4440 -14248
rect -4376 -14312 -4360 -14248
rect -4456 -14328 -4360 -14312
rect -4456 -14392 -4440 -14328
rect -4376 -14392 -4360 -14328
rect -4456 -14408 -4360 -14392
rect -4456 -14472 -4440 -14408
rect -4376 -14472 -4360 -14408
rect -4456 -14488 -4360 -14472
rect -4456 -14552 -4440 -14488
rect -4376 -14552 -4360 -14488
rect -4456 -14568 -4360 -14552
rect -4456 -14632 -4440 -14568
rect -4376 -14632 -4360 -14568
rect -4456 -14648 -4360 -14632
rect -4456 -14712 -4440 -14648
rect -4376 -14712 -4360 -14648
rect -4456 -14728 -4360 -14712
rect -4456 -14792 -4440 -14728
rect -4376 -14792 -4360 -14728
rect -4456 -14808 -4360 -14792
rect -4456 -14872 -4440 -14808
rect -4376 -14872 -4360 -14808
rect -4456 -14888 -4360 -14872
rect -5868 -14988 -5772 -14952
rect -4456 -14952 -4440 -14888
rect -4376 -14952 -4360 -14888
rect -4037 -14208 -3315 -14199
rect -4037 -14912 -4028 -14208
rect -3324 -14912 -3315 -14208
rect -4037 -14921 -3315 -14912
rect -3044 -14232 -3028 -14168
rect -2964 -14232 -2948 -14168
rect -1632 -14168 -1536 -14132
rect -3044 -14248 -2948 -14232
rect -3044 -14312 -3028 -14248
rect -2964 -14312 -2948 -14248
rect -3044 -14328 -2948 -14312
rect -3044 -14392 -3028 -14328
rect -2964 -14392 -2948 -14328
rect -3044 -14408 -2948 -14392
rect -3044 -14472 -3028 -14408
rect -2964 -14472 -2948 -14408
rect -3044 -14488 -2948 -14472
rect -3044 -14552 -3028 -14488
rect -2964 -14552 -2948 -14488
rect -3044 -14568 -2948 -14552
rect -3044 -14632 -3028 -14568
rect -2964 -14632 -2948 -14568
rect -3044 -14648 -2948 -14632
rect -3044 -14712 -3028 -14648
rect -2964 -14712 -2948 -14648
rect -3044 -14728 -2948 -14712
rect -3044 -14792 -3028 -14728
rect -2964 -14792 -2948 -14728
rect -3044 -14808 -2948 -14792
rect -3044 -14872 -3028 -14808
rect -2964 -14872 -2948 -14808
rect -3044 -14888 -2948 -14872
rect -4456 -14988 -4360 -14952
rect -3044 -14952 -3028 -14888
rect -2964 -14952 -2948 -14888
rect -2625 -14208 -1903 -14199
rect -2625 -14912 -2616 -14208
rect -1912 -14912 -1903 -14208
rect -2625 -14921 -1903 -14912
rect -1632 -14232 -1616 -14168
rect -1552 -14232 -1536 -14168
rect -220 -14168 -124 -14132
rect -1632 -14248 -1536 -14232
rect -1632 -14312 -1616 -14248
rect -1552 -14312 -1536 -14248
rect -1632 -14328 -1536 -14312
rect -1632 -14392 -1616 -14328
rect -1552 -14392 -1536 -14328
rect -1632 -14408 -1536 -14392
rect -1632 -14472 -1616 -14408
rect -1552 -14472 -1536 -14408
rect -1632 -14488 -1536 -14472
rect -1632 -14552 -1616 -14488
rect -1552 -14552 -1536 -14488
rect -1632 -14568 -1536 -14552
rect -1632 -14632 -1616 -14568
rect -1552 -14632 -1536 -14568
rect -1632 -14648 -1536 -14632
rect -1632 -14712 -1616 -14648
rect -1552 -14712 -1536 -14648
rect -1632 -14728 -1536 -14712
rect -1632 -14792 -1616 -14728
rect -1552 -14792 -1536 -14728
rect -1632 -14808 -1536 -14792
rect -1632 -14872 -1616 -14808
rect -1552 -14872 -1536 -14808
rect -1632 -14888 -1536 -14872
rect -3044 -14988 -2948 -14952
rect -1632 -14952 -1616 -14888
rect -1552 -14952 -1536 -14888
rect -1213 -14208 -491 -14199
rect -1213 -14912 -1204 -14208
rect -500 -14912 -491 -14208
rect -1213 -14921 -491 -14912
rect -220 -14232 -204 -14168
rect -140 -14232 -124 -14168
rect 1192 -14168 1288 -14132
rect -220 -14248 -124 -14232
rect -220 -14312 -204 -14248
rect -140 -14312 -124 -14248
rect -220 -14328 -124 -14312
rect -220 -14392 -204 -14328
rect -140 -14392 -124 -14328
rect -220 -14408 -124 -14392
rect -220 -14472 -204 -14408
rect -140 -14472 -124 -14408
rect -220 -14488 -124 -14472
rect -220 -14552 -204 -14488
rect -140 -14552 -124 -14488
rect -220 -14568 -124 -14552
rect -220 -14632 -204 -14568
rect -140 -14632 -124 -14568
rect -220 -14648 -124 -14632
rect -220 -14712 -204 -14648
rect -140 -14712 -124 -14648
rect -220 -14728 -124 -14712
rect -220 -14792 -204 -14728
rect -140 -14792 -124 -14728
rect -220 -14808 -124 -14792
rect -220 -14872 -204 -14808
rect -140 -14872 -124 -14808
rect -220 -14888 -124 -14872
rect -1632 -14988 -1536 -14952
rect -220 -14952 -204 -14888
rect -140 -14952 -124 -14888
rect 199 -14208 921 -14199
rect 199 -14912 208 -14208
rect 912 -14912 921 -14208
rect 199 -14921 921 -14912
rect 1192 -14232 1208 -14168
rect 1272 -14232 1288 -14168
rect 2604 -14168 2700 -14132
rect 1192 -14248 1288 -14232
rect 1192 -14312 1208 -14248
rect 1272 -14312 1288 -14248
rect 1192 -14328 1288 -14312
rect 1192 -14392 1208 -14328
rect 1272 -14392 1288 -14328
rect 1192 -14408 1288 -14392
rect 1192 -14472 1208 -14408
rect 1272 -14472 1288 -14408
rect 1192 -14488 1288 -14472
rect 1192 -14552 1208 -14488
rect 1272 -14552 1288 -14488
rect 1192 -14568 1288 -14552
rect 1192 -14632 1208 -14568
rect 1272 -14632 1288 -14568
rect 1192 -14648 1288 -14632
rect 1192 -14712 1208 -14648
rect 1272 -14712 1288 -14648
rect 1192 -14728 1288 -14712
rect 1192 -14792 1208 -14728
rect 1272 -14792 1288 -14728
rect 1192 -14808 1288 -14792
rect 1192 -14872 1208 -14808
rect 1272 -14872 1288 -14808
rect 1192 -14888 1288 -14872
rect -220 -14988 -124 -14952
rect 1192 -14952 1208 -14888
rect 1272 -14952 1288 -14888
rect 1611 -14208 2333 -14199
rect 1611 -14912 1620 -14208
rect 2324 -14912 2333 -14208
rect 1611 -14921 2333 -14912
rect 2604 -14232 2620 -14168
rect 2684 -14232 2700 -14168
rect 4016 -14168 4112 -14132
rect 2604 -14248 2700 -14232
rect 2604 -14312 2620 -14248
rect 2684 -14312 2700 -14248
rect 2604 -14328 2700 -14312
rect 2604 -14392 2620 -14328
rect 2684 -14392 2700 -14328
rect 2604 -14408 2700 -14392
rect 2604 -14472 2620 -14408
rect 2684 -14472 2700 -14408
rect 2604 -14488 2700 -14472
rect 2604 -14552 2620 -14488
rect 2684 -14552 2700 -14488
rect 2604 -14568 2700 -14552
rect 2604 -14632 2620 -14568
rect 2684 -14632 2700 -14568
rect 2604 -14648 2700 -14632
rect 2604 -14712 2620 -14648
rect 2684 -14712 2700 -14648
rect 2604 -14728 2700 -14712
rect 2604 -14792 2620 -14728
rect 2684 -14792 2700 -14728
rect 2604 -14808 2700 -14792
rect 2604 -14872 2620 -14808
rect 2684 -14872 2700 -14808
rect 2604 -14888 2700 -14872
rect 1192 -14988 1288 -14952
rect 2604 -14952 2620 -14888
rect 2684 -14952 2700 -14888
rect 3023 -14208 3745 -14199
rect 3023 -14912 3032 -14208
rect 3736 -14912 3745 -14208
rect 3023 -14921 3745 -14912
rect 4016 -14232 4032 -14168
rect 4096 -14232 4112 -14168
rect 5428 -14168 5524 -14132
rect 4016 -14248 4112 -14232
rect 4016 -14312 4032 -14248
rect 4096 -14312 4112 -14248
rect 4016 -14328 4112 -14312
rect 4016 -14392 4032 -14328
rect 4096 -14392 4112 -14328
rect 4016 -14408 4112 -14392
rect 4016 -14472 4032 -14408
rect 4096 -14472 4112 -14408
rect 4016 -14488 4112 -14472
rect 4016 -14552 4032 -14488
rect 4096 -14552 4112 -14488
rect 4016 -14568 4112 -14552
rect 4016 -14632 4032 -14568
rect 4096 -14632 4112 -14568
rect 4016 -14648 4112 -14632
rect 4016 -14712 4032 -14648
rect 4096 -14712 4112 -14648
rect 4016 -14728 4112 -14712
rect 4016 -14792 4032 -14728
rect 4096 -14792 4112 -14728
rect 4016 -14808 4112 -14792
rect 4016 -14872 4032 -14808
rect 4096 -14872 4112 -14808
rect 4016 -14888 4112 -14872
rect 2604 -14988 2700 -14952
rect 4016 -14952 4032 -14888
rect 4096 -14952 4112 -14888
rect 4435 -14208 5157 -14199
rect 4435 -14912 4444 -14208
rect 5148 -14912 5157 -14208
rect 4435 -14921 5157 -14912
rect 5428 -14232 5444 -14168
rect 5508 -14232 5524 -14168
rect 6840 -14168 6936 -14132
rect 5428 -14248 5524 -14232
rect 5428 -14312 5444 -14248
rect 5508 -14312 5524 -14248
rect 5428 -14328 5524 -14312
rect 5428 -14392 5444 -14328
rect 5508 -14392 5524 -14328
rect 5428 -14408 5524 -14392
rect 5428 -14472 5444 -14408
rect 5508 -14472 5524 -14408
rect 5428 -14488 5524 -14472
rect 5428 -14552 5444 -14488
rect 5508 -14552 5524 -14488
rect 5428 -14568 5524 -14552
rect 5428 -14632 5444 -14568
rect 5508 -14632 5524 -14568
rect 5428 -14648 5524 -14632
rect 5428 -14712 5444 -14648
rect 5508 -14712 5524 -14648
rect 5428 -14728 5524 -14712
rect 5428 -14792 5444 -14728
rect 5508 -14792 5524 -14728
rect 5428 -14808 5524 -14792
rect 5428 -14872 5444 -14808
rect 5508 -14872 5524 -14808
rect 5428 -14888 5524 -14872
rect 4016 -14988 4112 -14952
rect 5428 -14952 5444 -14888
rect 5508 -14952 5524 -14888
rect 5847 -14208 6569 -14199
rect 5847 -14912 5856 -14208
rect 6560 -14912 6569 -14208
rect 5847 -14921 6569 -14912
rect 6840 -14232 6856 -14168
rect 6920 -14232 6936 -14168
rect 8252 -14168 8348 -14132
rect 6840 -14248 6936 -14232
rect 6840 -14312 6856 -14248
rect 6920 -14312 6936 -14248
rect 6840 -14328 6936 -14312
rect 6840 -14392 6856 -14328
rect 6920 -14392 6936 -14328
rect 6840 -14408 6936 -14392
rect 6840 -14472 6856 -14408
rect 6920 -14472 6936 -14408
rect 6840 -14488 6936 -14472
rect 6840 -14552 6856 -14488
rect 6920 -14552 6936 -14488
rect 6840 -14568 6936 -14552
rect 6840 -14632 6856 -14568
rect 6920 -14632 6936 -14568
rect 6840 -14648 6936 -14632
rect 6840 -14712 6856 -14648
rect 6920 -14712 6936 -14648
rect 6840 -14728 6936 -14712
rect 6840 -14792 6856 -14728
rect 6920 -14792 6936 -14728
rect 6840 -14808 6936 -14792
rect 6840 -14872 6856 -14808
rect 6920 -14872 6936 -14808
rect 6840 -14888 6936 -14872
rect 5428 -14988 5524 -14952
rect 6840 -14952 6856 -14888
rect 6920 -14952 6936 -14888
rect 7259 -14208 7981 -14199
rect 7259 -14912 7268 -14208
rect 7972 -14912 7981 -14208
rect 7259 -14921 7981 -14912
rect 8252 -14232 8268 -14168
rect 8332 -14232 8348 -14168
rect 9664 -14168 9760 -14132
rect 8252 -14248 8348 -14232
rect 8252 -14312 8268 -14248
rect 8332 -14312 8348 -14248
rect 8252 -14328 8348 -14312
rect 8252 -14392 8268 -14328
rect 8332 -14392 8348 -14328
rect 8252 -14408 8348 -14392
rect 8252 -14472 8268 -14408
rect 8332 -14472 8348 -14408
rect 8252 -14488 8348 -14472
rect 8252 -14552 8268 -14488
rect 8332 -14552 8348 -14488
rect 8252 -14568 8348 -14552
rect 8252 -14632 8268 -14568
rect 8332 -14632 8348 -14568
rect 8252 -14648 8348 -14632
rect 8252 -14712 8268 -14648
rect 8332 -14712 8348 -14648
rect 8252 -14728 8348 -14712
rect 8252 -14792 8268 -14728
rect 8332 -14792 8348 -14728
rect 8252 -14808 8348 -14792
rect 8252 -14872 8268 -14808
rect 8332 -14872 8348 -14808
rect 8252 -14888 8348 -14872
rect 6840 -14988 6936 -14952
rect 8252 -14952 8268 -14888
rect 8332 -14952 8348 -14888
rect 8671 -14208 9393 -14199
rect 8671 -14912 8680 -14208
rect 9384 -14912 9393 -14208
rect 8671 -14921 9393 -14912
rect 9664 -14232 9680 -14168
rect 9744 -14232 9760 -14168
rect 11076 -14168 11172 -14132
rect 9664 -14248 9760 -14232
rect 9664 -14312 9680 -14248
rect 9744 -14312 9760 -14248
rect 9664 -14328 9760 -14312
rect 9664 -14392 9680 -14328
rect 9744 -14392 9760 -14328
rect 9664 -14408 9760 -14392
rect 9664 -14472 9680 -14408
rect 9744 -14472 9760 -14408
rect 9664 -14488 9760 -14472
rect 9664 -14552 9680 -14488
rect 9744 -14552 9760 -14488
rect 9664 -14568 9760 -14552
rect 9664 -14632 9680 -14568
rect 9744 -14632 9760 -14568
rect 9664 -14648 9760 -14632
rect 9664 -14712 9680 -14648
rect 9744 -14712 9760 -14648
rect 9664 -14728 9760 -14712
rect 9664 -14792 9680 -14728
rect 9744 -14792 9760 -14728
rect 9664 -14808 9760 -14792
rect 9664 -14872 9680 -14808
rect 9744 -14872 9760 -14808
rect 9664 -14888 9760 -14872
rect 8252 -14988 8348 -14952
rect 9664 -14952 9680 -14888
rect 9744 -14952 9760 -14888
rect 10083 -14208 10805 -14199
rect 10083 -14912 10092 -14208
rect 10796 -14912 10805 -14208
rect 10083 -14921 10805 -14912
rect 11076 -14232 11092 -14168
rect 11156 -14232 11172 -14168
rect 12488 -14168 12584 -14132
rect 11076 -14248 11172 -14232
rect 11076 -14312 11092 -14248
rect 11156 -14312 11172 -14248
rect 11076 -14328 11172 -14312
rect 11076 -14392 11092 -14328
rect 11156 -14392 11172 -14328
rect 11076 -14408 11172 -14392
rect 11076 -14472 11092 -14408
rect 11156 -14472 11172 -14408
rect 11076 -14488 11172 -14472
rect 11076 -14552 11092 -14488
rect 11156 -14552 11172 -14488
rect 11076 -14568 11172 -14552
rect 11076 -14632 11092 -14568
rect 11156 -14632 11172 -14568
rect 11076 -14648 11172 -14632
rect 11076 -14712 11092 -14648
rect 11156 -14712 11172 -14648
rect 11076 -14728 11172 -14712
rect 11076 -14792 11092 -14728
rect 11156 -14792 11172 -14728
rect 11076 -14808 11172 -14792
rect 11076 -14872 11092 -14808
rect 11156 -14872 11172 -14808
rect 11076 -14888 11172 -14872
rect 9664 -14988 9760 -14952
rect 11076 -14952 11092 -14888
rect 11156 -14952 11172 -14888
rect 11495 -14208 12217 -14199
rect 11495 -14912 11504 -14208
rect 12208 -14912 12217 -14208
rect 11495 -14921 12217 -14912
rect 12488 -14232 12504 -14168
rect 12568 -14232 12584 -14168
rect 13900 -14168 13996 -14132
rect 12488 -14248 12584 -14232
rect 12488 -14312 12504 -14248
rect 12568 -14312 12584 -14248
rect 12488 -14328 12584 -14312
rect 12488 -14392 12504 -14328
rect 12568 -14392 12584 -14328
rect 12488 -14408 12584 -14392
rect 12488 -14472 12504 -14408
rect 12568 -14472 12584 -14408
rect 12488 -14488 12584 -14472
rect 12488 -14552 12504 -14488
rect 12568 -14552 12584 -14488
rect 12488 -14568 12584 -14552
rect 12488 -14632 12504 -14568
rect 12568 -14632 12584 -14568
rect 12488 -14648 12584 -14632
rect 12488 -14712 12504 -14648
rect 12568 -14712 12584 -14648
rect 12488 -14728 12584 -14712
rect 12488 -14792 12504 -14728
rect 12568 -14792 12584 -14728
rect 12488 -14808 12584 -14792
rect 12488 -14872 12504 -14808
rect 12568 -14872 12584 -14808
rect 12488 -14888 12584 -14872
rect 11076 -14988 11172 -14952
rect 12488 -14952 12504 -14888
rect 12568 -14952 12584 -14888
rect 12907 -14208 13629 -14199
rect 12907 -14912 12916 -14208
rect 13620 -14912 13629 -14208
rect 12907 -14921 13629 -14912
rect 13900 -14232 13916 -14168
rect 13980 -14232 13996 -14168
rect 15312 -14168 15408 -14132
rect 13900 -14248 13996 -14232
rect 13900 -14312 13916 -14248
rect 13980 -14312 13996 -14248
rect 13900 -14328 13996 -14312
rect 13900 -14392 13916 -14328
rect 13980 -14392 13996 -14328
rect 13900 -14408 13996 -14392
rect 13900 -14472 13916 -14408
rect 13980 -14472 13996 -14408
rect 13900 -14488 13996 -14472
rect 13900 -14552 13916 -14488
rect 13980 -14552 13996 -14488
rect 13900 -14568 13996 -14552
rect 13900 -14632 13916 -14568
rect 13980 -14632 13996 -14568
rect 13900 -14648 13996 -14632
rect 13900 -14712 13916 -14648
rect 13980 -14712 13996 -14648
rect 13900 -14728 13996 -14712
rect 13900 -14792 13916 -14728
rect 13980 -14792 13996 -14728
rect 13900 -14808 13996 -14792
rect 13900 -14872 13916 -14808
rect 13980 -14872 13996 -14808
rect 13900 -14888 13996 -14872
rect 12488 -14988 12584 -14952
rect 13900 -14952 13916 -14888
rect 13980 -14952 13996 -14888
rect 14319 -14208 15041 -14199
rect 14319 -14912 14328 -14208
rect 15032 -14912 15041 -14208
rect 14319 -14921 15041 -14912
rect 15312 -14232 15328 -14168
rect 15392 -14232 15408 -14168
rect 16724 -14168 16820 -14132
rect 15312 -14248 15408 -14232
rect 15312 -14312 15328 -14248
rect 15392 -14312 15408 -14248
rect 15312 -14328 15408 -14312
rect 15312 -14392 15328 -14328
rect 15392 -14392 15408 -14328
rect 15312 -14408 15408 -14392
rect 15312 -14472 15328 -14408
rect 15392 -14472 15408 -14408
rect 15312 -14488 15408 -14472
rect 15312 -14552 15328 -14488
rect 15392 -14552 15408 -14488
rect 15312 -14568 15408 -14552
rect 15312 -14632 15328 -14568
rect 15392 -14632 15408 -14568
rect 15312 -14648 15408 -14632
rect 15312 -14712 15328 -14648
rect 15392 -14712 15408 -14648
rect 15312 -14728 15408 -14712
rect 15312 -14792 15328 -14728
rect 15392 -14792 15408 -14728
rect 15312 -14808 15408 -14792
rect 15312 -14872 15328 -14808
rect 15392 -14872 15408 -14808
rect 15312 -14888 15408 -14872
rect 13900 -14988 13996 -14952
rect 15312 -14952 15328 -14888
rect 15392 -14952 15408 -14888
rect 15731 -14208 16453 -14199
rect 15731 -14912 15740 -14208
rect 16444 -14912 16453 -14208
rect 15731 -14921 16453 -14912
rect 16724 -14232 16740 -14168
rect 16804 -14232 16820 -14168
rect 18136 -14168 18232 -14132
rect 16724 -14248 16820 -14232
rect 16724 -14312 16740 -14248
rect 16804 -14312 16820 -14248
rect 16724 -14328 16820 -14312
rect 16724 -14392 16740 -14328
rect 16804 -14392 16820 -14328
rect 16724 -14408 16820 -14392
rect 16724 -14472 16740 -14408
rect 16804 -14472 16820 -14408
rect 16724 -14488 16820 -14472
rect 16724 -14552 16740 -14488
rect 16804 -14552 16820 -14488
rect 16724 -14568 16820 -14552
rect 16724 -14632 16740 -14568
rect 16804 -14632 16820 -14568
rect 16724 -14648 16820 -14632
rect 16724 -14712 16740 -14648
rect 16804 -14712 16820 -14648
rect 16724 -14728 16820 -14712
rect 16724 -14792 16740 -14728
rect 16804 -14792 16820 -14728
rect 16724 -14808 16820 -14792
rect 16724 -14872 16740 -14808
rect 16804 -14872 16820 -14808
rect 16724 -14888 16820 -14872
rect 15312 -14988 15408 -14952
rect 16724 -14952 16740 -14888
rect 16804 -14952 16820 -14888
rect 17143 -14208 17865 -14199
rect 17143 -14912 17152 -14208
rect 17856 -14912 17865 -14208
rect 17143 -14921 17865 -14912
rect 18136 -14232 18152 -14168
rect 18216 -14232 18232 -14168
rect 19548 -14168 19644 -14132
rect 18136 -14248 18232 -14232
rect 18136 -14312 18152 -14248
rect 18216 -14312 18232 -14248
rect 18136 -14328 18232 -14312
rect 18136 -14392 18152 -14328
rect 18216 -14392 18232 -14328
rect 18136 -14408 18232 -14392
rect 18136 -14472 18152 -14408
rect 18216 -14472 18232 -14408
rect 18136 -14488 18232 -14472
rect 18136 -14552 18152 -14488
rect 18216 -14552 18232 -14488
rect 18136 -14568 18232 -14552
rect 18136 -14632 18152 -14568
rect 18216 -14632 18232 -14568
rect 18136 -14648 18232 -14632
rect 18136 -14712 18152 -14648
rect 18216 -14712 18232 -14648
rect 18136 -14728 18232 -14712
rect 18136 -14792 18152 -14728
rect 18216 -14792 18232 -14728
rect 18136 -14808 18232 -14792
rect 18136 -14872 18152 -14808
rect 18216 -14872 18232 -14808
rect 18136 -14888 18232 -14872
rect 16724 -14988 16820 -14952
rect 18136 -14952 18152 -14888
rect 18216 -14952 18232 -14888
rect 18555 -14208 19277 -14199
rect 18555 -14912 18564 -14208
rect 19268 -14912 19277 -14208
rect 18555 -14921 19277 -14912
rect 19548 -14232 19564 -14168
rect 19628 -14232 19644 -14168
rect 20960 -14168 21056 -14132
rect 19548 -14248 19644 -14232
rect 19548 -14312 19564 -14248
rect 19628 -14312 19644 -14248
rect 19548 -14328 19644 -14312
rect 19548 -14392 19564 -14328
rect 19628 -14392 19644 -14328
rect 19548 -14408 19644 -14392
rect 19548 -14472 19564 -14408
rect 19628 -14472 19644 -14408
rect 19548 -14488 19644 -14472
rect 19548 -14552 19564 -14488
rect 19628 -14552 19644 -14488
rect 19548 -14568 19644 -14552
rect 19548 -14632 19564 -14568
rect 19628 -14632 19644 -14568
rect 19548 -14648 19644 -14632
rect 19548 -14712 19564 -14648
rect 19628 -14712 19644 -14648
rect 19548 -14728 19644 -14712
rect 19548 -14792 19564 -14728
rect 19628 -14792 19644 -14728
rect 19548 -14808 19644 -14792
rect 19548 -14872 19564 -14808
rect 19628 -14872 19644 -14808
rect 19548 -14888 19644 -14872
rect 18136 -14988 18232 -14952
rect 19548 -14952 19564 -14888
rect 19628 -14952 19644 -14888
rect 19967 -14208 20689 -14199
rect 19967 -14912 19976 -14208
rect 20680 -14912 20689 -14208
rect 19967 -14921 20689 -14912
rect 20960 -14232 20976 -14168
rect 21040 -14232 21056 -14168
rect 22372 -14168 22468 -14132
rect 20960 -14248 21056 -14232
rect 20960 -14312 20976 -14248
rect 21040 -14312 21056 -14248
rect 20960 -14328 21056 -14312
rect 20960 -14392 20976 -14328
rect 21040 -14392 21056 -14328
rect 20960 -14408 21056 -14392
rect 20960 -14472 20976 -14408
rect 21040 -14472 21056 -14408
rect 20960 -14488 21056 -14472
rect 20960 -14552 20976 -14488
rect 21040 -14552 21056 -14488
rect 20960 -14568 21056 -14552
rect 20960 -14632 20976 -14568
rect 21040 -14632 21056 -14568
rect 20960 -14648 21056 -14632
rect 20960 -14712 20976 -14648
rect 21040 -14712 21056 -14648
rect 20960 -14728 21056 -14712
rect 20960 -14792 20976 -14728
rect 21040 -14792 21056 -14728
rect 20960 -14808 21056 -14792
rect 20960 -14872 20976 -14808
rect 21040 -14872 21056 -14808
rect 20960 -14888 21056 -14872
rect 19548 -14988 19644 -14952
rect 20960 -14952 20976 -14888
rect 21040 -14952 21056 -14888
rect 21379 -14208 22101 -14199
rect 21379 -14912 21388 -14208
rect 22092 -14912 22101 -14208
rect 21379 -14921 22101 -14912
rect 22372 -14232 22388 -14168
rect 22452 -14232 22468 -14168
rect 23784 -14168 23880 -14132
rect 22372 -14248 22468 -14232
rect 22372 -14312 22388 -14248
rect 22452 -14312 22468 -14248
rect 22372 -14328 22468 -14312
rect 22372 -14392 22388 -14328
rect 22452 -14392 22468 -14328
rect 22372 -14408 22468 -14392
rect 22372 -14472 22388 -14408
rect 22452 -14472 22468 -14408
rect 22372 -14488 22468 -14472
rect 22372 -14552 22388 -14488
rect 22452 -14552 22468 -14488
rect 22372 -14568 22468 -14552
rect 22372 -14632 22388 -14568
rect 22452 -14632 22468 -14568
rect 22372 -14648 22468 -14632
rect 22372 -14712 22388 -14648
rect 22452 -14712 22468 -14648
rect 22372 -14728 22468 -14712
rect 22372 -14792 22388 -14728
rect 22452 -14792 22468 -14728
rect 22372 -14808 22468 -14792
rect 22372 -14872 22388 -14808
rect 22452 -14872 22468 -14808
rect 22372 -14888 22468 -14872
rect 20960 -14988 21056 -14952
rect 22372 -14952 22388 -14888
rect 22452 -14952 22468 -14888
rect 22791 -14208 23513 -14199
rect 22791 -14912 22800 -14208
rect 23504 -14912 23513 -14208
rect 22791 -14921 23513 -14912
rect 23784 -14232 23800 -14168
rect 23864 -14232 23880 -14168
rect 23784 -14248 23880 -14232
rect 23784 -14312 23800 -14248
rect 23864 -14312 23880 -14248
rect 23784 -14328 23880 -14312
rect 23784 -14392 23800 -14328
rect 23864 -14392 23880 -14328
rect 23784 -14408 23880 -14392
rect 23784 -14472 23800 -14408
rect 23864 -14472 23880 -14408
rect 23784 -14488 23880 -14472
rect 23784 -14552 23800 -14488
rect 23864 -14552 23880 -14488
rect 23784 -14568 23880 -14552
rect 23784 -14632 23800 -14568
rect 23864 -14632 23880 -14568
rect 23784 -14648 23880 -14632
rect 23784 -14712 23800 -14648
rect 23864 -14712 23880 -14648
rect 23784 -14728 23880 -14712
rect 23784 -14792 23800 -14728
rect 23864 -14792 23880 -14728
rect 23784 -14808 23880 -14792
rect 23784 -14872 23800 -14808
rect 23864 -14872 23880 -14808
rect 23784 -14888 23880 -14872
rect 22372 -14988 22468 -14952
rect 23784 -14952 23800 -14888
rect 23864 -14952 23880 -14888
rect 23784 -14988 23880 -14952
rect -22812 -15288 -22716 -15252
rect -23805 -15328 -23083 -15319
rect -23805 -16032 -23796 -15328
rect -23092 -16032 -23083 -15328
rect -23805 -16041 -23083 -16032
rect -22812 -15352 -22796 -15288
rect -22732 -15352 -22716 -15288
rect -21400 -15288 -21304 -15252
rect -22812 -15368 -22716 -15352
rect -22812 -15432 -22796 -15368
rect -22732 -15432 -22716 -15368
rect -22812 -15448 -22716 -15432
rect -22812 -15512 -22796 -15448
rect -22732 -15512 -22716 -15448
rect -22812 -15528 -22716 -15512
rect -22812 -15592 -22796 -15528
rect -22732 -15592 -22716 -15528
rect -22812 -15608 -22716 -15592
rect -22812 -15672 -22796 -15608
rect -22732 -15672 -22716 -15608
rect -22812 -15688 -22716 -15672
rect -22812 -15752 -22796 -15688
rect -22732 -15752 -22716 -15688
rect -22812 -15768 -22716 -15752
rect -22812 -15832 -22796 -15768
rect -22732 -15832 -22716 -15768
rect -22812 -15848 -22716 -15832
rect -22812 -15912 -22796 -15848
rect -22732 -15912 -22716 -15848
rect -22812 -15928 -22716 -15912
rect -22812 -15992 -22796 -15928
rect -22732 -15992 -22716 -15928
rect -22812 -16008 -22716 -15992
rect -22812 -16072 -22796 -16008
rect -22732 -16072 -22716 -16008
rect -22393 -15328 -21671 -15319
rect -22393 -16032 -22384 -15328
rect -21680 -16032 -21671 -15328
rect -22393 -16041 -21671 -16032
rect -21400 -15352 -21384 -15288
rect -21320 -15352 -21304 -15288
rect -19988 -15288 -19892 -15252
rect -21400 -15368 -21304 -15352
rect -21400 -15432 -21384 -15368
rect -21320 -15432 -21304 -15368
rect -21400 -15448 -21304 -15432
rect -21400 -15512 -21384 -15448
rect -21320 -15512 -21304 -15448
rect -21400 -15528 -21304 -15512
rect -21400 -15592 -21384 -15528
rect -21320 -15592 -21304 -15528
rect -21400 -15608 -21304 -15592
rect -21400 -15672 -21384 -15608
rect -21320 -15672 -21304 -15608
rect -21400 -15688 -21304 -15672
rect -21400 -15752 -21384 -15688
rect -21320 -15752 -21304 -15688
rect -21400 -15768 -21304 -15752
rect -21400 -15832 -21384 -15768
rect -21320 -15832 -21304 -15768
rect -21400 -15848 -21304 -15832
rect -21400 -15912 -21384 -15848
rect -21320 -15912 -21304 -15848
rect -21400 -15928 -21304 -15912
rect -21400 -15992 -21384 -15928
rect -21320 -15992 -21304 -15928
rect -21400 -16008 -21304 -15992
rect -22812 -16108 -22716 -16072
rect -21400 -16072 -21384 -16008
rect -21320 -16072 -21304 -16008
rect -20981 -15328 -20259 -15319
rect -20981 -16032 -20972 -15328
rect -20268 -16032 -20259 -15328
rect -20981 -16041 -20259 -16032
rect -19988 -15352 -19972 -15288
rect -19908 -15352 -19892 -15288
rect -18576 -15288 -18480 -15252
rect -19988 -15368 -19892 -15352
rect -19988 -15432 -19972 -15368
rect -19908 -15432 -19892 -15368
rect -19988 -15448 -19892 -15432
rect -19988 -15512 -19972 -15448
rect -19908 -15512 -19892 -15448
rect -19988 -15528 -19892 -15512
rect -19988 -15592 -19972 -15528
rect -19908 -15592 -19892 -15528
rect -19988 -15608 -19892 -15592
rect -19988 -15672 -19972 -15608
rect -19908 -15672 -19892 -15608
rect -19988 -15688 -19892 -15672
rect -19988 -15752 -19972 -15688
rect -19908 -15752 -19892 -15688
rect -19988 -15768 -19892 -15752
rect -19988 -15832 -19972 -15768
rect -19908 -15832 -19892 -15768
rect -19988 -15848 -19892 -15832
rect -19988 -15912 -19972 -15848
rect -19908 -15912 -19892 -15848
rect -19988 -15928 -19892 -15912
rect -19988 -15992 -19972 -15928
rect -19908 -15992 -19892 -15928
rect -19988 -16008 -19892 -15992
rect -21400 -16108 -21304 -16072
rect -19988 -16072 -19972 -16008
rect -19908 -16072 -19892 -16008
rect -19569 -15328 -18847 -15319
rect -19569 -16032 -19560 -15328
rect -18856 -16032 -18847 -15328
rect -19569 -16041 -18847 -16032
rect -18576 -15352 -18560 -15288
rect -18496 -15352 -18480 -15288
rect -17164 -15288 -17068 -15252
rect -18576 -15368 -18480 -15352
rect -18576 -15432 -18560 -15368
rect -18496 -15432 -18480 -15368
rect -18576 -15448 -18480 -15432
rect -18576 -15512 -18560 -15448
rect -18496 -15512 -18480 -15448
rect -18576 -15528 -18480 -15512
rect -18576 -15592 -18560 -15528
rect -18496 -15592 -18480 -15528
rect -18576 -15608 -18480 -15592
rect -18576 -15672 -18560 -15608
rect -18496 -15672 -18480 -15608
rect -18576 -15688 -18480 -15672
rect -18576 -15752 -18560 -15688
rect -18496 -15752 -18480 -15688
rect -18576 -15768 -18480 -15752
rect -18576 -15832 -18560 -15768
rect -18496 -15832 -18480 -15768
rect -18576 -15848 -18480 -15832
rect -18576 -15912 -18560 -15848
rect -18496 -15912 -18480 -15848
rect -18576 -15928 -18480 -15912
rect -18576 -15992 -18560 -15928
rect -18496 -15992 -18480 -15928
rect -18576 -16008 -18480 -15992
rect -19988 -16108 -19892 -16072
rect -18576 -16072 -18560 -16008
rect -18496 -16072 -18480 -16008
rect -18157 -15328 -17435 -15319
rect -18157 -16032 -18148 -15328
rect -17444 -16032 -17435 -15328
rect -18157 -16041 -17435 -16032
rect -17164 -15352 -17148 -15288
rect -17084 -15352 -17068 -15288
rect -15752 -15288 -15656 -15252
rect -17164 -15368 -17068 -15352
rect -17164 -15432 -17148 -15368
rect -17084 -15432 -17068 -15368
rect -17164 -15448 -17068 -15432
rect -17164 -15512 -17148 -15448
rect -17084 -15512 -17068 -15448
rect -17164 -15528 -17068 -15512
rect -17164 -15592 -17148 -15528
rect -17084 -15592 -17068 -15528
rect -17164 -15608 -17068 -15592
rect -17164 -15672 -17148 -15608
rect -17084 -15672 -17068 -15608
rect -17164 -15688 -17068 -15672
rect -17164 -15752 -17148 -15688
rect -17084 -15752 -17068 -15688
rect -17164 -15768 -17068 -15752
rect -17164 -15832 -17148 -15768
rect -17084 -15832 -17068 -15768
rect -17164 -15848 -17068 -15832
rect -17164 -15912 -17148 -15848
rect -17084 -15912 -17068 -15848
rect -17164 -15928 -17068 -15912
rect -17164 -15992 -17148 -15928
rect -17084 -15992 -17068 -15928
rect -17164 -16008 -17068 -15992
rect -18576 -16108 -18480 -16072
rect -17164 -16072 -17148 -16008
rect -17084 -16072 -17068 -16008
rect -16745 -15328 -16023 -15319
rect -16745 -16032 -16736 -15328
rect -16032 -16032 -16023 -15328
rect -16745 -16041 -16023 -16032
rect -15752 -15352 -15736 -15288
rect -15672 -15352 -15656 -15288
rect -14340 -15288 -14244 -15252
rect -15752 -15368 -15656 -15352
rect -15752 -15432 -15736 -15368
rect -15672 -15432 -15656 -15368
rect -15752 -15448 -15656 -15432
rect -15752 -15512 -15736 -15448
rect -15672 -15512 -15656 -15448
rect -15752 -15528 -15656 -15512
rect -15752 -15592 -15736 -15528
rect -15672 -15592 -15656 -15528
rect -15752 -15608 -15656 -15592
rect -15752 -15672 -15736 -15608
rect -15672 -15672 -15656 -15608
rect -15752 -15688 -15656 -15672
rect -15752 -15752 -15736 -15688
rect -15672 -15752 -15656 -15688
rect -15752 -15768 -15656 -15752
rect -15752 -15832 -15736 -15768
rect -15672 -15832 -15656 -15768
rect -15752 -15848 -15656 -15832
rect -15752 -15912 -15736 -15848
rect -15672 -15912 -15656 -15848
rect -15752 -15928 -15656 -15912
rect -15752 -15992 -15736 -15928
rect -15672 -15992 -15656 -15928
rect -15752 -16008 -15656 -15992
rect -17164 -16108 -17068 -16072
rect -15752 -16072 -15736 -16008
rect -15672 -16072 -15656 -16008
rect -15333 -15328 -14611 -15319
rect -15333 -16032 -15324 -15328
rect -14620 -16032 -14611 -15328
rect -15333 -16041 -14611 -16032
rect -14340 -15352 -14324 -15288
rect -14260 -15352 -14244 -15288
rect -12928 -15288 -12832 -15252
rect -14340 -15368 -14244 -15352
rect -14340 -15432 -14324 -15368
rect -14260 -15432 -14244 -15368
rect -14340 -15448 -14244 -15432
rect -14340 -15512 -14324 -15448
rect -14260 -15512 -14244 -15448
rect -14340 -15528 -14244 -15512
rect -14340 -15592 -14324 -15528
rect -14260 -15592 -14244 -15528
rect -14340 -15608 -14244 -15592
rect -14340 -15672 -14324 -15608
rect -14260 -15672 -14244 -15608
rect -14340 -15688 -14244 -15672
rect -14340 -15752 -14324 -15688
rect -14260 -15752 -14244 -15688
rect -14340 -15768 -14244 -15752
rect -14340 -15832 -14324 -15768
rect -14260 -15832 -14244 -15768
rect -14340 -15848 -14244 -15832
rect -14340 -15912 -14324 -15848
rect -14260 -15912 -14244 -15848
rect -14340 -15928 -14244 -15912
rect -14340 -15992 -14324 -15928
rect -14260 -15992 -14244 -15928
rect -14340 -16008 -14244 -15992
rect -15752 -16108 -15656 -16072
rect -14340 -16072 -14324 -16008
rect -14260 -16072 -14244 -16008
rect -13921 -15328 -13199 -15319
rect -13921 -16032 -13912 -15328
rect -13208 -16032 -13199 -15328
rect -13921 -16041 -13199 -16032
rect -12928 -15352 -12912 -15288
rect -12848 -15352 -12832 -15288
rect -11516 -15288 -11420 -15252
rect -12928 -15368 -12832 -15352
rect -12928 -15432 -12912 -15368
rect -12848 -15432 -12832 -15368
rect -12928 -15448 -12832 -15432
rect -12928 -15512 -12912 -15448
rect -12848 -15512 -12832 -15448
rect -12928 -15528 -12832 -15512
rect -12928 -15592 -12912 -15528
rect -12848 -15592 -12832 -15528
rect -12928 -15608 -12832 -15592
rect -12928 -15672 -12912 -15608
rect -12848 -15672 -12832 -15608
rect -12928 -15688 -12832 -15672
rect -12928 -15752 -12912 -15688
rect -12848 -15752 -12832 -15688
rect -12928 -15768 -12832 -15752
rect -12928 -15832 -12912 -15768
rect -12848 -15832 -12832 -15768
rect -12928 -15848 -12832 -15832
rect -12928 -15912 -12912 -15848
rect -12848 -15912 -12832 -15848
rect -12928 -15928 -12832 -15912
rect -12928 -15992 -12912 -15928
rect -12848 -15992 -12832 -15928
rect -12928 -16008 -12832 -15992
rect -14340 -16108 -14244 -16072
rect -12928 -16072 -12912 -16008
rect -12848 -16072 -12832 -16008
rect -12509 -15328 -11787 -15319
rect -12509 -16032 -12500 -15328
rect -11796 -16032 -11787 -15328
rect -12509 -16041 -11787 -16032
rect -11516 -15352 -11500 -15288
rect -11436 -15352 -11420 -15288
rect -10104 -15288 -10008 -15252
rect -11516 -15368 -11420 -15352
rect -11516 -15432 -11500 -15368
rect -11436 -15432 -11420 -15368
rect -11516 -15448 -11420 -15432
rect -11516 -15512 -11500 -15448
rect -11436 -15512 -11420 -15448
rect -11516 -15528 -11420 -15512
rect -11516 -15592 -11500 -15528
rect -11436 -15592 -11420 -15528
rect -11516 -15608 -11420 -15592
rect -11516 -15672 -11500 -15608
rect -11436 -15672 -11420 -15608
rect -11516 -15688 -11420 -15672
rect -11516 -15752 -11500 -15688
rect -11436 -15752 -11420 -15688
rect -11516 -15768 -11420 -15752
rect -11516 -15832 -11500 -15768
rect -11436 -15832 -11420 -15768
rect -11516 -15848 -11420 -15832
rect -11516 -15912 -11500 -15848
rect -11436 -15912 -11420 -15848
rect -11516 -15928 -11420 -15912
rect -11516 -15992 -11500 -15928
rect -11436 -15992 -11420 -15928
rect -11516 -16008 -11420 -15992
rect -12928 -16108 -12832 -16072
rect -11516 -16072 -11500 -16008
rect -11436 -16072 -11420 -16008
rect -11097 -15328 -10375 -15319
rect -11097 -16032 -11088 -15328
rect -10384 -16032 -10375 -15328
rect -11097 -16041 -10375 -16032
rect -10104 -15352 -10088 -15288
rect -10024 -15352 -10008 -15288
rect -8692 -15288 -8596 -15252
rect -10104 -15368 -10008 -15352
rect -10104 -15432 -10088 -15368
rect -10024 -15432 -10008 -15368
rect -10104 -15448 -10008 -15432
rect -10104 -15512 -10088 -15448
rect -10024 -15512 -10008 -15448
rect -10104 -15528 -10008 -15512
rect -10104 -15592 -10088 -15528
rect -10024 -15592 -10008 -15528
rect -10104 -15608 -10008 -15592
rect -10104 -15672 -10088 -15608
rect -10024 -15672 -10008 -15608
rect -10104 -15688 -10008 -15672
rect -10104 -15752 -10088 -15688
rect -10024 -15752 -10008 -15688
rect -10104 -15768 -10008 -15752
rect -10104 -15832 -10088 -15768
rect -10024 -15832 -10008 -15768
rect -10104 -15848 -10008 -15832
rect -10104 -15912 -10088 -15848
rect -10024 -15912 -10008 -15848
rect -10104 -15928 -10008 -15912
rect -10104 -15992 -10088 -15928
rect -10024 -15992 -10008 -15928
rect -10104 -16008 -10008 -15992
rect -11516 -16108 -11420 -16072
rect -10104 -16072 -10088 -16008
rect -10024 -16072 -10008 -16008
rect -9685 -15328 -8963 -15319
rect -9685 -16032 -9676 -15328
rect -8972 -16032 -8963 -15328
rect -9685 -16041 -8963 -16032
rect -8692 -15352 -8676 -15288
rect -8612 -15352 -8596 -15288
rect -7280 -15288 -7184 -15252
rect -8692 -15368 -8596 -15352
rect -8692 -15432 -8676 -15368
rect -8612 -15432 -8596 -15368
rect -8692 -15448 -8596 -15432
rect -8692 -15512 -8676 -15448
rect -8612 -15512 -8596 -15448
rect -8692 -15528 -8596 -15512
rect -8692 -15592 -8676 -15528
rect -8612 -15592 -8596 -15528
rect -8692 -15608 -8596 -15592
rect -8692 -15672 -8676 -15608
rect -8612 -15672 -8596 -15608
rect -8692 -15688 -8596 -15672
rect -8692 -15752 -8676 -15688
rect -8612 -15752 -8596 -15688
rect -8692 -15768 -8596 -15752
rect -8692 -15832 -8676 -15768
rect -8612 -15832 -8596 -15768
rect -8692 -15848 -8596 -15832
rect -8692 -15912 -8676 -15848
rect -8612 -15912 -8596 -15848
rect -8692 -15928 -8596 -15912
rect -8692 -15992 -8676 -15928
rect -8612 -15992 -8596 -15928
rect -8692 -16008 -8596 -15992
rect -10104 -16108 -10008 -16072
rect -8692 -16072 -8676 -16008
rect -8612 -16072 -8596 -16008
rect -8273 -15328 -7551 -15319
rect -8273 -16032 -8264 -15328
rect -7560 -16032 -7551 -15328
rect -8273 -16041 -7551 -16032
rect -7280 -15352 -7264 -15288
rect -7200 -15352 -7184 -15288
rect -5868 -15288 -5772 -15252
rect -7280 -15368 -7184 -15352
rect -7280 -15432 -7264 -15368
rect -7200 -15432 -7184 -15368
rect -7280 -15448 -7184 -15432
rect -7280 -15512 -7264 -15448
rect -7200 -15512 -7184 -15448
rect -7280 -15528 -7184 -15512
rect -7280 -15592 -7264 -15528
rect -7200 -15592 -7184 -15528
rect -7280 -15608 -7184 -15592
rect -7280 -15672 -7264 -15608
rect -7200 -15672 -7184 -15608
rect -7280 -15688 -7184 -15672
rect -7280 -15752 -7264 -15688
rect -7200 -15752 -7184 -15688
rect -7280 -15768 -7184 -15752
rect -7280 -15832 -7264 -15768
rect -7200 -15832 -7184 -15768
rect -7280 -15848 -7184 -15832
rect -7280 -15912 -7264 -15848
rect -7200 -15912 -7184 -15848
rect -7280 -15928 -7184 -15912
rect -7280 -15992 -7264 -15928
rect -7200 -15992 -7184 -15928
rect -7280 -16008 -7184 -15992
rect -8692 -16108 -8596 -16072
rect -7280 -16072 -7264 -16008
rect -7200 -16072 -7184 -16008
rect -6861 -15328 -6139 -15319
rect -6861 -16032 -6852 -15328
rect -6148 -16032 -6139 -15328
rect -6861 -16041 -6139 -16032
rect -5868 -15352 -5852 -15288
rect -5788 -15352 -5772 -15288
rect -4456 -15288 -4360 -15252
rect -5868 -15368 -5772 -15352
rect -5868 -15432 -5852 -15368
rect -5788 -15432 -5772 -15368
rect -5868 -15448 -5772 -15432
rect -5868 -15512 -5852 -15448
rect -5788 -15512 -5772 -15448
rect -5868 -15528 -5772 -15512
rect -5868 -15592 -5852 -15528
rect -5788 -15592 -5772 -15528
rect -5868 -15608 -5772 -15592
rect -5868 -15672 -5852 -15608
rect -5788 -15672 -5772 -15608
rect -5868 -15688 -5772 -15672
rect -5868 -15752 -5852 -15688
rect -5788 -15752 -5772 -15688
rect -5868 -15768 -5772 -15752
rect -5868 -15832 -5852 -15768
rect -5788 -15832 -5772 -15768
rect -5868 -15848 -5772 -15832
rect -5868 -15912 -5852 -15848
rect -5788 -15912 -5772 -15848
rect -5868 -15928 -5772 -15912
rect -5868 -15992 -5852 -15928
rect -5788 -15992 -5772 -15928
rect -5868 -16008 -5772 -15992
rect -7280 -16108 -7184 -16072
rect -5868 -16072 -5852 -16008
rect -5788 -16072 -5772 -16008
rect -5449 -15328 -4727 -15319
rect -5449 -16032 -5440 -15328
rect -4736 -16032 -4727 -15328
rect -5449 -16041 -4727 -16032
rect -4456 -15352 -4440 -15288
rect -4376 -15352 -4360 -15288
rect -3044 -15288 -2948 -15252
rect -4456 -15368 -4360 -15352
rect -4456 -15432 -4440 -15368
rect -4376 -15432 -4360 -15368
rect -4456 -15448 -4360 -15432
rect -4456 -15512 -4440 -15448
rect -4376 -15512 -4360 -15448
rect -4456 -15528 -4360 -15512
rect -4456 -15592 -4440 -15528
rect -4376 -15592 -4360 -15528
rect -4456 -15608 -4360 -15592
rect -4456 -15672 -4440 -15608
rect -4376 -15672 -4360 -15608
rect -4456 -15688 -4360 -15672
rect -4456 -15752 -4440 -15688
rect -4376 -15752 -4360 -15688
rect -4456 -15768 -4360 -15752
rect -4456 -15832 -4440 -15768
rect -4376 -15832 -4360 -15768
rect -4456 -15848 -4360 -15832
rect -4456 -15912 -4440 -15848
rect -4376 -15912 -4360 -15848
rect -4456 -15928 -4360 -15912
rect -4456 -15992 -4440 -15928
rect -4376 -15992 -4360 -15928
rect -4456 -16008 -4360 -15992
rect -5868 -16108 -5772 -16072
rect -4456 -16072 -4440 -16008
rect -4376 -16072 -4360 -16008
rect -4037 -15328 -3315 -15319
rect -4037 -16032 -4028 -15328
rect -3324 -16032 -3315 -15328
rect -4037 -16041 -3315 -16032
rect -3044 -15352 -3028 -15288
rect -2964 -15352 -2948 -15288
rect -1632 -15288 -1536 -15252
rect -3044 -15368 -2948 -15352
rect -3044 -15432 -3028 -15368
rect -2964 -15432 -2948 -15368
rect -3044 -15448 -2948 -15432
rect -3044 -15512 -3028 -15448
rect -2964 -15512 -2948 -15448
rect -3044 -15528 -2948 -15512
rect -3044 -15592 -3028 -15528
rect -2964 -15592 -2948 -15528
rect -3044 -15608 -2948 -15592
rect -3044 -15672 -3028 -15608
rect -2964 -15672 -2948 -15608
rect -3044 -15688 -2948 -15672
rect -3044 -15752 -3028 -15688
rect -2964 -15752 -2948 -15688
rect -3044 -15768 -2948 -15752
rect -3044 -15832 -3028 -15768
rect -2964 -15832 -2948 -15768
rect -3044 -15848 -2948 -15832
rect -3044 -15912 -3028 -15848
rect -2964 -15912 -2948 -15848
rect -3044 -15928 -2948 -15912
rect -3044 -15992 -3028 -15928
rect -2964 -15992 -2948 -15928
rect -3044 -16008 -2948 -15992
rect -4456 -16108 -4360 -16072
rect -3044 -16072 -3028 -16008
rect -2964 -16072 -2948 -16008
rect -2625 -15328 -1903 -15319
rect -2625 -16032 -2616 -15328
rect -1912 -16032 -1903 -15328
rect -2625 -16041 -1903 -16032
rect -1632 -15352 -1616 -15288
rect -1552 -15352 -1536 -15288
rect -220 -15288 -124 -15252
rect -1632 -15368 -1536 -15352
rect -1632 -15432 -1616 -15368
rect -1552 -15432 -1536 -15368
rect -1632 -15448 -1536 -15432
rect -1632 -15512 -1616 -15448
rect -1552 -15512 -1536 -15448
rect -1632 -15528 -1536 -15512
rect -1632 -15592 -1616 -15528
rect -1552 -15592 -1536 -15528
rect -1632 -15608 -1536 -15592
rect -1632 -15672 -1616 -15608
rect -1552 -15672 -1536 -15608
rect -1632 -15688 -1536 -15672
rect -1632 -15752 -1616 -15688
rect -1552 -15752 -1536 -15688
rect -1632 -15768 -1536 -15752
rect -1632 -15832 -1616 -15768
rect -1552 -15832 -1536 -15768
rect -1632 -15848 -1536 -15832
rect -1632 -15912 -1616 -15848
rect -1552 -15912 -1536 -15848
rect -1632 -15928 -1536 -15912
rect -1632 -15992 -1616 -15928
rect -1552 -15992 -1536 -15928
rect -1632 -16008 -1536 -15992
rect -3044 -16108 -2948 -16072
rect -1632 -16072 -1616 -16008
rect -1552 -16072 -1536 -16008
rect -1213 -15328 -491 -15319
rect -1213 -16032 -1204 -15328
rect -500 -16032 -491 -15328
rect -1213 -16041 -491 -16032
rect -220 -15352 -204 -15288
rect -140 -15352 -124 -15288
rect 1192 -15288 1288 -15252
rect -220 -15368 -124 -15352
rect -220 -15432 -204 -15368
rect -140 -15432 -124 -15368
rect -220 -15448 -124 -15432
rect -220 -15512 -204 -15448
rect -140 -15512 -124 -15448
rect -220 -15528 -124 -15512
rect -220 -15592 -204 -15528
rect -140 -15592 -124 -15528
rect -220 -15608 -124 -15592
rect -220 -15672 -204 -15608
rect -140 -15672 -124 -15608
rect -220 -15688 -124 -15672
rect -220 -15752 -204 -15688
rect -140 -15752 -124 -15688
rect -220 -15768 -124 -15752
rect -220 -15832 -204 -15768
rect -140 -15832 -124 -15768
rect -220 -15848 -124 -15832
rect -220 -15912 -204 -15848
rect -140 -15912 -124 -15848
rect -220 -15928 -124 -15912
rect -220 -15992 -204 -15928
rect -140 -15992 -124 -15928
rect -220 -16008 -124 -15992
rect -1632 -16108 -1536 -16072
rect -220 -16072 -204 -16008
rect -140 -16072 -124 -16008
rect 199 -15328 921 -15319
rect 199 -16032 208 -15328
rect 912 -16032 921 -15328
rect 199 -16041 921 -16032
rect 1192 -15352 1208 -15288
rect 1272 -15352 1288 -15288
rect 2604 -15288 2700 -15252
rect 1192 -15368 1288 -15352
rect 1192 -15432 1208 -15368
rect 1272 -15432 1288 -15368
rect 1192 -15448 1288 -15432
rect 1192 -15512 1208 -15448
rect 1272 -15512 1288 -15448
rect 1192 -15528 1288 -15512
rect 1192 -15592 1208 -15528
rect 1272 -15592 1288 -15528
rect 1192 -15608 1288 -15592
rect 1192 -15672 1208 -15608
rect 1272 -15672 1288 -15608
rect 1192 -15688 1288 -15672
rect 1192 -15752 1208 -15688
rect 1272 -15752 1288 -15688
rect 1192 -15768 1288 -15752
rect 1192 -15832 1208 -15768
rect 1272 -15832 1288 -15768
rect 1192 -15848 1288 -15832
rect 1192 -15912 1208 -15848
rect 1272 -15912 1288 -15848
rect 1192 -15928 1288 -15912
rect 1192 -15992 1208 -15928
rect 1272 -15992 1288 -15928
rect 1192 -16008 1288 -15992
rect -220 -16108 -124 -16072
rect 1192 -16072 1208 -16008
rect 1272 -16072 1288 -16008
rect 1611 -15328 2333 -15319
rect 1611 -16032 1620 -15328
rect 2324 -16032 2333 -15328
rect 1611 -16041 2333 -16032
rect 2604 -15352 2620 -15288
rect 2684 -15352 2700 -15288
rect 4016 -15288 4112 -15252
rect 2604 -15368 2700 -15352
rect 2604 -15432 2620 -15368
rect 2684 -15432 2700 -15368
rect 2604 -15448 2700 -15432
rect 2604 -15512 2620 -15448
rect 2684 -15512 2700 -15448
rect 2604 -15528 2700 -15512
rect 2604 -15592 2620 -15528
rect 2684 -15592 2700 -15528
rect 2604 -15608 2700 -15592
rect 2604 -15672 2620 -15608
rect 2684 -15672 2700 -15608
rect 2604 -15688 2700 -15672
rect 2604 -15752 2620 -15688
rect 2684 -15752 2700 -15688
rect 2604 -15768 2700 -15752
rect 2604 -15832 2620 -15768
rect 2684 -15832 2700 -15768
rect 2604 -15848 2700 -15832
rect 2604 -15912 2620 -15848
rect 2684 -15912 2700 -15848
rect 2604 -15928 2700 -15912
rect 2604 -15992 2620 -15928
rect 2684 -15992 2700 -15928
rect 2604 -16008 2700 -15992
rect 1192 -16108 1288 -16072
rect 2604 -16072 2620 -16008
rect 2684 -16072 2700 -16008
rect 3023 -15328 3745 -15319
rect 3023 -16032 3032 -15328
rect 3736 -16032 3745 -15328
rect 3023 -16041 3745 -16032
rect 4016 -15352 4032 -15288
rect 4096 -15352 4112 -15288
rect 5428 -15288 5524 -15252
rect 4016 -15368 4112 -15352
rect 4016 -15432 4032 -15368
rect 4096 -15432 4112 -15368
rect 4016 -15448 4112 -15432
rect 4016 -15512 4032 -15448
rect 4096 -15512 4112 -15448
rect 4016 -15528 4112 -15512
rect 4016 -15592 4032 -15528
rect 4096 -15592 4112 -15528
rect 4016 -15608 4112 -15592
rect 4016 -15672 4032 -15608
rect 4096 -15672 4112 -15608
rect 4016 -15688 4112 -15672
rect 4016 -15752 4032 -15688
rect 4096 -15752 4112 -15688
rect 4016 -15768 4112 -15752
rect 4016 -15832 4032 -15768
rect 4096 -15832 4112 -15768
rect 4016 -15848 4112 -15832
rect 4016 -15912 4032 -15848
rect 4096 -15912 4112 -15848
rect 4016 -15928 4112 -15912
rect 4016 -15992 4032 -15928
rect 4096 -15992 4112 -15928
rect 4016 -16008 4112 -15992
rect 2604 -16108 2700 -16072
rect 4016 -16072 4032 -16008
rect 4096 -16072 4112 -16008
rect 4435 -15328 5157 -15319
rect 4435 -16032 4444 -15328
rect 5148 -16032 5157 -15328
rect 4435 -16041 5157 -16032
rect 5428 -15352 5444 -15288
rect 5508 -15352 5524 -15288
rect 6840 -15288 6936 -15252
rect 5428 -15368 5524 -15352
rect 5428 -15432 5444 -15368
rect 5508 -15432 5524 -15368
rect 5428 -15448 5524 -15432
rect 5428 -15512 5444 -15448
rect 5508 -15512 5524 -15448
rect 5428 -15528 5524 -15512
rect 5428 -15592 5444 -15528
rect 5508 -15592 5524 -15528
rect 5428 -15608 5524 -15592
rect 5428 -15672 5444 -15608
rect 5508 -15672 5524 -15608
rect 5428 -15688 5524 -15672
rect 5428 -15752 5444 -15688
rect 5508 -15752 5524 -15688
rect 5428 -15768 5524 -15752
rect 5428 -15832 5444 -15768
rect 5508 -15832 5524 -15768
rect 5428 -15848 5524 -15832
rect 5428 -15912 5444 -15848
rect 5508 -15912 5524 -15848
rect 5428 -15928 5524 -15912
rect 5428 -15992 5444 -15928
rect 5508 -15992 5524 -15928
rect 5428 -16008 5524 -15992
rect 4016 -16108 4112 -16072
rect 5428 -16072 5444 -16008
rect 5508 -16072 5524 -16008
rect 5847 -15328 6569 -15319
rect 5847 -16032 5856 -15328
rect 6560 -16032 6569 -15328
rect 5847 -16041 6569 -16032
rect 6840 -15352 6856 -15288
rect 6920 -15352 6936 -15288
rect 8252 -15288 8348 -15252
rect 6840 -15368 6936 -15352
rect 6840 -15432 6856 -15368
rect 6920 -15432 6936 -15368
rect 6840 -15448 6936 -15432
rect 6840 -15512 6856 -15448
rect 6920 -15512 6936 -15448
rect 6840 -15528 6936 -15512
rect 6840 -15592 6856 -15528
rect 6920 -15592 6936 -15528
rect 6840 -15608 6936 -15592
rect 6840 -15672 6856 -15608
rect 6920 -15672 6936 -15608
rect 6840 -15688 6936 -15672
rect 6840 -15752 6856 -15688
rect 6920 -15752 6936 -15688
rect 6840 -15768 6936 -15752
rect 6840 -15832 6856 -15768
rect 6920 -15832 6936 -15768
rect 6840 -15848 6936 -15832
rect 6840 -15912 6856 -15848
rect 6920 -15912 6936 -15848
rect 6840 -15928 6936 -15912
rect 6840 -15992 6856 -15928
rect 6920 -15992 6936 -15928
rect 6840 -16008 6936 -15992
rect 5428 -16108 5524 -16072
rect 6840 -16072 6856 -16008
rect 6920 -16072 6936 -16008
rect 7259 -15328 7981 -15319
rect 7259 -16032 7268 -15328
rect 7972 -16032 7981 -15328
rect 7259 -16041 7981 -16032
rect 8252 -15352 8268 -15288
rect 8332 -15352 8348 -15288
rect 9664 -15288 9760 -15252
rect 8252 -15368 8348 -15352
rect 8252 -15432 8268 -15368
rect 8332 -15432 8348 -15368
rect 8252 -15448 8348 -15432
rect 8252 -15512 8268 -15448
rect 8332 -15512 8348 -15448
rect 8252 -15528 8348 -15512
rect 8252 -15592 8268 -15528
rect 8332 -15592 8348 -15528
rect 8252 -15608 8348 -15592
rect 8252 -15672 8268 -15608
rect 8332 -15672 8348 -15608
rect 8252 -15688 8348 -15672
rect 8252 -15752 8268 -15688
rect 8332 -15752 8348 -15688
rect 8252 -15768 8348 -15752
rect 8252 -15832 8268 -15768
rect 8332 -15832 8348 -15768
rect 8252 -15848 8348 -15832
rect 8252 -15912 8268 -15848
rect 8332 -15912 8348 -15848
rect 8252 -15928 8348 -15912
rect 8252 -15992 8268 -15928
rect 8332 -15992 8348 -15928
rect 8252 -16008 8348 -15992
rect 6840 -16108 6936 -16072
rect 8252 -16072 8268 -16008
rect 8332 -16072 8348 -16008
rect 8671 -15328 9393 -15319
rect 8671 -16032 8680 -15328
rect 9384 -16032 9393 -15328
rect 8671 -16041 9393 -16032
rect 9664 -15352 9680 -15288
rect 9744 -15352 9760 -15288
rect 11076 -15288 11172 -15252
rect 9664 -15368 9760 -15352
rect 9664 -15432 9680 -15368
rect 9744 -15432 9760 -15368
rect 9664 -15448 9760 -15432
rect 9664 -15512 9680 -15448
rect 9744 -15512 9760 -15448
rect 9664 -15528 9760 -15512
rect 9664 -15592 9680 -15528
rect 9744 -15592 9760 -15528
rect 9664 -15608 9760 -15592
rect 9664 -15672 9680 -15608
rect 9744 -15672 9760 -15608
rect 9664 -15688 9760 -15672
rect 9664 -15752 9680 -15688
rect 9744 -15752 9760 -15688
rect 9664 -15768 9760 -15752
rect 9664 -15832 9680 -15768
rect 9744 -15832 9760 -15768
rect 9664 -15848 9760 -15832
rect 9664 -15912 9680 -15848
rect 9744 -15912 9760 -15848
rect 9664 -15928 9760 -15912
rect 9664 -15992 9680 -15928
rect 9744 -15992 9760 -15928
rect 9664 -16008 9760 -15992
rect 8252 -16108 8348 -16072
rect 9664 -16072 9680 -16008
rect 9744 -16072 9760 -16008
rect 10083 -15328 10805 -15319
rect 10083 -16032 10092 -15328
rect 10796 -16032 10805 -15328
rect 10083 -16041 10805 -16032
rect 11076 -15352 11092 -15288
rect 11156 -15352 11172 -15288
rect 12488 -15288 12584 -15252
rect 11076 -15368 11172 -15352
rect 11076 -15432 11092 -15368
rect 11156 -15432 11172 -15368
rect 11076 -15448 11172 -15432
rect 11076 -15512 11092 -15448
rect 11156 -15512 11172 -15448
rect 11076 -15528 11172 -15512
rect 11076 -15592 11092 -15528
rect 11156 -15592 11172 -15528
rect 11076 -15608 11172 -15592
rect 11076 -15672 11092 -15608
rect 11156 -15672 11172 -15608
rect 11076 -15688 11172 -15672
rect 11076 -15752 11092 -15688
rect 11156 -15752 11172 -15688
rect 11076 -15768 11172 -15752
rect 11076 -15832 11092 -15768
rect 11156 -15832 11172 -15768
rect 11076 -15848 11172 -15832
rect 11076 -15912 11092 -15848
rect 11156 -15912 11172 -15848
rect 11076 -15928 11172 -15912
rect 11076 -15992 11092 -15928
rect 11156 -15992 11172 -15928
rect 11076 -16008 11172 -15992
rect 9664 -16108 9760 -16072
rect 11076 -16072 11092 -16008
rect 11156 -16072 11172 -16008
rect 11495 -15328 12217 -15319
rect 11495 -16032 11504 -15328
rect 12208 -16032 12217 -15328
rect 11495 -16041 12217 -16032
rect 12488 -15352 12504 -15288
rect 12568 -15352 12584 -15288
rect 13900 -15288 13996 -15252
rect 12488 -15368 12584 -15352
rect 12488 -15432 12504 -15368
rect 12568 -15432 12584 -15368
rect 12488 -15448 12584 -15432
rect 12488 -15512 12504 -15448
rect 12568 -15512 12584 -15448
rect 12488 -15528 12584 -15512
rect 12488 -15592 12504 -15528
rect 12568 -15592 12584 -15528
rect 12488 -15608 12584 -15592
rect 12488 -15672 12504 -15608
rect 12568 -15672 12584 -15608
rect 12488 -15688 12584 -15672
rect 12488 -15752 12504 -15688
rect 12568 -15752 12584 -15688
rect 12488 -15768 12584 -15752
rect 12488 -15832 12504 -15768
rect 12568 -15832 12584 -15768
rect 12488 -15848 12584 -15832
rect 12488 -15912 12504 -15848
rect 12568 -15912 12584 -15848
rect 12488 -15928 12584 -15912
rect 12488 -15992 12504 -15928
rect 12568 -15992 12584 -15928
rect 12488 -16008 12584 -15992
rect 11076 -16108 11172 -16072
rect 12488 -16072 12504 -16008
rect 12568 -16072 12584 -16008
rect 12907 -15328 13629 -15319
rect 12907 -16032 12916 -15328
rect 13620 -16032 13629 -15328
rect 12907 -16041 13629 -16032
rect 13900 -15352 13916 -15288
rect 13980 -15352 13996 -15288
rect 15312 -15288 15408 -15252
rect 13900 -15368 13996 -15352
rect 13900 -15432 13916 -15368
rect 13980 -15432 13996 -15368
rect 13900 -15448 13996 -15432
rect 13900 -15512 13916 -15448
rect 13980 -15512 13996 -15448
rect 13900 -15528 13996 -15512
rect 13900 -15592 13916 -15528
rect 13980 -15592 13996 -15528
rect 13900 -15608 13996 -15592
rect 13900 -15672 13916 -15608
rect 13980 -15672 13996 -15608
rect 13900 -15688 13996 -15672
rect 13900 -15752 13916 -15688
rect 13980 -15752 13996 -15688
rect 13900 -15768 13996 -15752
rect 13900 -15832 13916 -15768
rect 13980 -15832 13996 -15768
rect 13900 -15848 13996 -15832
rect 13900 -15912 13916 -15848
rect 13980 -15912 13996 -15848
rect 13900 -15928 13996 -15912
rect 13900 -15992 13916 -15928
rect 13980 -15992 13996 -15928
rect 13900 -16008 13996 -15992
rect 12488 -16108 12584 -16072
rect 13900 -16072 13916 -16008
rect 13980 -16072 13996 -16008
rect 14319 -15328 15041 -15319
rect 14319 -16032 14328 -15328
rect 15032 -16032 15041 -15328
rect 14319 -16041 15041 -16032
rect 15312 -15352 15328 -15288
rect 15392 -15352 15408 -15288
rect 16724 -15288 16820 -15252
rect 15312 -15368 15408 -15352
rect 15312 -15432 15328 -15368
rect 15392 -15432 15408 -15368
rect 15312 -15448 15408 -15432
rect 15312 -15512 15328 -15448
rect 15392 -15512 15408 -15448
rect 15312 -15528 15408 -15512
rect 15312 -15592 15328 -15528
rect 15392 -15592 15408 -15528
rect 15312 -15608 15408 -15592
rect 15312 -15672 15328 -15608
rect 15392 -15672 15408 -15608
rect 15312 -15688 15408 -15672
rect 15312 -15752 15328 -15688
rect 15392 -15752 15408 -15688
rect 15312 -15768 15408 -15752
rect 15312 -15832 15328 -15768
rect 15392 -15832 15408 -15768
rect 15312 -15848 15408 -15832
rect 15312 -15912 15328 -15848
rect 15392 -15912 15408 -15848
rect 15312 -15928 15408 -15912
rect 15312 -15992 15328 -15928
rect 15392 -15992 15408 -15928
rect 15312 -16008 15408 -15992
rect 13900 -16108 13996 -16072
rect 15312 -16072 15328 -16008
rect 15392 -16072 15408 -16008
rect 15731 -15328 16453 -15319
rect 15731 -16032 15740 -15328
rect 16444 -16032 16453 -15328
rect 15731 -16041 16453 -16032
rect 16724 -15352 16740 -15288
rect 16804 -15352 16820 -15288
rect 18136 -15288 18232 -15252
rect 16724 -15368 16820 -15352
rect 16724 -15432 16740 -15368
rect 16804 -15432 16820 -15368
rect 16724 -15448 16820 -15432
rect 16724 -15512 16740 -15448
rect 16804 -15512 16820 -15448
rect 16724 -15528 16820 -15512
rect 16724 -15592 16740 -15528
rect 16804 -15592 16820 -15528
rect 16724 -15608 16820 -15592
rect 16724 -15672 16740 -15608
rect 16804 -15672 16820 -15608
rect 16724 -15688 16820 -15672
rect 16724 -15752 16740 -15688
rect 16804 -15752 16820 -15688
rect 16724 -15768 16820 -15752
rect 16724 -15832 16740 -15768
rect 16804 -15832 16820 -15768
rect 16724 -15848 16820 -15832
rect 16724 -15912 16740 -15848
rect 16804 -15912 16820 -15848
rect 16724 -15928 16820 -15912
rect 16724 -15992 16740 -15928
rect 16804 -15992 16820 -15928
rect 16724 -16008 16820 -15992
rect 15312 -16108 15408 -16072
rect 16724 -16072 16740 -16008
rect 16804 -16072 16820 -16008
rect 17143 -15328 17865 -15319
rect 17143 -16032 17152 -15328
rect 17856 -16032 17865 -15328
rect 17143 -16041 17865 -16032
rect 18136 -15352 18152 -15288
rect 18216 -15352 18232 -15288
rect 19548 -15288 19644 -15252
rect 18136 -15368 18232 -15352
rect 18136 -15432 18152 -15368
rect 18216 -15432 18232 -15368
rect 18136 -15448 18232 -15432
rect 18136 -15512 18152 -15448
rect 18216 -15512 18232 -15448
rect 18136 -15528 18232 -15512
rect 18136 -15592 18152 -15528
rect 18216 -15592 18232 -15528
rect 18136 -15608 18232 -15592
rect 18136 -15672 18152 -15608
rect 18216 -15672 18232 -15608
rect 18136 -15688 18232 -15672
rect 18136 -15752 18152 -15688
rect 18216 -15752 18232 -15688
rect 18136 -15768 18232 -15752
rect 18136 -15832 18152 -15768
rect 18216 -15832 18232 -15768
rect 18136 -15848 18232 -15832
rect 18136 -15912 18152 -15848
rect 18216 -15912 18232 -15848
rect 18136 -15928 18232 -15912
rect 18136 -15992 18152 -15928
rect 18216 -15992 18232 -15928
rect 18136 -16008 18232 -15992
rect 16724 -16108 16820 -16072
rect 18136 -16072 18152 -16008
rect 18216 -16072 18232 -16008
rect 18555 -15328 19277 -15319
rect 18555 -16032 18564 -15328
rect 19268 -16032 19277 -15328
rect 18555 -16041 19277 -16032
rect 19548 -15352 19564 -15288
rect 19628 -15352 19644 -15288
rect 20960 -15288 21056 -15252
rect 19548 -15368 19644 -15352
rect 19548 -15432 19564 -15368
rect 19628 -15432 19644 -15368
rect 19548 -15448 19644 -15432
rect 19548 -15512 19564 -15448
rect 19628 -15512 19644 -15448
rect 19548 -15528 19644 -15512
rect 19548 -15592 19564 -15528
rect 19628 -15592 19644 -15528
rect 19548 -15608 19644 -15592
rect 19548 -15672 19564 -15608
rect 19628 -15672 19644 -15608
rect 19548 -15688 19644 -15672
rect 19548 -15752 19564 -15688
rect 19628 -15752 19644 -15688
rect 19548 -15768 19644 -15752
rect 19548 -15832 19564 -15768
rect 19628 -15832 19644 -15768
rect 19548 -15848 19644 -15832
rect 19548 -15912 19564 -15848
rect 19628 -15912 19644 -15848
rect 19548 -15928 19644 -15912
rect 19548 -15992 19564 -15928
rect 19628 -15992 19644 -15928
rect 19548 -16008 19644 -15992
rect 18136 -16108 18232 -16072
rect 19548 -16072 19564 -16008
rect 19628 -16072 19644 -16008
rect 19967 -15328 20689 -15319
rect 19967 -16032 19976 -15328
rect 20680 -16032 20689 -15328
rect 19967 -16041 20689 -16032
rect 20960 -15352 20976 -15288
rect 21040 -15352 21056 -15288
rect 22372 -15288 22468 -15252
rect 20960 -15368 21056 -15352
rect 20960 -15432 20976 -15368
rect 21040 -15432 21056 -15368
rect 20960 -15448 21056 -15432
rect 20960 -15512 20976 -15448
rect 21040 -15512 21056 -15448
rect 20960 -15528 21056 -15512
rect 20960 -15592 20976 -15528
rect 21040 -15592 21056 -15528
rect 20960 -15608 21056 -15592
rect 20960 -15672 20976 -15608
rect 21040 -15672 21056 -15608
rect 20960 -15688 21056 -15672
rect 20960 -15752 20976 -15688
rect 21040 -15752 21056 -15688
rect 20960 -15768 21056 -15752
rect 20960 -15832 20976 -15768
rect 21040 -15832 21056 -15768
rect 20960 -15848 21056 -15832
rect 20960 -15912 20976 -15848
rect 21040 -15912 21056 -15848
rect 20960 -15928 21056 -15912
rect 20960 -15992 20976 -15928
rect 21040 -15992 21056 -15928
rect 20960 -16008 21056 -15992
rect 19548 -16108 19644 -16072
rect 20960 -16072 20976 -16008
rect 21040 -16072 21056 -16008
rect 21379 -15328 22101 -15319
rect 21379 -16032 21388 -15328
rect 22092 -16032 22101 -15328
rect 21379 -16041 22101 -16032
rect 22372 -15352 22388 -15288
rect 22452 -15352 22468 -15288
rect 23784 -15288 23880 -15252
rect 22372 -15368 22468 -15352
rect 22372 -15432 22388 -15368
rect 22452 -15432 22468 -15368
rect 22372 -15448 22468 -15432
rect 22372 -15512 22388 -15448
rect 22452 -15512 22468 -15448
rect 22372 -15528 22468 -15512
rect 22372 -15592 22388 -15528
rect 22452 -15592 22468 -15528
rect 22372 -15608 22468 -15592
rect 22372 -15672 22388 -15608
rect 22452 -15672 22468 -15608
rect 22372 -15688 22468 -15672
rect 22372 -15752 22388 -15688
rect 22452 -15752 22468 -15688
rect 22372 -15768 22468 -15752
rect 22372 -15832 22388 -15768
rect 22452 -15832 22468 -15768
rect 22372 -15848 22468 -15832
rect 22372 -15912 22388 -15848
rect 22452 -15912 22468 -15848
rect 22372 -15928 22468 -15912
rect 22372 -15992 22388 -15928
rect 22452 -15992 22468 -15928
rect 22372 -16008 22468 -15992
rect 20960 -16108 21056 -16072
rect 22372 -16072 22388 -16008
rect 22452 -16072 22468 -16008
rect 22791 -15328 23513 -15319
rect 22791 -16032 22800 -15328
rect 23504 -16032 23513 -15328
rect 22791 -16041 23513 -16032
rect 23784 -15352 23800 -15288
rect 23864 -15352 23880 -15288
rect 23784 -15368 23880 -15352
rect 23784 -15432 23800 -15368
rect 23864 -15432 23880 -15368
rect 23784 -15448 23880 -15432
rect 23784 -15512 23800 -15448
rect 23864 -15512 23880 -15448
rect 23784 -15528 23880 -15512
rect 23784 -15592 23800 -15528
rect 23864 -15592 23880 -15528
rect 23784 -15608 23880 -15592
rect 23784 -15672 23800 -15608
rect 23864 -15672 23880 -15608
rect 23784 -15688 23880 -15672
rect 23784 -15752 23800 -15688
rect 23864 -15752 23880 -15688
rect 23784 -15768 23880 -15752
rect 23784 -15832 23800 -15768
rect 23864 -15832 23880 -15768
rect 23784 -15848 23880 -15832
rect 23784 -15912 23800 -15848
rect 23864 -15912 23880 -15848
rect 23784 -15928 23880 -15912
rect 23784 -15992 23800 -15928
rect 23864 -15992 23880 -15928
rect 23784 -16008 23880 -15992
rect 22372 -16108 22468 -16072
rect 23784 -16072 23800 -16008
rect 23864 -16072 23880 -16008
rect 23784 -16108 23880 -16072
rect -22812 -16408 -22716 -16372
rect -23805 -16448 -23083 -16439
rect -23805 -17152 -23796 -16448
rect -23092 -17152 -23083 -16448
rect -23805 -17161 -23083 -17152
rect -22812 -16472 -22796 -16408
rect -22732 -16472 -22716 -16408
rect -21400 -16408 -21304 -16372
rect -22812 -16488 -22716 -16472
rect -22812 -16552 -22796 -16488
rect -22732 -16552 -22716 -16488
rect -22812 -16568 -22716 -16552
rect -22812 -16632 -22796 -16568
rect -22732 -16632 -22716 -16568
rect -22812 -16648 -22716 -16632
rect -22812 -16712 -22796 -16648
rect -22732 -16712 -22716 -16648
rect -22812 -16728 -22716 -16712
rect -22812 -16792 -22796 -16728
rect -22732 -16792 -22716 -16728
rect -22812 -16808 -22716 -16792
rect -22812 -16872 -22796 -16808
rect -22732 -16872 -22716 -16808
rect -22812 -16888 -22716 -16872
rect -22812 -16952 -22796 -16888
rect -22732 -16952 -22716 -16888
rect -22812 -16968 -22716 -16952
rect -22812 -17032 -22796 -16968
rect -22732 -17032 -22716 -16968
rect -22812 -17048 -22716 -17032
rect -22812 -17112 -22796 -17048
rect -22732 -17112 -22716 -17048
rect -22812 -17128 -22716 -17112
rect -22812 -17192 -22796 -17128
rect -22732 -17192 -22716 -17128
rect -22393 -16448 -21671 -16439
rect -22393 -17152 -22384 -16448
rect -21680 -17152 -21671 -16448
rect -22393 -17161 -21671 -17152
rect -21400 -16472 -21384 -16408
rect -21320 -16472 -21304 -16408
rect -19988 -16408 -19892 -16372
rect -21400 -16488 -21304 -16472
rect -21400 -16552 -21384 -16488
rect -21320 -16552 -21304 -16488
rect -21400 -16568 -21304 -16552
rect -21400 -16632 -21384 -16568
rect -21320 -16632 -21304 -16568
rect -21400 -16648 -21304 -16632
rect -21400 -16712 -21384 -16648
rect -21320 -16712 -21304 -16648
rect -21400 -16728 -21304 -16712
rect -21400 -16792 -21384 -16728
rect -21320 -16792 -21304 -16728
rect -21400 -16808 -21304 -16792
rect -21400 -16872 -21384 -16808
rect -21320 -16872 -21304 -16808
rect -21400 -16888 -21304 -16872
rect -21400 -16952 -21384 -16888
rect -21320 -16952 -21304 -16888
rect -21400 -16968 -21304 -16952
rect -21400 -17032 -21384 -16968
rect -21320 -17032 -21304 -16968
rect -21400 -17048 -21304 -17032
rect -21400 -17112 -21384 -17048
rect -21320 -17112 -21304 -17048
rect -21400 -17128 -21304 -17112
rect -22812 -17228 -22716 -17192
rect -21400 -17192 -21384 -17128
rect -21320 -17192 -21304 -17128
rect -20981 -16448 -20259 -16439
rect -20981 -17152 -20972 -16448
rect -20268 -17152 -20259 -16448
rect -20981 -17161 -20259 -17152
rect -19988 -16472 -19972 -16408
rect -19908 -16472 -19892 -16408
rect -18576 -16408 -18480 -16372
rect -19988 -16488 -19892 -16472
rect -19988 -16552 -19972 -16488
rect -19908 -16552 -19892 -16488
rect -19988 -16568 -19892 -16552
rect -19988 -16632 -19972 -16568
rect -19908 -16632 -19892 -16568
rect -19988 -16648 -19892 -16632
rect -19988 -16712 -19972 -16648
rect -19908 -16712 -19892 -16648
rect -19988 -16728 -19892 -16712
rect -19988 -16792 -19972 -16728
rect -19908 -16792 -19892 -16728
rect -19988 -16808 -19892 -16792
rect -19988 -16872 -19972 -16808
rect -19908 -16872 -19892 -16808
rect -19988 -16888 -19892 -16872
rect -19988 -16952 -19972 -16888
rect -19908 -16952 -19892 -16888
rect -19988 -16968 -19892 -16952
rect -19988 -17032 -19972 -16968
rect -19908 -17032 -19892 -16968
rect -19988 -17048 -19892 -17032
rect -19988 -17112 -19972 -17048
rect -19908 -17112 -19892 -17048
rect -19988 -17128 -19892 -17112
rect -21400 -17228 -21304 -17192
rect -19988 -17192 -19972 -17128
rect -19908 -17192 -19892 -17128
rect -19569 -16448 -18847 -16439
rect -19569 -17152 -19560 -16448
rect -18856 -17152 -18847 -16448
rect -19569 -17161 -18847 -17152
rect -18576 -16472 -18560 -16408
rect -18496 -16472 -18480 -16408
rect -17164 -16408 -17068 -16372
rect -18576 -16488 -18480 -16472
rect -18576 -16552 -18560 -16488
rect -18496 -16552 -18480 -16488
rect -18576 -16568 -18480 -16552
rect -18576 -16632 -18560 -16568
rect -18496 -16632 -18480 -16568
rect -18576 -16648 -18480 -16632
rect -18576 -16712 -18560 -16648
rect -18496 -16712 -18480 -16648
rect -18576 -16728 -18480 -16712
rect -18576 -16792 -18560 -16728
rect -18496 -16792 -18480 -16728
rect -18576 -16808 -18480 -16792
rect -18576 -16872 -18560 -16808
rect -18496 -16872 -18480 -16808
rect -18576 -16888 -18480 -16872
rect -18576 -16952 -18560 -16888
rect -18496 -16952 -18480 -16888
rect -18576 -16968 -18480 -16952
rect -18576 -17032 -18560 -16968
rect -18496 -17032 -18480 -16968
rect -18576 -17048 -18480 -17032
rect -18576 -17112 -18560 -17048
rect -18496 -17112 -18480 -17048
rect -18576 -17128 -18480 -17112
rect -19988 -17228 -19892 -17192
rect -18576 -17192 -18560 -17128
rect -18496 -17192 -18480 -17128
rect -18157 -16448 -17435 -16439
rect -18157 -17152 -18148 -16448
rect -17444 -17152 -17435 -16448
rect -18157 -17161 -17435 -17152
rect -17164 -16472 -17148 -16408
rect -17084 -16472 -17068 -16408
rect -15752 -16408 -15656 -16372
rect -17164 -16488 -17068 -16472
rect -17164 -16552 -17148 -16488
rect -17084 -16552 -17068 -16488
rect -17164 -16568 -17068 -16552
rect -17164 -16632 -17148 -16568
rect -17084 -16632 -17068 -16568
rect -17164 -16648 -17068 -16632
rect -17164 -16712 -17148 -16648
rect -17084 -16712 -17068 -16648
rect -17164 -16728 -17068 -16712
rect -17164 -16792 -17148 -16728
rect -17084 -16792 -17068 -16728
rect -17164 -16808 -17068 -16792
rect -17164 -16872 -17148 -16808
rect -17084 -16872 -17068 -16808
rect -17164 -16888 -17068 -16872
rect -17164 -16952 -17148 -16888
rect -17084 -16952 -17068 -16888
rect -17164 -16968 -17068 -16952
rect -17164 -17032 -17148 -16968
rect -17084 -17032 -17068 -16968
rect -17164 -17048 -17068 -17032
rect -17164 -17112 -17148 -17048
rect -17084 -17112 -17068 -17048
rect -17164 -17128 -17068 -17112
rect -18576 -17228 -18480 -17192
rect -17164 -17192 -17148 -17128
rect -17084 -17192 -17068 -17128
rect -16745 -16448 -16023 -16439
rect -16745 -17152 -16736 -16448
rect -16032 -17152 -16023 -16448
rect -16745 -17161 -16023 -17152
rect -15752 -16472 -15736 -16408
rect -15672 -16472 -15656 -16408
rect -14340 -16408 -14244 -16372
rect -15752 -16488 -15656 -16472
rect -15752 -16552 -15736 -16488
rect -15672 -16552 -15656 -16488
rect -15752 -16568 -15656 -16552
rect -15752 -16632 -15736 -16568
rect -15672 -16632 -15656 -16568
rect -15752 -16648 -15656 -16632
rect -15752 -16712 -15736 -16648
rect -15672 -16712 -15656 -16648
rect -15752 -16728 -15656 -16712
rect -15752 -16792 -15736 -16728
rect -15672 -16792 -15656 -16728
rect -15752 -16808 -15656 -16792
rect -15752 -16872 -15736 -16808
rect -15672 -16872 -15656 -16808
rect -15752 -16888 -15656 -16872
rect -15752 -16952 -15736 -16888
rect -15672 -16952 -15656 -16888
rect -15752 -16968 -15656 -16952
rect -15752 -17032 -15736 -16968
rect -15672 -17032 -15656 -16968
rect -15752 -17048 -15656 -17032
rect -15752 -17112 -15736 -17048
rect -15672 -17112 -15656 -17048
rect -15752 -17128 -15656 -17112
rect -17164 -17228 -17068 -17192
rect -15752 -17192 -15736 -17128
rect -15672 -17192 -15656 -17128
rect -15333 -16448 -14611 -16439
rect -15333 -17152 -15324 -16448
rect -14620 -17152 -14611 -16448
rect -15333 -17161 -14611 -17152
rect -14340 -16472 -14324 -16408
rect -14260 -16472 -14244 -16408
rect -12928 -16408 -12832 -16372
rect -14340 -16488 -14244 -16472
rect -14340 -16552 -14324 -16488
rect -14260 -16552 -14244 -16488
rect -14340 -16568 -14244 -16552
rect -14340 -16632 -14324 -16568
rect -14260 -16632 -14244 -16568
rect -14340 -16648 -14244 -16632
rect -14340 -16712 -14324 -16648
rect -14260 -16712 -14244 -16648
rect -14340 -16728 -14244 -16712
rect -14340 -16792 -14324 -16728
rect -14260 -16792 -14244 -16728
rect -14340 -16808 -14244 -16792
rect -14340 -16872 -14324 -16808
rect -14260 -16872 -14244 -16808
rect -14340 -16888 -14244 -16872
rect -14340 -16952 -14324 -16888
rect -14260 -16952 -14244 -16888
rect -14340 -16968 -14244 -16952
rect -14340 -17032 -14324 -16968
rect -14260 -17032 -14244 -16968
rect -14340 -17048 -14244 -17032
rect -14340 -17112 -14324 -17048
rect -14260 -17112 -14244 -17048
rect -14340 -17128 -14244 -17112
rect -15752 -17228 -15656 -17192
rect -14340 -17192 -14324 -17128
rect -14260 -17192 -14244 -17128
rect -13921 -16448 -13199 -16439
rect -13921 -17152 -13912 -16448
rect -13208 -17152 -13199 -16448
rect -13921 -17161 -13199 -17152
rect -12928 -16472 -12912 -16408
rect -12848 -16472 -12832 -16408
rect -11516 -16408 -11420 -16372
rect -12928 -16488 -12832 -16472
rect -12928 -16552 -12912 -16488
rect -12848 -16552 -12832 -16488
rect -12928 -16568 -12832 -16552
rect -12928 -16632 -12912 -16568
rect -12848 -16632 -12832 -16568
rect -12928 -16648 -12832 -16632
rect -12928 -16712 -12912 -16648
rect -12848 -16712 -12832 -16648
rect -12928 -16728 -12832 -16712
rect -12928 -16792 -12912 -16728
rect -12848 -16792 -12832 -16728
rect -12928 -16808 -12832 -16792
rect -12928 -16872 -12912 -16808
rect -12848 -16872 -12832 -16808
rect -12928 -16888 -12832 -16872
rect -12928 -16952 -12912 -16888
rect -12848 -16952 -12832 -16888
rect -12928 -16968 -12832 -16952
rect -12928 -17032 -12912 -16968
rect -12848 -17032 -12832 -16968
rect -12928 -17048 -12832 -17032
rect -12928 -17112 -12912 -17048
rect -12848 -17112 -12832 -17048
rect -12928 -17128 -12832 -17112
rect -14340 -17228 -14244 -17192
rect -12928 -17192 -12912 -17128
rect -12848 -17192 -12832 -17128
rect -12509 -16448 -11787 -16439
rect -12509 -17152 -12500 -16448
rect -11796 -17152 -11787 -16448
rect -12509 -17161 -11787 -17152
rect -11516 -16472 -11500 -16408
rect -11436 -16472 -11420 -16408
rect -10104 -16408 -10008 -16372
rect -11516 -16488 -11420 -16472
rect -11516 -16552 -11500 -16488
rect -11436 -16552 -11420 -16488
rect -11516 -16568 -11420 -16552
rect -11516 -16632 -11500 -16568
rect -11436 -16632 -11420 -16568
rect -11516 -16648 -11420 -16632
rect -11516 -16712 -11500 -16648
rect -11436 -16712 -11420 -16648
rect -11516 -16728 -11420 -16712
rect -11516 -16792 -11500 -16728
rect -11436 -16792 -11420 -16728
rect -11516 -16808 -11420 -16792
rect -11516 -16872 -11500 -16808
rect -11436 -16872 -11420 -16808
rect -11516 -16888 -11420 -16872
rect -11516 -16952 -11500 -16888
rect -11436 -16952 -11420 -16888
rect -11516 -16968 -11420 -16952
rect -11516 -17032 -11500 -16968
rect -11436 -17032 -11420 -16968
rect -11516 -17048 -11420 -17032
rect -11516 -17112 -11500 -17048
rect -11436 -17112 -11420 -17048
rect -11516 -17128 -11420 -17112
rect -12928 -17228 -12832 -17192
rect -11516 -17192 -11500 -17128
rect -11436 -17192 -11420 -17128
rect -11097 -16448 -10375 -16439
rect -11097 -17152 -11088 -16448
rect -10384 -17152 -10375 -16448
rect -11097 -17161 -10375 -17152
rect -10104 -16472 -10088 -16408
rect -10024 -16472 -10008 -16408
rect -8692 -16408 -8596 -16372
rect -10104 -16488 -10008 -16472
rect -10104 -16552 -10088 -16488
rect -10024 -16552 -10008 -16488
rect -10104 -16568 -10008 -16552
rect -10104 -16632 -10088 -16568
rect -10024 -16632 -10008 -16568
rect -10104 -16648 -10008 -16632
rect -10104 -16712 -10088 -16648
rect -10024 -16712 -10008 -16648
rect -10104 -16728 -10008 -16712
rect -10104 -16792 -10088 -16728
rect -10024 -16792 -10008 -16728
rect -10104 -16808 -10008 -16792
rect -10104 -16872 -10088 -16808
rect -10024 -16872 -10008 -16808
rect -10104 -16888 -10008 -16872
rect -10104 -16952 -10088 -16888
rect -10024 -16952 -10008 -16888
rect -10104 -16968 -10008 -16952
rect -10104 -17032 -10088 -16968
rect -10024 -17032 -10008 -16968
rect -10104 -17048 -10008 -17032
rect -10104 -17112 -10088 -17048
rect -10024 -17112 -10008 -17048
rect -10104 -17128 -10008 -17112
rect -11516 -17228 -11420 -17192
rect -10104 -17192 -10088 -17128
rect -10024 -17192 -10008 -17128
rect -9685 -16448 -8963 -16439
rect -9685 -17152 -9676 -16448
rect -8972 -17152 -8963 -16448
rect -9685 -17161 -8963 -17152
rect -8692 -16472 -8676 -16408
rect -8612 -16472 -8596 -16408
rect -7280 -16408 -7184 -16372
rect -8692 -16488 -8596 -16472
rect -8692 -16552 -8676 -16488
rect -8612 -16552 -8596 -16488
rect -8692 -16568 -8596 -16552
rect -8692 -16632 -8676 -16568
rect -8612 -16632 -8596 -16568
rect -8692 -16648 -8596 -16632
rect -8692 -16712 -8676 -16648
rect -8612 -16712 -8596 -16648
rect -8692 -16728 -8596 -16712
rect -8692 -16792 -8676 -16728
rect -8612 -16792 -8596 -16728
rect -8692 -16808 -8596 -16792
rect -8692 -16872 -8676 -16808
rect -8612 -16872 -8596 -16808
rect -8692 -16888 -8596 -16872
rect -8692 -16952 -8676 -16888
rect -8612 -16952 -8596 -16888
rect -8692 -16968 -8596 -16952
rect -8692 -17032 -8676 -16968
rect -8612 -17032 -8596 -16968
rect -8692 -17048 -8596 -17032
rect -8692 -17112 -8676 -17048
rect -8612 -17112 -8596 -17048
rect -8692 -17128 -8596 -17112
rect -10104 -17228 -10008 -17192
rect -8692 -17192 -8676 -17128
rect -8612 -17192 -8596 -17128
rect -8273 -16448 -7551 -16439
rect -8273 -17152 -8264 -16448
rect -7560 -17152 -7551 -16448
rect -8273 -17161 -7551 -17152
rect -7280 -16472 -7264 -16408
rect -7200 -16472 -7184 -16408
rect -5868 -16408 -5772 -16372
rect -7280 -16488 -7184 -16472
rect -7280 -16552 -7264 -16488
rect -7200 -16552 -7184 -16488
rect -7280 -16568 -7184 -16552
rect -7280 -16632 -7264 -16568
rect -7200 -16632 -7184 -16568
rect -7280 -16648 -7184 -16632
rect -7280 -16712 -7264 -16648
rect -7200 -16712 -7184 -16648
rect -7280 -16728 -7184 -16712
rect -7280 -16792 -7264 -16728
rect -7200 -16792 -7184 -16728
rect -7280 -16808 -7184 -16792
rect -7280 -16872 -7264 -16808
rect -7200 -16872 -7184 -16808
rect -7280 -16888 -7184 -16872
rect -7280 -16952 -7264 -16888
rect -7200 -16952 -7184 -16888
rect -7280 -16968 -7184 -16952
rect -7280 -17032 -7264 -16968
rect -7200 -17032 -7184 -16968
rect -7280 -17048 -7184 -17032
rect -7280 -17112 -7264 -17048
rect -7200 -17112 -7184 -17048
rect -7280 -17128 -7184 -17112
rect -8692 -17228 -8596 -17192
rect -7280 -17192 -7264 -17128
rect -7200 -17192 -7184 -17128
rect -6861 -16448 -6139 -16439
rect -6861 -17152 -6852 -16448
rect -6148 -17152 -6139 -16448
rect -6861 -17161 -6139 -17152
rect -5868 -16472 -5852 -16408
rect -5788 -16472 -5772 -16408
rect -4456 -16408 -4360 -16372
rect -5868 -16488 -5772 -16472
rect -5868 -16552 -5852 -16488
rect -5788 -16552 -5772 -16488
rect -5868 -16568 -5772 -16552
rect -5868 -16632 -5852 -16568
rect -5788 -16632 -5772 -16568
rect -5868 -16648 -5772 -16632
rect -5868 -16712 -5852 -16648
rect -5788 -16712 -5772 -16648
rect -5868 -16728 -5772 -16712
rect -5868 -16792 -5852 -16728
rect -5788 -16792 -5772 -16728
rect -5868 -16808 -5772 -16792
rect -5868 -16872 -5852 -16808
rect -5788 -16872 -5772 -16808
rect -5868 -16888 -5772 -16872
rect -5868 -16952 -5852 -16888
rect -5788 -16952 -5772 -16888
rect -5868 -16968 -5772 -16952
rect -5868 -17032 -5852 -16968
rect -5788 -17032 -5772 -16968
rect -5868 -17048 -5772 -17032
rect -5868 -17112 -5852 -17048
rect -5788 -17112 -5772 -17048
rect -5868 -17128 -5772 -17112
rect -7280 -17228 -7184 -17192
rect -5868 -17192 -5852 -17128
rect -5788 -17192 -5772 -17128
rect -5449 -16448 -4727 -16439
rect -5449 -17152 -5440 -16448
rect -4736 -17152 -4727 -16448
rect -5449 -17161 -4727 -17152
rect -4456 -16472 -4440 -16408
rect -4376 -16472 -4360 -16408
rect -3044 -16408 -2948 -16372
rect -4456 -16488 -4360 -16472
rect -4456 -16552 -4440 -16488
rect -4376 -16552 -4360 -16488
rect -4456 -16568 -4360 -16552
rect -4456 -16632 -4440 -16568
rect -4376 -16632 -4360 -16568
rect -4456 -16648 -4360 -16632
rect -4456 -16712 -4440 -16648
rect -4376 -16712 -4360 -16648
rect -4456 -16728 -4360 -16712
rect -4456 -16792 -4440 -16728
rect -4376 -16792 -4360 -16728
rect -4456 -16808 -4360 -16792
rect -4456 -16872 -4440 -16808
rect -4376 -16872 -4360 -16808
rect -4456 -16888 -4360 -16872
rect -4456 -16952 -4440 -16888
rect -4376 -16952 -4360 -16888
rect -4456 -16968 -4360 -16952
rect -4456 -17032 -4440 -16968
rect -4376 -17032 -4360 -16968
rect -4456 -17048 -4360 -17032
rect -4456 -17112 -4440 -17048
rect -4376 -17112 -4360 -17048
rect -4456 -17128 -4360 -17112
rect -5868 -17228 -5772 -17192
rect -4456 -17192 -4440 -17128
rect -4376 -17192 -4360 -17128
rect -4037 -16448 -3315 -16439
rect -4037 -17152 -4028 -16448
rect -3324 -17152 -3315 -16448
rect -4037 -17161 -3315 -17152
rect -3044 -16472 -3028 -16408
rect -2964 -16472 -2948 -16408
rect -1632 -16408 -1536 -16372
rect -3044 -16488 -2948 -16472
rect -3044 -16552 -3028 -16488
rect -2964 -16552 -2948 -16488
rect -3044 -16568 -2948 -16552
rect -3044 -16632 -3028 -16568
rect -2964 -16632 -2948 -16568
rect -3044 -16648 -2948 -16632
rect -3044 -16712 -3028 -16648
rect -2964 -16712 -2948 -16648
rect -3044 -16728 -2948 -16712
rect -3044 -16792 -3028 -16728
rect -2964 -16792 -2948 -16728
rect -3044 -16808 -2948 -16792
rect -3044 -16872 -3028 -16808
rect -2964 -16872 -2948 -16808
rect -3044 -16888 -2948 -16872
rect -3044 -16952 -3028 -16888
rect -2964 -16952 -2948 -16888
rect -3044 -16968 -2948 -16952
rect -3044 -17032 -3028 -16968
rect -2964 -17032 -2948 -16968
rect -3044 -17048 -2948 -17032
rect -3044 -17112 -3028 -17048
rect -2964 -17112 -2948 -17048
rect -3044 -17128 -2948 -17112
rect -4456 -17228 -4360 -17192
rect -3044 -17192 -3028 -17128
rect -2964 -17192 -2948 -17128
rect -2625 -16448 -1903 -16439
rect -2625 -17152 -2616 -16448
rect -1912 -17152 -1903 -16448
rect -2625 -17161 -1903 -17152
rect -1632 -16472 -1616 -16408
rect -1552 -16472 -1536 -16408
rect -220 -16408 -124 -16372
rect -1632 -16488 -1536 -16472
rect -1632 -16552 -1616 -16488
rect -1552 -16552 -1536 -16488
rect -1632 -16568 -1536 -16552
rect -1632 -16632 -1616 -16568
rect -1552 -16632 -1536 -16568
rect -1632 -16648 -1536 -16632
rect -1632 -16712 -1616 -16648
rect -1552 -16712 -1536 -16648
rect -1632 -16728 -1536 -16712
rect -1632 -16792 -1616 -16728
rect -1552 -16792 -1536 -16728
rect -1632 -16808 -1536 -16792
rect -1632 -16872 -1616 -16808
rect -1552 -16872 -1536 -16808
rect -1632 -16888 -1536 -16872
rect -1632 -16952 -1616 -16888
rect -1552 -16952 -1536 -16888
rect -1632 -16968 -1536 -16952
rect -1632 -17032 -1616 -16968
rect -1552 -17032 -1536 -16968
rect -1632 -17048 -1536 -17032
rect -1632 -17112 -1616 -17048
rect -1552 -17112 -1536 -17048
rect -1632 -17128 -1536 -17112
rect -3044 -17228 -2948 -17192
rect -1632 -17192 -1616 -17128
rect -1552 -17192 -1536 -17128
rect -1213 -16448 -491 -16439
rect -1213 -17152 -1204 -16448
rect -500 -17152 -491 -16448
rect -1213 -17161 -491 -17152
rect -220 -16472 -204 -16408
rect -140 -16472 -124 -16408
rect 1192 -16408 1288 -16372
rect -220 -16488 -124 -16472
rect -220 -16552 -204 -16488
rect -140 -16552 -124 -16488
rect -220 -16568 -124 -16552
rect -220 -16632 -204 -16568
rect -140 -16632 -124 -16568
rect -220 -16648 -124 -16632
rect -220 -16712 -204 -16648
rect -140 -16712 -124 -16648
rect -220 -16728 -124 -16712
rect -220 -16792 -204 -16728
rect -140 -16792 -124 -16728
rect -220 -16808 -124 -16792
rect -220 -16872 -204 -16808
rect -140 -16872 -124 -16808
rect -220 -16888 -124 -16872
rect -220 -16952 -204 -16888
rect -140 -16952 -124 -16888
rect -220 -16968 -124 -16952
rect -220 -17032 -204 -16968
rect -140 -17032 -124 -16968
rect -220 -17048 -124 -17032
rect -220 -17112 -204 -17048
rect -140 -17112 -124 -17048
rect -220 -17128 -124 -17112
rect -1632 -17228 -1536 -17192
rect -220 -17192 -204 -17128
rect -140 -17192 -124 -17128
rect 199 -16448 921 -16439
rect 199 -17152 208 -16448
rect 912 -17152 921 -16448
rect 199 -17161 921 -17152
rect 1192 -16472 1208 -16408
rect 1272 -16472 1288 -16408
rect 2604 -16408 2700 -16372
rect 1192 -16488 1288 -16472
rect 1192 -16552 1208 -16488
rect 1272 -16552 1288 -16488
rect 1192 -16568 1288 -16552
rect 1192 -16632 1208 -16568
rect 1272 -16632 1288 -16568
rect 1192 -16648 1288 -16632
rect 1192 -16712 1208 -16648
rect 1272 -16712 1288 -16648
rect 1192 -16728 1288 -16712
rect 1192 -16792 1208 -16728
rect 1272 -16792 1288 -16728
rect 1192 -16808 1288 -16792
rect 1192 -16872 1208 -16808
rect 1272 -16872 1288 -16808
rect 1192 -16888 1288 -16872
rect 1192 -16952 1208 -16888
rect 1272 -16952 1288 -16888
rect 1192 -16968 1288 -16952
rect 1192 -17032 1208 -16968
rect 1272 -17032 1288 -16968
rect 1192 -17048 1288 -17032
rect 1192 -17112 1208 -17048
rect 1272 -17112 1288 -17048
rect 1192 -17128 1288 -17112
rect -220 -17228 -124 -17192
rect 1192 -17192 1208 -17128
rect 1272 -17192 1288 -17128
rect 1611 -16448 2333 -16439
rect 1611 -17152 1620 -16448
rect 2324 -17152 2333 -16448
rect 1611 -17161 2333 -17152
rect 2604 -16472 2620 -16408
rect 2684 -16472 2700 -16408
rect 4016 -16408 4112 -16372
rect 2604 -16488 2700 -16472
rect 2604 -16552 2620 -16488
rect 2684 -16552 2700 -16488
rect 2604 -16568 2700 -16552
rect 2604 -16632 2620 -16568
rect 2684 -16632 2700 -16568
rect 2604 -16648 2700 -16632
rect 2604 -16712 2620 -16648
rect 2684 -16712 2700 -16648
rect 2604 -16728 2700 -16712
rect 2604 -16792 2620 -16728
rect 2684 -16792 2700 -16728
rect 2604 -16808 2700 -16792
rect 2604 -16872 2620 -16808
rect 2684 -16872 2700 -16808
rect 2604 -16888 2700 -16872
rect 2604 -16952 2620 -16888
rect 2684 -16952 2700 -16888
rect 2604 -16968 2700 -16952
rect 2604 -17032 2620 -16968
rect 2684 -17032 2700 -16968
rect 2604 -17048 2700 -17032
rect 2604 -17112 2620 -17048
rect 2684 -17112 2700 -17048
rect 2604 -17128 2700 -17112
rect 1192 -17228 1288 -17192
rect 2604 -17192 2620 -17128
rect 2684 -17192 2700 -17128
rect 3023 -16448 3745 -16439
rect 3023 -17152 3032 -16448
rect 3736 -17152 3745 -16448
rect 3023 -17161 3745 -17152
rect 4016 -16472 4032 -16408
rect 4096 -16472 4112 -16408
rect 5428 -16408 5524 -16372
rect 4016 -16488 4112 -16472
rect 4016 -16552 4032 -16488
rect 4096 -16552 4112 -16488
rect 4016 -16568 4112 -16552
rect 4016 -16632 4032 -16568
rect 4096 -16632 4112 -16568
rect 4016 -16648 4112 -16632
rect 4016 -16712 4032 -16648
rect 4096 -16712 4112 -16648
rect 4016 -16728 4112 -16712
rect 4016 -16792 4032 -16728
rect 4096 -16792 4112 -16728
rect 4016 -16808 4112 -16792
rect 4016 -16872 4032 -16808
rect 4096 -16872 4112 -16808
rect 4016 -16888 4112 -16872
rect 4016 -16952 4032 -16888
rect 4096 -16952 4112 -16888
rect 4016 -16968 4112 -16952
rect 4016 -17032 4032 -16968
rect 4096 -17032 4112 -16968
rect 4016 -17048 4112 -17032
rect 4016 -17112 4032 -17048
rect 4096 -17112 4112 -17048
rect 4016 -17128 4112 -17112
rect 2604 -17228 2700 -17192
rect 4016 -17192 4032 -17128
rect 4096 -17192 4112 -17128
rect 4435 -16448 5157 -16439
rect 4435 -17152 4444 -16448
rect 5148 -17152 5157 -16448
rect 4435 -17161 5157 -17152
rect 5428 -16472 5444 -16408
rect 5508 -16472 5524 -16408
rect 6840 -16408 6936 -16372
rect 5428 -16488 5524 -16472
rect 5428 -16552 5444 -16488
rect 5508 -16552 5524 -16488
rect 5428 -16568 5524 -16552
rect 5428 -16632 5444 -16568
rect 5508 -16632 5524 -16568
rect 5428 -16648 5524 -16632
rect 5428 -16712 5444 -16648
rect 5508 -16712 5524 -16648
rect 5428 -16728 5524 -16712
rect 5428 -16792 5444 -16728
rect 5508 -16792 5524 -16728
rect 5428 -16808 5524 -16792
rect 5428 -16872 5444 -16808
rect 5508 -16872 5524 -16808
rect 5428 -16888 5524 -16872
rect 5428 -16952 5444 -16888
rect 5508 -16952 5524 -16888
rect 5428 -16968 5524 -16952
rect 5428 -17032 5444 -16968
rect 5508 -17032 5524 -16968
rect 5428 -17048 5524 -17032
rect 5428 -17112 5444 -17048
rect 5508 -17112 5524 -17048
rect 5428 -17128 5524 -17112
rect 4016 -17228 4112 -17192
rect 5428 -17192 5444 -17128
rect 5508 -17192 5524 -17128
rect 5847 -16448 6569 -16439
rect 5847 -17152 5856 -16448
rect 6560 -17152 6569 -16448
rect 5847 -17161 6569 -17152
rect 6840 -16472 6856 -16408
rect 6920 -16472 6936 -16408
rect 8252 -16408 8348 -16372
rect 6840 -16488 6936 -16472
rect 6840 -16552 6856 -16488
rect 6920 -16552 6936 -16488
rect 6840 -16568 6936 -16552
rect 6840 -16632 6856 -16568
rect 6920 -16632 6936 -16568
rect 6840 -16648 6936 -16632
rect 6840 -16712 6856 -16648
rect 6920 -16712 6936 -16648
rect 6840 -16728 6936 -16712
rect 6840 -16792 6856 -16728
rect 6920 -16792 6936 -16728
rect 6840 -16808 6936 -16792
rect 6840 -16872 6856 -16808
rect 6920 -16872 6936 -16808
rect 6840 -16888 6936 -16872
rect 6840 -16952 6856 -16888
rect 6920 -16952 6936 -16888
rect 6840 -16968 6936 -16952
rect 6840 -17032 6856 -16968
rect 6920 -17032 6936 -16968
rect 6840 -17048 6936 -17032
rect 6840 -17112 6856 -17048
rect 6920 -17112 6936 -17048
rect 6840 -17128 6936 -17112
rect 5428 -17228 5524 -17192
rect 6840 -17192 6856 -17128
rect 6920 -17192 6936 -17128
rect 7259 -16448 7981 -16439
rect 7259 -17152 7268 -16448
rect 7972 -17152 7981 -16448
rect 7259 -17161 7981 -17152
rect 8252 -16472 8268 -16408
rect 8332 -16472 8348 -16408
rect 9664 -16408 9760 -16372
rect 8252 -16488 8348 -16472
rect 8252 -16552 8268 -16488
rect 8332 -16552 8348 -16488
rect 8252 -16568 8348 -16552
rect 8252 -16632 8268 -16568
rect 8332 -16632 8348 -16568
rect 8252 -16648 8348 -16632
rect 8252 -16712 8268 -16648
rect 8332 -16712 8348 -16648
rect 8252 -16728 8348 -16712
rect 8252 -16792 8268 -16728
rect 8332 -16792 8348 -16728
rect 8252 -16808 8348 -16792
rect 8252 -16872 8268 -16808
rect 8332 -16872 8348 -16808
rect 8252 -16888 8348 -16872
rect 8252 -16952 8268 -16888
rect 8332 -16952 8348 -16888
rect 8252 -16968 8348 -16952
rect 8252 -17032 8268 -16968
rect 8332 -17032 8348 -16968
rect 8252 -17048 8348 -17032
rect 8252 -17112 8268 -17048
rect 8332 -17112 8348 -17048
rect 8252 -17128 8348 -17112
rect 6840 -17228 6936 -17192
rect 8252 -17192 8268 -17128
rect 8332 -17192 8348 -17128
rect 8671 -16448 9393 -16439
rect 8671 -17152 8680 -16448
rect 9384 -17152 9393 -16448
rect 8671 -17161 9393 -17152
rect 9664 -16472 9680 -16408
rect 9744 -16472 9760 -16408
rect 11076 -16408 11172 -16372
rect 9664 -16488 9760 -16472
rect 9664 -16552 9680 -16488
rect 9744 -16552 9760 -16488
rect 9664 -16568 9760 -16552
rect 9664 -16632 9680 -16568
rect 9744 -16632 9760 -16568
rect 9664 -16648 9760 -16632
rect 9664 -16712 9680 -16648
rect 9744 -16712 9760 -16648
rect 9664 -16728 9760 -16712
rect 9664 -16792 9680 -16728
rect 9744 -16792 9760 -16728
rect 9664 -16808 9760 -16792
rect 9664 -16872 9680 -16808
rect 9744 -16872 9760 -16808
rect 9664 -16888 9760 -16872
rect 9664 -16952 9680 -16888
rect 9744 -16952 9760 -16888
rect 9664 -16968 9760 -16952
rect 9664 -17032 9680 -16968
rect 9744 -17032 9760 -16968
rect 9664 -17048 9760 -17032
rect 9664 -17112 9680 -17048
rect 9744 -17112 9760 -17048
rect 9664 -17128 9760 -17112
rect 8252 -17228 8348 -17192
rect 9664 -17192 9680 -17128
rect 9744 -17192 9760 -17128
rect 10083 -16448 10805 -16439
rect 10083 -17152 10092 -16448
rect 10796 -17152 10805 -16448
rect 10083 -17161 10805 -17152
rect 11076 -16472 11092 -16408
rect 11156 -16472 11172 -16408
rect 12488 -16408 12584 -16372
rect 11076 -16488 11172 -16472
rect 11076 -16552 11092 -16488
rect 11156 -16552 11172 -16488
rect 11076 -16568 11172 -16552
rect 11076 -16632 11092 -16568
rect 11156 -16632 11172 -16568
rect 11076 -16648 11172 -16632
rect 11076 -16712 11092 -16648
rect 11156 -16712 11172 -16648
rect 11076 -16728 11172 -16712
rect 11076 -16792 11092 -16728
rect 11156 -16792 11172 -16728
rect 11076 -16808 11172 -16792
rect 11076 -16872 11092 -16808
rect 11156 -16872 11172 -16808
rect 11076 -16888 11172 -16872
rect 11076 -16952 11092 -16888
rect 11156 -16952 11172 -16888
rect 11076 -16968 11172 -16952
rect 11076 -17032 11092 -16968
rect 11156 -17032 11172 -16968
rect 11076 -17048 11172 -17032
rect 11076 -17112 11092 -17048
rect 11156 -17112 11172 -17048
rect 11076 -17128 11172 -17112
rect 9664 -17228 9760 -17192
rect 11076 -17192 11092 -17128
rect 11156 -17192 11172 -17128
rect 11495 -16448 12217 -16439
rect 11495 -17152 11504 -16448
rect 12208 -17152 12217 -16448
rect 11495 -17161 12217 -17152
rect 12488 -16472 12504 -16408
rect 12568 -16472 12584 -16408
rect 13900 -16408 13996 -16372
rect 12488 -16488 12584 -16472
rect 12488 -16552 12504 -16488
rect 12568 -16552 12584 -16488
rect 12488 -16568 12584 -16552
rect 12488 -16632 12504 -16568
rect 12568 -16632 12584 -16568
rect 12488 -16648 12584 -16632
rect 12488 -16712 12504 -16648
rect 12568 -16712 12584 -16648
rect 12488 -16728 12584 -16712
rect 12488 -16792 12504 -16728
rect 12568 -16792 12584 -16728
rect 12488 -16808 12584 -16792
rect 12488 -16872 12504 -16808
rect 12568 -16872 12584 -16808
rect 12488 -16888 12584 -16872
rect 12488 -16952 12504 -16888
rect 12568 -16952 12584 -16888
rect 12488 -16968 12584 -16952
rect 12488 -17032 12504 -16968
rect 12568 -17032 12584 -16968
rect 12488 -17048 12584 -17032
rect 12488 -17112 12504 -17048
rect 12568 -17112 12584 -17048
rect 12488 -17128 12584 -17112
rect 11076 -17228 11172 -17192
rect 12488 -17192 12504 -17128
rect 12568 -17192 12584 -17128
rect 12907 -16448 13629 -16439
rect 12907 -17152 12916 -16448
rect 13620 -17152 13629 -16448
rect 12907 -17161 13629 -17152
rect 13900 -16472 13916 -16408
rect 13980 -16472 13996 -16408
rect 15312 -16408 15408 -16372
rect 13900 -16488 13996 -16472
rect 13900 -16552 13916 -16488
rect 13980 -16552 13996 -16488
rect 13900 -16568 13996 -16552
rect 13900 -16632 13916 -16568
rect 13980 -16632 13996 -16568
rect 13900 -16648 13996 -16632
rect 13900 -16712 13916 -16648
rect 13980 -16712 13996 -16648
rect 13900 -16728 13996 -16712
rect 13900 -16792 13916 -16728
rect 13980 -16792 13996 -16728
rect 13900 -16808 13996 -16792
rect 13900 -16872 13916 -16808
rect 13980 -16872 13996 -16808
rect 13900 -16888 13996 -16872
rect 13900 -16952 13916 -16888
rect 13980 -16952 13996 -16888
rect 13900 -16968 13996 -16952
rect 13900 -17032 13916 -16968
rect 13980 -17032 13996 -16968
rect 13900 -17048 13996 -17032
rect 13900 -17112 13916 -17048
rect 13980 -17112 13996 -17048
rect 13900 -17128 13996 -17112
rect 12488 -17228 12584 -17192
rect 13900 -17192 13916 -17128
rect 13980 -17192 13996 -17128
rect 14319 -16448 15041 -16439
rect 14319 -17152 14328 -16448
rect 15032 -17152 15041 -16448
rect 14319 -17161 15041 -17152
rect 15312 -16472 15328 -16408
rect 15392 -16472 15408 -16408
rect 16724 -16408 16820 -16372
rect 15312 -16488 15408 -16472
rect 15312 -16552 15328 -16488
rect 15392 -16552 15408 -16488
rect 15312 -16568 15408 -16552
rect 15312 -16632 15328 -16568
rect 15392 -16632 15408 -16568
rect 15312 -16648 15408 -16632
rect 15312 -16712 15328 -16648
rect 15392 -16712 15408 -16648
rect 15312 -16728 15408 -16712
rect 15312 -16792 15328 -16728
rect 15392 -16792 15408 -16728
rect 15312 -16808 15408 -16792
rect 15312 -16872 15328 -16808
rect 15392 -16872 15408 -16808
rect 15312 -16888 15408 -16872
rect 15312 -16952 15328 -16888
rect 15392 -16952 15408 -16888
rect 15312 -16968 15408 -16952
rect 15312 -17032 15328 -16968
rect 15392 -17032 15408 -16968
rect 15312 -17048 15408 -17032
rect 15312 -17112 15328 -17048
rect 15392 -17112 15408 -17048
rect 15312 -17128 15408 -17112
rect 13900 -17228 13996 -17192
rect 15312 -17192 15328 -17128
rect 15392 -17192 15408 -17128
rect 15731 -16448 16453 -16439
rect 15731 -17152 15740 -16448
rect 16444 -17152 16453 -16448
rect 15731 -17161 16453 -17152
rect 16724 -16472 16740 -16408
rect 16804 -16472 16820 -16408
rect 18136 -16408 18232 -16372
rect 16724 -16488 16820 -16472
rect 16724 -16552 16740 -16488
rect 16804 -16552 16820 -16488
rect 16724 -16568 16820 -16552
rect 16724 -16632 16740 -16568
rect 16804 -16632 16820 -16568
rect 16724 -16648 16820 -16632
rect 16724 -16712 16740 -16648
rect 16804 -16712 16820 -16648
rect 16724 -16728 16820 -16712
rect 16724 -16792 16740 -16728
rect 16804 -16792 16820 -16728
rect 16724 -16808 16820 -16792
rect 16724 -16872 16740 -16808
rect 16804 -16872 16820 -16808
rect 16724 -16888 16820 -16872
rect 16724 -16952 16740 -16888
rect 16804 -16952 16820 -16888
rect 16724 -16968 16820 -16952
rect 16724 -17032 16740 -16968
rect 16804 -17032 16820 -16968
rect 16724 -17048 16820 -17032
rect 16724 -17112 16740 -17048
rect 16804 -17112 16820 -17048
rect 16724 -17128 16820 -17112
rect 15312 -17228 15408 -17192
rect 16724 -17192 16740 -17128
rect 16804 -17192 16820 -17128
rect 17143 -16448 17865 -16439
rect 17143 -17152 17152 -16448
rect 17856 -17152 17865 -16448
rect 17143 -17161 17865 -17152
rect 18136 -16472 18152 -16408
rect 18216 -16472 18232 -16408
rect 19548 -16408 19644 -16372
rect 18136 -16488 18232 -16472
rect 18136 -16552 18152 -16488
rect 18216 -16552 18232 -16488
rect 18136 -16568 18232 -16552
rect 18136 -16632 18152 -16568
rect 18216 -16632 18232 -16568
rect 18136 -16648 18232 -16632
rect 18136 -16712 18152 -16648
rect 18216 -16712 18232 -16648
rect 18136 -16728 18232 -16712
rect 18136 -16792 18152 -16728
rect 18216 -16792 18232 -16728
rect 18136 -16808 18232 -16792
rect 18136 -16872 18152 -16808
rect 18216 -16872 18232 -16808
rect 18136 -16888 18232 -16872
rect 18136 -16952 18152 -16888
rect 18216 -16952 18232 -16888
rect 18136 -16968 18232 -16952
rect 18136 -17032 18152 -16968
rect 18216 -17032 18232 -16968
rect 18136 -17048 18232 -17032
rect 18136 -17112 18152 -17048
rect 18216 -17112 18232 -17048
rect 18136 -17128 18232 -17112
rect 16724 -17228 16820 -17192
rect 18136 -17192 18152 -17128
rect 18216 -17192 18232 -17128
rect 18555 -16448 19277 -16439
rect 18555 -17152 18564 -16448
rect 19268 -17152 19277 -16448
rect 18555 -17161 19277 -17152
rect 19548 -16472 19564 -16408
rect 19628 -16472 19644 -16408
rect 20960 -16408 21056 -16372
rect 19548 -16488 19644 -16472
rect 19548 -16552 19564 -16488
rect 19628 -16552 19644 -16488
rect 19548 -16568 19644 -16552
rect 19548 -16632 19564 -16568
rect 19628 -16632 19644 -16568
rect 19548 -16648 19644 -16632
rect 19548 -16712 19564 -16648
rect 19628 -16712 19644 -16648
rect 19548 -16728 19644 -16712
rect 19548 -16792 19564 -16728
rect 19628 -16792 19644 -16728
rect 19548 -16808 19644 -16792
rect 19548 -16872 19564 -16808
rect 19628 -16872 19644 -16808
rect 19548 -16888 19644 -16872
rect 19548 -16952 19564 -16888
rect 19628 -16952 19644 -16888
rect 19548 -16968 19644 -16952
rect 19548 -17032 19564 -16968
rect 19628 -17032 19644 -16968
rect 19548 -17048 19644 -17032
rect 19548 -17112 19564 -17048
rect 19628 -17112 19644 -17048
rect 19548 -17128 19644 -17112
rect 18136 -17228 18232 -17192
rect 19548 -17192 19564 -17128
rect 19628 -17192 19644 -17128
rect 19967 -16448 20689 -16439
rect 19967 -17152 19976 -16448
rect 20680 -17152 20689 -16448
rect 19967 -17161 20689 -17152
rect 20960 -16472 20976 -16408
rect 21040 -16472 21056 -16408
rect 22372 -16408 22468 -16372
rect 20960 -16488 21056 -16472
rect 20960 -16552 20976 -16488
rect 21040 -16552 21056 -16488
rect 20960 -16568 21056 -16552
rect 20960 -16632 20976 -16568
rect 21040 -16632 21056 -16568
rect 20960 -16648 21056 -16632
rect 20960 -16712 20976 -16648
rect 21040 -16712 21056 -16648
rect 20960 -16728 21056 -16712
rect 20960 -16792 20976 -16728
rect 21040 -16792 21056 -16728
rect 20960 -16808 21056 -16792
rect 20960 -16872 20976 -16808
rect 21040 -16872 21056 -16808
rect 20960 -16888 21056 -16872
rect 20960 -16952 20976 -16888
rect 21040 -16952 21056 -16888
rect 20960 -16968 21056 -16952
rect 20960 -17032 20976 -16968
rect 21040 -17032 21056 -16968
rect 20960 -17048 21056 -17032
rect 20960 -17112 20976 -17048
rect 21040 -17112 21056 -17048
rect 20960 -17128 21056 -17112
rect 19548 -17228 19644 -17192
rect 20960 -17192 20976 -17128
rect 21040 -17192 21056 -17128
rect 21379 -16448 22101 -16439
rect 21379 -17152 21388 -16448
rect 22092 -17152 22101 -16448
rect 21379 -17161 22101 -17152
rect 22372 -16472 22388 -16408
rect 22452 -16472 22468 -16408
rect 23784 -16408 23880 -16372
rect 22372 -16488 22468 -16472
rect 22372 -16552 22388 -16488
rect 22452 -16552 22468 -16488
rect 22372 -16568 22468 -16552
rect 22372 -16632 22388 -16568
rect 22452 -16632 22468 -16568
rect 22372 -16648 22468 -16632
rect 22372 -16712 22388 -16648
rect 22452 -16712 22468 -16648
rect 22372 -16728 22468 -16712
rect 22372 -16792 22388 -16728
rect 22452 -16792 22468 -16728
rect 22372 -16808 22468 -16792
rect 22372 -16872 22388 -16808
rect 22452 -16872 22468 -16808
rect 22372 -16888 22468 -16872
rect 22372 -16952 22388 -16888
rect 22452 -16952 22468 -16888
rect 22372 -16968 22468 -16952
rect 22372 -17032 22388 -16968
rect 22452 -17032 22468 -16968
rect 22372 -17048 22468 -17032
rect 22372 -17112 22388 -17048
rect 22452 -17112 22468 -17048
rect 22372 -17128 22468 -17112
rect 20960 -17228 21056 -17192
rect 22372 -17192 22388 -17128
rect 22452 -17192 22468 -17128
rect 22791 -16448 23513 -16439
rect 22791 -17152 22800 -16448
rect 23504 -17152 23513 -16448
rect 22791 -17161 23513 -17152
rect 23784 -16472 23800 -16408
rect 23864 -16472 23880 -16408
rect 23784 -16488 23880 -16472
rect 23784 -16552 23800 -16488
rect 23864 -16552 23880 -16488
rect 23784 -16568 23880 -16552
rect 23784 -16632 23800 -16568
rect 23864 -16632 23880 -16568
rect 23784 -16648 23880 -16632
rect 23784 -16712 23800 -16648
rect 23864 -16712 23880 -16648
rect 23784 -16728 23880 -16712
rect 23784 -16792 23800 -16728
rect 23864 -16792 23880 -16728
rect 23784 -16808 23880 -16792
rect 23784 -16872 23800 -16808
rect 23864 -16872 23880 -16808
rect 23784 -16888 23880 -16872
rect 23784 -16952 23800 -16888
rect 23864 -16952 23880 -16888
rect 23784 -16968 23880 -16952
rect 23784 -17032 23800 -16968
rect 23864 -17032 23880 -16968
rect 23784 -17048 23880 -17032
rect 23784 -17112 23800 -17048
rect 23864 -17112 23880 -17048
rect 23784 -17128 23880 -17112
rect 22372 -17228 22468 -17192
rect 23784 -17192 23800 -17128
rect 23864 -17192 23880 -17128
rect 23784 -17228 23880 -17192
rect -22812 -17528 -22716 -17492
rect -23805 -17568 -23083 -17559
rect -23805 -18272 -23796 -17568
rect -23092 -18272 -23083 -17568
rect -23805 -18281 -23083 -18272
rect -22812 -17592 -22796 -17528
rect -22732 -17592 -22716 -17528
rect -21400 -17528 -21304 -17492
rect -22812 -17608 -22716 -17592
rect -22812 -17672 -22796 -17608
rect -22732 -17672 -22716 -17608
rect -22812 -17688 -22716 -17672
rect -22812 -17752 -22796 -17688
rect -22732 -17752 -22716 -17688
rect -22812 -17768 -22716 -17752
rect -22812 -17832 -22796 -17768
rect -22732 -17832 -22716 -17768
rect -22812 -17848 -22716 -17832
rect -22812 -17912 -22796 -17848
rect -22732 -17912 -22716 -17848
rect -22812 -17928 -22716 -17912
rect -22812 -17992 -22796 -17928
rect -22732 -17992 -22716 -17928
rect -22812 -18008 -22716 -17992
rect -22812 -18072 -22796 -18008
rect -22732 -18072 -22716 -18008
rect -22812 -18088 -22716 -18072
rect -22812 -18152 -22796 -18088
rect -22732 -18152 -22716 -18088
rect -22812 -18168 -22716 -18152
rect -22812 -18232 -22796 -18168
rect -22732 -18232 -22716 -18168
rect -22812 -18248 -22716 -18232
rect -22812 -18312 -22796 -18248
rect -22732 -18312 -22716 -18248
rect -22393 -17568 -21671 -17559
rect -22393 -18272 -22384 -17568
rect -21680 -18272 -21671 -17568
rect -22393 -18281 -21671 -18272
rect -21400 -17592 -21384 -17528
rect -21320 -17592 -21304 -17528
rect -19988 -17528 -19892 -17492
rect -21400 -17608 -21304 -17592
rect -21400 -17672 -21384 -17608
rect -21320 -17672 -21304 -17608
rect -21400 -17688 -21304 -17672
rect -21400 -17752 -21384 -17688
rect -21320 -17752 -21304 -17688
rect -21400 -17768 -21304 -17752
rect -21400 -17832 -21384 -17768
rect -21320 -17832 -21304 -17768
rect -21400 -17848 -21304 -17832
rect -21400 -17912 -21384 -17848
rect -21320 -17912 -21304 -17848
rect -21400 -17928 -21304 -17912
rect -21400 -17992 -21384 -17928
rect -21320 -17992 -21304 -17928
rect -21400 -18008 -21304 -17992
rect -21400 -18072 -21384 -18008
rect -21320 -18072 -21304 -18008
rect -21400 -18088 -21304 -18072
rect -21400 -18152 -21384 -18088
rect -21320 -18152 -21304 -18088
rect -21400 -18168 -21304 -18152
rect -21400 -18232 -21384 -18168
rect -21320 -18232 -21304 -18168
rect -21400 -18248 -21304 -18232
rect -22812 -18348 -22716 -18312
rect -21400 -18312 -21384 -18248
rect -21320 -18312 -21304 -18248
rect -20981 -17568 -20259 -17559
rect -20981 -18272 -20972 -17568
rect -20268 -18272 -20259 -17568
rect -20981 -18281 -20259 -18272
rect -19988 -17592 -19972 -17528
rect -19908 -17592 -19892 -17528
rect -18576 -17528 -18480 -17492
rect -19988 -17608 -19892 -17592
rect -19988 -17672 -19972 -17608
rect -19908 -17672 -19892 -17608
rect -19988 -17688 -19892 -17672
rect -19988 -17752 -19972 -17688
rect -19908 -17752 -19892 -17688
rect -19988 -17768 -19892 -17752
rect -19988 -17832 -19972 -17768
rect -19908 -17832 -19892 -17768
rect -19988 -17848 -19892 -17832
rect -19988 -17912 -19972 -17848
rect -19908 -17912 -19892 -17848
rect -19988 -17928 -19892 -17912
rect -19988 -17992 -19972 -17928
rect -19908 -17992 -19892 -17928
rect -19988 -18008 -19892 -17992
rect -19988 -18072 -19972 -18008
rect -19908 -18072 -19892 -18008
rect -19988 -18088 -19892 -18072
rect -19988 -18152 -19972 -18088
rect -19908 -18152 -19892 -18088
rect -19988 -18168 -19892 -18152
rect -19988 -18232 -19972 -18168
rect -19908 -18232 -19892 -18168
rect -19988 -18248 -19892 -18232
rect -21400 -18348 -21304 -18312
rect -19988 -18312 -19972 -18248
rect -19908 -18312 -19892 -18248
rect -19569 -17568 -18847 -17559
rect -19569 -18272 -19560 -17568
rect -18856 -18272 -18847 -17568
rect -19569 -18281 -18847 -18272
rect -18576 -17592 -18560 -17528
rect -18496 -17592 -18480 -17528
rect -17164 -17528 -17068 -17492
rect -18576 -17608 -18480 -17592
rect -18576 -17672 -18560 -17608
rect -18496 -17672 -18480 -17608
rect -18576 -17688 -18480 -17672
rect -18576 -17752 -18560 -17688
rect -18496 -17752 -18480 -17688
rect -18576 -17768 -18480 -17752
rect -18576 -17832 -18560 -17768
rect -18496 -17832 -18480 -17768
rect -18576 -17848 -18480 -17832
rect -18576 -17912 -18560 -17848
rect -18496 -17912 -18480 -17848
rect -18576 -17928 -18480 -17912
rect -18576 -17992 -18560 -17928
rect -18496 -17992 -18480 -17928
rect -18576 -18008 -18480 -17992
rect -18576 -18072 -18560 -18008
rect -18496 -18072 -18480 -18008
rect -18576 -18088 -18480 -18072
rect -18576 -18152 -18560 -18088
rect -18496 -18152 -18480 -18088
rect -18576 -18168 -18480 -18152
rect -18576 -18232 -18560 -18168
rect -18496 -18232 -18480 -18168
rect -18576 -18248 -18480 -18232
rect -19988 -18348 -19892 -18312
rect -18576 -18312 -18560 -18248
rect -18496 -18312 -18480 -18248
rect -18157 -17568 -17435 -17559
rect -18157 -18272 -18148 -17568
rect -17444 -18272 -17435 -17568
rect -18157 -18281 -17435 -18272
rect -17164 -17592 -17148 -17528
rect -17084 -17592 -17068 -17528
rect -15752 -17528 -15656 -17492
rect -17164 -17608 -17068 -17592
rect -17164 -17672 -17148 -17608
rect -17084 -17672 -17068 -17608
rect -17164 -17688 -17068 -17672
rect -17164 -17752 -17148 -17688
rect -17084 -17752 -17068 -17688
rect -17164 -17768 -17068 -17752
rect -17164 -17832 -17148 -17768
rect -17084 -17832 -17068 -17768
rect -17164 -17848 -17068 -17832
rect -17164 -17912 -17148 -17848
rect -17084 -17912 -17068 -17848
rect -17164 -17928 -17068 -17912
rect -17164 -17992 -17148 -17928
rect -17084 -17992 -17068 -17928
rect -17164 -18008 -17068 -17992
rect -17164 -18072 -17148 -18008
rect -17084 -18072 -17068 -18008
rect -17164 -18088 -17068 -18072
rect -17164 -18152 -17148 -18088
rect -17084 -18152 -17068 -18088
rect -17164 -18168 -17068 -18152
rect -17164 -18232 -17148 -18168
rect -17084 -18232 -17068 -18168
rect -17164 -18248 -17068 -18232
rect -18576 -18348 -18480 -18312
rect -17164 -18312 -17148 -18248
rect -17084 -18312 -17068 -18248
rect -16745 -17568 -16023 -17559
rect -16745 -18272 -16736 -17568
rect -16032 -18272 -16023 -17568
rect -16745 -18281 -16023 -18272
rect -15752 -17592 -15736 -17528
rect -15672 -17592 -15656 -17528
rect -14340 -17528 -14244 -17492
rect -15752 -17608 -15656 -17592
rect -15752 -17672 -15736 -17608
rect -15672 -17672 -15656 -17608
rect -15752 -17688 -15656 -17672
rect -15752 -17752 -15736 -17688
rect -15672 -17752 -15656 -17688
rect -15752 -17768 -15656 -17752
rect -15752 -17832 -15736 -17768
rect -15672 -17832 -15656 -17768
rect -15752 -17848 -15656 -17832
rect -15752 -17912 -15736 -17848
rect -15672 -17912 -15656 -17848
rect -15752 -17928 -15656 -17912
rect -15752 -17992 -15736 -17928
rect -15672 -17992 -15656 -17928
rect -15752 -18008 -15656 -17992
rect -15752 -18072 -15736 -18008
rect -15672 -18072 -15656 -18008
rect -15752 -18088 -15656 -18072
rect -15752 -18152 -15736 -18088
rect -15672 -18152 -15656 -18088
rect -15752 -18168 -15656 -18152
rect -15752 -18232 -15736 -18168
rect -15672 -18232 -15656 -18168
rect -15752 -18248 -15656 -18232
rect -17164 -18348 -17068 -18312
rect -15752 -18312 -15736 -18248
rect -15672 -18312 -15656 -18248
rect -15333 -17568 -14611 -17559
rect -15333 -18272 -15324 -17568
rect -14620 -18272 -14611 -17568
rect -15333 -18281 -14611 -18272
rect -14340 -17592 -14324 -17528
rect -14260 -17592 -14244 -17528
rect -12928 -17528 -12832 -17492
rect -14340 -17608 -14244 -17592
rect -14340 -17672 -14324 -17608
rect -14260 -17672 -14244 -17608
rect -14340 -17688 -14244 -17672
rect -14340 -17752 -14324 -17688
rect -14260 -17752 -14244 -17688
rect -14340 -17768 -14244 -17752
rect -14340 -17832 -14324 -17768
rect -14260 -17832 -14244 -17768
rect -14340 -17848 -14244 -17832
rect -14340 -17912 -14324 -17848
rect -14260 -17912 -14244 -17848
rect -14340 -17928 -14244 -17912
rect -14340 -17992 -14324 -17928
rect -14260 -17992 -14244 -17928
rect -14340 -18008 -14244 -17992
rect -14340 -18072 -14324 -18008
rect -14260 -18072 -14244 -18008
rect -14340 -18088 -14244 -18072
rect -14340 -18152 -14324 -18088
rect -14260 -18152 -14244 -18088
rect -14340 -18168 -14244 -18152
rect -14340 -18232 -14324 -18168
rect -14260 -18232 -14244 -18168
rect -14340 -18248 -14244 -18232
rect -15752 -18348 -15656 -18312
rect -14340 -18312 -14324 -18248
rect -14260 -18312 -14244 -18248
rect -13921 -17568 -13199 -17559
rect -13921 -18272 -13912 -17568
rect -13208 -18272 -13199 -17568
rect -13921 -18281 -13199 -18272
rect -12928 -17592 -12912 -17528
rect -12848 -17592 -12832 -17528
rect -11516 -17528 -11420 -17492
rect -12928 -17608 -12832 -17592
rect -12928 -17672 -12912 -17608
rect -12848 -17672 -12832 -17608
rect -12928 -17688 -12832 -17672
rect -12928 -17752 -12912 -17688
rect -12848 -17752 -12832 -17688
rect -12928 -17768 -12832 -17752
rect -12928 -17832 -12912 -17768
rect -12848 -17832 -12832 -17768
rect -12928 -17848 -12832 -17832
rect -12928 -17912 -12912 -17848
rect -12848 -17912 -12832 -17848
rect -12928 -17928 -12832 -17912
rect -12928 -17992 -12912 -17928
rect -12848 -17992 -12832 -17928
rect -12928 -18008 -12832 -17992
rect -12928 -18072 -12912 -18008
rect -12848 -18072 -12832 -18008
rect -12928 -18088 -12832 -18072
rect -12928 -18152 -12912 -18088
rect -12848 -18152 -12832 -18088
rect -12928 -18168 -12832 -18152
rect -12928 -18232 -12912 -18168
rect -12848 -18232 -12832 -18168
rect -12928 -18248 -12832 -18232
rect -14340 -18348 -14244 -18312
rect -12928 -18312 -12912 -18248
rect -12848 -18312 -12832 -18248
rect -12509 -17568 -11787 -17559
rect -12509 -18272 -12500 -17568
rect -11796 -18272 -11787 -17568
rect -12509 -18281 -11787 -18272
rect -11516 -17592 -11500 -17528
rect -11436 -17592 -11420 -17528
rect -10104 -17528 -10008 -17492
rect -11516 -17608 -11420 -17592
rect -11516 -17672 -11500 -17608
rect -11436 -17672 -11420 -17608
rect -11516 -17688 -11420 -17672
rect -11516 -17752 -11500 -17688
rect -11436 -17752 -11420 -17688
rect -11516 -17768 -11420 -17752
rect -11516 -17832 -11500 -17768
rect -11436 -17832 -11420 -17768
rect -11516 -17848 -11420 -17832
rect -11516 -17912 -11500 -17848
rect -11436 -17912 -11420 -17848
rect -11516 -17928 -11420 -17912
rect -11516 -17992 -11500 -17928
rect -11436 -17992 -11420 -17928
rect -11516 -18008 -11420 -17992
rect -11516 -18072 -11500 -18008
rect -11436 -18072 -11420 -18008
rect -11516 -18088 -11420 -18072
rect -11516 -18152 -11500 -18088
rect -11436 -18152 -11420 -18088
rect -11516 -18168 -11420 -18152
rect -11516 -18232 -11500 -18168
rect -11436 -18232 -11420 -18168
rect -11516 -18248 -11420 -18232
rect -12928 -18348 -12832 -18312
rect -11516 -18312 -11500 -18248
rect -11436 -18312 -11420 -18248
rect -11097 -17568 -10375 -17559
rect -11097 -18272 -11088 -17568
rect -10384 -18272 -10375 -17568
rect -11097 -18281 -10375 -18272
rect -10104 -17592 -10088 -17528
rect -10024 -17592 -10008 -17528
rect -8692 -17528 -8596 -17492
rect -10104 -17608 -10008 -17592
rect -10104 -17672 -10088 -17608
rect -10024 -17672 -10008 -17608
rect -10104 -17688 -10008 -17672
rect -10104 -17752 -10088 -17688
rect -10024 -17752 -10008 -17688
rect -10104 -17768 -10008 -17752
rect -10104 -17832 -10088 -17768
rect -10024 -17832 -10008 -17768
rect -10104 -17848 -10008 -17832
rect -10104 -17912 -10088 -17848
rect -10024 -17912 -10008 -17848
rect -10104 -17928 -10008 -17912
rect -10104 -17992 -10088 -17928
rect -10024 -17992 -10008 -17928
rect -10104 -18008 -10008 -17992
rect -10104 -18072 -10088 -18008
rect -10024 -18072 -10008 -18008
rect -10104 -18088 -10008 -18072
rect -10104 -18152 -10088 -18088
rect -10024 -18152 -10008 -18088
rect -10104 -18168 -10008 -18152
rect -10104 -18232 -10088 -18168
rect -10024 -18232 -10008 -18168
rect -10104 -18248 -10008 -18232
rect -11516 -18348 -11420 -18312
rect -10104 -18312 -10088 -18248
rect -10024 -18312 -10008 -18248
rect -9685 -17568 -8963 -17559
rect -9685 -18272 -9676 -17568
rect -8972 -18272 -8963 -17568
rect -9685 -18281 -8963 -18272
rect -8692 -17592 -8676 -17528
rect -8612 -17592 -8596 -17528
rect -7280 -17528 -7184 -17492
rect -8692 -17608 -8596 -17592
rect -8692 -17672 -8676 -17608
rect -8612 -17672 -8596 -17608
rect -8692 -17688 -8596 -17672
rect -8692 -17752 -8676 -17688
rect -8612 -17752 -8596 -17688
rect -8692 -17768 -8596 -17752
rect -8692 -17832 -8676 -17768
rect -8612 -17832 -8596 -17768
rect -8692 -17848 -8596 -17832
rect -8692 -17912 -8676 -17848
rect -8612 -17912 -8596 -17848
rect -8692 -17928 -8596 -17912
rect -8692 -17992 -8676 -17928
rect -8612 -17992 -8596 -17928
rect -8692 -18008 -8596 -17992
rect -8692 -18072 -8676 -18008
rect -8612 -18072 -8596 -18008
rect -8692 -18088 -8596 -18072
rect -8692 -18152 -8676 -18088
rect -8612 -18152 -8596 -18088
rect -8692 -18168 -8596 -18152
rect -8692 -18232 -8676 -18168
rect -8612 -18232 -8596 -18168
rect -8692 -18248 -8596 -18232
rect -10104 -18348 -10008 -18312
rect -8692 -18312 -8676 -18248
rect -8612 -18312 -8596 -18248
rect -8273 -17568 -7551 -17559
rect -8273 -18272 -8264 -17568
rect -7560 -18272 -7551 -17568
rect -8273 -18281 -7551 -18272
rect -7280 -17592 -7264 -17528
rect -7200 -17592 -7184 -17528
rect -5868 -17528 -5772 -17492
rect -7280 -17608 -7184 -17592
rect -7280 -17672 -7264 -17608
rect -7200 -17672 -7184 -17608
rect -7280 -17688 -7184 -17672
rect -7280 -17752 -7264 -17688
rect -7200 -17752 -7184 -17688
rect -7280 -17768 -7184 -17752
rect -7280 -17832 -7264 -17768
rect -7200 -17832 -7184 -17768
rect -7280 -17848 -7184 -17832
rect -7280 -17912 -7264 -17848
rect -7200 -17912 -7184 -17848
rect -7280 -17928 -7184 -17912
rect -7280 -17992 -7264 -17928
rect -7200 -17992 -7184 -17928
rect -7280 -18008 -7184 -17992
rect -7280 -18072 -7264 -18008
rect -7200 -18072 -7184 -18008
rect -7280 -18088 -7184 -18072
rect -7280 -18152 -7264 -18088
rect -7200 -18152 -7184 -18088
rect -7280 -18168 -7184 -18152
rect -7280 -18232 -7264 -18168
rect -7200 -18232 -7184 -18168
rect -7280 -18248 -7184 -18232
rect -8692 -18348 -8596 -18312
rect -7280 -18312 -7264 -18248
rect -7200 -18312 -7184 -18248
rect -6861 -17568 -6139 -17559
rect -6861 -18272 -6852 -17568
rect -6148 -18272 -6139 -17568
rect -6861 -18281 -6139 -18272
rect -5868 -17592 -5852 -17528
rect -5788 -17592 -5772 -17528
rect -4456 -17528 -4360 -17492
rect -5868 -17608 -5772 -17592
rect -5868 -17672 -5852 -17608
rect -5788 -17672 -5772 -17608
rect -5868 -17688 -5772 -17672
rect -5868 -17752 -5852 -17688
rect -5788 -17752 -5772 -17688
rect -5868 -17768 -5772 -17752
rect -5868 -17832 -5852 -17768
rect -5788 -17832 -5772 -17768
rect -5868 -17848 -5772 -17832
rect -5868 -17912 -5852 -17848
rect -5788 -17912 -5772 -17848
rect -5868 -17928 -5772 -17912
rect -5868 -17992 -5852 -17928
rect -5788 -17992 -5772 -17928
rect -5868 -18008 -5772 -17992
rect -5868 -18072 -5852 -18008
rect -5788 -18072 -5772 -18008
rect -5868 -18088 -5772 -18072
rect -5868 -18152 -5852 -18088
rect -5788 -18152 -5772 -18088
rect -5868 -18168 -5772 -18152
rect -5868 -18232 -5852 -18168
rect -5788 -18232 -5772 -18168
rect -5868 -18248 -5772 -18232
rect -7280 -18348 -7184 -18312
rect -5868 -18312 -5852 -18248
rect -5788 -18312 -5772 -18248
rect -5449 -17568 -4727 -17559
rect -5449 -18272 -5440 -17568
rect -4736 -18272 -4727 -17568
rect -5449 -18281 -4727 -18272
rect -4456 -17592 -4440 -17528
rect -4376 -17592 -4360 -17528
rect -3044 -17528 -2948 -17492
rect -4456 -17608 -4360 -17592
rect -4456 -17672 -4440 -17608
rect -4376 -17672 -4360 -17608
rect -4456 -17688 -4360 -17672
rect -4456 -17752 -4440 -17688
rect -4376 -17752 -4360 -17688
rect -4456 -17768 -4360 -17752
rect -4456 -17832 -4440 -17768
rect -4376 -17832 -4360 -17768
rect -4456 -17848 -4360 -17832
rect -4456 -17912 -4440 -17848
rect -4376 -17912 -4360 -17848
rect -4456 -17928 -4360 -17912
rect -4456 -17992 -4440 -17928
rect -4376 -17992 -4360 -17928
rect -4456 -18008 -4360 -17992
rect -4456 -18072 -4440 -18008
rect -4376 -18072 -4360 -18008
rect -4456 -18088 -4360 -18072
rect -4456 -18152 -4440 -18088
rect -4376 -18152 -4360 -18088
rect -4456 -18168 -4360 -18152
rect -4456 -18232 -4440 -18168
rect -4376 -18232 -4360 -18168
rect -4456 -18248 -4360 -18232
rect -5868 -18348 -5772 -18312
rect -4456 -18312 -4440 -18248
rect -4376 -18312 -4360 -18248
rect -4037 -17568 -3315 -17559
rect -4037 -18272 -4028 -17568
rect -3324 -18272 -3315 -17568
rect -4037 -18281 -3315 -18272
rect -3044 -17592 -3028 -17528
rect -2964 -17592 -2948 -17528
rect -1632 -17528 -1536 -17492
rect -3044 -17608 -2948 -17592
rect -3044 -17672 -3028 -17608
rect -2964 -17672 -2948 -17608
rect -3044 -17688 -2948 -17672
rect -3044 -17752 -3028 -17688
rect -2964 -17752 -2948 -17688
rect -3044 -17768 -2948 -17752
rect -3044 -17832 -3028 -17768
rect -2964 -17832 -2948 -17768
rect -3044 -17848 -2948 -17832
rect -3044 -17912 -3028 -17848
rect -2964 -17912 -2948 -17848
rect -3044 -17928 -2948 -17912
rect -3044 -17992 -3028 -17928
rect -2964 -17992 -2948 -17928
rect -3044 -18008 -2948 -17992
rect -3044 -18072 -3028 -18008
rect -2964 -18072 -2948 -18008
rect -3044 -18088 -2948 -18072
rect -3044 -18152 -3028 -18088
rect -2964 -18152 -2948 -18088
rect -3044 -18168 -2948 -18152
rect -3044 -18232 -3028 -18168
rect -2964 -18232 -2948 -18168
rect -3044 -18248 -2948 -18232
rect -4456 -18348 -4360 -18312
rect -3044 -18312 -3028 -18248
rect -2964 -18312 -2948 -18248
rect -2625 -17568 -1903 -17559
rect -2625 -18272 -2616 -17568
rect -1912 -18272 -1903 -17568
rect -2625 -18281 -1903 -18272
rect -1632 -17592 -1616 -17528
rect -1552 -17592 -1536 -17528
rect -220 -17528 -124 -17492
rect -1632 -17608 -1536 -17592
rect -1632 -17672 -1616 -17608
rect -1552 -17672 -1536 -17608
rect -1632 -17688 -1536 -17672
rect -1632 -17752 -1616 -17688
rect -1552 -17752 -1536 -17688
rect -1632 -17768 -1536 -17752
rect -1632 -17832 -1616 -17768
rect -1552 -17832 -1536 -17768
rect -1632 -17848 -1536 -17832
rect -1632 -17912 -1616 -17848
rect -1552 -17912 -1536 -17848
rect -1632 -17928 -1536 -17912
rect -1632 -17992 -1616 -17928
rect -1552 -17992 -1536 -17928
rect -1632 -18008 -1536 -17992
rect -1632 -18072 -1616 -18008
rect -1552 -18072 -1536 -18008
rect -1632 -18088 -1536 -18072
rect -1632 -18152 -1616 -18088
rect -1552 -18152 -1536 -18088
rect -1632 -18168 -1536 -18152
rect -1632 -18232 -1616 -18168
rect -1552 -18232 -1536 -18168
rect -1632 -18248 -1536 -18232
rect -3044 -18348 -2948 -18312
rect -1632 -18312 -1616 -18248
rect -1552 -18312 -1536 -18248
rect -1213 -17568 -491 -17559
rect -1213 -18272 -1204 -17568
rect -500 -18272 -491 -17568
rect -1213 -18281 -491 -18272
rect -220 -17592 -204 -17528
rect -140 -17592 -124 -17528
rect 1192 -17528 1288 -17492
rect -220 -17608 -124 -17592
rect -220 -17672 -204 -17608
rect -140 -17672 -124 -17608
rect -220 -17688 -124 -17672
rect -220 -17752 -204 -17688
rect -140 -17752 -124 -17688
rect -220 -17768 -124 -17752
rect -220 -17832 -204 -17768
rect -140 -17832 -124 -17768
rect -220 -17848 -124 -17832
rect -220 -17912 -204 -17848
rect -140 -17912 -124 -17848
rect -220 -17928 -124 -17912
rect -220 -17992 -204 -17928
rect -140 -17992 -124 -17928
rect -220 -18008 -124 -17992
rect -220 -18072 -204 -18008
rect -140 -18072 -124 -18008
rect -220 -18088 -124 -18072
rect -220 -18152 -204 -18088
rect -140 -18152 -124 -18088
rect -220 -18168 -124 -18152
rect -220 -18232 -204 -18168
rect -140 -18232 -124 -18168
rect -220 -18248 -124 -18232
rect -1632 -18348 -1536 -18312
rect -220 -18312 -204 -18248
rect -140 -18312 -124 -18248
rect 199 -17568 921 -17559
rect 199 -18272 208 -17568
rect 912 -18272 921 -17568
rect 199 -18281 921 -18272
rect 1192 -17592 1208 -17528
rect 1272 -17592 1288 -17528
rect 2604 -17528 2700 -17492
rect 1192 -17608 1288 -17592
rect 1192 -17672 1208 -17608
rect 1272 -17672 1288 -17608
rect 1192 -17688 1288 -17672
rect 1192 -17752 1208 -17688
rect 1272 -17752 1288 -17688
rect 1192 -17768 1288 -17752
rect 1192 -17832 1208 -17768
rect 1272 -17832 1288 -17768
rect 1192 -17848 1288 -17832
rect 1192 -17912 1208 -17848
rect 1272 -17912 1288 -17848
rect 1192 -17928 1288 -17912
rect 1192 -17992 1208 -17928
rect 1272 -17992 1288 -17928
rect 1192 -18008 1288 -17992
rect 1192 -18072 1208 -18008
rect 1272 -18072 1288 -18008
rect 1192 -18088 1288 -18072
rect 1192 -18152 1208 -18088
rect 1272 -18152 1288 -18088
rect 1192 -18168 1288 -18152
rect 1192 -18232 1208 -18168
rect 1272 -18232 1288 -18168
rect 1192 -18248 1288 -18232
rect -220 -18348 -124 -18312
rect 1192 -18312 1208 -18248
rect 1272 -18312 1288 -18248
rect 1611 -17568 2333 -17559
rect 1611 -18272 1620 -17568
rect 2324 -18272 2333 -17568
rect 1611 -18281 2333 -18272
rect 2604 -17592 2620 -17528
rect 2684 -17592 2700 -17528
rect 4016 -17528 4112 -17492
rect 2604 -17608 2700 -17592
rect 2604 -17672 2620 -17608
rect 2684 -17672 2700 -17608
rect 2604 -17688 2700 -17672
rect 2604 -17752 2620 -17688
rect 2684 -17752 2700 -17688
rect 2604 -17768 2700 -17752
rect 2604 -17832 2620 -17768
rect 2684 -17832 2700 -17768
rect 2604 -17848 2700 -17832
rect 2604 -17912 2620 -17848
rect 2684 -17912 2700 -17848
rect 2604 -17928 2700 -17912
rect 2604 -17992 2620 -17928
rect 2684 -17992 2700 -17928
rect 2604 -18008 2700 -17992
rect 2604 -18072 2620 -18008
rect 2684 -18072 2700 -18008
rect 2604 -18088 2700 -18072
rect 2604 -18152 2620 -18088
rect 2684 -18152 2700 -18088
rect 2604 -18168 2700 -18152
rect 2604 -18232 2620 -18168
rect 2684 -18232 2700 -18168
rect 2604 -18248 2700 -18232
rect 1192 -18348 1288 -18312
rect 2604 -18312 2620 -18248
rect 2684 -18312 2700 -18248
rect 3023 -17568 3745 -17559
rect 3023 -18272 3032 -17568
rect 3736 -18272 3745 -17568
rect 3023 -18281 3745 -18272
rect 4016 -17592 4032 -17528
rect 4096 -17592 4112 -17528
rect 5428 -17528 5524 -17492
rect 4016 -17608 4112 -17592
rect 4016 -17672 4032 -17608
rect 4096 -17672 4112 -17608
rect 4016 -17688 4112 -17672
rect 4016 -17752 4032 -17688
rect 4096 -17752 4112 -17688
rect 4016 -17768 4112 -17752
rect 4016 -17832 4032 -17768
rect 4096 -17832 4112 -17768
rect 4016 -17848 4112 -17832
rect 4016 -17912 4032 -17848
rect 4096 -17912 4112 -17848
rect 4016 -17928 4112 -17912
rect 4016 -17992 4032 -17928
rect 4096 -17992 4112 -17928
rect 4016 -18008 4112 -17992
rect 4016 -18072 4032 -18008
rect 4096 -18072 4112 -18008
rect 4016 -18088 4112 -18072
rect 4016 -18152 4032 -18088
rect 4096 -18152 4112 -18088
rect 4016 -18168 4112 -18152
rect 4016 -18232 4032 -18168
rect 4096 -18232 4112 -18168
rect 4016 -18248 4112 -18232
rect 2604 -18348 2700 -18312
rect 4016 -18312 4032 -18248
rect 4096 -18312 4112 -18248
rect 4435 -17568 5157 -17559
rect 4435 -18272 4444 -17568
rect 5148 -18272 5157 -17568
rect 4435 -18281 5157 -18272
rect 5428 -17592 5444 -17528
rect 5508 -17592 5524 -17528
rect 6840 -17528 6936 -17492
rect 5428 -17608 5524 -17592
rect 5428 -17672 5444 -17608
rect 5508 -17672 5524 -17608
rect 5428 -17688 5524 -17672
rect 5428 -17752 5444 -17688
rect 5508 -17752 5524 -17688
rect 5428 -17768 5524 -17752
rect 5428 -17832 5444 -17768
rect 5508 -17832 5524 -17768
rect 5428 -17848 5524 -17832
rect 5428 -17912 5444 -17848
rect 5508 -17912 5524 -17848
rect 5428 -17928 5524 -17912
rect 5428 -17992 5444 -17928
rect 5508 -17992 5524 -17928
rect 5428 -18008 5524 -17992
rect 5428 -18072 5444 -18008
rect 5508 -18072 5524 -18008
rect 5428 -18088 5524 -18072
rect 5428 -18152 5444 -18088
rect 5508 -18152 5524 -18088
rect 5428 -18168 5524 -18152
rect 5428 -18232 5444 -18168
rect 5508 -18232 5524 -18168
rect 5428 -18248 5524 -18232
rect 4016 -18348 4112 -18312
rect 5428 -18312 5444 -18248
rect 5508 -18312 5524 -18248
rect 5847 -17568 6569 -17559
rect 5847 -18272 5856 -17568
rect 6560 -18272 6569 -17568
rect 5847 -18281 6569 -18272
rect 6840 -17592 6856 -17528
rect 6920 -17592 6936 -17528
rect 8252 -17528 8348 -17492
rect 6840 -17608 6936 -17592
rect 6840 -17672 6856 -17608
rect 6920 -17672 6936 -17608
rect 6840 -17688 6936 -17672
rect 6840 -17752 6856 -17688
rect 6920 -17752 6936 -17688
rect 6840 -17768 6936 -17752
rect 6840 -17832 6856 -17768
rect 6920 -17832 6936 -17768
rect 6840 -17848 6936 -17832
rect 6840 -17912 6856 -17848
rect 6920 -17912 6936 -17848
rect 6840 -17928 6936 -17912
rect 6840 -17992 6856 -17928
rect 6920 -17992 6936 -17928
rect 6840 -18008 6936 -17992
rect 6840 -18072 6856 -18008
rect 6920 -18072 6936 -18008
rect 6840 -18088 6936 -18072
rect 6840 -18152 6856 -18088
rect 6920 -18152 6936 -18088
rect 6840 -18168 6936 -18152
rect 6840 -18232 6856 -18168
rect 6920 -18232 6936 -18168
rect 6840 -18248 6936 -18232
rect 5428 -18348 5524 -18312
rect 6840 -18312 6856 -18248
rect 6920 -18312 6936 -18248
rect 7259 -17568 7981 -17559
rect 7259 -18272 7268 -17568
rect 7972 -18272 7981 -17568
rect 7259 -18281 7981 -18272
rect 8252 -17592 8268 -17528
rect 8332 -17592 8348 -17528
rect 9664 -17528 9760 -17492
rect 8252 -17608 8348 -17592
rect 8252 -17672 8268 -17608
rect 8332 -17672 8348 -17608
rect 8252 -17688 8348 -17672
rect 8252 -17752 8268 -17688
rect 8332 -17752 8348 -17688
rect 8252 -17768 8348 -17752
rect 8252 -17832 8268 -17768
rect 8332 -17832 8348 -17768
rect 8252 -17848 8348 -17832
rect 8252 -17912 8268 -17848
rect 8332 -17912 8348 -17848
rect 8252 -17928 8348 -17912
rect 8252 -17992 8268 -17928
rect 8332 -17992 8348 -17928
rect 8252 -18008 8348 -17992
rect 8252 -18072 8268 -18008
rect 8332 -18072 8348 -18008
rect 8252 -18088 8348 -18072
rect 8252 -18152 8268 -18088
rect 8332 -18152 8348 -18088
rect 8252 -18168 8348 -18152
rect 8252 -18232 8268 -18168
rect 8332 -18232 8348 -18168
rect 8252 -18248 8348 -18232
rect 6840 -18348 6936 -18312
rect 8252 -18312 8268 -18248
rect 8332 -18312 8348 -18248
rect 8671 -17568 9393 -17559
rect 8671 -18272 8680 -17568
rect 9384 -18272 9393 -17568
rect 8671 -18281 9393 -18272
rect 9664 -17592 9680 -17528
rect 9744 -17592 9760 -17528
rect 11076 -17528 11172 -17492
rect 9664 -17608 9760 -17592
rect 9664 -17672 9680 -17608
rect 9744 -17672 9760 -17608
rect 9664 -17688 9760 -17672
rect 9664 -17752 9680 -17688
rect 9744 -17752 9760 -17688
rect 9664 -17768 9760 -17752
rect 9664 -17832 9680 -17768
rect 9744 -17832 9760 -17768
rect 9664 -17848 9760 -17832
rect 9664 -17912 9680 -17848
rect 9744 -17912 9760 -17848
rect 9664 -17928 9760 -17912
rect 9664 -17992 9680 -17928
rect 9744 -17992 9760 -17928
rect 9664 -18008 9760 -17992
rect 9664 -18072 9680 -18008
rect 9744 -18072 9760 -18008
rect 9664 -18088 9760 -18072
rect 9664 -18152 9680 -18088
rect 9744 -18152 9760 -18088
rect 9664 -18168 9760 -18152
rect 9664 -18232 9680 -18168
rect 9744 -18232 9760 -18168
rect 9664 -18248 9760 -18232
rect 8252 -18348 8348 -18312
rect 9664 -18312 9680 -18248
rect 9744 -18312 9760 -18248
rect 10083 -17568 10805 -17559
rect 10083 -18272 10092 -17568
rect 10796 -18272 10805 -17568
rect 10083 -18281 10805 -18272
rect 11076 -17592 11092 -17528
rect 11156 -17592 11172 -17528
rect 12488 -17528 12584 -17492
rect 11076 -17608 11172 -17592
rect 11076 -17672 11092 -17608
rect 11156 -17672 11172 -17608
rect 11076 -17688 11172 -17672
rect 11076 -17752 11092 -17688
rect 11156 -17752 11172 -17688
rect 11076 -17768 11172 -17752
rect 11076 -17832 11092 -17768
rect 11156 -17832 11172 -17768
rect 11076 -17848 11172 -17832
rect 11076 -17912 11092 -17848
rect 11156 -17912 11172 -17848
rect 11076 -17928 11172 -17912
rect 11076 -17992 11092 -17928
rect 11156 -17992 11172 -17928
rect 11076 -18008 11172 -17992
rect 11076 -18072 11092 -18008
rect 11156 -18072 11172 -18008
rect 11076 -18088 11172 -18072
rect 11076 -18152 11092 -18088
rect 11156 -18152 11172 -18088
rect 11076 -18168 11172 -18152
rect 11076 -18232 11092 -18168
rect 11156 -18232 11172 -18168
rect 11076 -18248 11172 -18232
rect 9664 -18348 9760 -18312
rect 11076 -18312 11092 -18248
rect 11156 -18312 11172 -18248
rect 11495 -17568 12217 -17559
rect 11495 -18272 11504 -17568
rect 12208 -18272 12217 -17568
rect 11495 -18281 12217 -18272
rect 12488 -17592 12504 -17528
rect 12568 -17592 12584 -17528
rect 13900 -17528 13996 -17492
rect 12488 -17608 12584 -17592
rect 12488 -17672 12504 -17608
rect 12568 -17672 12584 -17608
rect 12488 -17688 12584 -17672
rect 12488 -17752 12504 -17688
rect 12568 -17752 12584 -17688
rect 12488 -17768 12584 -17752
rect 12488 -17832 12504 -17768
rect 12568 -17832 12584 -17768
rect 12488 -17848 12584 -17832
rect 12488 -17912 12504 -17848
rect 12568 -17912 12584 -17848
rect 12488 -17928 12584 -17912
rect 12488 -17992 12504 -17928
rect 12568 -17992 12584 -17928
rect 12488 -18008 12584 -17992
rect 12488 -18072 12504 -18008
rect 12568 -18072 12584 -18008
rect 12488 -18088 12584 -18072
rect 12488 -18152 12504 -18088
rect 12568 -18152 12584 -18088
rect 12488 -18168 12584 -18152
rect 12488 -18232 12504 -18168
rect 12568 -18232 12584 -18168
rect 12488 -18248 12584 -18232
rect 11076 -18348 11172 -18312
rect 12488 -18312 12504 -18248
rect 12568 -18312 12584 -18248
rect 12907 -17568 13629 -17559
rect 12907 -18272 12916 -17568
rect 13620 -18272 13629 -17568
rect 12907 -18281 13629 -18272
rect 13900 -17592 13916 -17528
rect 13980 -17592 13996 -17528
rect 15312 -17528 15408 -17492
rect 13900 -17608 13996 -17592
rect 13900 -17672 13916 -17608
rect 13980 -17672 13996 -17608
rect 13900 -17688 13996 -17672
rect 13900 -17752 13916 -17688
rect 13980 -17752 13996 -17688
rect 13900 -17768 13996 -17752
rect 13900 -17832 13916 -17768
rect 13980 -17832 13996 -17768
rect 13900 -17848 13996 -17832
rect 13900 -17912 13916 -17848
rect 13980 -17912 13996 -17848
rect 13900 -17928 13996 -17912
rect 13900 -17992 13916 -17928
rect 13980 -17992 13996 -17928
rect 13900 -18008 13996 -17992
rect 13900 -18072 13916 -18008
rect 13980 -18072 13996 -18008
rect 13900 -18088 13996 -18072
rect 13900 -18152 13916 -18088
rect 13980 -18152 13996 -18088
rect 13900 -18168 13996 -18152
rect 13900 -18232 13916 -18168
rect 13980 -18232 13996 -18168
rect 13900 -18248 13996 -18232
rect 12488 -18348 12584 -18312
rect 13900 -18312 13916 -18248
rect 13980 -18312 13996 -18248
rect 14319 -17568 15041 -17559
rect 14319 -18272 14328 -17568
rect 15032 -18272 15041 -17568
rect 14319 -18281 15041 -18272
rect 15312 -17592 15328 -17528
rect 15392 -17592 15408 -17528
rect 16724 -17528 16820 -17492
rect 15312 -17608 15408 -17592
rect 15312 -17672 15328 -17608
rect 15392 -17672 15408 -17608
rect 15312 -17688 15408 -17672
rect 15312 -17752 15328 -17688
rect 15392 -17752 15408 -17688
rect 15312 -17768 15408 -17752
rect 15312 -17832 15328 -17768
rect 15392 -17832 15408 -17768
rect 15312 -17848 15408 -17832
rect 15312 -17912 15328 -17848
rect 15392 -17912 15408 -17848
rect 15312 -17928 15408 -17912
rect 15312 -17992 15328 -17928
rect 15392 -17992 15408 -17928
rect 15312 -18008 15408 -17992
rect 15312 -18072 15328 -18008
rect 15392 -18072 15408 -18008
rect 15312 -18088 15408 -18072
rect 15312 -18152 15328 -18088
rect 15392 -18152 15408 -18088
rect 15312 -18168 15408 -18152
rect 15312 -18232 15328 -18168
rect 15392 -18232 15408 -18168
rect 15312 -18248 15408 -18232
rect 13900 -18348 13996 -18312
rect 15312 -18312 15328 -18248
rect 15392 -18312 15408 -18248
rect 15731 -17568 16453 -17559
rect 15731 -18272 15740 -17568
rect 16444 -18272 16453 -17568
rect 15731 -18281 16453 -18272
rect 16724 -17592 16740 -17528
rect 16804 -17592 16820 -17528
rect 18136 -17528 18232 -17492
rect 16724 -17608 16820 -17592
rect 16724 -17672 16740 -17608
rect 16804 -17672 16820 -17608
rect 16724 -17688 16820 -17672
rect 16724 -17752 16740 -17688
rect 16804 -17752 16820 -17688
rect 16724 -17768 16820 -17752
rect 16724 -17832 16740 -17768
rect 16804 -17832 16820 -17768
rect 16724 -17848 16820 -17832
rect 16724 -17912 16740 -17848
rect 16804 -17912 16820 -17848
rect 16724 -17928 16820 -17912
rect 16724 -17992 16740 -17928
rect 16804 -17992 16820 -17928
rect 16724 -18008 16820 -17992
rect 16724 -18072 16740 -18008
rect 16804 -18072 16820 -18008
rect 16724 -18088 16820 -18072
rect 16724 -18152 16740 -18088
rect 16804 -18152 16820 -18088
rect 16724 -18168 16820 -18152
rect 16724 -18232 16740 -18168
rect 16804 -18232 16820 -18168
rect 16724 -18248 16820 -18232
rect 15312 -18348 15408 -18312
rect 16724 -18312 16740 -18248
rect 16804 -18312 16820 -18248
rect 17143 -17568 17865 -17559
rect 17143 -18272 17152 -17568
rect 17856 -18272 17865 -17568
rect 17143 -18281 17865 -18272
rect 18136 -17592 18152 -17528
rect 18216 -17592 18232 -17528
rect 19548 -17528 19644 -17492
rect 18136 -17608 18232 -17592
rect 18136 -17672 18152 -17608
rect 18216 -17672 18232 -17608
rect 18136 -17688 18232 -17672
rect 18136 -17752 18152 -17688
rect 18216 -17752 18232 -17688
rect 18136 -17768 18232 -17752
rect 18136 -17832 18152 -17768
rect 18216 -17832 18232 -17768
rect 18136 -17848 18232 -17832
rect 18136 -17912 18152 -17848
rect 18216 -17912 18232 -17848
rect 18136 -17928 18232 -17912
rect 18136 -17992 18152 -17928
rect 18216 -17992 18232 -17928
rect 18136 -18008 18232 -17992
rect 18136 -18072 18152 -18008
rect 18216 -18072 18232 -18008
rect 18136 -18088 18232 -18072
rect 18136 -18152 18152 -18088
rect 18216 -18152 18232 -18088
rect 18136 -18168 18232 -18152
rect 18136 -18232 18152 -18168
rect 18216 -18232 18232 -18168
rect 18136 -18248 18232 -18232
rect 16724 -18348 16820 -18312
rect 18136 -18312 18152 -18248
rect 18216 -18312 18232 -18248
rect 18555 -17568 19277 -17559
rect 18555 -18272 18564 -17568
rect 19268 -18272 19277 -17568
rect 18555 -18281 19277 -18272
rect 19548 -17592 19564 -17528
rect 19628 -17592 19644 -17528
rect 20960 -17528 21056 -17492
rect 19548 -17608 19644 -17592
rect 19548 -17672 19564 -17608
rect 19628 -17672 19644 -17608
rect 19548 -17688 19644 -17672
rect 19548 -17752 19564 -17688
rect 19628 -17752 19644 -17688
rect 19548 -17768 19644 -17752
rect 19548 -17832 19564 -17768
rect 19628 -17832 19644 -17768
rect 19548 -17848 19644 -17832
rect 19548 -17912 19564 -17848
rect 19628 -17912 19644 -17848
rect 19548 -17928 19644 -17912
rect 19548 -17992 19564 -17928
rect 19628 -17992 19644 -17928
rect 19548 -18008 19644 -17992
rect 19548 -18072 19564 -18008
rect 19628 -18072 19644 -18008
rect 19548 -18088 19644 -18072
rect 19548 -18152 19564 -18088
rect 19628 -18152 19644 -18088
rect 19548 -18168 19644 -18152
rect 19548 -18232 19564 -18168
rect 19628 -18232 19644 -18168
rect 19548 -18248 19644 -18232
rect 18136 -18348 18232 -18312
rect 19548 -18312 19564 -18248
rect 19628 -18312 19644 -18248
rect 19967 -17568 20689 -17559
rect 19967 -18272 19976 -17568
rect 20680 -18272 20689 -17568
rect 19967 -18281 20689 -18272
rect 20960 -17592 20976 -17528
rect 21040 -17592 21056 -17528
rect 22372 -17528 22468 -17492
rect 20960 -17608 21056 -17592
rect 20960 -17672 20976 -17608
rect 21040 -17672 21056 -17608
rect 20960 -17688 21056 -17672
rect 20960 -17752 20976 -17688
rect 21040 -17752 21056 -17688
rect 20960 -17768 21056 -17752
rect 20960 -17832 20976 -17768
rect 21040 -17832 21056 -17768
rect 20960 -17848 21056 -17832
rect 20960 -17912 20976 -17848
rect 21040 -17912 21056 -17848
rect 20960 -17928 21056 -17912
rect 20960 -17992 20976 -17928
rect 21040 -17992 21056 -17928
rect 20960 -18008 21056 -17992
rect 20960 -18072 20976 -18008
rect 21040 -18072 21056 -18008
rect 20960 -18088 21056 -18072
rect 20960 -18152 20976 -18088
rect 21040 -18152 21056 -18088
rect 20960 -18168 21056 -18152
rect 20960 -18232 20976 -18168
rect 21040 -18232 21056 -18168
rect 20960 -18248 21056 -18232
rect 19548 -18348 19644 -18312
rect 20960 -18312 20976 -18248
rect 21040 -18312 21056 -18248
rect 21379 -17568 22101 -17559
rect 21379 -18272 21388 -17568
rect 22092 -18272 22101 -17568
rect 21379 -18281 22101 -18272
rect 22372 -17592 22388 -17528
rect 22452 -17592 22468 -17528
rect 23784 -17528 23880 -17492
rect 22372 -17608 22468 -17592
rect 22372 -17672 22388 -17608
rect 22452 -17672 22468 -17608
rect 22372 -17688 22468 -17672
rect 22372 -17752 22388 -17688
rect 22452 -17752 22468 -17688
rect 22372 -17768 22468 -17752
rect 22372 -17832 22388 -17768
rect 22452 -17832 22468 -17768
rect 22372 -17848 22468 -17832
rect 22372 -17912 22388 -17848
rect 22452 -17912 22468 -17848
rect 22372 -17928 22468 -17912
rect 22372 -17992 22388 -17928
rect 22452 -17992 22468 -17928
rect 22372 -18008 22468 -17992
rect 22372 -18072 22388 -18008
rect 22452 -18072 22468 -18008
rect 22372 -18088 22468 -18072
rect 22372 -18152 22388 -18088
rect 22452 -18152 22468 -18088
rect 22372 -18168 22468 -18152
rect 22372 -18232 22388 -18168
rect 22452 -18232 22468 -18168
rect 22372 -18248 22468 -18232
rect 20960 -18348 21056 -18312
rect 22372 -18312 22388 -18248
rect 22452 -18312 22468 -18248
rect 22791 -17568 23513 -17559
rect 22791 -18272 22800 -17568
rect 23504 -18272 23513 -17568
rect 22791 -18281 23513 -18272
rect 23784 -17592 23800 -17528
rect 23864 -17592 23880 -17528
rect 23784 -17608 23880 -17592
rect 23784 -17672 23800 -17608
rect 23864 -17672 23880 -17608
rect 23784 -17688 23880 -17672
rect 23784 -17752 23800 -17688
rect 23864 -17752 23880 -17688
rect 23784 -17768 23880 -17752
rect 23784 -17832 23800 -17768
rect 23864 -17832 23880 -17768
rect 23784 -17848 23880 -17832
rect 23784 -17912 23800 -17848
rect 23864 -17912 23880 -17848
rect 23784 -17928 23880 -17912
rect 23784 -17992 23800 -17928
rect 23864 -17992 23880 -17928
rect 23784 -18008 23880 -17992
rect 23784 -18072 23800 -18008
rect 23864 -18072 23880 -18008
rect 23784 -18088 23880 -18072
rect 23784 -18152 23800 -18088
rect 23864 -18152 23880 -18088
rect 23784 -18168 23880 -18152
rect 23784 -18232 23800 -18168
rect 23864 -18232 23880 -18168
rect 23784 -18248 23880 -18232
rect 22372 -18348 22468 -18312
rect 23784 -18312 23800 -18248
rect 23864 -18312 23880 -18248
rect 23784 -18348 23880 -18312
<< properties >>
string FIXED_BBOX 22712 17480 23592 18360
<< end >>
