magic
tech sky130A
magscale 1 2
timestamp 1757830127
<< metal1 >>
rect -32202 -960 -32192 -864
rect -32096 -960 -31492 -864
rect -31412 -960 -31180 -864
rect -31084 -960 -31074 -864
rect -32202 -3120 -32192 -3024
rect -32096 -3120 -31652 -3024
rect -31572 -3120 -31180 -3024
rect -31084 -3120 -31074 -3024
rect -32202 -3840 -32192 -3744
rect -32096 -3840 -31812 -3744
rect -31732 -3840 -31180 -3744
rect -31084 -3840 -31074 -3744
rect -32834 -4668 -32824 -4572
rect -32744 -4668 -32192 -4572
rect -32096 -4668 -32086 -4572
rect -32514 -5028 -32504 -4932
rect -32424 -5028 -31180 -4932
rect -31084 -5028 -31074 -4932
rect -32674 -5388 -32664 -5292
rect -32584 -5388 -31180 -5292
rect -31084 -5388 -31074 -5292
rect -32514 -5748 -32504 -5652
rect -32424 -5748 -32192 -5652
rect -32096 -5748 -32086 -5652
rect -32202 -6000 -32192 -5904
rect -32096 -6000 -31812 -5904
rect -31732 -6000 -31180 -5904
rect -31084 -6000 -31074 -5904
rect -32202 -7440 -32192 -7344
rect -32096 -7440 -31652 -7344
rect -31572 -7440 -31180 -7344
rect -31084 -7440 -31074 -7344
rect -32202 -9600 -32192 -9504
rect -32096 -9600 -31492 -9504
rect -31412 -9600 -31180 -9504
rect -31084 -9600 -31074 -9504
rect -63568 -11336 -48388 -11232
rect -48284 -11336 -14992 -11232
rect -14888 -11336 292 -11232
rect -63568 -11544 -40292 -11440
rect -40188 -11544 -23088 -11440
rect -22984 -11544 292 -11440
rect -63568 -11752 -36244 -11648
rect -36140 -11752 -27136 -11648
rect -27032 -11752 292 -11648
rect -63568 -11960 -34220 -11856
rect -34116 -11960 -29160 -11856
rect -29056 -11960 292 -11856
rect -63568 -12168 -33208 -12064
rect -33104 -12168 -30172 -12064
rect -30068 -12168 292 -12064
rect -63568 -12376 -31492 -12272
rect -31412 -12376 292 -12272
rect -63568 -12584 -31652 -12480
rect -31572 -12584 292 -12480
rect -63568 -12792 -31812 -12688
rect -31732 -12792 292 -12688
rect -63568 -13000 -32504 -12896
rect -32424 -13000 292 -12896
rect -63568 -13208 -32664 -13104
rect -32584 -13208 292 -13104
rect -63568 -13416 -32824 -13312
rect -32744 -13416 292 -13312
<< via1 >>
rect -32192 -960 -32096 -864
rect -31492 -960 -31412 -864
rect -31180 -960 -31084 -864
rect -32192 -3120 -32096 -3024
rect -31652 -3120 -31572 -3024
rect -31180 -3120 -31084 -3024
rect -32192 -3840 -32096 -3744
rect -31812 -3840 -31732 -3744
rect -31180 -3840 -31084 -3744
rect -32824 -4668 -32744 -4572
rect -32192 -4668 -32096 -4572
rect -32504 -5028 -32424 -4932
rect -31180 -5028 -31084 -4932
rect -32664 -5388 -32584 -5292
rect -31180 -5388 -31084 -5292
rect -32504 -5748 -32424 -5652
rect -32192 -5748 -32096 -5652
rect -32192 -6000 -32096 -5904
rect -31812 -6000 -31732 -5904
rect -31180 -6000 -31084 -5904
rect -32192 -7440 -32096 -7344
rect -31652 -7440 -31572 -7344
rect -31180 -7440 -31084 -7344
rect -32192 -9600 -32096 -9504
rect -31492 -9600 -31412 -9504
rect -31180 -9600 -31084 -9504
rect -48388 -11336 -48284 -11232
rect -14992 -11336 -14888 -11232
rect -40292 -11544 -40188 -11440
rect -23088 -11544 -22984 -11440
rect -36244 -11752 -36140 -11648
rect -27136 -11752 -27032 -11648
rect -34220 -11960 -34116 -11856
rect -29160 -11960 -29056 -11856
rect -33208 -12168 -33104 -12064
rect -30172 -12168 -30068 -12064
rect -31492 -12376 -31412 -12272
rect -31652 -12584 -31572 -12480
rect -31812 -12792 -31732 -12688
rect -32504 -13000 -32424 -12896
rect -32664 -13208 -32584 -13104
rect -32824 -13416 -32744 -13312
<< metal2 >>
rect -32192 -864 -32096 -854
rect -32192 -970 -32096 -960
rect -31492 -864 -31412 -858
rect -32192 -3024 -32096 -3014
rect -32192 -3130 -32096 -3120
rect -31652 -3024 -31572 -3018
rect -32192 -3744 -32096 -3734
rect -32192 -3850 -32096 -3840
rect -31812 -3744 -31732 -3738
rect -32824 -4572 -32744 -4566
rect -48388 -11232 -48284 -11222
rect -48388 -11346 -48284 -11336
rect -40292 -11440 -40188 -11430
rect -40292 -11554 -40188 -11544
rect -36244 -11648 -36140 -11638
rect -36244 -11762 -36140 -11752
rect -34220 -11856 -34116 -11846
rect -34220 -11970 -34116 -11960
rect -33208 -12064 -33104 -12054
rect -33208 -12178 -33104 -12168
rect -32824 -13312 -32744 -4668
rect -32192 -4572 -32096 -4562
rect -32192 -4678 -32096 -4668
rect -32504 -4932 -32424 -4926
rect -32664 -5292 -32584 -5286
rect -32664 -13104 -32584 -5388
rect -32504 -5652 -32424 -5028
rect -32504 -12896 -32424 -5748
rect -32192 -5652 -32096 -5642
rect -32192 -5758 -32096 -5748
rect -32192 -5904 -32096 -5894
rect -32192 -6010 -32096 -6000
rect -31812 -5904 -31732 -3840
rect -32192 -7344 -32096 -7334
rect -32192 -7450 -32096 -7440
rect -32192 -9504 -32096 -9494
rect -32192 -9610 -32096 -9600
rect -31812 -12688 -31732 -6000
rect -31652 -7344 -31572 -3120
rect -31652 -12480 -31572 -7440
rect -31492 -9504 -31412 -960
rect -31180 -864 -31084 -854
rect -31180 -970 -31084 -960
rect -31180 -3024 -31084 -3014
rect -31180 -3130 -31084 -3120
rect -31180 -3744 -31084 -3734
rect -31180 -3850 -31084 -3840
rect -31180 -4932 -31084 -4922
rect -31180 -5038 -31084 -5028
rect -31180 -5292 -31084 -5282
rect -31180 -5398 -31084 -5388
rect -31180 -5904 -31084 -5894
rect -31180 -6010 -31084 -6000
rect -31180 -7344 -31084 -7334
rect -31180 -7450 -31084 -7440
rect -31492 -12272 -31412 -9600
rect -31180 -9504 -31084 -9494
rect -31180 -9610 -31084 -9600
rect -14992 -11232 -14888 -11222
rect -14992 -11346 -14888 -11336
rect -23088 -11440 -22984 -11430
rect -23088 -11554 -22984 -11544
rect -27136 -11648 -27032 -11638
rect -27136 -11762 -27032 -11752
rect -29160 -11856 -29056 -11846
rect -29160 -11970 -29056 -11960
rect -30172 -12064 -30068 -12054
rect -30172 -12178 -30068 -12168
rect -31492 -12386 -31412 -12376
rect -31652 -12594 -31572 -12584
rect -31812 -12802 -31732 -12792
rect -32504 -13010 -32424 -13000
rect -32664 -13218 -32584 -13208
rect -32824 -13426 -32744 -13416
<< via2 >>
rect -32192 -960 -32096 -864
rect -32192 -3120 -32096 -3024
rect -32192 -3840 -32096 -3744
rect -48388 -11336 -48284 -11232
rect -40292 -11544 -40188 -11440
rect -36244 -11752 -36140 -11648
rect -34220 -11960 -34116 -11856
rect -33208 -12168 -33104 -12064
rect -32192 -4668 -32096 -4572
rect -32192 -5748 -32096 -5652
rect -32192 -6000 -32096 -5904
rect -32192 -7440 -32096 -7344
rect -32192 -9600 -32096 -9504
rect -31180 -960 -31084 -864
rect -31180 -3120 -31084 -3024
rect -31180 -3840 -31084 -3744
rect -31180 -5028 -31084 -4932
rect -31180 -5388 -31084 -5292
rect -31180 -6000 -31084 -5904
rect -31180 -7440 -31084 -7344
rect -31180 -9600 -31084 -9504
rect -14992 -11336 -14888 -11232
rect -23088 -11544 -22984 -11440
rect -27136 -11752 -27032 -11648
rect -29160 -11960 -29056 -11856
rect -30172 -12168 -30068 -12064
<< metal3 >>
rect -32202 -864 -32086 -859
rect -32202 -960 -32192 -864
rect -32096 -960 -32086 -864
rect -32202 -965 -32086 -960
rect -31190 -864 -31074 -859
rect -31190 -960 -31180 -864
rect -31084 -960 -31074 -864
rect -31190 -965 -31074 -960
rect -32202 -3024 -32086 -3019
rect -32202 -3120 -32192 -3024
rect -32096 -3120 -32086 -3024
rect -32202 -3125 -32086 -3120
rect -31190 -3024 -31074 -3019
rect -31190 -3120 -31180 -3024
rect -31084 -3120 -31074 -3024
rect -31190 -3125 -31074 -3120
rect -32202 -3744 -32086 -3739
rect -32202 -3840 -32192 -3744
rect -32096 -3840 -32086 -3744
rect -32202 -3845 -32086 -3840
rect -31190 -3744 -31074 -3739
rect -31190 -3840 -31180 -3744
rect -31084 -3840 -31074 -3744
rect -31190 -3845 -31074 -3840
rect -32202 -4572 -32086 -4567
rect -32202 -4668 -32192 -4572
rect -32096 -4668 -32086 -4572
rect -32202 -4673 -32086 -4668
rect -31190 -4932 -31074 -4927
rect -31190 -5028 -31180 -4932
rect -31084 -5028 -31074 -4932
rect -31190 -5033 -31074 -5028
rect -31190 -5292 -31074 -5287
rect -31190 -5388 -31180 -5292
rect -31084 -5388 -31074 -5292
rect -31190 -5393 -31074 -5388
rect -32202 -5652 -32086 -5647
rect -32202 -5748 -32192 -5652
rect -32096 -5748 -32086 -5652
rect -32202 -5753 -32086 -5748
rect -32202 -5904 -32086 -5899
rect -32202 -6000 -32192 -5904
rect -32096 -6000 -32086 -5904
rect -32202 -6005 -32086 -6000
rect -31190 -5904 -31074 -5899
rect -31190 -6000 -31180 -5904
rect -31084 -6000 -31074 -5904
rect -31190 -6005 -31074 -6000
rect -32202 -7344 -32086 -7339
rect -32202 -7440 -32192 -7344
rect -32096 -7440 -32086 -7344
rect -32202 -7445 -32086 -7440
rect -31190 -7344 -31074 -7339
rect -31190 -7440 -31180 -7344
rect -31084 -7440 -31074 -7344
rect -31190 -7445 -31074 -7440
rect -32202 -9504 -32086 -9499
rect -32202 -9600 -32192 -9504
rect -32096 -9600 -32086 -9504
rect -32202 -9605 -32086 -9600
rect -31190 -9504 -31074 -9499
rect -31190 -9600 -31180 -9504
rect -31084 -9600 -31074 -9504
rect -31190 -9605 -31074 -9600
rect -48398 -11232 -48274 -11227
rect -48398 -11336 -48388 -11232
rect -48284 -11336 -48274 -11232
rect -48398 -11341 -48274 -11336
rect -15002 -11232 -14878 -11227
rect -15002 -11336 -14992 -11232
rect -14888 -11336 -14878 -11232
rect -15002 -11341 -14878 -11336
rect -40302 -11440 -40178 -11435
rect -40302 -11544 -40292 -11440
rect -40188 -11544 -40178 -11440
rect -40302 -11549 -40178 -11544
rect -23098 -11440 -22974 -11435
rect -23098 -11544 -23088 -11440
rect -22984 -11544 -22974 -11440
rect -23098 -11549 -22974 -11544
rect -36254 -11648 -36130 -11643
rect -36254 -11752 -36244 -11648
rect -36140 -11752 -36130 -11648
rect -36254 -11757 -36130 -11752
rect -27146 -11648 -27022 -11643
rect -27146 -11752 -27136 -11648
rect -27032 -11752 -27022 -11648
rect -27146 -11757 -27022 -11752
rect -34230 -11856 -34106 -11851
rect -34230 -11960 -34220 -11856
rect -34116 -11960 -34106 -11856
rect -34230 -11965 -34106 -11960
rect -29170 -11856 -29046 -11851
rect -29170 -11960 -29160 -11856
rect -29056 -11960 -29046 -11856
rect -29170 -11965 -29046 -11960
rect -33218 -12064 -33094 -12059
rect -33218 -12168 -33208 -12064
rect -33104 -12168 -33094 -12064
rect -33218 -12173 -33094 -12168
rect -30182 -12064 -30058 -12059
rect -30182 -12168 -30172 -12064
rect -30068 -12168 -30058 -12064
rect -30182 -12173 -30058 -12168
<< via3 >>
rect -32192 -960 -32096 -864
rect -31180 -960 -31084 -864
rect -32192 -3120 -32096 -3024
rect -31180 -3120 -31084 -3024
rect -32192 -3840 -32096 -3744
rect -31180 -3840 -31084 -3744
rect -32192 -6000 -32096 -5904
rect -31180 -6000 -31084 -5904
rect -32192 -7440 -32096 -7344
rect -31180 -7440 -31084 -7344
rect -32192 -9600 -32096 -9504
rect -31180 -9600 -31084 -9504
rect -48388 -11336 -48284 -11232
rect -14992 -11336 -14888 -11232
rect -40292 -11544 -40188 -11440
rect -23088 -11544 -22984 -11440
rect -36244 -11752 -36140 -11648
rect -27136 -11752 -27032 -11648
rect -34220 -11960 -34116 -11856
rect -29160 -11960 -29056 -11856
rect -33208 -12168 -33104 -12064
rect -30172 -12168 -30068 -12064
<< metal4 >>
rect -64048 704 -188 808
rect -64048 600 -63944 704
rect -63036 600 -62932 704
rect -62024 600 -61920 704
rect -61012 600 -60908 704
rect -60000 600 -59896 704
rect -58988 600 -58884 704
rect -57976 600 -57872 704
rect -56964 600 -56860 704
rect -55952 600 -55848 704
rect -54940 600 -54836 704
rect -53928 600 -53824 704
rect -52916 600 -52812 704
rect -51904 600 -51800 704
rect -50892 600 -50788 704
rect -49880 600 -49776 704
rect -48868 600 -48764 704
rect -47856 600 -47752 704
rect -46844 600 -46740 704
rect -45832 600 -45728 704
rect -44820 600 -44716 704
rect -43808 600 -43704 704
rect -42796 600 -42692 704
rect -41784 600 -41680 704
rect -40772 600 -40668 704
rect -39760 600 -39656 704
rect -38748 600 -38644 704
rect -37736 600 -37632 704
rect -36724 600 -36620 704
rect -35712 600 -35608 704
rect -34700 600 -34596 704
rect -33688 600 -33584 704
rect -32676 600 -32572 704
rect -31664 600 -31560 704
rect -30652 600 -30548 704
rect -29640 600 -29536 704
rect -28628 600 -28524 704
rect -27616 600 -27512 704
rect -26604 600 -26500 704
rect -25592 600 -25488 704
rect -24580 600 -24476 704
rect -23568 600 -23464 704
rect -22556 600 -22452 704
rect -21544 600 -21440 704
rect -20532 600 -20428 704
rect -19520 600 -19416 704
rect -18508 600 -18404 704
rect -17496 600 -17392 704
rect -16484 600 -16380 704
rect -15472 600 -15368 704
rect -14460 600 -14356 704
rect -13448 600 -13344 704
rect -12436 600 -12332 704
rect -11424 600 -11320 704
rect -10412 600 -10308 704
rect -9400 600 -9296 704
rect -8388 600 -8284 704
rect -7376 600 -7272 704
rect -6364 600 -6260 704
rect -5352 600 -5248 704
rect -4340 600 -4236 704
rect -3328 600 -3224 704
rect -2316 600 -2212 704
rect -1304 600 -1200 704
rect -292 600 -188 704
rect -32192 -863 -32096 12
rect -31180 -863 -31084 12
rect -32193 -864 -32095 -863
rect -32193 -960 -32192 -864
rect -32096 -960 -32095 -864
rect -32193 -961 -32095 -960
rect -31181 -864 -31083 -863
rect -31181 -960 -31180 -864
rect -31084 -960 -31083 -864
rect -31181 -961 -31083 -960
rect -32192 -1692 -32096 -961
rect -31180 -1692 -31084 -961
rect -32192 -3023 -32096 -2868
rect -31180 -3023 -31084 -2868
rect -32193 -3024 -32095 -3023
rect -32193 -3120 -32192 -3024
rect -32096 -3120 -32095 -3024
rect -32193 -3121 -32095 -3120
rect -31181 -3024 -31083 -3023
rect -31181 -3120 -31180 -3024
rect -31084 -3120 -31083 -3024
rect -31181 -3121 -31083 -3120
rect -32192 -3132 -32096 -3121
rect -31180 -3132 -31084 -3121
rect -32193 -3744 -32095 -3743
rect -32193 -3840 -32192 -3744
rect -32096 -3840 -32095 -3744
rect -32193 -3841 -32095 -3840
rect -31181 -3744 -31083 -3743
rect -31181 -3840 -31180 -3744
rect -31084 -3840 -31083 -3744
rect -31181 -3841 -31083 -3840
rect -32192 -3854 -32096 -3841
rect -31180 -3852 -31084 -3841
rect -32193 -5904 -32095 -5903
rect -32193 -6000 -32192 -5904
rect -32096 -6000 -32095 -5904
rect -32193 -6001 -32095 -6000
rect -31181 -5904 -31083 -5903
rect -31181 -6000 -31180 -5904
rect -31084 -6000 -31083 -5904
rect -31181 -6001 -31083 -6000
rect -32192 -6012 -32096 -6001
rect -31180 -6012 -31084 -6001
rect -32192 -7343 -32096 -7188
rect -31180 -7343 -31084 -7188
rect -32193 -7344 -32095 -7343
rect -32193 -7440 -32192 -7344
rect -32096 -7440 -32095 -7344
rect -32193 -7441 -32095 -7440
rect -31181 -7344 -31083 -7343
rect -31181 -7440 -31180 -7344
rect -31084 -7440 -31083 -7344
rect -31181 -7441 -31083 -7440
rect -32192 -7452 -32096 -7441
rect -31180 -7452 -31084 -7441
rect -32192 -9503 -32096 -8628
rect -31180 -9503 -31084 -8628
rect -32193 -9504 -32095 -9503
rect -32193 -9600 -32192 -9504
rect -32096 -9600 -32095 -9504
rect -32193 -9601 -32095 -9600
rect -31181 -9504 -31083 -9503
rect -31181 -9600 -31180 -9504
rect -31084 -9600 -31083 -9504
rect -31181 -9601 -31083 -9600
rect -32192 -10332 -32096 -9601
rect -31180 -10332 -31084 -9601
rect -63568 -11024 -63464 -10920
rect -62556 -11024 -62452 -10920
rect -61544 -11024 -61440 -10920
rect -60532 -11024 -60428 -10920
rect -59520 -11024 -59416 -10920
rect -58508 -11024 -58404 -10920
rect -57496 -11024 -57392 -10920
rect -56484 -11024 -56380 -10920
rect -55472 -11024 -55368 -10920
rect -54460 -11024 -54356 -10920
rect -53448 -11024 -53344 -10920
rect -52436 -11024 -52332 -10920
rect -51424 -11024 -51320 -10920
rect -50412 -11024 -50308 -10920
rect -49400 -11024 -49296 -10920
rect -48388 -11024 -48284 -10920
rect -63568 -11128 -48284 -11024
rect -47376 -11024 -47272 -10920
rect -46364 -11024 -46260 -10920
rect -45352 -11024 -45248 -10920
rect -44340 -11024 -44236 -10920
rect -43328 -11024 -43224 -10920
rect -42316 -11024 -42212 -10920
rect -41304 -11024 -41200 -10920
rect -40292 -11024 -40188 -10920
rect -47376 -11128 -40188 -11024
rect -39280 -11024 -39176 -10920
rect -38268 -11024 -38164 -10920
rect -37256 -11024 -37152 -10920
rect -36244 -11024 -36140 -10920
rect -39280 -11128 -36140 -11024
rect -35232 -11024 -35128 -10920
rect -34220 -11024 -34116 -10920
rect -35232 -11128 -34116 -11024
rect -48388 -11231 -48284 -11128
rect -48389 -11232 -48283 -11231
rect -48389 -11336 -48388 -11232
rect -48284 -11336 -48283 -11232
rect -48389 -11337 -48283 -11336
rect -40292 -11439 -40188 -11128
rect -40293 -11440 -40187 -11439
rect -40293 -11544 -40292 -11440
rect -40188 -11544 -40187 -11440
rect -40293 -11545 -40187 -11544
rect -36244 -11647 -36140 -11128
rect -36245 -11648 -36139 -11647
rect -36245 -11752 -36244 -11648
rect -36140 -11752 -36139 -11648
rect -36245 -11753 -36139 -11752
rect -34220 -11855 -34116 -11128
rect -34221 -11856 -34115 -11855
rect -34221 -11960 -34220 -11856
rect -34116 -11960 -34115 -11856
rect -34221 -11961 -34115 -11960
rect -33208 -12063 -33104 -10920
rect -30172 -12063 -30068 -10920
rect -29160 -11024 -29056 -10920
rect -28148 -11024 -28044 -10816
rect -29160 -11128 -28044 -11024
rect -27136 -11024 -27032 -10920
rect -26124 -11024 -26020 -10816
rect -25112 -11024 -25008 -10810
rect -24100 -11024 -23996 -10816
rect -27136 -11128 -23996 -11024
rect -23088 -11024 -22984 -10920
rect -22076 -11024 -21972 -10816
rect -21064 -11024 -20960 -10816
rect -20052 -11024 -19948 -10811
rect -19040 -11024 -18936 -10816
rect -18028 -11024 -17924 -10811
rect -17016 -11024 -16912 -10816
rect -16004 -11024 -15900 -10816
rect -23088 -11128 -15900 -11024
rect -14992 -11024 -14888 -10920
rect -13980 -11024 -13876 -10812
rect -12968 -11024 -12864 -10815
rect -11956 -11024 -11852 -10816
rect -10944 -11024 -10840 -10816
rect -9932 -11024 -9828 -10816
rect -8920 -11024 -8816 -10816
rect -7908 -11024 -7804 -10816
rect -6896 -11024 -6792 -10816
rect -5884 -11024 -5780 -10816
rect -4872 -11024 -4768 -10807
rect -3860 -11024 -3756 -10816
rect -2848 -11024 -2744 -10807
rect -1836 -11024 -1732 -10805
rect -824 -11024 -720 -10815
rect 188 -11024 292 -10816
rect -14992 -11128 292 -11024
rect -29160 -11855 -29056 -11128
rect -27136 -11647 -27032 -11128
rect -23088 -11439 -22984 -11128
rect -14992 -11231 -14888 -11128
rect -14993 -11232 -14887 -11231
rect -14993 -11336 -14992 -11232
rect -14888 -11336 -14887 -11232
rect -14993 -11337 -14887 -11336
rect -23089 -11440 -22983 -11439
rect -23089 -11544 -23088 -11440
rect -22984 -11544 -22983 -11440
rect -23089 -11545 -22983 -11544
rect -27137 -11648 -27031 -11647
rect -27137 -11752 -27136 -11648
rect -27032 -11752 -27031 -11648
rect -27137 -11753 -27031 -11752
rect -29161 -11856 -29055 -11855
rect -29161 -11960 -29160 -11856
rect -29056 -11960 -29055 -11856
rect -29161 -11961 -29055 -11960
rect -33209 -12064 -33103 -12063
rect -33209 -12168 -33208 -12064
rect -33104 -12168 -33103 -12064
rect -33209 -12169 -33103 -12168
rect -30173 -12064 -30067 -12063
rect -30173 -12168 -30172 -12064
rect -30068 -12168 -30067 -12064
rect -30173 -12169 -30067 -12168
use sky130_fd_pr__cap_mim_m3_1_NLQ4WR  sky130_fd_pr__cap_mim_m3_1_NLQ4WR_0
timestamp 1757810374
transform 1 0 -31972 0 1 -5160
box -892 -5760 892 5760
use sky130_fd_pr__cap_mim_m3_1_TE2AE4  sky130_fd_pr__cap_mim_m3_1_TE2AE4_0
timestamp 1757383169
transform 1 0 -15274 0 1 -5160
box -15566 -5760 15566 5760
use sky130_fd_pr__cap_mim_m3_1_TE2AE4  sky130_fd_pr__cap_mim_m3_1_TE2AE4_1
timestamp 1757383169
transform 1 0 -48670 0 1 -5160
box -15566 -5760 15566 5760
<< labels >>
flabel metal1 188 -13416 292 -13312 0 FreeSans 320 0 0 0 VCM
port 10 nsew
flabel metal4 -414 704 -310 808 0 FreeSans 320 0 0 0 VC
port 12 nsew
flabel metal1 188 -13208 292 -13104 0 FreeSans 320 0 0 0 S[9]
port 0 nsew
flabel metal1 188 -13000 292 -12896 0 FreeSans 320 0 0 0 S[8]
port 1 nsew
flabel metal1 188 -12792 292 -12688 0 FreeSans 320 0 0 0 S[7]
port 2 nsew
flabel metal1 188 -12584 292 -12480 0 FreeSans 320 0 0 0 S[6]
port 3 nsew
flabel metal1 188 -12376 292 -12272 0 FreeSans 320 0 0 0 S[5]
port 4 nsew
flabel metal1 188 -12168 292 -12064 0 FreeSans 320 0 0 0 S[4]
port 5 nsew
flabel metal1 188 -11960 292 -11856 0 FreeSans 320 0 0 0 S[3]
port 6 nsew
flabel metal1 188 -11752 292 -11648 0 FreeSans 320 0 0 0 S[2]
port 7 nsew
flabel metal1 188 -11544 292 -11440 0 FreeSans 320 0 0 0 S[1]
port 8 nsew
flabel metal1 188 -11336 292 -11232 0 FreeSans 320 0 0 0 S[0]
port 9 nsew
<< end >>
