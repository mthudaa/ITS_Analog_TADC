magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< metal3 >>
rect -2704 2092 -1532 2120
rect -2704 1268 -1616 2092
rect -1552 1268 -1532 2092
rect -2704 1240 -1532 1268
rect -1292 2092 -120 2120
rect -1292 1268 -204 2092
rect -140 1268 -120 2092
rect -1292 1240 -120 1268
rect 120 2092 1292 2120
rect 120 1268 1208 2092
rect 1272 1268 1292 2092
rect 120 1240 1292 1268
rect 1532 2092 2704 2120
rect 1532 1268 2620 2092
rect 2684 1268 2704 2092
rect 1532 1240 2704 1268
rect -2704 972 -1532 1000
rect -2704 148 -1616 972
rect -1552 148 -1532 972
rect -2704 120 -1532 148
rect -1292 972 -120 1000
rect -1292 148 -204 972
rect -140 148 -120 972
rect -1292 120 -120 148
rect 120 972 1292 1000
rect 120 148 1208 972
rect 1272 148 1292 972
rect 120 120 1292 148
rect 1532 972 2704 1000
rect 1532 148 2620 972
rect 2684 148 2704 972
rect 1532 120 2704 148
rect -2704 -148 -1532 -120
rect -2704 -972 -1616 -148
rect -1552 -972 -1532 -148
rect -2704 -1000 -1532 -972
rect -1292 -148 -120 -120
rect -1292 -972 -204 -148
rect -140 -972 -120 -148
rect -1292 -1000 -120 -972
rect 120 -148 1292 -120
rect 120 -972 1208 -148
rect 1272 -972 1292 -148
rect 120 -1000 1292 -972
rect 1532 -148 2704 -120
rect 1532 -972 2620 -148
rect 2684 -972 2704 -148
rect 1532 -1000 2704 -972
rect -2704 -1268 -1532 -1240
rect -2704 -2092 -1616 -1268
rect -1552 -2092 -1532 -1268
rect -2704 -2120 -1532 -2092
rect -1292 -1268 -120 -1240
rect -1292 -2092 -204 -1268
rect -140 -2092 -120 -1268
rect -1292 -2120 -120 -2092
rect 120 -1268 1292 -1240
rect 120 -2092 1208 -1268
rect 1272 -2092 1292 -1268
rect 120 -2120 1292 -2092
rect 1532 -1268 2704 -1240
rect 1532 -2092 2620 -1268
rect 2684 -2092 2704 -1268
rect 1532 -2120 2704 -2092
<< via3 >>
rect -1616 1268 -1552 2092
rect -204 1268 -140 2092
rect 1208 1268 1272 2092
rect 2620 1268 2684 2092
rect -1616 148 -1552 972
rect -204 148 -140 972
rect 1208 148 1272 972
rect 2620 148 2684 972
rect -1616 -972 -1552 -148
rect -204 -972 -140 -148
rect 1208 -972 1272 -148
rect 2620 -972 2684 -148
rect -1616 -2092 -1552 -1268
rect -204 -2092 -140 -1268
rect 1208 -2092 1272 -1268
rect 2620 -2092 2684 -1268
<< mimcap >>
rect -2664 2040 -1864 2080
rect -2664 1320 -2624 2040
rect -1904 1320 -1864 2040
rect -2664 1280 -1864 1320
rect -1252 2040 -452 2080
rect -1252 1320 -1212 2040
rect -492 1320 -452 2040
rect -1252 1280 -452 1320
rect 160 2040 960 2080
rect 160 1320 200 2040
rect 920 1320 960 2040
rect 160 1280 960 1320
rect 1572 2040 2372 2080
rect 1572 1320 1612 2040
rect 2332 1320 2372 2040
rect 1572 1280 2372 1320
rect -2664 920 -1864 960
rect -2664 200 -2624 920
rect -1904 200 -1864 920
rect -2664 160 -1864 200
rect -1252 920 -452 960
rect -1252 200 -1212 920
rect -492 200 -452 920
rect -1252 160 -452 200
rect 160 920 960 960
rect 160 200 200 920
rect 920 200 960 920
rect 160 160 960 200
rect 1572 920 2372 960
rect 1572 200 1612 920
rect 2332 200 2372 920
rect 1572 160 2372 200
rect -2664 -200 -1864 -160
rect -2664 -920 -2624 -200
rect -1904 -920 -1864 -200
rect -2664 -960 -1864 -920
rect -1252 -200 -452 -160
rect -1252 -920 -1212 -200
rect -492 -920 -452 -200
rect -1252 -960 -452 -920
rect 160 -200 960 -160
rect 160 -920 200 -200
rect 920 -920 960 -200
rect 160 -960 960 -920
rect 1572 -200 2372 -160
rect 1572 -920 1612 -200
rect 2332 -920 2372 -200
rect 1572 -960 2372 -920
rect -2664 -1320 -1864 -1280
rect -2664 -2040 -2624 -1320
rect -1904 -2040 -1864 -1320
rect -2664 -2080 -1864 -2040
rect -1252 -1320 -452 -1280
rect -1252 -2040 -1212 -1320
rect -492 -2040 -452 -1320
rect -1252 -2080 -452 -2040
rect 160 -1320 960 -1280
rect 160 -2040 200 -1320
rect 920 -2040 960 -1320
rect 160 -2080 960 -2040
rect 1572 -1320 2372 -1280
rect 1572 -2040 1612 -1320
rect 2332 -2040 2372 -1320
rect 1572 -2080 2372 -2040
<< mimcapcontact >>
rect -2624 1320 -1904 2040
rect -1212 1320 -492 2040
rect 200 1320 920 2040
rect 1612 1320 2332 2040
rect -2624 200 -1904 920
rect -1212 200 -492 920
rect 200 200 920 920
rect 1612 200 2332 920
rect -2624 -920 -1904 -200
rect -1212 -920 -492 -200
rect 200 -920 920 -200
rect 1612 -920 2332 -200
rect -2624 -2040 -1904 -1320
rect -1212 -2040 -492 -1320
rect 200 -2040 920 -1320
rect 1612 -2040 2332 -1320
<< metal4 >>
rect -2316 2041 -2212 2240
rect -1636 2092 -1532 2240
rect -2625 2040 -1903 2041
rect -2625 1320 -2624 2040
rect -1904 1320 -1903 2040
rect -2625 1319 -1903 1320
rect -2316 921 -2212 1319
rect -1636 1268 -1616 2092
rect -1552 1268 -1532 2092
rect -904 2041 -800 2240
rect -224 2092 -120 2240
rect -1213 2040 -491 2041
rect -1213 1320 -1212 2040
rect -492 1320 -491 2040
rect -1213 1319 -491 1320
rect -1636 972 -1532 1268
rect -2625 920 -1903 921
rect -2625 200 -2624 920
rect -1904 200 -1903 920
rect -2625 199 -1903 200
rect -2316 -199 -2212 199
rect -1636 148 -1616 972
rect -1552 148 -1532 972
rect -904 921 -800 1319
rect -224 1268 -204 2092
rect -140 1268 -120 2092
rect 508 2041 612 2240
rect 1188 2092 1292 2240
rect 199 2040 921 2041
rect 199 1320 200 2040
rect 920 1320 921 2040
rect 199 1319 921 1320
rect -224 972 -120 1268
rect -1213 920 -491 921
rect -1213 200 -1212 920
rect -492 200 -491 920
rect -1213 199 -491 200
rect -1636 -148 -1532 148
rect -2625 -200 -1903 -199
rect -2625 -920 -2624 -200
rect -1904 -920 -1903 -200
rect -2625 -921 -1903 -920
rect -2316 -1319 -2212 -921
rect -1636 -972 -1616 -148
rect -1552 -972 -1532 -148
rect -904 -199 -800 199
rect -224 148 -204 972
rect -140 148 -120 972
rect 508 921 612 1319
rect 1188 1268 1208 2092
rect 1272 1268 1292 2092
rect 1920 2041 2024 2240
rect 2600 2092 2704 2240
rect 1611 2040 2333 2041
rect 1611 1320 1612 2040
rect 2332 1320 2333 2040
rect 1611 1319 2333 1320
rect 1188 972 1292 1268
rect 199 920 921 921
rect 199 200 200 920
rect 920 200 921 920
rect 199 199 921 200
rect -224 -148 -120 148
rect -1213 -200 -491 -199
rect -1213 -920 -1212 -200
rect -492 -920 -491 -200
rect -1213 -921 -491 -920
rect -1636 -1268 -1532 -972
rect -2625 -1320 -1903 -1319
rect -2625 -2040 -2624 -1320
rect -1904 -2040 -1903 -1320
rect -2625 -2041 -1903 -2040
rect -2316 -2240 -2212 -2041
rect -1636 -2092 -1616 -1268
rect -1552 -2092 -1532 -1268
rect -904 -1319 -800 -921
rect -224 -972 -204 -148
rect -140 -972 -120 -148
rect 508 -199 612 199
rect 1188 148 1208 972
rect 1272 148 1292 972
rect 1920 921 2024 1319
rect 2600 1268 2620 2092
rect 2684 1268 2704 2092
rect 2600 972 2704 1268
rect 1611 920 2333 921
rect 1611 200 1612 920
rect 2332 200 2333 920
rect 1611 199 2333 200
rect 1188 -148 1292 148
rect 199 -200 921 -199
rect 199 -920 200 -200
rect 920 -920 921 -200
rect 199 -921 921 -920
rect -224 -1268 -120 -972
rect -1213 -1320 -491 -1319
rect -1213 -2040 -1212 -1320
rect -492 -2040 -491 -1320
rect -1213 -2041 -491 -2040
rect -1636 -2240 -1532 -2092
rect -904 -2240 -800 -2041
rect -224 -2092 -204 -1268
rect -140 -2092 -120 -1268
rect 508 -1319 612 -921
rect 1188 -972 1208 -148
rect 1272 -972 1292 -148
rect 1920 -199 2024 199
rect 2600 148 2620 972
rect 2684 148 2704 972
rect 2600 -148 2704 148
rect 1611 -200 2333 -199
rect 1611 -920 1612 -200
rect 2332 -920 2333 -200
rect 1611 -921 2333 -920
rect 1188 -1268 1292 -972
rect 199 -1320 921 -1319
rect 199 -2040 200 -1320
rect 920 -2040 921 -1320
rect 199 -2041 921 -2040
rect -224 -2240 -120 -2092
rect 508 -2240 612 -2041
rect 1188 -2092 1208 -1268
rect 1272 -2092 1292 -1268
rect 1920 -1319 2024 -921
rect 2600 -972 2620 -148
rect 2684 -972 2704 -148
rect 2600 -1268 2704 -972
rect 1611 -1320 2333 -1319
rect 1611 -2040 1612 -1320
rect 2332 -2040 2333 -1320
rect 1611 -2041 2333 -2040
rect 1188 -2240 1292 -2092
rect 1920 -2240 2024 -2041
rect 2600 -2092 2620 -1268
rect 2684 -2092 2704 -1268
rect 2600 -2240 2704 -2092
<< properties >>
string FIXED_BBOX 1532 1240 2412 2120
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
