magic
tech sky130A
magscale 1 2
timestamp 1757961500
<< metal1 >>
rect -9429 2654 -9419 2750
rect -9323 2654 -9313 2750
rect -32230 -960 -32220 -864
rect -32124 -960 -31492 -864
rect -31412 -960 -30808 -864
rect -30712 -960 -30702 -864
rect -32230 -3120 -32220 -3024
rect -32124 -3120 -31652 -3024
rect -31572 -3120 -30808 -3024
rect -30712 -3120 -30702 -3024
rect -32230 -3840 -32220 -3744
rect -32124 -3840 -31812 -3744
rect -31732 -3840 -30808 -3744
rect -30712 -3840 -30702 -3744
rect -33234 -4668 -33224 -4572
rect -33144 -4668 -32220 -4572
rect -32124 -4668 -32114 -4572
rect -32914 -5028 -32904 -4932
rect -32824 -5028 -30808 -4932
rect -30712 -5028 -30702 -4932
rect -33074 -5388 -33064 -5292
rect -32984 -5388 -30808 -5292
rect -30712 -5388 -30702 -5292
rect -32914 -5748 -32904 -5652
rect -32824 -5748 -32220 -5652
rect -32124 -5748 -32114 -5652
rect -32230 -6000 -32220 -5904
rect -32124 -6000 -31812 -5904
rect -31732 -6000 -30808 -5904
rect -30712 -6000 -30702 -5904
rect -32230 -7440 -32220 -7344
rect -32124 -7440 -31652 -7344
rect -31572 -7440 -30808 -7344
rect -30712 -7440 -30702 -7344
rect -32230 -9600 -32220 -9504
rect -32124 -9600 -31492 -9504
rect -31412 -9600 -30808 -9504
rect -30712 -9600 -30702 -9504
rect -48444 -11304 -40692 -11200
rect -40588 -11304 -22688 -11200
rect -22584 -11304 -15500 -11200
rect -48444 -11512 -36644 -11408
rect -36540 -11512 -26736 -11408
rect -26632 -11512 -15500 -11408
rect -48444 -11720 -34620 -11616
rect -34516 -11720 -28760 -11616
rect -28656 -11720 -15500 -11616
rect -48444 -11928 -33608 -11824
rect -33504 -11928 -29772 -11824
rect -29668 -11928 -15500 -11824
rect -48444 -12136 -31492 -12032
rect -31412 -12136 -15500 -12032
rect -48444 -12344 -31652 -12240
rect -31572 -12344 -15500 -12240
rect -48444 -12552 -31812 -12448
rect -31732 -12552 -15500 -12448
rect -48444 -12760 -32904 -12656
rect -32824 -12760 -15500 -12656
rect -48444 -12968 -33064 -12864
rect -32984 -12968 -15500 -12864
rect -48444 -13176 -33224 -13072
rect -33144 -13176 -15500 -13072
<< via1 >>
rect -9419 2654 -9323 2750
rect -32220 -960 -32124 -864
rect -31492 -960 -31412 -864
rect -30808 -960 -30712 -864
rect -32220 -3120 -32124 -3024
rect -31652 -3120 -31572 -3024
rect -30808 -3120 -30712 -3024
rect -32220 -3840 -32124 -3744
rect -31812 -3840 -31732 -3744
rect -30808 -3840 -30712 -3744
rect -33224 -4668 -33144 -4572
rect -32220 -4668 -32124 -4572
rect -32904 -5028 -32824 -4932
rect -30808 -5028 -30712 -4932
rect -33064 -5388 -32984 -5292
rect -30808 -5388 -30712 -5292
rect -32904 -5748 -32824 -5652
rect -32220 -5748 -32124 -5652
rect -32220 -6000 -32124 -5904
rect -31812 -6000 -31732 -5904
rect -30808 -6000 -30712 -5904
rect -32220 -7440 -32124 -7344
rect -31652 -7440 -31572 -7344
rect -30808 -7440 -30712 -7344
rect -32220 -9600 -32124 -9504
rect -31492 -9600 -31412 -9504
rect -30808 -9600 -30712 -9504
rect -40692 -11304 -40588 -11200
rect -22688 -11304 -22584 -11200
rect -36644 -11512 -36540 -11408
rect -26736 -11512 -26632 -11408
rect -34620 -11720 -34516 -11616
rect -28760 -11720 -28656 -11616
rect -33608 -11928 -33504 -11824
rect -29772 -11928 -29668 -11824
rect -31492 -12136 -31412 -12032
rect -31652 -12344 -31572 -12240
rect -31812 -12552 -31732 -12448
rect -32904 -12760 -32824 -12656
rect -33064 -12968 -32984 -12864
rect -33224 -13176 -33144 -13072
<< metal2 >>
rect -9419 2750 -9323 2760
rect -9419 2644 -9323 2654
rect -32220 -864 -32124 -854
rect -32220 -970 -32124 -960
rect -31492 -864 -31412 -858
rect -32220 -3024 -32124 -3014
rect -32220 -3130 -32124 -3120
rect -31652 -3024 -31572 -3018
rect -32220 -3744 -32124 -3734
rect -32220 -3850 -32124 -3840
rect -31812 -3744 -31732 -3738
rect -33224 -4572 -33144 -4566
rect -40692 -11200 -40588 -11190
rect -40692 -11314 -40588 -11304
rect -36644 -11408 -36540 -11398
rect -36644 -11522 -36540 -11512
rect -34620 -11616 -34516 -11606
rect -34620 -11730 -34516 -11720
rect -33608 -11824 -33504 -11814
rect -33608 -11938 -33504 -11928
rect -33224 -13072 -33144 -4668
rect -32220 -4572 -32124 -4562
rect -32220 -4678 -32124 -4668
rect -32904 -4932 -32824 -4926
rect -33064 -5292 -32984 -5286
rect -33064 -12864 -32984 -5388
rect -32904 -5652 -32824 -5028
rect -32904 -12656 -32824 -5748
rect -32220 -5652 -32124 -5642
rect -32220 -5758 -32124 -5748
rect -32220 -5904 -32124 -5894
rect -32220 -6010 -32124 -6000
rect -31812 -5904 -31732 -3840
rect -32220 -7344 -32124 -7334
rect -32220 -7450 -32124 -7440
rect -32220 -9504 -32124 -9494
rect -32220 -9610 -32124 -9600
rect -31812 -12448 -31732 -6000
rect -31652 -7344 -31572 -3120
rect -31652 -12240 -31572 -7440
rect -31492 -9504 -31412 -960
rect -30808 -864 -30712 -854
rect -30808 -970 -30712 -960
rect -30808 -3024 -30712 -3014
rect -30808 -3130 -30712 -3120
rect -30808 -3744 -30712 -3734
rect -30808 -3850 -30712 -3840
rect -30808 -4932 -30712 -4922
rect -30808 -5038 -30712 -5028
rect -30808 -5292 -30712 -5282
rect -30808 -5398 -30712 -5388
rect -30808 -5904 -30712 -5894
rect -30808 -6010 -30712 -6000
rect -30808 -7344 -30712 -7334
rect -30808 -7450 -30712 -7440
rect -31492 -12032 -31412 -9600
rect -30808 -9504 -30712 -9494
rect -30808 -9610 -30712 -9600
rect -22688 -11200 -22584 -11190
rect -22688 -11314 -22584 -11304
rect -26736 -11408 -26632 -11398
rect -26736 -11522 -26632 -11512
rect -28760 -11616 -28656 -11606
rect -28760 -11730 -28656 -11720
rect -29772 -11824 -29668 -11814
rect -29772 -11938 -29668 -11928
rect -31492 -12146 -31412 -12136
rect -31652 -12354 -31572 -12344
rect -31812 -12562 -31732 -12552
rect -32904 -12770 -32824 -12760
rect -33064 -12978 -32984 -12968
rect -33224 -13186 -33144 -13176
<< via2 >>
rect -9419 2654 -9323 2750
rect -32220 -960 -32124 -864
rect -32220 -3120 -32124 -3024
rect -32220 -3840 -32124 -3744
rect -40692 -11304 -40588 -11200
rect -36644 -11512 -36540 -11408
rect -34620 -11720 -34516 -11616
rect -33608 -11928 -33504 -11824
rect -32220 -4668 -32124 -4572
rect -32220 -5748 -32124 -5652
rect -32220 -6000 -32124 -5904
rect -32220 -7440 -32124 -7344
rect -32220 -9600 -32124 -9504
rect -30808 -960 -30712 -864
rect -30808 -3120 -30712 -3024
rect -30808 -3840 -30712 -3744
rect -30808 -5028 -30712 -4932
rect -30808 -5388 -30712 -5292
rect -30808 -6000 -30712 -5904
rect -30808 -7440 -30712 -7344
rect -30808 -9600 -30712 -9504
rect -22688 -11304 -22584 -11200
rect -26736 -11512 -26632 -11408
rect -28760 -11720 -28656 -11616
rect -29772 -11928 -29668 -11824
<< metal3 >>
rect -9429 2750 -9313 2755
rect -9429 2654 -9419 2750
rect -9323 2654 -9313 2750
rect -9429 2649 -9313 2654
rect -32230 -864 -32114 -859
rect -32230 -960 -32220 -864
rect -32124 -960 -32114 -864
rect -32230 -965 -32114 -960
rect -30818 -864 -30702 -859
rect -30818 -960 -30808 -864
rect -30712 -960 -30702 -864
rect -30818 -965 -30702 -960
rect -32230 -3024 -32114 -3019
rect -32230 -3120 -32220 -3024
rect -32124 -3120 -32114 -3024
rect -32230 -3125 -32114 -3120
rect -30818 -3024 -30702 -3019
rect -30818 -3120 -30808 -3024
rect -30712 -3120 -30702 -3024
rect -30818 -3125 -30702 -3120
rect -32230 -3744 -32114 -3739
rect -32230 -3840 -32220 -3744
rect -32124 -3840 -32114 -3744
rect -32230 -3845 -32114 -3840
rect -30818 -3744 -30702 -3739
rect -30818 -3840 -30808 -3744
rect -30712 -3840 -30702 -3744
rect -30818 -3845 -30702 -3840
rect -32230 -4572 -32114 -4567
rect -32230 -4668 -32220 -4572
rect -32124 -4668 -32114 -4572
rect -32230 -4673 -32114 -4668
rect -30818 -4932 -30702 -4927
rect -30818 -5028 -30808 -4932
rect -30712 -5028 -30702 -4932
rect -30818 -5033 -30702 -5028
rect -30818 -5292 -30702 -5287
rect -30818 -5388 -30808 -5292
rect -30712 -5388 -30702 -5292
rect -30818 -5393 -30702 -5388
rect -32230 -5652 -32114 -5647
rect -32230 -5748 -32220 -5652
rect -32124 -5748 -32114 -5652
rect -32230 -5753 -32114 -5748
rect -32230 -5904 -32114 -5899
rect -32230 -6000 -32220 -5904
rect -32124 -6000 -32114 -5904
rect -32230 -6005 -32114 -6000
rect -30818 -5904 -30702 -5899
rect -30818 -6000 -30808 -5904
rect -30712 -6000 -30702 -5904
rect -30818 -6005 -30702 -6000
rect -32230 -7344 -32114 -7339
rect -32230 -7440 -32220 -7344
rect -32124 -7440 -32114 -7344
rect -32230 -7445 -32114 -7440
rect -30818 -7344 -30702 -7339
rect -30818 -7440 -30808 -7344
rect -30712 -7440 -30702 -7344
rect -30818 -7445 -30702 -7440
rect -32230 -9504 -32114 -9499
rect -32230 -9600 -32220 -9504
rect -32124 -9600 -32114 -9504
rect -32230 -9605 -32114 -9600
rect -30818 -9504 -30702 -9499
rect -30818 -9600 -30808 -9504
rect -30712 -9600 -30702 -9504
rect -30818 -9605 -30702 -9600
rect -40702 -11200 -40578 -11195
rect -40702 -11304 -40692 -11200
rect -40588 -11304 -40578 -11200
rect -40702 -11309 -40578 -11304
rect -22698 -11200 -22574 -11195
rect -22698 -11304 -22688 -11200
rect -22584 -11304 -22574 -11200
rect -22698 -11309 -22574 -11304
rect -36654 -11408 -36530 -11403
rect -36654 -11512 -36644 -11408
rect -36540 -11512 -36530 -11408
rect -36654 -11517 -36530 -11512
rect -26746 -11408 -26622 -11403
rect -26746 -11512 -26736 -11408
rect -26632 -11512 -26622 -11408
rect -26746 -11517 -26622 -11512
rect -34630 -11616 -34506 -11611
rect -34630 -11720 -34620 -11616
rect -34516 -11720 -34506 -11616
rect -34630 -11725 -34506 -11720
rect -28770 -11616 -28646 -11611
rect -28770 -11720 -28760 -11616
rect -28656 -11720 -28646 -11616
rect -28770 -11725 -28646 -11720
rect -33618 -11824 -33494 -11819
rect -33618 -11928 -33608 -11824
rect -33504 -11928 -33494 -11824
rect -33618 -11933 -33494 -11928
rect -29782 -11824 -29658 -11819
rect -29782 -11928 -29772 -11824
rect -29668 -11928 -29658 -11824
rect -29782 -11933 -29658 -11928
<< via3 >>
rect -9419 2654 -9323 2750
rect -32220 -960 -32124 -864
rect -30808 -960 -30712 -864
rect -32220 -3120 -32124 -3024
rect -30808 -3120 -30712 -3024
rect -32220 -3840 -32124 -3744
rect -30808 -3840 -30712 -3744
rect -32220 -4668 -32124 -4572
rect -30808 -5028 -30712 -4932
rect -30808 -5388 -30712 -5292
rect -32220 -5748 -32124 -5652
rect -32220 -6000 -32124 -5904
rect -30808 -6000 -30712 -5904
rect -32220 -7440 -32124 -7344
rect -30808 -7440 -30712 -7344
rect -32220 -9600 -32124 -9504
rect -30808 -9600 -30712 -9504
rect -40692 -11304 -40588 -11200
rect -22688 -11304 -22584 -11200
rect -36644 -11512 -36540 -11408
rect -26736 -11512 -26632 -11408
rect -34620 -11720 -34516 -11616
rect -28760 -11720 -28656 -11616
rect -33608 -11928 -33504 -11824
rect -29772 -11928 -29668 -11824
<< metal4 >>
rect -9420 2750 -9322 2751
rect -9695 2654 -9419 2750
rect -9323 2654 -9322 2750
rect -9420 2653 -9322 2654
rect -48444 704 -15450 808
rect -48256 600 -48152 704
rect -47244 600 -47140 704
rect -46232 600 -46128 704
rect -45220 600 -45116 704
rect -44208 600 -44104 704
rect -43196 600 -43092 704
rect -42184 600 -42080 704
rect -41172 600 -41068 704
rect -40160 600 -40056 704
rect -39148 600 -39044 704
rect -38136 600 -38032 704
rect -37124 600 -37020 704
rect -36112 600 -36008 704
rect -35100 600 -34996 704
rect -34088 600 -33984 704
rect -33076 600 -32972 704
rect -31664 600 -31560 704
rect -30252 455 -30148 704
rect -29240 463 -29136 704
rect -28228 600 -28124 704
rect -27216 600 -27112 704
rect -26204 600 -26100 704
rect -25192 600 -25088 704
rect -24180 600 -24076 704
rect -23168 600 -23064 704
rect -22156 600 -22052 704
rect -21144 600 -21040 704
rect -20132 600 -20028 704
rect -19120 600 -19016 704
rect -18108 600 -18004 704
rect -17096 600 -16992 704
rect -16084 600 -15980 704
rect -32592 -864 -32496 12
rect -32221 -864 -32123 -863
rect -32592 -960 -32220 -864
rect -32124 -960 -32123 -864
rect -32592 -1692 -32496 -960
rect -32221 -961 -32123 -960
rect -31180 -864 -31084 12
rect -30809 -864 -30711 -863
rect -31180 -960 -30808 -864
rect -30712 -960 -30711 -864
rect -31180 -1692 -31084 -960
rect -30809 -961 -30711 -960
rect -32592 -3024 -32496 -2868
rect -32221 -3024 -32123 -3023
rect -32592 -3120 -32220 -3024
rect -32124 -3120 -32123 -3024
rect -32592 -3177 -32496 -3120
rect -32221 -3121 -32123 -3120
rect -31180 -3024 -31084 -2868
rect -30809 -3024 -30711 -3023
rect -31180 -3120 -30808 -3024
rect -30712 -3120 -30711 -3024
rect -31180 -3186 -31084 -3120
rect -30809 -3121 -30711 -3120
rect -32221 -3744 -32123 -3743
rect -30809 -3744 -30711 -3743
rect -32592 -3840 -32220 -3744
rect -32124 -3840 -32123 -3744
rect -32592 -3923 -32496 -3840
rect -32221 -3841 -32123 -3840
rect -31180 -3840 -30808 -3744
rect -30712 -3840 -30711 -3744
rect -31180 -3949 -31084 -3840
rect -30809 -3841 -30711 -3840
rect -32221 -4572 -32123 -4571
rect -32496 -4668 -32220 -4572
rect -32124 -4668 -32123 -4572
rect -32221 -4669 -32123 -4668
rect -30809 -4932 -30711 -4931
rect -31084 -5028 -30808 -4932
rect -30712 -5028 -30711 -4932
rect -30809 -5029 -30711 -5028
rect -30809 -5292 -30711 -5291
rect -31155 -5388 -30808 -5292
rect -30712 -5388 -30711 -5292
rect -30809 -5389 -30711 -5388
rect -32221 -5652 -32123 -5651
rect -32565 -5748 -32220 -5652
rect -32124 -5748 -32123 -5652
rect -32221 -5749 -32123 -5748
rect -32221 -5904 -32123 -5903
rect -30809 -5904 -30711 -5903
rect -32592 -6000 -32220 -5904
rect -32124 -6000 -32123 -5904
rect -32592 -6070 -32496 -6000
rect -32221 -6001 -32123 -6000
rect -31180 -6000 -30808 -5904
rect -30712 -6000 -30711 -5904
rect -31180 -6089 -31084 -6000
rect -30809 -6001 -30711 -6000
rect -32592 -7344 -32496 -7188
rect -32221 -7344 -32123 -7343
rect -32592 -7440 -32220 -7344
rect -32124 -7440 -32123 -7344
rect -32592 -7503 -32496 -7440
rect -32221 -7441 -32123 -7440
rect -31180 -7344 -31084 -7188
rect -30809 -7344 -30711 -7343
rect -31180 -7440 -30808 -7344
rect -30712 -7440 -30711 -7344
rect -31180 -7492 -31084 -7440
rect -30809 -7441 -30711 -7440
rect -32592 -9504 -32496 -8628
rect -32221 -9504 -32123 -9503
rect -32592 -9600 -32220 -9504
rect -32124 -9600 -32123 -9504
rect -32592 -10332 -32496 -9600
rect -32221 -9601 -32123 -9600
rect -31180 -9504 -31084 -8628
rect -30809 -9504 -30711 -9503
rect -31180 -9600 -30808 -9504
rect -30712 -9600 -30711 -9504
rect -31180 -10332 -31084 -9600
rect -30809 -9601 -30711 -9600
rect -47776 -11024 -47672 -10920
rect -46764 -11024 -46660 -10920
rect -45752 -11024 -45648 -10920
rect -44740 -11024 -44636 -10920
rect -43728 -11024 -43624 -10920
rect -42716 -11024 -42612 -10920
rect -41704 -11024 -41600 -10920
rect -40692 -11024 -40588 -10920
rect -47776 -11128 -40588 -11024
rect -39680 -11024 -39576 -10920
rect -38668 -11024 -38564 -10920
rect -37656 -11024 -37552 -10920
rect -36644 -11024 -36540 -10920
rect -39680 -11128 -36540 -11024
rect -35632 -11024 -35528 -10920
rect -34620 -11024 -34516 -10920
rect -35632 -11128 -34516 -11024
rect -40692 -11199 -40588 -11128
rect -40693 -11200 -40587 -11199
rect -40693 -11304 -40692 -11200
rect -40588 -11304 -40587 -11200
rect -40693 -11305 -40587 -11304
rect -36644 -11407 -36540 -11128
rect -36645 -11408 -36539 -11407
rect -36645 -11512 -36644 -11408
rect -36540 -11512 -36539 -11408
rect -36645 -11513 -36539 -11512
rect -34620 -11615 -34516 -11128
rect -34621 -11616 -34515 -11615
rect -34621 -11720 -34620 -11616
rect -34516 -11720 -34515 -11616
rect -34621 -11721 -34515 -11720
rect -33608 -11823 -33504 -10920
rect -29772 -11823 -29668 -10857
rect -28760 -11024 -28656 -10920
rect -27748 -11024 -27644 -10816
rect -28760 -11128 -27644 -11024
rect -26736 -11024 -26632 -10920
rect -25724 -11024 -25620 -10816
rect -24712 -11024 -24608 -10810
rect -23700 -11024 -23596 -10816
rect -26736 -11128 -23596 -11024
rect -22688 -11024 -22584 -10920
rect -21676 -11024 -21572 -10816
rect -20664 -11024 -20560 -10816
rect -19652 -11024 -19548 -10811
rect -18640 -11024 -18536 -10816
rect -17628 -11024 -17524 -10811
rect -16616 -11024 -16512 -10816
rect -15604 -11024 -15500 -10816
rect -22688 -11128 -15500 -11024
rect -28760 -11615 -28656 -11128
rect -26736 -11407 -26632 -11128
rect -22688 -11199 -22584 -11128
rect -22689 -11200 -22583 -11199
rect -22689 -11304 -22688 -11200
rect -22584 -11304 -22583 -11200
rect -22689 -11305 -22583 -11304
rect -26737 -11408 -26631 -11407
rect -26737 -11512 -26736 -11408
rect -26632 -11512 -26631 -11408
rect -26737 -11513 -26631 -11512
rect -28761 -11616 -28655 -11615
rect -28761 -11720 -28760 -11616
rect -28656 -11720 -28655 -11616
rect -28761 -11721 -28655 -11720
rect -33609 -11824 -33503 -11823
rect -33609 -11928 -33608 -11824
rect -33504 -11928 -33503 -11824
rect -33609 -11929 -33503 -11928
rect -29773 -11824 -29667 -11823
rect -29773 -11928 -29772 -11824
rect -29668 -11928 -29667 -11824
rect -29773 -11929 -29667 -11928
use sky130_fd_pr__cap_mim_m3_1_NL85WR  sky130_fd_pr__cap_mim_m3_1_NL85WR_0
timestamp 1757961500
transform 1 0 -31466 0 1 -5160
box -386 -5760 386 5760
use sky130_fd_pr__cap_mim_m3_1_NL85WR  sky130_fd_pr__cap_mim_m3_1_NL85WR_1
timestamp 1757961500
transform 1 0 -32878 0 1 -5160
box -386 -5760 386 5760
use sky130_fd_pr__cap_mim_m3_1_TE2UD4  sky130_fd_pr__cap_mim_m3_1_TE2UD4_0
timestamp 1757858808
transform 1 0 -40974 0 1 -5160
box -7470 -5760 7470 5760
use sky130_fd_pr__cap_mim_m3_1_TE2UD4  sky130_fd_pr__cap_mim_m3_1_TE2UD4_1
timestamp 1757858808
transform 1 0 -22970 0 1 -5160
box -7470 -5760 7470 5760
<< labels >>
flabel metal1 -15604 -13176 -15500 -13072 0 FreeSans 320 0 0 0 VCM
port 10 nsew
flabel metal1 -15604 -11304 -15500 -11200 0 FreeSans 320 0 0 0 S[0]
port 9 nsew
flabel metal1 -15604 -11512 -15500 -11408 0 FreeSans 320 0 0 0 S[1]
port 8 nsew
flabel metal1 -15604 -11720 -15500 -11616 0 FreeSans 320 0 0 0 S[2]
port 7 nsew
flabel metal1 -15604 -11928 -15500 -11824 0 FreeSans 320 0 0 0 S[3]
port 6 nsew
flabel metal1 -15604 -12136 -15500 -12032 0 FreeSans 320 0 0 0 S[4]
port 5 nsew
flabel metal1 -15604 -12344 -15500 -12240 0 FreeSans 320 0 0 0 S[5]
port 4 nsew
flabel metal1 -15604 -12552 -15500 -12448 0 FreeSans 320 0 0 0 S[6]
port 3 nsew
flabel metal1 -15604 -12760 -15500 -12656 0 FreeSans 320 0 0 0 S[7]
port 2 nsew
flabel metal1 -15604 -12968 -15500 -12864 0 FreeSans 320 0 0 0 S[8]
port 1 nsew
<< end >>
