magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< pwell >>
rect -236 -565 236 565
<< nmos >>
rect -50 265 50 365
rect -50 55 50 155
rect -50 -155 50 -55
rect -50 -365 50 -265
<< ndiff >>
rect -108 332 -50 365
rect -108 298 -96 332
rect -62 298 -50 332
rect -108 265 -50 298
rect 50 332 108 365
rect 50 298 62 332
rect 96 298 108 332
rect 50 265 108 298
rect -108 122 -50 155
rect -108 88 -96 122
rect -62 88 -50 122
rect -108 55 -50 88
rect 50 122 108 155
rect 50 88 62 122
rect 96 88 108 122
rect 50 55 108 88
rect -108 -88 -50 -55
rect -108 -122 -96 -88
rect -62 -122 -50 -88
rect -108 -155 -50 -122
rect 50 -88 108 -55
rect 50 -122 62 -88
rect 96 -122 108 -88
rect 50 -155 108 -122
rect -108 -298 -50 -265
rect -108 -332 -96 -298
rect -62 -332 -50 -298
rect -108 -365 -50 -332
rect 50 -298 108 -265
rect 50 -332 62 -298
rect 96 -332 108 -298
rect 50 -365 108 -332
<< ndiffc >>
rect -96 298 -62 332
rect 62 298 96 332
rect -96 88 -62 122
rect 62 88 96 122
rect -96 -122 -62 -88
rect 62 -122 96 -88
rect -96 -332 -62 -298
rect 62 -332 96 -298
<< psubdiff >>
rect -210 505 -85 539
rect -51 505 -17 539
rect 17 505 51 539
rect 85 505 210 539
rect -210 425 -176 505
rect -210 357 -176 391
rect 176 425 210 505
rect -210 289 -176 323
rect 176 357 210 391
rect 176 289 210 323
rect -210 221 -176 255
rect -210 153 -176 187
rect 176 221 210 255
rect -210 85 -176 119
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect 176 -119 210 -85
rect -210 -255 -176 -221
rect 176 -187 210 -153
rect 176 -255 210 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect 176 -323 210 -289
rect -210 -505 -176 -425
rect 176 -391 210 -357
rect 176 -505 210 -425
rect -210 -539 -85 -505
rect -51 -539 -17 -505
rect 17 -539 51 -505
rect 85 -539 210 -505
<< psubdiffcont >>
rect -85 505 -51 539
rect -17 505 17 539
rect 51 505 85 539
rect -210 391 -176 425
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect 176 323 210 357
rect -210 187 -176 221
rect 176 255 210 289
rect 176 187 210 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect 176 -85 210 -51
rect 176 -153 210 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect 176 -221 210 -187
rect -210 -357 -176 -323
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect 176 -425 210 -391
rect -85 -539 -51 -505
rect -17 -539 17 -505
rect 51 -539 85 -505
<< poly >>
rect -50 437 50 453
rect -50 403 -17 437
rect 17 403 50 437
rect -50 365 50 403
rect -50 227 50 265
rect -50 193 -17 227
rect 17 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect -50 -265 50 -227
rect -50 -403 50 -365
rect -50 -437 -17 -403
rect 17 -437 50 -403
rect -50 -453 50 -437
<< polycont >>
rect -17 403 17 437
rect -17 193 17 227
rect -17 -17 17 17
rect -17 -227 17 -193
rect -17 -437 17 -403
<< locali >>
rect -210 505 -85 539
rect -51 505 -17 539
rect 17 505 51 539
rect 85 505 210 539
rect -210 425 -176 505
rect -50 403 -17 437
rect 17 403 50 437
rect 176 425 210 505
rect -210 357 -176 391
rect -210 289 -176 323
rect -96 332 -62 369
rect -96 261 -62 298
rect 62 332 96 369
rect 62 261 96 298
rect 176 357 210 391
rect 176 289 210 323
rect -210 221 -176 255
rect -50 193 -17 227
rect 17 193 50 227
rect 176 221 210 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -96 122 -62 159
rect -96 51 -62 88
rect 62 122 96 159
rect 62 51 96 88
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect 176 17 210 51
rect -50 -17 -17 17
rect 17 -17 50 17
rect -210 -51 -176 -17
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -96 -88 -62 -51
rect -96 -159 -62 -122
rect 62 -88 96 -51
rect 62 -159 96 -122
rect 176 -119 210 -85
rect 176 -187 210 -153
rect -210 -255 -176 -221
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect 176 -255 210 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -96 -298 -62 -261
rect -96 -369 -62 -332
rect 62 -298 96 -261
rect 62 -369 96 -332
rect 176 -323 210 -289
rect 176 -391 210 -357
rect -210 -505 -176 -425
rect -50 -437 -17 -403
rect 17 -437 50 -403
rect 176 -505 210 -425
rect -210 -539 -85 -505
rect -51 -539 -17 -505
rect 17 -539 51 -505
rect 85 -539 210 -505
<< viali >>
rect -17 403 17 437
rect -96 298 -62 332
rect 62 298 96 332
rect -17 193 17 227
rect -96 88 -62 122
rect 62 88 96 122
rect -17 -17 17 17
rect -96 -122 -62 -88
rect 62 -122 96 -88
rect -17 -227 17 -193
rect -96 -332 -62 -298
rect 62 -332 96 -298
rect -17 -437 17 -403
<< metal1 >>
rect -46 437 46 443
rect -46 403 -17 437
rect 17 403 46 437
rect -46 397 46 403
rect -102 332 -56 365
rect -102 298 -96 332
rect -62 298 -56 332
rect -102 265 -56 298
rect 56 332 102 365
rect 56 298 62 332
rect 96 298 102 332
rect 56 265 102 298
rect -46 227 46 233
rect -46 193 -17 227
rect 17 193 46 227
rect -46 187 46 193
rect -102 122 -56 155
rect -102 88 -96 122
rect -62 88 -56 122
rect -102 55 -56 88
rect 56 122 102 155
rect 56 88 62 122
rect 96 88 102 122
rect 56 55 102 88
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -88 -56 -55
rect -102 -122 -96 -88
rect -62 -122 -56 -88
rect -102 -155 -56 -122
rect 56 -88 102 -55
rect 56 -122 62 -88
rect 96 -122 102 -88
rect 56 -155 102 -122
rect -46 -193 46 -187
rect -46 -227 -17 -193
rect 17 -227 46 -193
rect -46 -233 46 -227
rect -102 -298 -56 -265
rect -102 -332 -96 -298
rect -62 -332 -56 -298
rect -102 -365 -56 -332
rect 56 -298 102 -265
rect 56 -332 62 -298
rect 96 -332 102 -298
rect 56 -365 102 -332
rect -46 -403 46 -397
rect -46 -437 -17 -403
rect 17 -437 46 -403
rect -46 -443 46 -437
<< properties >>
string FIXED_BBOX -193 -522 193 522
<< end >>
