magic
tech sky130A
magscale 1 2
timestamp 1757961947
<< viali >>
rect 46770 20680 46870 20780
<< metal1 >>
rect 22350 19550 22450 25770
rect 22560 23580 22660 24940
rect 22550 23480 22560 23580
rect 22660 23480 22670 23580
rect 22560 20459 22660 23480
rect 22750 21680 22760 21780
rect 22860 21680 22870 21780
rect 22760 20520 22860 21680
rect 21880 19370 21890 19550
rect 22070 19530 22450 19550
rect 22070 19370 22372 19530
rect 23960 18884 24112 26836
rect 25716 18593 25890 26767
rect 27362 23380 27462 24968
rect 27352 23280 27362 23380
rect 27462 23280 27472 23380
rect 27362 20519 27462 23280
rect 27552 21480 27562 21580
rect 27662 21480 27672 21580
rect 27562 20518 27662 21480
rect 28762 18664 28914 26836
rect 30518 18630 30692 26847
rect 32164 23180 32264 24940
rect 32154 23080 32164 23180
rect 32264 23080 32274 23180
rect 32164 20544 32264 23080
rect 32354 21280 32364 21380
rect 32464 21280 32474 21380
rect 32364 20515 32464 21280
rect 33564 18684 33716 26836
rect 35320 18613 35494 27047
rect 36966 22980 37066 24970
rect 37166 24780 37266 24940
rect 37156 24680 37166 24780
rect 37266 24680 37276 24780
rect 36956 22880 36966 22980
rect 37066 22880 37076 22980
rect 36966 20479 37066 22880
rect 37156 21080 37166 21180
rect 37266 21080 37276 21180
rect 37166 20520 37266 21080
rect 38366 18744 38518 26796
rect 40122 18673 40296 26847
rect 41768 22780 41868 24941
rect 41968 24580 42068 24940
rect 41958 24480 41968 24580
rect 42068 24480 42078 24580
rect 41758 22680 41768 22780
rect 41868 22680 41878 22780
rect 41768 20541 41868 22680
rect 41958 20880 41968 20980
rect 42068 20880 42078 20980
rect 41968 20520 42068 20880
rect 43168 18644 43320 26796
rect 44924 18653 45098 26830
rect 46570 22580 46670 24911
rect 46770 24380 46870 24940
rect 46760 24280 46770 24380
rect 46870 24280 46880 24380
rect 46560 22480 46570 22580
rect 46670 22480 46680 22580
rect 46570 20516 46670 22480
rect 46758 20780 46882 20786
rect 46758 20680 46770 20780
rect 46870 20680 46882 20780
rect 46758 20674 46882 20680
rect 46770 20520 46870 20674
rect 47971 18804 48123 26816
rect 49727 18673 49901 26847
rect 51372 22380 51472 24909
rect 51572 24180 51672 24940
rect 51562 24080 51572 24180
rect 51672 24080 51682 24180
rect 51362 22280 51372 22380
rect 51472 22280 51482 22380
rect 51372 20520 51472 22280
rect 51562 20480 51572 20580
rect 51672 20480 51682 20580
rect 52782 18764 52934 26796
rect 54538 18630 54712 26787
rect 56174 22180 56274 24937
rect 56374 23980 56474 24943
rect 56364 23880 56374 23980
rect 56474 23880 56484 23980
rect 56164 22080 56174 22180
rect 56274 22080 56284 22180
rect 56174 20520 56274 22080
rect 57574 18804 57726 26616
rect 59330 18630 59504 26787
rect 60976 21980 61076 24902
rect 61176 23780 61276 24940
rect 61166 23680 61176 23780
rect 61276 23680 61286 23780
rect 60966 21880 60976 21980
rect 61076 21880 61086 21980
rect 60976 20510 61076 21880
rect 62376 18764 62528 26836
rect 64132 18630 64306 26747
rect 16623 14220 16633 14300
rect 16713 14220 16723 14300
rect 5218 14072 5228 14128
rect 5284 14072 5294 14128
rect 10786 14090 10796 14152
rect 10852 14141 10862 14152
rect 10852 14101 16615 14141
rect 10852 14090 10862 14101
rect 5234 14001 5274 14072
rect 5234 13961 16403 14001
rect 16363 13717 16403 13961
rect 16575 13711 16615 14101
rect 16654 13708 16694 14220
rect 18727 13980 18737 14080
rect 18837 13980 20699 14080
rect 20599 8800 20699 13980
rect 20599 8700 23888 8800
rect 12701 7984 12711 8088
rect 12815 7984 12825 8088
rect 8465 7470 8475 7530
rect 8531 7470 8541 7530
rect 791 7149 801 7245
rect 1200 7149 3374 7245
rect 12711 7048 12815 7984
rect 15986 7245 16020 8406
rect 14717 6989 16020 7245
rect 16202 7245 16236 8423
rect 19429 8250 19439 8354
rect 19543 8250 19553 8354
rect 16202 6989 17451 7245
rect 19439 7059 19543 8250
rect 23788 7486 23888 8700
rect 190 1135 200 1231
rect 600 1135 11763 1231
<< via1 >>
rect 22560 23480 22660 23580
rect 22760 21680 22860 21780
rect 21890 19370 22070 19550
rect 27362 23280 27462 23380
rect 27562 21480 27662 21580
rect 32164 23080 32264 23180
rect 32364 21280 32464 21380
rect 37166 24680 37266 24780
rect 36966 22880 37066 22980
rect 37166 21080 37266 21180
rect 41968 24480 42068 24580
rect 41768 22680 41868 22780
rect 41968 20880 42068 20980
rect 46770 24280 46870 24380
rect 46570 22480 46670 22580
rect 46770 20680 46870 20780
rect 51572 24080 51672 24180
rect 51372 22280 51472 22380
rect 51572 20480 51672 20580
rect 56374 23880 56474 23980
rect 56174 22080 56274 22180
rect 61176 23680 61276 23780
rect 60976 21880 61076 21980
rect 16633 14220 16713 14300
rect 5228 14072 5284 14128
rect 10796 14090 10852 14152
rect 18737 13980 18837 14080
rect 12711 7984 12815 8088
rect 8475 7470 8531 7530
rect 801 7149 1200 7245
rect 19439 8250 19543 8354
rect 200 1135 600 1231
<< metal2 >>
rect 27620 42240 27760 42250
rect 19131 42220 19231 42230
rect 19231 42141 27620 42201
rect 19131 42110 19231 42120
rect 27620 42090 27760 42100
rect 17020 33160 17420 33170
rect 17420 32760 21420 33160
rect 17020 32750 17420 32760
rect 17020 32360 17420 32370
rect 17420 31960 20540 32360
rect 17020 31950 17420 31960
rect 1640 31400 1760 31410
rect 1640 30570 1760 30580
rect 2800 31400 2920 31410
rect 2800 30570 2920 30580
rect 3940 31400 4060 31410
rect 3940 30570 4060 30580
rect 5100 31400 5220 31410
rect 5100 30570 5220 30580
rect 6240 31400 6360 31410
rect 6240 30570 6360 30580
rect 7400 31400 7520 31410
rect 7400 30570 7520 30580
rect 8560 31400 8680 31410
rect 8560 30570 8680 30580
rect 9700 31400 9820 31410
rect 9700 30570 9820 30580
rect 10860 31400 10980 31410
rect 10860 30570 10980 30580
rect 12020 31400 12140 31410
rect 12020 30570 12140 30580
rect 13160 31400 13280 31410
rect 13160 30570 13280 30580
rect 14320 31400 14440 31410
rect 18340 31045 18420 31055
rect 14440 30965 18340 31045
rect 18340 30955 18420 30965
rect 14320 30570 14440 30580
rect 20140 18880 20540 31960
rect 21020 26480 21420 32760
rect 21020 26380 22850 26480
rect 65150 25380 65890 25480
rect 22760 25080 22860 25090
rect 22760 24970 22860 24980
rect 27562 25080 27662 25090
rect 27562 24970 27662 24980
rect 32364 25080 32464 25090
rect 32364 24970 32464 24980
rect 37166 24780 37266 24790
rect 37166 24670 37266 24680
rect 41968 24580 42068 24590
rect 41968 24470 42068 24480
rect 46770 24380 46870 24390
rect 46770 24270 46870 24280
rect 51572 24180 51672 24190
rect 51572 24070 51672 24080
rect 56374 23980 56474 23990
rect 56374 23870 56474 23880
rect 61176 23780 61276 23790
rect 61176 23670 61276 23680
rect 22560 23580 22660 23590
rect 22560 23470 22660 23480
rect 27362 23380 27462 23390
rect 27362 23270 27462 23280
rect 32164 23180 32264 23190
rect 32164 23070 32264 23080
rect 36966 22980 37066 22990
rect 36966 22870 37066 22880
rect 41768 22780 41868 22790
rect 41768 22670 41868 22680
rect 46570 22580 46670 22590
rect 46570 22470 46670 22480
rect 51372 22380 51472 22390
rect 51372 22270 51472 22280
rect 56174 22180 56274 22190
rect 56174 22070 56274 22080
rect 60976 21980 61076 21990
rect 60976 21870 61076 21880
rect 22760 21780 22860 21790
rect 22760 21670 22860 21680
rect 27562 21580 27662 21590
rect 27562 21470 27662 21480
rect 32364 21380 32464 21390
rect 32364 21270 32464 21280
rect 37166 21180 37266 21190
rect 37166 21070 37266 21080
rect 41968 20980 42068 20990
rect 41968 20870 42068 20880
rect 46770 20780 46870 20790
rect 46770 20670 46870 20680
rect 51572 20580 51672 20590
rect 51572 20470 51672 20480
rect 56374 20480 56474 20490
rect 56374 20370 56474 20380
rect 61176 20480 61276 20490
rect 61176 20370 61276 20380
rect 65790 20080 65890 25380
rect 65450 19980 65890 20080
rect 21890 19550 22070 19560
rect 21890 19360 22070 19370
rect 20140 18780 22850 18880
rect 18340 14600 18420 14610
rect 18340 14510 18420 14520
rect 8000 14300 8080 14310
rect 8000 14210 8080 14220
rect 16633 14300 16713 14310
rect 16633 14210 16713 14220
rect 10796 14152 10852 14162
rect 5228 14128 5284 14138
rect 2420 14080 2520 14090
rect 10796 14080 10852 14090
rect 5228 14062 5284 14072
rect 2420 13970 2520 13980
rect 13580 8648 13636 14154
rect 14460 13700 14620 13710
rect 14460 13530 14620 13540
rect 18354 8677 18406 14510
rect 18737 14080 18837 14090
rect 18737 13970 18837 13980
rect 8475 8592 13636 8648
rect 16150 8625 18406 8677
rect 8475 7530 8531 8592
rect 14260 8360 14420 8370
rect 19439 8354 19543 8364
rect 19439 8240 19543 8250
rect 14260 8190 14420 8200
rect 12711 8088 12815 8098
rect 12711 7974 12815 7984
rect 8475 7460 8531 7470
rect 801 7245 1200 7255
rect 801 7139 1200 7149
rect 200 1231 600 1241
rect 200 1125 600 1135
<< via2 >>
rect 19131 42120 19231 42220
rect 27620 42100 27760 42240
rect 17020 32760 17420 33160
rect 17020 31960 17420 32360
rect 1640 30580 1760 31400
rect 2800 30580 2920 31400
rect 3940 30580 4060 31400
rect 5100 30580 5220 31400
rect 6240 30580 6360 31400
rect 7400 30580 7520 31400
rect 8560 30580 8680 31400
rect 9700 30580 9820 31400
rect 10860 30580 10980 31400
rect 12020 30580 12140 31400
rect 13160 30580 13280 31400
rect 14320 30580 14440 31400
rect 18340 30965 18420 31045
rect 22760 24980 22860 25080
rect 27562 24980 27662 25080
rect 32364 24980 32464 25080
rect 37166 24680 37266 24780
rect 41968 24480 42068 24580
rect 46770 24280 46870 24380
rect 51572 24080 51672 24180
rect 56374 23880 56474 23980
rect 61176 23680 61276 23780
rect 22560 23480 22660 23580
rect 27362 23280 27462 23380
rect 32164 23080 32264 23180
rect 36966 22880 37066 22980
rect 41768 22680 41868 22780
rect 46570 22480 46670 22580
rect 51372 22280 51472 22380
rect 56174 22080 56274 22180
rect 60976 21880 61076 21980
rect 22760 21680 22860 21780
rect 27562 21480 27662 21580
rect 32364 21280 32464 21380
rect 37166 21080 37266 21180
rect 41968 20880 42068 20980
rect 46770 20680 46870 20780
rect 51572 20480 51672 20580
rect 56374 20380 56474 20480
rect 61176 20380 61276 20480
rect 21890 19370 22070 19550
rect 18340 14520 18420 14600
rect 8000 14220 8080 14300
rect 16633 14220 16713 14300
rect 2420 13980 2520 14080
rect 14460 13540 14620 13700
rect 18737 13980 18837 14080
rect 14260 8200 14420 8360
rect 19439 8250 19543 8354
rect 12711 7984 12815 8088
rect 801 7149 1200 7245
rect 200 1135 600 1231
<< metal3 >>
rect 19439 44544 33043 44648
rect 33147 44544 33157 44648
rect 9410 44360 9420 44460
rect 9520 44360 9530 44460
rect 9970 44360 9980 44460
rect 10080 44360 10090 44460
rect 9420 43025 9520 44360
rect 9980 43025 10080 44360
rect 190 42625 200 43025
rect 600 42625 10080 43025
rect 19121 42220 19241 42225
rect 1644 42120 1654 42220
rect 1754 42201 1764 42220
rect 19121 42201 19131 42220
rect 1754 42141 19131 42201
rect 1754 42120 1764 42141
rect 19121 42120 19131 42141
rect 19231 42120 19241 42220
rect 19121 42115 19241 42120
rect 17010 33160 17430 33165
rect 190 32760 200 33160
rect 600 32760 17020 33160
rect 17420 32760 17430 33160
rect 17010 32755 17430 32760
rect 17010 32360 17430 32365
rect 790 31960 800 32360
rect 1200 31960 17020 32360
rect 17420 31960 17430 32360
rect 17010 31955 17430 31960
rect 1630 31400 1770 31405
rect 1630 30580 1640 31400
rect 1760 30580 1770 31400
rect 1630 30575 1770 30580
rect 2790 31400 2930 31405
rect 2790 30580 2800 31400
rect 2920 30580 2930 31400
rect 2790 30575 2930 30580
rect 3930 31400 4070 31405
rect 3930 30580 3940 31400
rect 4060 30580 4070 31400
rect 3930 30575 4070 30580
rect 5090 31400 5230 31405
rect 5090 30580 5100 31400
rect 5220 30580 5230 31400
rect 5090 30575 5230 30580
rect 6230 31400 6370 31405
rect 6230 30580 6240 31400
rect 6360 30580 6370 31400
rect 6230 30575 6370 30580
rect 7390 31400 7530 31405
rect 7390 30580 7400 31400
rect 7520 30580 7530 31400
rect 7390 30575 7530 30580
rect 8550 31400 8690 31405
rect 8550 30580 8560 31400
rect 8680 30580 8690 31400
rect 8550 30575 8690 30580
rect 9690 31400 9830 31405
rect 9690 30580 9700 31400
rect 9820 30580 9830 31400
rect 9690 30575 9830 30580
rect 10850 31400 10990 31405
rect 10850 30580 10860 31400
rect 10980 30580 10990 31400
rect 10850 30575 10990 30580
rect 12010 31400 12150 31405
rect 12010 30580 12020 31400
rect 12140 30580 12150 31400
rect 12010 30575 12150 30580
rect 13150 31400 13290 31405
rect 13150 30580 13160 31400
rect 13280 30580 13290 31400
rect 13150 30575 13290 30580
rect 14310 31400 14450 31405
rect 14310 30580 14320 31400
rect 14440 30580 14450 31400
rect 18330 31045 18430 31050
rect 18330 30965 18340 31045
rect 18420 30965 18430 31045
rect 18330 30960 18430 30965
rect 14310 30575 14450 30580
rect 14376 30366 14386 30486
rect 15186 30366 15196 30486
rect 190 29380 200 29780
rect 600 29380 2840 29780
rect 3240 29380 3250 29780
rect 14376 29774 14386 29894
rect 15186 29774 15196 29894
rect 14376 29182 14386 29302
rect 15186 29182 15196 29302
rect 14376 28590 14386 28710
rect 15186 28590 15196 28710
rect 14376 27998 14386 28118
rect 15186 27998 15196 28118
rect 14376 27406 14386 27526
rect 15186 27406 15196 27526
rect 14376 26814 14386 26934
rect 15186 26814 15196 26934
rect 14376 26222 14386 26342
rect 15186 26222 15196 26342
rect 14376 25630 14386 25750
rect 15186 25630 15196 25750
rect 14376 25038 14386 25158
rect 15186 25038 15196 25158
rect 14376 24446 14386 24566
rect 15186 24446 15196 24566
rect 14376 23854 14386 23974
rect 15186 23854 15196 23974
rect 14376 23262 14386 23382
rect 15186 23262 15196 23382
rect 14376 22670 14386 22790
rect 15186 22670 15196 22790
rect 14376 22078 14386 22198
rect 15186 22078 15196 22198
rect 14376 21486 14386 21606
rect 15186 21486 15196 21606
rect 14376 20894 14386 21014
rect 15186 20894 15196 21014
rect 14376 20302 14386 20422
rect 15186 20302 15196 20422
rect 14376 19710 14386 19830
rect 15186 19710 15196 19830
rect 14376 19118 14386 19238
rect 15186 19118 15196 19238
rect 14376 18526 14386 18646
rect 15186 18526 15196 18646
rect 14376 17934 14386 18054
rect 15186 17934 15196 18054
rect 14376 17342 14386 17462
rect 15186 17342 15196 17462
rect 14376 16750 14386 16870
rect 15186 16750 15196 16870
rect 14376 16158 14386 16278
rect 15186 16158 15196 16278
rect 14376 15566 14386 15686
rect 15186 15566 15196 15686
rect 14376 14974 14386 15094
rect 15186 14974 15196 15094
rect 18340 14605 18420 30960
rect 18330 14600 18430 14605
rect 18330 14520 18340 14600
rect 18420 14520 18430 14600
rect 18330 14515 18430 14520
rect 7990 14300 8090 14305
rect 16623 14300 16723 14305
rect 7990 14220 8000 14300
rect 8080 14220 16633 14300
rect 16713 14220 16723 14300
rect 7990 14215 8090 14220
rect 16623 14215 16723 14220
rect 2410 14080 2530 14085
rect 18727 14080 18847 14085
rect 2410 13980 2420 14080
rect 2520 13980 18737 14080
rect 18837 13980 18847 14080
rect 2410 13975 2530 13980
rect 18727 13975 18847 13980
rect 14450 13700 14630 13705
rect 790 13540 800 13700
rect 1200 13540 14460 13700
rect 14620 13540 14630 13700
rect 14450 13535 14630 13540
rect 14250 8360 14430 8365
rect 190 8200 200 8360
rect 600 8200 14260 8360
rect 14420 8200 14430 8360
rect 19439 8359 19543 44544
rect 27610 42240 27770 42245
rect 27610 42100 27620 42240
rect 27760 42100 27770 42240
rect 27610 42095 27770 42100
rect 22750 25280 22760 25380
rect 22860 25280 22870 25380
rect 22760 25085 22860 25280
rect 22750 25080 22870 25085
rect 22750 24980 22760 25080
rect 22860 24980 22870 25080
rect 22750 24975 22870 24980
rect 27552 24980 27562 25180
rect 27662 24980 27672 25180
rect 27552 24975 27672 24980
rect 32354 25080 32474 25085
rect 32354 24980 32364 25080
rect 32464 24980 32474 25080
rect 32354 24975 32474 24980
rect 37156 24780 37276 24785
rect 37156 24680 37166 24780
rect 37266 24680 37276 24780
rect 37156 24675 37276 24680
rect 41958 24580 42078 24585
rect 41958 24480 41968 24580
rect 42068 24480 42078 24580
rect 41958 24475 42078 24480
rect 46760 24380 46880 24385
rect 46760 24280 46770 24380
rect 46870 24280 46880 24380
rect 46760 24275 46880 24280
rect 51562 24180 51682 24185
rect 51562 24080 51572 24180
rect 51672 24080 51682 24180
rect 51562 24075 51682 24080
rect 56364 23980 56484 23985
rect 56364 23880 56374 23980
rect 56474 23880 56484 23980
rect 56364 23875 56484 23880
rect 61166 23780 61286 23785
rect 61166 23680 61176 23780
rect 61276 23680 61286 23780
rect 61166 23675 61286 23680
rect 22550 23580 22670 23585
rect 22550 23480 22560 23580
rect 22660 23480 22670 23580
rect 22550 23475 22670 23480
rect 27352 23380 27472 23385
rect 27352 23280 27362 23380
rect 27462 23280 27472 23380
rect 27352 23275 27472 23280
rect 32154 23180 32274 23185
rect 32154 23080 32164 23180
rect 32264 23080 32274 23180
rect 32154 23075 32274 23080
rect 36956 22980 37076 22985
rect 36956 22880 36966 22980
rect 37066 22880 37076 22980
rect 36956 22875 37076 22880
rect 41758 22780 41878 22785
rect 41758 22680 41768 22780
rect 41868 22680 41878 22780
rect 41758 22675 41878 22680
rect 46560 22580 46680 22585
rect 46560 22480 46570 22580
rect 46670 22480 46680 22580
rect 46560 22475 46680 22480
rect 51362 22380 51482 22385
rect 51362 22280 51372 22380
rect 51472 22280 51482 22380
rect 51362 22275 51482 22280
rect 56164 22180 56284 22185
rect 56164 22080 56174 22180
rect 56274 22080 56284 22180
rect 56164 22075 56284 22080
rect 60966 21980 61086 21985
rect 60966 21880 60976 21980
rect 61076 21880 61086 21980
rect 60966 21875 61086 21880
rect 22750 21780 22870 21785
rect 22750 21680 22760 21780
rect 22860 21680 22870 21780
rect 22750 21675 22870 21680
rect 27552 21580 27672 21585
rect 27552 21480 27562 21580
rect 27662 21480 27672 21580
rect 27552 21475 27672 21480
rect 32354 21380 32474 21385
rect 32354 21280 32364 21380
rect 32464 21280 32474 21380
rect 32354 21275 32474 21280
rect 37156 21180 37276 21185
rect 37156 21080 37166 21180
rect 37266 21080 37276 21180
rect 37156 21075 37276 21080
rect 41958 20980 42078 20985
rect 41958 20880 41968 20980
rect 42068 20880 42078 20980
rect 41958 20875 42078 20880
rect 46760 20780 46880 20785
rect 46760 20680 46770 20780
rect 46870 20680 46880 20780
rect 46760 20675 46880 20680
rect 51562 20580 51682 20585
rect 51562 20480 51572 20580
rect 51672 20480 51682 20580
rect 51562 20475 51682 20480
rect 56364 20480 56484 20485
rect 56364 20380 56374 20480
rect 56474 20380 56484 20480
rect 56364 20375 56484 20380
rect 61166 20480 61286 20485
rect 61166 20380 61176 20480
rect 61276 20380 61286 20480
rect 61166 20375 61286 20380
rect 21880 19550 22080 19555
rect 21880 19370 21890 19550
rect 22070 19370 22080 19550
rect 21880 19365 22080 19370
rect 19429 8354 19553 8359
rect 19429 8250 19439 8354
rect 19543 8250 19553 8354
rect 19429 8245 19553 8250
rect 14250 8195 14430 8200
rect 12701 8088 12825 8093
rect 12701 7984 12711 8088
rect 12815 7984 32586 8088
rect 12701 7979 12825 7984
rect 791 7245 1210 7250
rect 791 7149 801 7245
rect 1200 7149 1210 7245
rect 791 7144 1210 7149
rect 190 1231 610 1236
rect 190 1135 200 1231
rect 600 1135 610 1231
rect 13482 1154 13492 1370
rect 15228 1154 15238 1370
rect 16986 1154 16996 1370
rect 18732 1154 18742 1370
rect 190 1130 610 1135
rect 32482 916 32586 7984
rect 32482 812 33043 916
rect 33147 812 33157 916
<< via3 >>
rect 33043 44544 33147 44648
rect 9420 44360 9520 44460
rect 9980 44360 10080 44460
rect 200 42625 600 43025
rect 1654 42120 1754 42220
rect 200 32760 600 33160
rect 800 31960 1200 32360
rect 1640 30580 1760 31400
rect 2800 30580 2920 31400
rect 3940 30580 4060 31400
rect 5100 30580 5220 31400
rect 6240 30580 6360 31400
rect 7400 30580 7520 31400
rect 8560 30580 8680 31400
rect 9700 30580 9820 31400
rect 10860 30580 10980 31400
rect 12020 30580 12140 31400
rect 13160 30580 13280 31400
rect 14320 30580 14440 31400
rect 14386 30366 15186 30486
rect 200 29380 600 29780
rect 2840 29380 3240 29780
rect 14386 29774 15186 29894
rect 14386 29182 15186 29302
rect 14386 28590 15186 28710
rect 14386 27998 15186 28118
rect 14386 27406 15186 27526
rect 14386 26814 15186 26934
rect 14386 26222 15186 26342
rect 14386 25630 15186 25750
rect 14386 25038 15186 25158
rect 14386 24446 15186 24566
rect 14386 23854 15186 23974
rect 14386 23262 15186 23382
rect 14386 22670 15186 22790
rect 14386 22078 15186 22198
rect 14386 21486 15186 21606
rect 14386 20894 15186 21014
rect 14386 20302 15186 20422
rect 14386 19710 15186 19830
rect 14386 19118 15186 19238
rect 14386 18526 15186 18646
rect 14386 17934 15186 18054
rect 14386 17342 15186 17462
rect 14386 16750 15186 16870
rect 14386 16158 15186 16278
rect 14386 15566 15186 15686
rect 14386 14974 15186 15094
rect 800 13540 1200 13700
rect 200 8200 600 8360
rect 27620 42100 27760 42240
rect 22760 25280 22860 25380
rect 27562 25080 27662 25180
rect 32364 24980 32464 25080
rect 37166 24680 37266 24780
rect 41968 24480 42068 24580
rect 46770 24280 46870 24380
rect 51572 24080 51672 24180
rect 56374 23880 56474 23980
rect 61176 23680 61276 23780
rect 22560 23480 22660 23580
rect 27362 23280 27462 23380
rect 32164 23080 32264 23180
rect 36966 22880 37066 22980
rect 41768 22680 41868 22780
rect 46570 22480 46670 22580
rect 51372 22280 51472 22380
rect 56174 22080 56274 22180
rect 60976 21880 61076 21980
rect 22760 21680 22860 21780
rect 27562 21480 27662 21580
rect 32364 21280 32464 21380
rect 37166 21080 37266 21180
rect 41968 20880 42068 20980
rect 46770 20680 46870 20780
rect 51572 20480 51672 20580
rect 56374 20380 56474 20480
rect 61176 20380 61276 20480
rect 21890 19370 22070 19550
rect 801 7149 1200 7245
rect 200 1135 600 1231
rect 13492 1154 15228 1370
rect 16996 1154 18732 1370
rect 33043 812 33147 916
<< metal4 >>
rect 200 43026 600 44152
rect 800 43843 1200 44152
rect 6134 43843 6194 45152
rect 6686 43843 6746 45152
rect 7238 43843 7298 45152
rect 7790 43843 7850 45152
rect 8342 43843 8402 45152
rect 8894 43843 8954 45152
rect 9446 44461 9506 45152
rect 9998 44461 10058 45152
rect 9419 44460 9521 44461
rect 9419 44360 9420 44460
rect 9520 44360 9521 44460
rect 9419 44359 9521 44360
rect 9979 44460 10081 44461
rect 9979 44360 9980 44460
rect 10080 44360 10081 44460
rect 9979 44359 10081 44360
rect 10550 43843 10610 45152
rect 11102 43843 11162 45152
rect 11654 43843 11714 45152
rect 12206 43843 12266 45152
rect 12758 43843 12818 45152
rect 13310 43843 13370 45152
rect 800 43443 13370 43843
rect 199 43025 601 43026
rect 199 42625 200 43025
rect 600 42625 601 43025
rect 199 42624 601 42625
rect 200 33161 600 42624
rect 199 33160 601 33161
rect 199 32760 200 33160
rect 600 32760 601 33160
rect 199 32759 601 32760
rect 200 29781 600 32759
rect 800 32361 1200 43443
rect 1653 42220 1755 42221
rect 1653 42120 1654 42220
rect 1754 42120 1755 42220
rect 1653 42119 1755 42120
rect 799 32360 1201 32361
rect 799 31960 800 32360
rect 1200 31960 1201 32360
rect 799 31959 1201 31960
rect 199 29780 601 29781
rect 199 29380 200 29780
rect 600 29380 601 29780
rect 199 29379 601 29380
rect 200 8361 600 29379
rect 800 16100 1200 31959
rect 1674 31401 1734 42119
rect 13862 41180 13922 45152
rect 2825 41120 13922 41180
rect 2825 31401 2885 41120
rect 14414 40491 14474 45152
rect 3978 40431 14474 40491
rect 3978 31401 4038 40431
rect 14966 39832 15026 45152
rect 5130 39772 15026 39832
rect 5130 31401 5190 39772
rect 15518 39240 15578 45152
rect 6282 39180 15578 39240
rect 6282 31401 6342 39180
rect 16070 38633 16130 45152
rect 7434 38573 16130 38633
rect 7434 31401 7494 38573
rect 16622 38060 16682 45152
rect 8586 38000 16682 38060
rect 8586 31401 8646 38000
rect 17174 37556 17234 45152
rect 9738 37496 17234 37556
rect 9738 31401 9798 37496
rect 17726 37171 17786 45152
rect 10890 37111 17786 37171
rect 10890 31401 10950 37111
rect 18278 36758 18338 45152
rect 12042 36698 18338 36758
rect 12042 31401 12102 36698
rect 18830 36440 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 42241 27722 45152
rect 28214 44952 28274 45152
rect 27619 42240 27761 42241
rect 27619 42100 27620 42240
rect 27760 42100 27761 42240
rect 27619 42099 27761 42100
rect 13194 36380 18890 36440
rect 13194 31401 13254 36380
rect 28766 33967 28826 45152
rect 29318 44952 29378 45152
rect 33042 44648 33148 44649
rect 33042 44544 33043 44648
rect 33147 44544 33148 44648
rect 33042 44543 33148 44544
rect 14346 33907 28826 33967
rect 14346 31401 14406 33907
rect 1639 31400 1761 31401
rect 1639 30580 1640 31400
rect 1760 30580 1761 31400
rect 1639 30579 1761 30580
rect 2799 31400 2921 31401
rect 2799 30580 2800 31400
rect 2920 30580 2921 31400
rect 2799 30579 2921 30580
rect 3939 31400 4061 31401
rect 3939 30580 3940 31400
rect 4060 30580 4061 31400
rect 3939 30579 4061 30580
rect 5099 31400 5221 31401
rect 5099 30580 5100 31400
rect 5220 30580 5221 31400
rect 5099 30579 5221 30580
rect 6239 31400 6361 31401
rect 6239 30580 6240 31400
rect 6360 30580 6361 31400
rect 6239 30579 6361 30580
rect 7399 31400 7521 31401
rect 7399 30580 7400 31400
rect 7520 30580 7521 31400
rect 7399 30579 7521 30580
rect 8559 31400 8681 31401
rect 8559 30580 8560 31400
rect 8680 30580 8681 31400
rect 8559 30579 8681 30580
rect 9699 31400 9821 31401
rect 9699 30580 9700 31400
rect 9820 30580 9821 31400
rect 9699 30579 9821 30580
rect 10859 31400 10981 31401
rect 10859 30580 10860 31400
rect 10980 30580 10981 31400
rect 10859 30579 10981 30580
rect 12019 31400 12141 31401
rect 12019 30580 12020 31400
rect 12140 30580 12141 31400
rect 12019 30579 12141 30580
rect 13159 31400 13281 31401
rect 13159 30580 13160 31400
rect 13280 30580 13281 31400
rect 13159 30579 13281 30580
rect 14319 31400 14441 31401
rect 14319 30580 14320 31400
rect 14440 30580 14441 31400
rect 14319 30579 14441 30580
rect 14385 30486 15187 30487
rect 14385 30366 14386 30486
rect 15186 30476 15187 30486
rect 15186 30376 18750 30476
rect 15186 30366 15187 30376
rect 14385 30365 15187 30366
rect 14385 29894 15187 29895
rect 2839 29780 3241 29781
rect 2839 29380 2840 29780
rect 3240 29380 3241 29780
rect 14385 29774 14386 29894
rect 15186 29885 15187 29894
rect 15186 29785 18430 29885
rect 15186 29774 15187 29785
rect 14385 29773 15187 29774
rect 2839 29379 3241 29380
rect 2840 28300 3240 29379
rect 14385 29302 15187 29303
rect 14385 29182 14386 29302
rect 15186 29291 15187 29302
rect 15186 29191 18130 29291
rect 15186 29182 15187 29191
rect 14385 29181 15187 29182
rect 14385 28710 15187 28711
rect 14385 28590 14386 28710
rect 15186 28700 15187 28710
rect 15186 28600 17850 28700
rect 15186 28590 15187 28600
rect 14385 28589 15187 28590
rect 14385 28118 15187 28119
rect 14385 27998 14386 28118
rect 15186 28108 15187 28118
rect 15186 28008 17550 28108
rect 15186 27998 15187 28008
rect 14385 27997 15187 27998
rect 14385 27526 15187 27527
rect 14385 27406 14386 27526
rect 15186 27516 15187 27526
rect 15186 27416 17290 27516
rect 15186 27406 15187 27416
rect 14385 27405 15187 27406
rect 14385 26934 15187 26935
rect 14385 26814 14386 26934
rect 15186 26926 15187 26934
rect 15186 26826 17030 26926
rect 15186 26814 15187 26826
rect 14385 26813 15187 26814
rect 14385 26342 15187 26343
rect 14385 26222 14386 26342
rect 15186 26331 15187 26342
rect 15186 26231 16790 26331
rect 15186 26222 15187 26231
rect 14385 26221 15187 26222
rect 14385 25750 15187 25751
rect 14385 25630 14386 25750
rect 15186 25740 15187 25750
rect 15186 25640 16530 25740
rect 15186 25630 15187 25640
rect 14385 25629 15187 25630
rect 14385 25158 15187 25159
rect 14385 25038 14386 25158
rect 15186 25149 15187 25158
rect 15186 25049 16270 25149
rect 15186 25038 15187 25049
rect 14385 25037 15187 25038
rect 14385 24566 15187 24567
rect 14385 24446 14386 24566
rect 15186 24554 15187 24566
rect 15186 24454 16030 24554
rect 15186 24446 15187 24454
rect 14385 24445 15187 24446
rect 14385 23974 15187 23975
rect 14385 23854 14386 23974
rect 15186 23964 15187 23974
rect 15186 23864 15810 23964
rect 15186 23854 15187 23864
rect 14385 23853 15187 23854
rect 14385 23382 15187 23383
rect 14385 23262 14386 23382
rect 15186 23370 15187 23382
rect 15186 23270 15580 23370
rect 15186 23262 15187 23270
rect 14385 23261 15187 23262
rect 15480 22980 15580 23270
rect 15710 23180 15810 23864
rect 15930 23380 16030 24454
rect 16170 23580 16270 25049
rect 16430 23780 16530 25640
rect 16690 23980 16790 26231
rect 16930 24180 17030 26826
rect 17190 24380 17290 27416
rect 17450 24580 17550 28008
rect 17750 24780 17850 28600
rect 18030 24980 18130 29191
rect 18330 25180 18430 29785
rect 18650 25380 18750 30376
rect 22759 25380 22861 25381
rect 18650 25280 22760 25380
rect 22860 25280 22861 25380
rect 22759 25279 22861 25280
rect 27561 25180 27663 25181
rect 18330 25080 27562 25180
rect 27662 25080 27663 25180
rect 27561 25079 27663 25080
rect 32363 25080 32465 25081
rect 32363 24980 32364 25080
rect 32464 24980 32465 25080
rect 18030 24979 32465 24980
rect 18030 24880 32464 24979
rect 37165 24780 37267 24781
rect 17750 24680 37166 24780
rect 37266 24680 37267 24780
rect 37165 24679 37267 24680
rect 41967 24580 42069 24581
rect 17450 24480 41968 24580
rect 42068 24480 42069 24580
rect 41967 24479 42069 24480
rect 46769 24380 46871 24381
rect 17190 24280 46770 24380
rect 46870 24280 46871 24380
rect 46769 24279 46871 24280
rect 51571 24180 51673 24181
rect 16930 24080 51572 24180
rect 51672 24080 51673 24180
rect 51571 24079 51673 24080
rect 56373 23980 56475 23981
rect 16690 23880 56374 23980
rect 56474 23880 56475 23980
rect 56373 23879 56475 23880
rect 61175 23780 61277 23781
rect 16430 23680 61176 23780
rect 61276 23680 61277 23780
rect 61175 23679 61277 23680
rect 22559 23580 22661 23581
rect 16170 23480 22560 23580
rect 22660 23480 22661 23580
rect 22559 23479 22661 23480
rect 27361 23380 27463 23381
rect 15930 23280 27362 23380
rect 27462 23280 27463 23380
rect 27361 23279 27463 23280
rect 32163 23180 32265 23181
rect 15710 23080 32164 23180
rect 32264 23080 32265 23180
rect 32163 23079 32265 23080
rect 36965 22980 37067 22981
rect 15480 22880 36966 22980
rect 37066 22880 37067 22980
rect 36965 22879 37067 22880
rect 14385 22790 15187 22791
rect 14385 22670 14386 22790
rect 15186 22780 15187 22790
rect 41767 22780 41869 22781
rect 15186 22680 41768 22780
rect 41868 22680 41869 22780
rect 15186 22670 15187 22680
rect 41767 22679 41869 22680
rect 14385 22669 15187 22670
rect 46569 22580 46671 22581
rect 15480 22480 46570 22580
rect 46670 22480 46671 22580
rect 14385 22198 15187 22199
rect 14385 22078 14386 22198
rect 15186 22190 15187 22198
rect 15480 22190 15580 22480
rect 46569 22479 46671 22480
rect 51371 22380 51473 22381
rect 15186 22090 15580 22190
rect 15710 22280 51372 22380
rect 51472 22280 51473 22380
rect 15186 22078 15187 22090
rect 14385 22077 15187 22078
rect 14385 21606 15187 21607
rect 14385 21486 14386 21606
rect 15186 21596 15187 21606
rect 15710 21596 15810 22280
rect 51371 22279 51473 22280
rect 56173 22180 56275 22181
rect 15186 21496 15810 21596
rect 15930 22080 56174 22180
rect 56274 22080 56275 22180
rect 15186 21486 15187 21496
rect 14385 21485 15187 21486
rect 14385 21014 15187 21015
rect 14385 20894 14386 21014
rect 15186 21006 15187 21014
rect 15930 21006 16030 22080
rect 56173 22079 56275 22080
rect 60975 21980 61077 21981
rect 15186 20906 16030 21006
rect 16170 21880 60976 21980
rect 61076 21880 61077 21980
rect 15186 20894 15187 20906
rect 14385 20893 15187 20894
rect 14385 20422 15187 20423
rect 14385 20302 14386 20422
rect 15186 20411 15187 20422
rect 16170 20411 16270 21880
rect 60975 21879 61077 21880
rect 22759 21780 22861 21781
rect 15186 20311 16270 20411
rect 16430 21680 22760 21780
rect 22860 21680 22861 21780
rect 15186 20302 15187 20311
rect 14385 20301 15187 20302
rect 14385 19830 15187 19831
rect 14385 19710 14386 19830
rect 15186 19820 15187 19830
rect 16430 19820 16530 21680
rect 22759 21679 22861 21680
rect 27561 21580 27663 21581
rect 15186 19720 16530 19820
rect 16690 21480 27562 21580
rect 27662 21480 27663 21580
rect 15186 19710 15187 19720
rect 14385 19709 15187 19710
rect 14385 19238 15187 19239
rect 14385 19118 14386 19238
rect 15186 19229 15187 19238
rect 16690 19229 16790 21480
rect 27561 21479 27663 21480
rect 32363 21380 32465 21381
rect 15186 19129 16790 19229
rect 16930 21280 32364 21380
rect 32464 21280 32465 21380
rect 15186 19118 15187 19129
rect 14385 19117 15187 19118
rect 14385 18646 15187 18647
rect 14385 18526 14386 18646
rect 15186 18634 15187 18646
rect 16930 18634 17030 21280
rect 32363 21279 32465 21280
rect 37165 21180 37267 21181
rect 15186 18534 17030 18634
rect 17190 21080 37166 21180
rect 37266 21080 37267 21180
rect 15186 18526 15187 18534
rect 14385 18525 15187 18526
rect 14385 18054 15187 18055
rect 14385 17934 14386 18054
rect 15186 18044 15187 18054
rect 17190 18044 17290 21080
rect 37165 21079 37267 21080
rect 41967 20980 42069 20981
rect 15186 17944 17290 18044
rect 17450 20880 41968 20980
rect 42068 20880 42069 20980
rect 15186 17934 15187 17944
rect 14385 17933 15187 17934
rect 14385 17462 15187 17463
rect 14385 17342 14386 17462
rect 15186 17452 15187 17462
rect 17450 17452 17550 20880
rect 41967 20879 42069 20880
rect 46769 20780 46871 20781
rect 15186 17352 17550 17452
rect 17750 20680 46770 20780
rect 46870 20680 46871 20780
rect 15186 17342 15187 17352
rect 14385 17341 15187 17342
rect 5840 16100 6240 17240
rect 14385 16870 15187 16871
rect 14385 16750 14386 16870
rect 15186 16860 15187 16870
rect 17750 16860 17850 20680
rect 46769 20679 46871 20680
rect 51571 20580 51673 20581
rect 15186 16760 17850 16860
rect 18030 20480 51572 20580
rect 51672 20480 51673 20580
rect 15186 16750 15187 16760
rect 14385 16749 15187 16750
rect 14385 16278 15187 16279
rect 14385 16158 14386 16278
rect 15186 16269 15187 16278
rect 18030 16269 18130 20480
rect 51571 20479 51673 20480
rect 56373 20480 56475 20481
rect 56373 20380 56374 20480
rect 56474 20380 56475 20480
rect 15186 16169 18130 16269
rect 18330 20379 56475 20380
rect 61175 20480 61277 20481
rect 61175 20380 61176 20480
rect 61276 20380 61277 20480
rect 61175 20379 61277 20380
rect 18330 20280 56474 20379
rect 15186 16158 15187 16169
rect 14385 16157 15187 16158
rect 800 15700 6240 16100
rect 800 13701 1200 15700
rect 14385 15686 15187 15687
rect 14385 15566 14386 15686
rect 15186 15675 15187 15686
rect 18330 15675 18430 20280
rect 61176 20180 61276 20379
rect 15186 15575 18430 15675
rect 18650 20080 61276 20180
rect 15186 15566 15187 15575
rect 14385 15565 15187 15566
rect 14385 15094 15187 15095
rect 14385 14974 14386 15094
rect 15186 15084 15187 15094
rect 18650 15084 18750 20080
rect 21889 19550 22071 19551
rect 21889 19370 21890 19550
rect 22070 19370 22071 19550
rect 21889 19369 22071 19370
rect 15186 14984 18750 15084
rect 15186 14974 15187 14984
rect 14385 14973 15187 14974
rect 799 13700 1201 13701
rect 799 13540 800 13700
rect 1200 13540 1201 13700
rect 799 13539 1201 13540
rect 199 8360 601 8361
rect 199 8200 200 8360
rect 600 8200 601 8360
rect 199 8199 601 8200
rect 200 1232 600 8199
rect 800 7246 1200 13539
rect 21890 11150 22070 19369
rect 21890 10970 30542 11150
rect 800 7245 1201 7246
rect 800 7149 801 7245
rect 1200 7149 1201 7245
rect 800 7148 1201 7149
rect 199 1231 601 1232
rect 199 1135 200 1231
rect 600 1135 601 1231
rect 199 1134 601 1135
rect 200 1000 600 1134
rect 800 1000 1200 7148
rect 13491 1370 15229 1371
rect 13491 1154 13492 1370
rect 15228 1154 15229 1370
rect 13491 1153 15229 1154
rect 16995 1370 18733 1371
rect 16995 1154 16996 1370
rect 18732 1154 18733 1370
rect 16995 1153 18733 1154
rect 14250 531 14430 1153
rect 17790 840 17970 1153
rect 17790 660 26678 840
rect 22634 531 22814 532
rect 14250 351 22814 531
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 351
rect 26498 0 26678 660
rect 30362 0 30542 10970
rect 33042 916 33148 917
rect 33042 812 33043 916
rect 33147 812 33148 916
rect 33042 811 33148 812
use sar9b  sar9b_0
timestamp 1757911661
transform 1 0 888 0 1 14072
box 784 0 14298 17322
use single_9b_cdac  single_9b_cdac_0
timestamp 1757961500
transform -1 0 64504 0 1 61688
box -1533 -36848 42164 -15088
use single_9b_cdac  single_9b_cdac_1
timestamp 1757961500
transform -1 0 64504 0 -1 -16228
box -1533 -36848 42164 -15088
use tdc  tdc_0
timestamp 1757893939
transform 0 -1 17291 1 0 8455
box -224 -646 5424 3006
use th_dif_sw  th_dif_sw_0
timestamp 1757961904
transform -1 0 31942 0 -1 7509
box 3069 -413 28591 6385
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
