magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 238 1527 240 1561
rect 274 1527 312 1561
rect 346 1527 384 1561
rect 418 1527 456 1561
rect 490 1527 528 1561
rect 562 1527 600 1561
rect 634 1527 672 1561
rect 706 1527 744 1561
rect 778 1527 816 1561
rect 850 1527 888 1561
rect 922 1527 960 1561
rect 994 1527 1032 1561
rect 1066 1527 1104 1561
rect 1138 1527 1140 1561
rect 272 -123 310 -89
rect 344 -123 382 -89
rect 416 -123 454 -89
rect 488 -123 526 -89
rect 560 -123 598 -89
rect 632 -123 670 -89
<< viali >>
rect 240 1527 274 1561
rect 312 1527 346 1561
rect 384 1527 418 1561
rect 456 1527 490 1561
rect 528 1527 562 1561
rect 600 1527 634 1561
rect 672 1527 706 1561
rect 744 1527 778 1561
rect 816 1527 850 1561
rect 888 1527 922 1561
rect 960 1527 994 1561
rect 1032 1527 1066 1561
rect 1104 1527 1138 1561
rect 238 -123 272 -89
rect 310 -123 344 -89
rect 382 -123 416 -89
rect 454 -123 488 -89
rect 526 -123 560 -89
rect 598 -123 632 -89
rect 670 -123 704 -89
<< metal1 >>
rect 106 1561 1272 1597
rect 106 1527 240 1561
rect 274 1527 312 1561
rect 346 1527 384 1561
rect 418 1527 456 1561
rect 490 1527 528 1561
rect 562 1527 600 1561
rect 634 1527 672 1561
rect 706 1527 744 1561
rect 778 1527 816 1561
rect 850 1527 888 1561
rect 922 1527 960 1561
rect 994 1527 1032 1561
rect 1066 1527 1104 1561
rect 1138 1527 1272 1561
rect 106 1521 1272 1527
rect 325 1447 1053 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 1053 1255
rect 106 915 284 1015
rect 106 570 1272 869
rect 106 423 284 523
rect 316 183 626 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 626 -9
rect 106 -89 1272 -83
rect 106 -123 238 -89
rect 272 -123 310 -89
rect 344 -123 382 -89
rect 416 -123 454 -89
rect 488 -123 526 -89
rect 560 -123 598 -89
rect 632 -123 670 -89
rect 704 -123 1272 -89
rect 106 -159 1272 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_RXFLWN  sky130_fd_pr__nfet_01v8_RXFLWN_0
timestamp 1750100919
transform 0 1 471 -1 0 87
box -236 -355 236 355
use sky130_fd_pr__pfet_01v8_NMYYUH  sky130_fd_pr__pfet_01v8_NMYYUH_0
timestamp 1750100919
transform 0 1 689 -1 0 965
box -246 -583 246 583
use sky130_fd_pr__pfet_01v8_NMYYUH  XM1
timestamp 1750100919
transform 0 1 689 -1 0 1351
box -246 -583 246 583
use sky130_fd_pr__nfet_01v8_RXFLWN  XM3
timestamp 1750100919
transform 0 1 471 -1 0 473
box -236 -355 236 355
<< labels >>
flabel metal1 s 106 1521 238 1597 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 106 1301 176 1401 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 106 915 284 1015 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 106 423 284 523 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 106 -159 238 -83 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 106 570 1272 869 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
