magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< error_p >>
rect -29 -86 29 -80
rect -29 -120 -17 -86
rect -29 -126 29 -120
<< nwell >>
rect -211 -259 211 259
<< pmos >>
rect -15 -39 15 111
<< pdiff >>
rect -73 87 -15 111
rect -73 53 -61 87
rect -27 53 -15 87
rect -73 19 -15 53
rect -73 -15 -61 19
rect -27 -15 -15 19
rect -73 -39 -15 -15
rect 15 87 73 111
rect 15 53 27 87
rect 61 53 73 87
rect 15 19 73 53
rect 15 -15 27 19
rect 61 -15 73 19
rect 15 -39 73 -15
<< pdiffc >>
rect -61 53 -27 87
rect -61 -15 -27 19
rect 27 53 61 87
rect 27 -15 61 19
<< nsubdiff >>
rect -175 189 -51 223
rect -17 189 17 223
rect 51 189 175 223
rect -175 119 -141 189
rect 141 119 175 189
rect -175 51 -141 85
rect -175 -17 -141 17
rect 141 51 175 85
rect 141 -17 175 17
rect -175 -85 -141 -51
rect -175 -189 -141 -119
rect 141 -85 175 -51
rect 141 -189 175 -119
rect -175 -223 -51 -189
rect -17 -223 17 -189
rect 51 -223 175 -189
<< nsubdiffcont >>
rect -51 189 -17 223
rect 17 189 51 223
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect 141 -119 175 -85
rect -51 -223 -17 -189
rect 17 -223 51 -189
<< poly >>
rect -15 111 15 137
rect -15 -70 15 -39
rect -33 -86 33 -70
rect -33 -120 -17 -86
rect 17 -120 33 -86
rect -33 -136 33 -120
<< polycont >>
rect -17 -120 17 -86
<< locali >>
rect -175 189 -51 223
rect -17 189 17 223
rect 51 189 175 223
rect -175 119 -141 189
rect 141 119 175 189
rect -175 51 -141 85
rect -175 -17 -141 17
rect -61 89 -27 115
rect -61 19 -27 53
rect -61 -43 -27 -17
rect 27 89 61 115
rect 27 19 61 53
rect 27 -43 61 -17
rect 141 51 175 85
rect 141 -17 175 17
rect -175 -85 -141 -51
rect 141 -85 175 -51
rect -175 -189 -141 -119
rect -33 -120 -17 -86
rect 17 -120 33 -86
rect 141 -189 175 -119
rect -175 -223 -51 -189
rect -17 -223 17 -189
rect 51 -223 175 -189
<< viali >>
rect -61 87 -27 89
rect -61 55 -27 87
rect -61 -15 -27 17
rect -61 -17 -27 -15
rect 27 87 61 89
rect 27 55 61 87
rect 27 -15 61 17
rect 27 -17 61 -15
rect -17 -120 17 -86
<< metal1 >>
rect -67 89 -21 111
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -39 -21 -17
rect 21 89 67 111
rect 21 55 27 89
rect 61 55 67 89
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -39 67 -17
rect -29 -86 29 -80
rect -29 -120 -17 -86
rect 17 -120 29 -86
rect -29 -126 29 -120
<< properties >>
string FIXED_BBOX -158 -206 158 206
<< end >>
