magic
tech sky130A
magscale 1 2
timestamp 1757832914
<< error_p >>
rect -29 -211 29 -205
rect -29 -245 -17 -211
rect -29 -251 29 -245
<< nwell >>
rect -211 -384 211 384
<< pmos >>
rect -15 -164 15 236
<< pdiff >>
rect -73 223 -15 236
rect -73 189 -61 223
rect -27 189 -15 223
rect -73 155 -15 189
rect -73 121 -61 155
rect -27 121 -15 155
rect -73 87 -15 121
rect -73 53 -61 87
rect -27 53 -15 87
rect -73 19 -15 53
rect -73 -15 -61 19
rect -27 -15 -15 19
rect -73 -49 -15 -15
rect -73 -83 -61 -49
rect -27 -83 -15 -49
rect -73 -117 -15 -83
rect -73 -151 -61 -117
rect -27 -151 -15 -117
rect -73 -164 -15 -151
rect 15 223 73 236
rect 15 189 27 223
rect 61 189 73 223
rect 15 155 73 189
rect 15 121 27 155
rect 61 121 73 155
rect 15 87 73 121
rect 15 53 27 87
rect 61 53 73 87
rect 15 19 73 53
rect 15 -15 27 19
rect 61 -15 73 19
rect 15 -49 73 -15
rect 15 -83 27 -49
rect 61 -83 73 -49
rect 15 -117 73 -83
rect 15 -151 27 -117
rect 61 -151 73 -117
rect 15 -164 73 -151
<< pdiffc >>
rect -61 189 -27 223
rect -61 121 -27 155
rect -61 53 -27 87
rect -61 -15 -27 19
rect -61 -83 -27 -49
rect -61 -151 -27 -117
rect 27 189 61 223
rect 27 121 61 155
rect 27 53 61 87
rect 27 -15 61 19
rect 27 -83 61 -49
rect 27 -151 61 -117
<< nsubdiff >>
rect -175 314 -51 348
rect -17 314 17 348
rect 51 314 175 348
rect -175 -314 -141 314
rect 141 221 175 314
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -314 175 -221
rect -175 -348 -51 -314
rect -17 -348 17 -314
rect 51 -348 175 -314
<< nsubdiffcont >>
rect -51 314 -17 348
rect 17 314 51 348
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect -51 -348 -17 -314
rect 17 -348 51 -314
<< poly >>
rect -15 236 15 262
rect -15 -195 15 -164
rect -33 -211 33 -195
rect -33 -245 -17 -211
rect 17 -245 33 -211
rect -33 -261 33 -245
<< polycont >>
rect -17 -245 17 -211
<< locali >>
rect -175 314 -51 348
rect -17 314 17 348
rect 51 314 175 348
rect -175 -314 -141 314
rect -61 223 -27 240
rect -61 155 -27 163
rect -61 87 -27 91
rect -61 -19 -27 -15
rect -61 -91 -27 -83
rect -61 -168 -27 -151
rect 27 223 61 240
rect 27 155 61 163
rect 27 87 61 91
rect 27 -19 61 -15
rect 27 -91 61 -83
rect 27 -168 61 -151
rect 141 221 175 314
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect -33 -245 -17 -211
rect 17 -245 33 -211
rect 141 -314 175 -221
rect -175 -348 -51 -314
rect -17 -348 17 -314
rect 51 -348 175 -314
<< viali >>
rect -61 189 -27 197
rect -61 163 -27 189
rect -61 121 -27 125
rect -61 91 -27 121
rect -61 19 -27 53
rect -61 -49 -27 -19
rect -61 -53 -27 -49
rect -61 -117 -27 -91
rect -61 -125 -27 -117
rect 27 189 61 197
rect 27 163 61 189
rect 27 121 61 125
rect 27 91 61 121
rect 27 19 61 53
rect 27 -49 61 -19
rect 27 -53 61 -49
rect 27 -117 61 -91
rect 27 -125 61 -117
rect -17 -245 17 -211
<< metal1 >>
rect -67 197 -21 236
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -164 -21 -125
rect 21 197 67 236
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -164 67 -125
rect -29 -211 29 -205
rect -29 -245 -17 -211
rect 17 -245 29 -211
rect -29 -251 29 -245
<< properties >>
string FIXED_BBOX -158 -331 158 331
<< end >>
