magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 -3 403
rect 31 369 69 403
rect 103 369 141 403
rect 175 369 213 403
rect 247 369 285 403
rect 319 369 357 403
rect 391 369 429 403
rect 463 369 501 403
rect 535 369 573 403
rect 607 369 645 403
rect 679 369 717 403
rect 751 369 789 403
rect 823 369 861 403
rect 895 369 933 403
rect 967 369 1005 403
rect 1039 369 1077 403
rect 1111 369 1149 403
rect 1183 369 1221 403
rect 1255 369 1293 403
rect 1327 369 1365 403
rect 1399 369 1437 403
rect 1471 369 1509 403
rect 1543 369 1581 403
rect 1615 369 1653 403
rect 1687 369 1725 403
rect 1759 369 1797 403
rect 1831 369 1869 403
rect 1903 369 1941 403
rect 1975 369 2013 403
rect 2047 369 2085 403
rect 2119 369 2157 403
rect 2191 369 2229 403
rect 2263 369 2301 403
rect 2335 369 2373 403
rect 2407 369 2445 403
rect 2479 369 2517 403
rect 2551 369 2589 403
rect 2623 369 2661 403
rect 2695 369 2733 403
rect 2767 369 2805 403
rect 2839 369 2877 403
rect 2911 369 2949 403
rect 2983 369 3021 403
rect 3055 369 3093 403
rect 3127 369 3165 403
rect 3199 369 3237 403
rect 3271 369 3309 403
rect 3343 369 3381 403
rect 3415 369 3453 403
rect 3487 369 3525 403
rect 3559 369 3597 403
rect 3631 369 3645 403
rect 3717 -17 3723 17
rect 3757 -17 3795 17
rect 3829 -17 3867 17
rect 3901 -17 3939 17
rect 3973 -17 4011 17
rect 4045 -17 4083 17
rect 4117 -17 4155 17
rect 4189 -17 4227 17
rect 4261 -17 4299 17
rect 4333 -17 4371 17
rect 4405 -17 4443 17
rect 4477 -17 4515 17
rect 4549 -17 4587 17
rect 4621 -17 4659 17
rect 4693 -17 4731 17
rect 4765 -17 4803 17
rect 4837 -17 4875 17
rect 4909 -17 4947 17
rect 4981 -17 5019 17
rect 5053 -17 5091 17
rect 5125 -17 5163 17
rect 5197 -17 5235 17
rect 5269 -17 5307 17
rect 5341 -17 5379 17
rect 5413 -17 5451 17
rect 5485 -17 5523 17
rect 5557 -17 5595 17
rect 5629 -17 5635 17
<< viali >>
rect -3 369 31 403
rect 69 369 103 403
rect 141 369 175 403
rect 213 369 247 403
rect 285 369 319 403
rect 357 369 391 403
rect 429 369 463 403
rect 501 369 535 403
rect 573 369 607 403
rect 645 369 679 403
rect 717 369 751 403
rect 789 369 823 403
rect 861 369 895 403
rect 933 369 967 403
rect 1005 369 1039 403
rect 1077 369 1111 403
rect 1149 369 1183 403
rect 1221 369 1255 403
rect 1293 369 1327 403
rect 1365 369 1399 403
rect 1437 369 1471 403
rect 1509 369 1543 403
rect 1581 369 1615 403
rect 1653 369 1687 403
rect 1725 369 1759 403
rect 1797 369 1831 403
rect 1869 369 1903 403
rect 1941 369 1975 403
rect 2013 369 2047 403
rect 2085 369 2119 403
rect 2157 369 2191 403
rect 2229 369 2263 403
rect 2301 369 2335 403
rect 2373 369 2407 403
rect 2445 369 2479 403
rect 2517 369 2551 403
rect 2589 369 2623 403
rect 2661 369 2695 403
rect 2733 369 2767 403
rect 2805 369 2839 403
rect 2877 369 2911 403
rect 2949 369 2983 403
rect 3021 369 3055 403
rect 3093 369 3127 403
rect 3165 369 3199 403
rect 3237 369 3271 403
rect 3309 369 3343 403
rect 3381 369 3415 403
rect 3453 369 3487 403
rect 3525 369 3559 403
rect 3597 369 3631 403
rect 3723 -17 3757 17
rect 3795 -17 3829 17
rect 3867 -17 3901 17
rect 3939 -17 3973 17
rect 4011 -17 4045 17
rect 4083 -17 4117 17
rect 4155 -17 4189 17
rect 4227 -17 4261 17
rect 4299 -17 4333 17
rect 4371 -17 4405 17
rect 4443 -17 4477 17
rect 4515 -17 4549 17
rect 4587 -17 4621 17
rect 4659 -17 4693 17
rect 4731 -17 4765 17
rect 4803 -17 4837 17
rect 4875 -17 4909 17
rect 4947 -17 4981 17
rect 5019 -17 5053 17
rect 5091 -17 5125 17
rect 5163 -17 5197 17
rect 5235 -17 5269 17
rect 5307 -17 5341 17
rect 5379 -17 5413 17
rect 5451 -17 5485 17
rect 5523 -17 5557 17
rect 5595 -17 5629 17
<< metal1 >>
rect -53 403 5671 439
rect -53 369 -3 403
rect 31 369 69 403
rect 103 369 141 403
rect 175 369 213 403
rect 247 369 285 403
rect 319 369 357 403
rect 391 369 429 403
rect 463 369 501 403
rect 535 369 573 403
rect 607 369 645 403
rect 679 369 717 403
rect 751 369 789 403
rect 823 369 861 403
rect 895 369 933 403
rect 967 369 1005 403
rect 1039 369 1077 403
rect 1111 369 1149 403
rect 1183 369 1221 403
rect 1255 369 1293 403
rect 1327 369 1365 403
rect 1399 369 1437 403
rect 1471 369 1509 403
rect 1543 369 1581 403
rect 1615 369 1653 403
rect 1687 369 1725 403
rect 1759 369 1797 403
rect 1831 369 1869 403
rect 1903 369 1941 403
rect 1975 369 2013 403
rect 2047 369 2085 403
rect 2119 369 2157 403
rect 2191 369 2229 403
rect 2263 369 2301 403
rect 2335 369 2373 403
rect 2407 369 2445 403
rect 2479 369 2517 403
rect 2551 369 2589 403
rect 2623 369 2661 403
rect 2695 369 2733 403
rect 2767 369 2805 403
rect 2839 369 2877 403
rect 2911 369 2949 403
rect 2983 369 3021 403
rect 3055 369 3093 403
rect 3127 369 3165 403
rect 3199 369 3237 403
rect 3271 369 3309 403
rect 3343 369 3381 403
rect 3415 369 3453 403
rect 3487 369 3525 403
rect 3559 369 3597 403
rect 3631 369 5671 403
rect -53 363 5671 369
rect -53 289 5461 323
rect -53 143 125 243
rect 5493 143 5671 243
rect 166 63 5671 97
rect -53 17 5671 23
rect -53 -17 3723 17
rect 3757 -17 3795 17
rect 3829 -17 3867 17
rect 3901 -17 3939 17
rect 3973 -17 4011 17
rect 4045 -17 4083 17
rect 4117 -17 4155 17
rect 4189 -17 4227 17
rect 4261 -17 4299 17
rect 4333 -17 4371 17
rect 4405 -17 4443 17
rect 4477 -17 4515 17
rect 4549 -17 4587 17
rect 4621 -17 4659 17
rect 4693 -17 4731 17
rect 4765 -17 4803 17
rect 4837 -17 4875 17
rect 4909 -17 4947 17
rect 4981 -17 5019 17
rect 5053 -17 5091 17
rect 5125 -17 5163 17
rect 5197 -17 5235 17
rect 5269 -17 5307 17
rect 5341 -17 5379 17
rect 5413 -17 5451 17
rect 5485 -17 5523 17
rect 5557 -17 5595 17
rect 5629 -17 5671 17
rect -53 -53 5671 -17
use sky130_fd_pr__pfet_01v8_FFQTRC  XM1
timestamp 1750100919
transform 0 1 1814 -1 0 193
box -246 -1867 246 1867
use sky130_fd_pr__nfet_01v8_4SAWNX  XM2
timestamp 1750100919
transform 0 1 4676 -1 0 193
box -236 -985 236 985
<< labels >>
flabel metal1 s -40 398 -28 407 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -36 -19 -24 -10 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -47 302 -35 311 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -41 189 -29 198 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 5649 188 5661 197 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 5649 76 5661 85 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
