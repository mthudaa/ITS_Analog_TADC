magic
tech sky130A
magscale 1 2
timestamp 1749307785
<< metal3 >>
rect -586 17772 586 17800
rect -586 16948 502 17772
rect 566 16948 586 17772
rect -586 16920 586 16948
rect -586 16652 586 16680
rect -586 15828 502 16652
rect 566 15828 586 16652
rect -586 15800 586 15828
rect -586 15532 586 15560
rect -586 14708 502 15532
rect 566 14708 586 15532
rect -586 14680 586 14708
rect -586 14412 586 14440
rect -586 13588 502 14412
rect 566 13588 586 14412
rect -586 13560 586 13588
rect -586 13292 586 13320
rect -586 12468 502 13292
rect 566 12468 586 13292
rect -586 12440 586 12468
rect -586 12172 586 12200
rect -586 11348 502 12172
rect 566 11348 586 12172
rect -586 11320 586 11348
rect -586 11052 586 11080
rect -586 10228 502 11052
rect 566 10228 586 11052
rect -586 10200 586 10228
rect -586 9932 586 9960
rect -586 9108 502 9932
rect 566 9108 586 9932
rect -586 9080 586 9108
rect -586 8812 586 8840
rect -586 7988 502 8812
rect 566 7988 586 8812
rect -586 7960 586 7988
rect -586 7692 586 7720
rect -586 6868 502 7692
rect 566 6868 586 7692
rect -586 6840 586 6868
rect -586 6572 586 6600
rect -586 5748 502 6572
rect 566 5748 586 6572
rect -586 5720 586 5748
rect -586 5452 586 5480
rect -586 4628 502 5452
rect 566 4628 586 5452
rect -586 4600 586 4628
rect -586 4332 586 4360
rect -586 3508 502 4332
rect 566 3508 586 4332
rect -586 3480 586 3508
rect -586 3212 586 3240
rect -586 2388 502 3212
rect 566 2388 586 3212
rect -586 2360 586 2388
rect -586 2092 586 2120
rect -586 1268 502 2092
rect 566 1268 586 2092
rect -586 1240 586 1268
rect -586 972 586 1000
rect -586 148 502 972
rect 566 148 586 972
rect -586 120 586 148
rect -586 -148 586 -120
rect -586 -972 502 -148
rect 566 -972 586 -148
rect -586 -1000 586 -972
rect -586 -1268 586 -1240
rect -586 -2092 502 -1268
rect 566 -2092 586 -1268
rect -586 -2120 586 -2092
rect -586 -2388 586 -2360
rect -586 -3212 502 -2388
rect 566 -3212 586 -2388
rect -586 -3240 586 -3212
rect -586 -3508 586 -3480
rect -586 -4332 502 -3508
rect 566 -4332 586 -3508
rect -586 -4360 586 -4332
rect -586 -4628 586 -4600
rect -586 -5452 502 -4628
rect 566 -5452 586 -4628
rect -586 -5480 586 -5452
rect -586 -5748 586 -5720
rect -586 -6572 502 -5748
rect 566 -6572 586 -5748
rect -586 -6600 586 -6572
rect -586 -6868 586 -6840
rect -586 -7692 502 -6868
rect 566 -7692 586 -6868
rect -586 -7720 586 -7692
rect -586 -7988 586 -7960
rect -586 -8812 502 -7988
rect 566 -8812 586 -7988
rect -586 -8840 586 -8812
rect -586 -9108 586 -9080
rect -586 -9932 502 -9108
rect 566 -9932 586 -9108
rect -586 -9960 586 -9932
rect -586 -10228 586 -10200
rect -586 -11052 502 -10228
rect 566 -11052 586 -10228
rect -586 -11080 586 -11052
rect -586 -11348 586 -11320
rect -586 -12172 502 -11348
rect 566 -12172 586 -11348
rect -586 -12200 586 -12172
rect -586 -12468 586 -12440
rect -586 -13292 502 -12468
rect 566 -13292 586 -12468
rect -586 -13320 586 -13292
rect -586 -13588 586 -13560
rect -586 -14412 502 -13588
rect 566 -14412 586 -13588
rect -586 -14440 586 -14412
rect -586 -14708 586 -14680
rect -586 -15532 502 -14708
rect 566 -15532 586 -14708
rect -586 -15560 586 -15532
rect -586 -15828 586 -15800
rect -586 -16652 502 -15828
rect 566 -16652 586 -15828
rect -586 -16680 586 -16652
rect -586 -16948 586 -16920
rect -586 -17772 502 -16948
rect 566 -17772 586 -16948
rect -586 -17800 586 -17772
<< via3 >>
rect 502 16948 566 17772
rect 502 15828 566 16652
rect 502 14708 566 15532
rect 502 13588 566 14412
rect 502 12468 566 13292
rect 502 11348 566 12172
rect 502 10228 566 11052
rect 502 9108 566 9932
rect 502 7988 566 8812
rect 502 6868 566 7692
rect 502 5748 566 6572
rect 502 4628 566 5452
rect 502 3508 566 4332
rect 502 2388 566 3212
rect 502 1268 566 2092
rect 502 148 566 972
rect 502 -972 566 -148
rect 502 -2092 566 -1268
rect 502 -3212 566 -2388
rect 502 -4332 566 -3508
rect 502 -5452 566 -4628
rect 502 -6572 566 -5748
rect 502 -7692 566 -6868
rect 502 -8812 566 -7988
rect 502 -9932 566 -9108
rect 502 -11052 566 -10228
rect 502 -12172 566 -11348
rect 502 -13292 566 -12468
rect 502 -14412 566 -13588
rect 502 -15532 566 -14708
rect 502 -16652 566 -15828
rect 502 -17772 566 -16948
<< mimcap >>
rect -546 17720 254 17760
rect -546 17000 -506 17720
rect 214 17000 254 17720
rect -546 16960 254 17000
rect -546 16600 254 16640
rect -546 15880 -506 16600
rect 214 15880 254 16600
rect -546 15840 254 15880
rect -546 15480 254 15520
rect -546 14760 -506 15480
rect 214 14760 254 15480
rect -546 14720 254 14760
rect -546 14360 254 14400
rect -546 13640 -506 14360
rect 214 13640 254 14360
rect -546 13600 254 13640
rect -546 13240 254 13280
rect -546 12520 -506 13240
rect 214 12520 254 13240
rect -546 12480 254 12520
rect -546 12120 254 12160
rect -546 11400 -506 12120
rect 214 11400 254 12120
rect -546 11360 254 11400
rect -546 11000 254 11040
rect -546 10280 -506 11000
rect 214 10280 254 11000
rect -546 10240 254 10280
rect -546 9880 254 9920
rect -546 9160 -506 9880
rect 214 9160 254 9880
rect -546 9120 254 9160
rect -546 8760 254 8800
rect -546 8040 -506 8760
rect 214 8040 254 8760
rect -546 8000 254 8040
rect -546 7640 254 7680
rect -546 6920 -506 7640
rect 214 6920 254 7640
rect -546 6880 254 6920
rect -546 6520 254 6560
rect -546 5800 -506 6520
rect 214 5800 254 6520
rect -546 5760 254 5800
rect -546 5400 254 5440
rect -546 4680 -506 5400
rect 214 4680 254 5400
rect -546 4640 254 4680
rect -546 4280 254 4320
rect -546 3560 -506 4280
rect 214 3560 254 4280
rect -546 3520 254 3560
rect -546 3160 254 3200
rect -546 2440 -506 3160
rect 214 2440 254 3160
rect -546 2400 254 2440
rect -546 2040 254 2080
rect -546 1320 -506 2040
rect 214 1320 254 2040
rect -546 1280 254 1320
rect -546 920 254 960
rect -546 200 -506 920
rect 214 200 254 920
rect -546 160 254 200
rect -546 -200 254 -160
rect -546 -920 -506 -200
rect 214 -920 254 -200
rect -546 -960 254 -920
rect -546 -1320 254 -1280
rect -546 -2040 -506 -1320
rect 214 -2040 254 -1320
rect -546 -2080 254 -2040
rect -546 -2440 254 -2400
rect -546 -3160 -506 -2440
rect 214 -3160 254 -2440
rect -546 -3200 254 -3160
rect -546 -3560 254 -3520
rect -546 -4280 -506 -3560
rect 214 -4280 254 -3560
rect -546 -4320 254 -4280
rect -546 -4680 254 -4640
rect -546 -5400 -506 -4680
rect 214 -5400 254 -4680
rect -546 -5440 254 -5400
rect -546 -5800 254 -5760
rect -546 -6520 -506 -5800
rect 214 -6520 254 -5800
rect -546 -6560 254 -6520
rect -546 -6920 254 -6880
rect -546 -7640 -506 -6920
rect 214 -7640 254 -6920
rect -546 -7680 254 -7640
rect -546 -8040 254 -8000
rect -546 -8760 -506 -8040
rect 214 -8760 254 -8040
rect -546 -8800 254 -8760
rect -546 -9160 254 -9120
rect -546 -9880 -506 -9160
rect 214 -9880 254 -9160
rect -546 -9920 254 -9880
rect -546 -10280 254 -10240
rect -546 -11000 -506 -10280
rect 214 -11000 254 -10280
rect -546 -11040 254 -11000
rect -546 -11400 254 -11360
rect -546 -12120 -506 -11400
rect 214 -12120 254 -11400
rect -546 -12160 254 -12120
rect -546 -12520 254 -12480
rect -546 -13240 -506 -12520
rect 214 -13240 254 -12520
rect -546 -13280 254 -13240
rect -546 -13640 254 -13600
rect -546 -14360 -506 -13640
rect 214 -14360 254 -13640
rect -546 -14400 254 -14360
rect -546 -14760 254 -14720
rect -546 -15480 -506 -14760
rect 214 -15480 254 -14760
rect -546 -15520 254 -15480
rect -546 -15880 254 -15840
rect -546 -16600 -506 -15880
rect 214 -16600 254 -15880
rect -546 -16640 254 -16600
rect -546 -17000 254 -16960
rect -546 -17720 -506 -17000
rect 214 -17720 254 -17000
rect -546 -17760 254 -17720
<< mimcapcontact >>
rect -506 17000 214 17720
rect -506 15880 214 16600
rect -506 14760 214 15480
rect -506 13640 214 14360
rect -506 12520 214 13240
rect -506 11400 214 12120
rect -506 10280 214 11000
rect -506 9160 214 9880
rect -506 8040 214 8760
rect -506 6920 214 7640
rect -506 5800 214 6520
rect -506 4680 214 5400
rect -506 3560 214 4280
rect -506 2440 214 3160
rect -506 1320 214 2040
rect -506 200 214 920
rect -506 -920 214 -200
rect -506 -2040 214 -1320
rect -506 -3160 214 -2440
rect -506 -4280 214 -3560
rect -506 -5400 214 -4680
rect -506 -6520 214 -5800
rect -506 -7640 214 -6920
rect -506 -8760 214 -8040
rect -506 -9880 214 -9160
rect -506 -11000 214 -10280
rect -506 -12120 214 -11400
rect -506 -13240 214 -12520
rect -506 -14360 214 -13640
rect -506 -15480 214 -14760
rect -506 -16600 214 -15880
rect -506 -17720 214 -17000
<< metal4 >>
rect -198 17721 -94 17920
rect 482 17772 586 17920
rect -507 17720 215 17721
rect -507 17000 -506 17720
rect 214 17000 215 17720
rect -507 16999 215 17000
rect -198 16601 -94 16999
rect 482 16948 502 17772
rect 566 16948 586 17772
rect 482 16652 586 16948
rect -507 16600 215 16601
rect -507 15880 -506 16600
rect 214 15880 215 16600
rect -507 15879 215 15880
rect -198 15481 -94 15879
rect 482 15828 502 16652
rect 566 15828 586 16652
rect 482 15532 586 15828
rect -507 15480 215 15481
rect -507 14760 -506 15480
rect 214 14760 215 15480
rect -507 14759 215 14760
rect -198 14361 -94 14759
rect 482 14708 502 15532
rect 566 14708 586 15532
rect 482 14412 586 14708
rect -507 14360 215 14361
rect -507 13640 -506 14360
rect 214 13640 215 14360
rect -507 13639 215 13640
rect -198 13241 -94 13639
rect 482 13588 502 14412
rect 566 13588 586 14412
rect 482 13292 586 13588
rect -507 13240 215 13241
rect -507 12520 -506 13240
rect 214 12520 215 13240
rect -507 12519 215 12520
rect -198 12121 -94 12519
rect 482 12468 502 13292
rect 566 12468 586 13292
rect 482 12172 586 12468
rect -507 12120 215 12121
rect -507 11400 -506 12120
rect 214 11400 215 12120
rect -507 11399 215 11400
rect -198 11001 -94 11399
rect 482 11348 502 12172
rect 566 11348 586 12172
rect 482 11052 586 11348
rect -507 11000 215 11001
rect -507 10280 -506 11000
rect 214 10280 215 11000
rect -507 10279 215 10280
rect -198 9881 -94 10279
rect 482 10228 502 11052
rect 566 10228 586 11052
rect 482 9932 586 10228
rect -507 9880 215 9881
rect -507 9160 -506 9880
rect 214 9160 215 9880
rect -507 9159 215 9160
rect -198 8761 -94 9159
rect 482 9108 502 9932
rect 566 9108 586 9932
rect 482 8812 586 9108
rect -507 8760 215 8761
rect -507 8040 -506 8760
rect 214 8040 215 8760
rect -507 8039 215 8040
rect -198 7641 -94 8039
rect 482 7988 502 8812
rect 566 7988 586 8812
rect 482 7692 586 7988
rect -507 7640 215 7641
rect -507 6920 -506 7640
rect 214 6920 215 7640
rect -507 6919 215 6920
rect -198 6521 -94 6919
rect 482 6868 502 7692
rect 566 6868 586 7692
rect 482 6572 586 6868
rect -507 6520 215 6521
rect -507 5800 -506 6520
rect 214 5800 215 6520
rect -507 5799 215 5800
rect -198 5401 -94 5799
rect 482 5748 502 6572
rect 566 5748 586 6572
rect 482 5452 586 5748
rect -507 5400 215 5401
rect -507 4680 -506 5400
rect 214 4680 215 5400
rect -507 4679 215 4680
rect -198 4281 -94 4679
rect 482 4628 502 5452
rect 566 4628 586 5452
rect 482 4332 586 4628
rect -507 4280 215 4281
rect -507 3560 -506 4280
rect 214 3560 215 4280
rect -507 3559 215 3560
rect -198 3161 -94 3559
rect 482 3508 502 4332
rect 566 3508 586 4332
rect 482 3212 586 3508
rect -507 3160 215 3161
rect -507 2440 -506 3160
rect 214 2440 215 3160
rect -507 2439 215 2440
rect -198 2041 -94 2439
rect 482 2388 502 3212
rect 566 2388 586 3212
rect 482 2092 586 2388
rect -507 2040 215 2041
rect -507 1320 -506 2040
rect 214 1320 215 2040
rect -507 1319 215 1320
rect -198 921 -94 1319
rect 482 1268 502 2092
rect 566 1268 586 2092
rect 482 972 586 1268
rect -507 920 215 921
rect -507 200 -506 920
rect 214 200 215 920
rect -507 199 215 200
rect -198 -199 -94 199
rect 482 148 502 972
rect 566 148 586 972
rect 482 -148 586 148
rect -507 -200 215 -199
rect -507 -920 -506 -200
rect 214 -920 215 -200
rect -507 -921 215 -920
rect -198 -1319 -94 -921
rect 482 -972 502 -148
rect 566 -972 586 -148
rect 482 -1268 586 -972
rect -507 -1320 215 -1319
rect -507 -2040 -506 -1320
rect 214 -2040 215 -1320
rect -507 -2041 215 -2040
rect -198 -2439 -94 -2041
rect 482 -2092 502 -1268
rect 566 -2092 586 -1268
rect 482 -2388 586 -2092
rect -507 -2440 215 -2439
rect -507 -3160 -506 -2440
rect 214 -3160 215 -2440
rect -507 -3161 215 -3160
rect -198 -3559 -94 -3161
rect 482 -3212 502 -2388
rect 566 -3212 586 -2388
rect 482 -3508 586 -3212
rect -507 -3560 215 -3559
rect -507 -4280 -506 -3560
rect 214 -4280 215 -3560
rect -507 -4281 215 -4280
rect -198 -4679 -94 -4281
rect 482 -4332 502 -3508
rect 566 -4332 586 -3508
rect 482 -4628 586 -4332
rect -507 -4680 215 -4679
rect -507 -5400 -506 -4680
rect 214 -5400 215 -4680
rect -507 -5401 215 -5400
rect -198 -5799 -94 -5401
rect 482 -5452 502 -4628
rect 566 -5452 586 -4628
rect 482 -5748 586 -5452
rect -507 -5800 215 -5799
rect -507 -6520 -506 -5800
rect 214 -6520 215 -5800
rect -507 -6521 215 -6520
rect -198 -6919 -94 -6521
rect 482 -6572 502 -5748
rect 566 -6572 586 -5748
rect 482 -6868 586 -6572
rect -507 -6920 215 -6919
rect -507 -7640 -506 -6920
rect 214 -7640 215 -6920
rect -507 -7641 215 -7640
rect -198 -8039 -94 -7641
rect 482 -7692 502 -6868
rect 566 -7692 586 -6868
rect 482 -7988 586 -7692
rect -507 -8040 215 -8039
rect -507 -8760 -506 -8040
rect 214 -8760 215 -8040
rect -507 -8761 215 -8760
rect -198 -9159 -94 -8761
rect 482 -8812 502 -7988
rect 566 -8812 586 -7988
rect 482 -9108 586 -8812
rect -507 -9160 215 -9159
rect -507 -9880 -506 -9160
rect 214 -9880 215 -9160
rect -507 -9881 215 -9880
rect -198 -10279 -94 -9881
rect 482 -9932 502 -9108
rect 566 -9932 586 -9108
rect 482 -10228 586 -9932
rect -507 -10280 215 -10279
rect -507 -11000 -506 -10280
rect 214 -11000 215 -10280
rect -507 -11001 215 -11000
rect -198 -11399 -94 -11001
rect 482 -11052 502 -10228
rect 566 -11052 586 -10228
rect 482 -11348 586 -11052
rect -507 -11400 215 -11399
rect -507 -12120 -506 -11400
rect 214 -12120 215 -11400
rect -507 -12121 215 -12120
rect -198 -12519 -94 -12121
rect 482 -12172 502 -11348
rect 566 -12172 586 -11348
rect 482 -12468 586 -12172
rect -507 -12520 215 -12519
rect -507 -13240 -506 -12520
rect 214 -13240 215 -12520
rect -507 -13241 215 -13240
rect -198 -13639 -94 -13241
rect 482 -13292 502 -12468
rect 566 -13292 586 -12468
rect 482 -13588 586 -13292
rect -507 -13640 215 -13639
rect -507 -14360 -506 -13640
rect 214 -14360 215 -13640
rect -507 -14361 215 -14360
rect -198 -14759 -94 -14361
rect 482 -14412 502 -13588
rect 566 -14412 586 -13588
rect 482 -14708 586 -14412
rect -507 -14760 215 -14759
rect -507 -15480 -506 -14760
rect 214 -15480 215 -14760
rect -507 -15481 215 -15480
rect -198 -15879 -94 -15481
rect 482 -15532 502 -14708
rect 566 -15532 586 -14708
rect 482 -15828 586 -15532
rect -507 -15880 215 -15879
rect -507 -16600 -506 -15880
rect 214 -16600 215 -15880
rect -507 -16601 215 -16600
rect -198 -16999 -94 -16601
rect 482 -16652 502 -15828
rect 566 -16652 586 -15828
rect 482 -16948 586 -16652
rect -507 -17000 215 -16999
rect -507 -17720 -506 -17000
rect 214 -17720 215 -17000
rect -507 -17721 215 -17720
rect -198 -17920 -94 -17721
rect 482 -17772 502 -16948
rect 566 -17772 586 -16948
rect 482 -17920 586 -17772
<< properties >>
string FIXED_BBOX -586 16920 294 17800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 1 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
