magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -194 -364 194 398
<< pmos >>
rect -100 -264 100 336
<< pdiff >>
rect -158 291 -100 336
rect -158 257 -146 291
rect -112 257 -100 291
rect -158 223 -100 257
rect -158 189 -146 223
rect -112 189 -100 223
rect -158 155 -100 189
rect -158 121 -146 155
rect -112 121 -100 155
rect -158 87 -100 121
rect -158 53 -146 87
rect -112 53 -100 87
rect -158 19 -100 53
rect -158 -15 -146 19
rect -112 -15 -100 19
rect -158 -49 -100 -15
rect -158 -83 -146 -49
rect -112 -83 -100 -49
rect -158 -117 -100 -83
rect -158 -151 -146 -117
rect -112 -151 -100 -117
rect -158 -185 -100 -151
rect -158 -219 -146 -185
rect -112 -219 -100 -185
rect -158 -264 -100 -219
rect 100 291 158 336
rect 100 257 112 291
rect 146 257 158 291
rect 100 223 158 257
rect 100 189 112 223
rect 146 189 158 223
rect 100 155 158 189
rect 100 121 112 155
rect 146 121 158 155
rect 100 87 158 121
rect 100 53 112 87
rect 146 53 158 87
rect 100 19 158 53
rect 100 -15 112 19
rect 146 -15 158 19
rect 100 -49 158 -15
rect 100 -83 112 -49
rect 146 -83 158 -49
rect 100 -117 158 -83
rect 100 -151 112 -117
rect 146 -151 158 -117
rect 100 -185 158 -151
rect 100 -219 112 -185
rect 146 -219 158 -185
rect 100 -264 158 -219
<< pdiffc >>
rect -146 257 -112 291
rect -146 189 -112 223
rect -146 121 -112 155
rect -146 53 -112 87
rect -146 -15 -112 19
rect -146 -83 -112 -49
rect -146 -151 -112 -117
rect -146 -219 -112 -185
rect 112 257 146 291
rect 112 189 146 223
rect 112 121 146 155
rect 112 53 146 87
rect 112 -15 146 19
rect 112 -83 146 -49
rect 112 -151 146 -117
rect 112 -219 146 -185
<< poly >>
rect -100 336 100 362
rect -100 -311 100 -264
rect -100 -328 -17 -311
rect -58 -345 -17 -328
rect 17 -328 100 -311
rect 17 -345 58 -328
rect -58 -361 58 -345
<< polycont >>
rect -17 -345 17 -311
<< locali >>
rect -146 305 -112 340
rect -146 233 -112 257
rect -146 161 -112 189
rect -146 89 -112 121
rect -146 19 -112 53
rect -146 -49 -112 -17
rect -146 -117 -112 -89
rect -146 -185 -112 -161
rect -146 -268 -112 -233
rect 112 305 146 340
rect 112 233 146 257
rect 112 161 146 189
rect 112 89 146 121
rect 112 19 146 53
rect 112 -49 146 -17
rect 112 -117 146 -89
rect 112 -185 146 -161
rect 112 -268 146 -233
rect -58 -345 -17 -311
rect 17 -345 58 -311
<< viali >>
rect -146 291 -112 305
rect -146 271 -112 291
rect -146 223 -112 233
rect -146 199 -112 223
rect -146 155 -112 161
rect -146 127 -112 155
rect -146 87 -112 89
rect -146 55 -112 87
rect -146 -15 -112 17
rect -146 -17 -112 -15
rect -146 -83 -112 -55
rect -146 -89 -112 -83
rect -146 -151 -112 -127
rect -146 -161 -112 -151
rect -146 -219 -112 -199
rect -146 -233 -112 -219
rect 112 291 146 305
rect 112 271 146 291
rect 112 223 146 233
rect 112 199 146 223
rect 112 155 146 161
rect 112 127 146 155
rect 112 87 146 89
rect 112 55 146 87
rect 112 -15 146 17
rect 112 -17 146 -15
rect 112 -83 146 -55
rect 112 -89 146 -83
rect 112 -151 146 -127
rect 112 -161 146 -151
rect 112 -219 146 -199
rect 112 -233 146 -219
rect -17 -345 17 -311
<< metal1 >>
rect -152 305 -106 336
rect -152 271 -146 305
rect -112 271 -106 305
rect -152 233 -106 271
rect -152 199 -146 233
rect -112 199 -106 233
rect -152 161 -106 199
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -199 -106 -161
rect -152 -233 -146 -199
rect -112 -233 -106 -199
rect -152 -264 -106 -233
rect 106 305 152 336
rect 106 271 112 305
rect 146 271 152 305
rect 106 233 152 271
rect 106 199 112 233
rect 146 199 152 233
rect 106 161 152 199
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -199 152 -161
rect 106 -233 112 -199
rect 146 -233 152 -199
rect 106 -264 152 -233
rect -54 -311 54 -305
rect -54 -345 -17 -311
rect 17 -345 54 -311
rect -54 -351 54 -345
<< end >>
