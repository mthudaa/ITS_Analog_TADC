magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 17 403
rect 51 369 89 403
rect 123 369 161 403
rect 195 369 233 403
rect 267 369 305 403
rect 339 369 377 403
rect 411 369 449 403
rect 483 369 521 403
rect 555 369 593 403
rect 627 369 665 403
rect 699 369 737 403
rect 771 369 809 403
rect 843 369 881 403
rect 915 369 953 403
rect 987 369 1025 403
rect 1059 369 1097 403
rect 1131 369 1169 403
rect 1203 369 1241 403
rect 1275 369 1313 403
rect 1347 369 1385 403
rect 1419 369 1457 403
rect 1491 369 1529 403
rect 1563 369 1601 403
rect 1635 369 1673 403
rect 1707 369 1745 403
rect 1779 369 1817 403
rect 1851 369 1889 403
rect 1923 369 1961 403
rect 1995 369 2033 403
rect 2067 369 2105 403
rect 2139 369 2177 403
rect 2211 369 2249 403
rect 2283 369 2321 403
rect 2355 369 2393 403
rect 2427 369 2465 403
rect 2499 369 2537 403
rect 2571 369 2609 403
rect 2643 369 2681 403
rect 2715 369 2753 403
rect 2787 369 2825 403
rect 2859 369 2897 403
rect 2931 369 2969 403
rect 3003 369 3041 403
rect 3075 369 3113 403
rect 3147 369 3185 403
rect 3219 369 3257 403
rect 3291 369 3329 403
rect 3363 369 3401 403
rect 3435 369 3473 403
rect 3507 369 3545 403
rect 3579 369 3617 403
rect 3651 369 3689 403
rect 3723 369 3761 403
rect 3795 369 3833 403
rect 3867 369 3905 403
rect 3939 369 3977 403
rect 4011 369 4049 403
rect 4083 369 4121 403
rect 4155 369 4193 403
rect 4227 369 4265 403
rect 4299 369 4337 403
rect 4371 369 4409 403
rect 4443 369 4481 403
rect 4515 369 4553 403
rect 4587 369 4625 403
rect 4659 369 4697 403
rect 4731 369 4769 403
rect 4803 369 4841 403
rect 4875 369 4913 403
rect 4947 369 4985 403
rect 5019 369 5057 403
rect 5091 369 5129 403
rect 5163 369 5201 403
rect 5235 369 5273 403
rect 5307 369 5345 403
rect 5379 369 5417 403
rect 5451 369 5489 403
rect 5523 369 5561 403
rect 5595 369 5633 403
rect 5667 369 5705 403
rect 5739 369 5777 403
rect 5811 369 5849 403
rect 5883 369 5921 403
rect 5955 369 5993 403
rect 6027 369 6065 403
rect 6099 369 6137 403
rect 6171 369 6209 403
rect 6243 369 6281 403
rect 6315 369 6353 403
rect 6387 369 6425 403
rect 6459 369 6497 403
rect 6531 369 6569 403
rect 6603 369 6641 403
rect 6675 369 6713 403
rect 6747 369 6785 403
rect 6819 369 6857 403
rect 6891 369 6929 403
rect 6963 369 7001 403
rect 7035 369 7069 403
rect 7141 -17 7159 17
rect 7193 -17 7231 17
rect 7265 -17 7303 17
rect 7337 -17 7375 17
rect 7409 -17 7447 17
rect 7481 -17 7519 17
rect 7553 -17 7591 17
rect 7625 -17 7663 17
rect 7697 -17 7735 17
rect 7769 -17 7807 17
rect 7841 -17 7879 17
rect 7913 -17 7951 17
rect 7985 -17 8023 17
rect 8057 -17 8095 17
rect 8129 -17 8167 17
rect 8201 -17 8239 17
rect 8273 -17 8311 17
rect 8345 -17 8383 17
rect 8417 -17 8455 17
rect 8489 -17 8527 17
rect 8561 -17 8599 17
rect 8633 -17 8671 17
rect 8705 -17 8743 17
rect 8777 -17 8815 17
rect 8849 -17 8887 17
rect 8921 -17 8959 17
rect 8993 -17 9031 17
rect 9065 -17 9103 17
rect 9137 -17 9175 17
rect 9209 -17 9247 17
rect 9281 -17 9319 17
rect 9353 -17 9391 17
rect 9425 -17 9463 17
rect 9497 -17 9535 17
rect 9569 -17 9607 17
rect 9641 -17 9679 17
rect 9713 -17 9751 17
rect 9785 -17 9823 17
rect 9857 -17 9895 17
rect 9929 -17 9967 17
rect 10001 -17 10039 17
rect 10073 -17 10111 17
rect 10145 -17 10183 17
rect 10217 -17 10255 17
rect 10289 -17 10327 17
rect 10361 -17 10399 17
rect 10433 -17 10471 17
rect 10505 -17 10543 17
rect 10577 -17 10615 17
rect 10649 -17 10687 17
rect 10721 -17 10739 17
<< viali >>
rect 17 369 51 403
rect 89 369 123 403
rect 161 369 195 403
rect 233 369 267 403
rect 305 369 339 403
rect 377 369 411 403
rect 449 369 483 403
rect 521 369 555 403
rect 593 369 627 403
rect 665 369 699 403
rect 737 369 771 403
rect 809 369 843 403
rect 881 369 915 403
rect 953 369 987 403
rect 1025 369 1059 403
rect 1097 369 1131 403
rect 1169 369 1203 403
rect 1241 369 1275 403
rect 1313 369 1347 403
rect 1385 369 1419 403
rect 1457 369 1491 403
rect 1529 369 1563 403
rect 1601 369 1635 403
rect 1673 369 1707 403
rect 1745 369 1779 403
rect 1817 369 1851 403
rect 1889 369 1923 403
rect 1961 369 1995 403
rect 2033 369 2067 403
rect 2105 369 2139 403
rect 2177 369 2211 403
rect 2249 369 2283 403
rect 2321 369 2355 403
rect 2393 369 2427 403
rect 2465 369 2499 403
rect 2537 369 2571 403
rect 2609 369 2643 403
rect 2681 369 2715 403
rect 2753 369 2787 403
rect 2825 369 2859 403
rect 2897 369 2931 403
rect 2969 369 3003 403
rect 3041 369 3075 403
rect 3113 369 3147 403
rect 3185 369 3219 403
rect 3257 369 3291 403
rect 3329 369 3363 403
rect 3401 369 3435 403
rect 3473 369 3507 403
rect 3545 369 3579 403
rect 3617 369 3651 403
rect 3689 369 3723 403
rect 3761 369 3795 403
rect 3833 369 3867 403
rect 3905 369 3939 403
rect 3977 369 4011 403
rect 4049 369 4083 403
rect 4121 369 4155 403
rect 4193 369 4227 403
rect 4265 369 4299 403
rect 4337 369 4371 403
rect 4409 369 4443 403
rect 4481 369 4515 403
rect 4553 369 4587 403
rect 4625 369 4659 403
rect 4697 369 4731 403
rect 4769 369 4803 403
rect 4841 369 4875 403
rect 4913 369 4947 403
rect 4985 369 5019 403
rect 5057 369 5091 403
rect 5129 369 5163 403
rect 5201 369 5235 403
rect 5273 369 5307 403
rect 5345 369 5379 403
rect 5417 369 5451 403
rect 5489 369 5523 403
rect 5561 369 5595 403
rect 5633 369 5667 403
rect 5705 369 5739 403
rect 5777 369 5811 403
rect 5849 369 5883 403
rect 5921 369 5955 403
rect 5993 369 6027 403
rect 6065 369 6099 403
rect 6137 369 6171 403
rect 6209 369 6243 403
rect 6281 369 6315 403
rect 6353 369 6387 403
rect 6425 369 6459 403
rect 6497 369 6531 403
rect 6569 369 6603 403
rect 6641 369 6675 403
rect 6713 369 6747 403
rect 6785 369 6819 403
rect 6857 369 6891 403
rect 6929 369 6963 403
rect 7001 369 7035 403
rect 7159 -17 7193 17
rect 7231 -17 7265 17
rect 7303 -17 7337 17
rect 7375 -17 7409 17
rect 7447 -17 7481 17
rect 7519 -17 7553 17
rect 7591 -17 7625 17
rect 7663 -17 7697 17
rect 7735 -17 7769 17
rect 7807 -17 7841 17
rect 7879 -17 7913 17
rect 7951 -17 7985 17
rect 8023 -17 8057 17
rect 8095 -17 8129 17
rect 8167 -17 8201 17
rect 8239 -17 8273 17
rect 8311 -17 8345 17
rect 8383 -17 8417 17
rect 8455 -17 8489 17
rect 8527 -17 8561 17
rect 8599 -17 8633 17
rect 8671 -17 8705 17
rect 8743 -17 8777 17
rect 8815 -17 8849 17
rect 8887 -17 8921 17
rect 8959 -17 8993 17
rect 9031 -17 9065 17
rect 9103 -17 9137 17
rect 9175 -17 9209 17
rect 9247 -17 9281 17
rect 9319 -17 9353 17
rect 9391 -17 9425 17
rect 9463 -17 9497 17
rect 9535 -17 9569 17
rect 9607 -17 9641 17
rect 9679 -17 9713 17
rect 9751 -17 9785 17
rect 9823 -17 9857 17
rect 9895 -17 9929 17
rect 9967 -17 10001 17
rect 10039 -17 10073 17
rect 10111 -17 10145 17
rect 10183 -17 10217 17
rect 10255 -17 10289 17
rect 10327 -17 10361 17
rect 10399 -17 10433 17
rect 10471 -17 10505 17
rect 10543 -17 10577 17
rect 10615 -17 10649 17
rect 10687 -17 10721 17
<< metal1 >>
rect -53 403 10775 439
rect -53 369 17 403
rect 51 369 89 403
rect 123 369 161 403
rect 195 369 233 403
rect 267 369 305 403
rect 339 369 377 403
rect 411 369 449 403
rect 483 369 521 403
rect 555 369 593 403
rect 627 369 665 403
rect 699 369 737 403
rect 771 369 809 403
rect 843 369 881 403
rect 915 369 953 403
rect 987 369 1025 403
rect 1059 369 1097 403
rect 1131 369 1169 403
rect 1203 369 1241 403
rect 1275 369 1313 403
rect 1347 369 1385 403
rect 1419 369 1457 403
rect 1491 369 1529 403
rect 1563 369 1601 403
rect 1635 369 1673 403
rect 1707 369 1745 403
rect 1779 369 1817 403
rect 1851 369 1889 403
rect 1923 369 1961 403
rect 1995 369 2033 403
rect 2067 369 2105 403
rect 2139 369 2177 403
rect 2211 369 2249 403
rect 2283 369 2321 403
rect 2355 369 2393 403
rect 2427 369 2465 403
rect 2499 369 2537 403
rect 2571 369 2609 403
rect 2643 369 2681 403
rect 2715 369 2753 403
rect 2787 369 2825 403
rect 2859 369 2897 403
rect 2931 369 2969 403
rect 3003 369 3041 403
rect 3075 369 3113 403
rect 3147 369 3185 403
rect 3219 369 3257 403
rect 3291 369 3329 403
rect 3363 369 3401 403
rect 3435 369 3473 403
rect 3507 369 3545 403
rect 3579 369 3617 403
rect 3651 369 3689 403
rect 3723 369 3761 403
rect 3795 369 3833 403
rect 3867 369 3905 403
rect 3939 369 3977 403
rect 4011 369 4049 403
rect 4083 369 4121 403
rect 4155 369 4193 403
rect 4227 369 4265 403
rect 4299 369 4337 403
rect 4371 369 4409 403
rect 4443 369 4481 403
rect 4515 369 4553 403
rect 4587 369 4625 403
rect 4659 369 4697 403
rect 4731 369 4769 403
rect 4803 369 4841 403
rect 4875 369 4913 403
rect 4947 369 4985 403
rect 5019 369 5057 403
rect 5091 369 5129 403
rect 5163 369 5201 403
rect 5235 369 5273 403
rect 5307 369 5345 403
rect 5379 369 5417 403
rect 5451 369 5489 403
rect 5523 369 5561 403
rect 5595 369 5633 403
rect 5667 369 5705 403
rect 5739 369 5777 403
rect 5811 369 5849 403
rect 5883 369 5921 403
rect 5955 369 5993 403
rect 6027 369 6065 403
rect 6099 369 6137 403
rect 6171 369 6209 403
rect 6243 369 6281 403
rect 6315 369 6353 403
rect 6387 369 6425 403
rect 6459 369 6497 403
rect 6531 369 6569 403
rect 6603 369 6641 403
rect 6675 369 6713 403
rect 6747 369 6785 403
rect 6819 369 6857 403
rect 6891 369 6929 403
rect 6963 369 7001 403
rect 7035 369 10775 403
rect -53 363 10775 369
rect -53 289 10565 323
rect -53 147 125 239
rect 10597 147 10775 239
rect 166 63 10775 97
rect -53 17 10775 23
rect -53 -17 7159 17
rect 7193 -17 7231 17
rect 7265 -17 7303 17
rect 7337 -17 7375 17
rect 7409 -17 7447 17
rect 7481 -17 7519 17
rect 7553 -17 7591 17
rect 7625 -17 7663 17
rect 7697 -17 7735 17
rect 7769 -17 7807 17
rect 7841 -17 7879 17
rect 7913 -17 7951 17
rect 7985 -17 8023 17
rect 8057 -17 8095 17
rect 8129 -17 8167 17
rect 8201 -17 8239 17
rect 8273 -17 8311 17
rect 8345 -17 8383 17
rect 8417 -17 8455 17
rect 8489 -17 8527 17
rect 8561 -17 8599 17
rect 8633 -17 8671 17
rect 8705 -17 8743 17
rect 8777 -17 8815 17
rect 8849 -17 8887 17
rect 8921 -17 8959 17
rect 8993 -17 9031 17
rect 9065 -17 9103 17
rect 9137 -17 9175 17
rect 9209 -17 9247 17
rect 9281 -17 9319 17
rect 9353 -17 9391 17
rect 9425 -17 9463 17
rect 9497 -17 9535 17
rect 9569 -17 9607 17
rect 9641 -17 9679 17
rect 9713 -17 9751 17
rect 9785 -17 9823 17
rect 9857 -17 9895 17
rect 9929 -17 9967 17
rect 10001 -17 10039 17
rect 10073 -17 10111 17
rect 10145 -17 10183 17
rect 10217 -17 10255 17
rect 10289 -17 10327 17
rect 10361 -17 10399 17
rect 10433 -17 10471 17
rect 10505 -17 10543 17
rect 10577 -17 10615 17
rect 10649 -17 10687 17
rect 10721 -17 10775 17
rect -53 -53 10775 -17
use sky130_fd_pr__pfet_01v8_D9Q5W2  XM1
timestamp 1750100919
transform 0 1 3526 -1 0 193
box -246 -3579 246 3579
use sky130_fd_pr__nfet_01v8_K9ZN2D  XM2
timestamp 1750100919
transform 0 1 8940 -1 0 193
box -236 -1825 236 1825
<< labels >>
flabel metal1 s -38 405 -26 413 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -44 -31 -32 -23 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -39 303 -27 311 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -42 186 -30 194 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 10751 187 10763 195 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 10756 76 10768 84 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
