magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< metal3 >>
rect -586 8812 586 8840
rect -586 7988 502 8812
rect 566 7988 586 8812
rect -586 7960 586 7988
rect -586 7692 586 7720
rect -586 6868 502 7692
rect 566 6868 586 7692
rect -586 6840 586 6868
rect -586 6572 586 6600
rect -586 5748 502 6572
rect 566 5748 586 6572
rect -586 5720 586 5748
rect -586 5452 586 5480
rect -586 4628 502 5452
rect 566 4628 586 5452
rect -586 4600 586 4628
rect -586 4332 586 4360
rect -586 3508 502 4332
rect 566 3508 586 4332
rect -586 3480 586 3508
rect -586 3212 586 3240
rect -586 2388 502 3212
rect 566 2388 586 3212
rect -586 2360 586 2388
rect -586 2092 586 2120
rect -586 1268 502 2092
rect 566 1268 586 2092
rect -586 1240 586 1268
rect -586 972 586 1000
rect -586 148 502 972
rect 566 148 586 972
rect -586 120 586 148
rect -586 -148 586 -120
rect -586 -972 502 -148
rect 566 -972 586 -148
rect -586 -1000 586 -972
rect -586 -1268 586 -1240
rect -586 -2092 502 -1268
rect 566 -2092 586 -1268
rect -586 -2120 586 -2092
rect -586 -2388 586 -2360
rect -586 -3212 502 -2388
rect 566 -3212 586 -2388
rect -586 -3240 586 -3212
rect -586 -3508 586 -3480
rect -586 -4332 502 -3508
rect 566 -4332 586 -3508
rect -586 -4360 586 -4332
rect -586 -4628 586 -4600
rect -586 -5452 502 -4628
rect 566 -5452 586 -4628
rect -586 -5480 586 -5452
rect -586 -5748 586 -5720
rect -586 -6572 502 -5748
rect 566 -6572 586 -5748
rect -586 -6600 586 -6572
rect -586 -6868 586 -6840
rect -586 -7692 502 -6868
rect 566 -7692 586 -6868
rect -586 -7720 586 -7692
rect -586 -7988 586 -7960
rect -586 -8812 502 -7988
rect 566 -8812 586 -7988
rect -586 -8840 586 -8812
<< via3 >>
rect 502 7988 566 8812
rect 502 6868 566 7692
rect 502 5748 566 6572
rect 502 4628 566 5452
rect 502 3508 566 4332
rect 502 2388 566 3212
rect 502 1268 566 2092
rect 502 148 566 972
rect 502 -972 566 -148
rect 502 -2092 566 -1268
rect 502 -3212 566 -2388
rect 502 -4332 566 -3508
rect 502 -5452 566 -4628
rect 502 -6572 566 -5748
rect 502 -7692 566 -6868
rect 502 -8812 566 -7988
<< mimcap >>
rect -546 8760 254 8800
rect -546 8040 -506 8760
rect 214 8040 254 8760
rect -546 8000 254 8040
rect -546 7640 254 7680
rect -546 6920 -506 7640
rect 214 6920 254 7640
rect -546 6880 254 6920
rect -546 6520 254 6560
rect -546 5800 -506 6520
rect 214 5800 254 6520
rect -546 5760 254 5800
rect -546 5400 254 5440
rect -546 4680 -506 5400
rect 214 4680 254 5400
rect -546 4640 254 4680
rect -546 4280 254 4320
rect -546 3560 -506 4280
rect 214 3560 254 4280
rect -546 3520 254 3560
rect -546 3160 254 3200
rect -546 2440 -506 3160
rect 214 2440 254 3160
rect -546 2400 254 2440
rect -546 2040 254 2080
rect -546 1320 -506 2040
rect 214 1320 254 2040
rect -546 1280 254 1320
rect -546 920 254 960
rect -546 200 -506 920
rect 214 200 254 920
rect -546 160 254 200
rect -546 -200 254 -160
rect -546 -920 -506 -200
rect 214 -920 254 -200
rect -546 -960 254 -920
rect -546 -1320 254 -1280
rect -546 -2040 -506 -1320
rect 214 -2040 254 -1320
rect -546 -2080 254 -2040
rect -546 -2440 254 -2400
rect -546 -3160 -506 -2440
rect 214 -3160 254 -2440
rect -546 -3200 254 -3160
rect -546 -3560 254 -3520
rect -546 -4280 -506 -3560
rect 214 -4280 254 -3560
rect -546 -4320 254 -4280
rect -546 -4680 254 -4640
rect -546 -5400 -506 -4680
rect 214 -5400 254 -4680
rect -546 -5440 254 -5400
rect -546 -5800 254 -5760
rect -546 -6520 -506 -5800
rect 214 -6520 254 -5800
rect -546 -6560 254 -6520
rect -546 -6920 254 -6880
rect -546 -7640 -506 -6920
rect 214 -7640 254 -6920
rect -546 -7680 254 -7640
rect -546 -8040 254 -8000
rect -546 -8760 -506 -8040
rect 214 -8760 254 -8040
rect -546 -8800 254 -8760
<< mimcapcontact >>
rect -506 8040 214 8760
rect -506 6920 214 7640
rect -506 5800 214 6520
rect -506 4680 214 5400
rect -506 3560 214 4280
rect -506 2440 214 3160
rect -506 1320 214 2040
rect -506 200 214 920
rect -506 -920 214 -200
rect -506 -2040 214 -1320
rect -506 -3160 214 -2440
rect -506 -4280 214 -3560
rect -506 -5400 214 -4680
rect -506 -6520 214 -5800
rect -506 -7640 214 -6920
rect -506 -8760 214 -8040
<< metal4 >>
rect -198 8761 -94 8960
rect 482 8812 586 8960
rect -507 8760 215 8761
rect -507 8040 -506 8760
rect 214 8040 215 8760
rect -507 8039 215 8040
rect -198 7641 -94 8039
rect 482 7988 502 8812
rect 566 7988 586 8812
rect 482 7692 586 7988
rect -507 7640 215 7641
rect -507 6920 -506 7640
rect 214 6920 215 7640
rect -507 6919 215 6920
rect -198 6521 -94 6919
rect 482 6868 502 7692
rect 566 6868 586 7692
rect 482 6572 586 6868
rect -507 6520 215 6521
rect -507 5800 -506 6520
rect 214 5800 215 6520
rect -507 5799 215 5800
rect -198 5401 -94 5799
rect 482 5748 502 6572
rect 566 5748 586 6572
rect 482 5452 586 5748
rect -507 5400 215 5401
rect -507 4680 -506 5400
rect 214 4680 215 5400
rect -507 4679 215 4680
rect -198 4281 -94 4679
rect 482 4628 502 5452
rect 566 4628 586 5452
rect 482 4332 586 4628
rect -507 4280 215 4281
rect -507 3560 -506 4280
rect 214 3560 215 4280
rect -507 3559 215 3560
rect -198 3161 -94 3559
rect 482 3508 502 4332
rect 566 3508 586 4332
rect 482 3212 586 3508
rect -507 3160 215 3161
rect -507 2440 -506 3160
rect 214 2440 215 3160
rect -507 2439 215 2440
rect -198 2041 -94 2439
rect 482 2388 502 3212
rect 566 2388 586 3212
rect 482 2092 586 2388
rect -507 2040 215 2041
rect -507 1320 -506 2040
rect 214 1320 215 2040
rect -507 1319 215 1320
rect -198 921 -94 1319
rect 482 1268 502 2092
rect 566 1268 586 2092
rect 482 972 586 1268
rect -507 920 215 921
rect -507 200 -506 920
rect 214 200 215 920
rect -507 199 215 200
rect -198 -199 -94 199
rect 482 148 502 972
rect 566 148 586 972
rect 482 -148 586 148
rect -507 -200 215 -199
rect -507 -920 -506 -200
rect 214 -920 215 -200
rect -507 -921 215 -920
rect -198 -1319 -94 -921
rect 482 -972 502 -148
rect 566 -972 586 -148
rect 482 -1268 586 -972
rect -507 -1320 215 -1319
rect -507 -2040 -506 -1320
rect 214 -2040 215 -1320
rect -507 -2041 215 -2040
rect -198 -2439 -94 -2041
rect 482 -2092 502 -1268
rect 566 -2092 586 -1268
rect 482 -2388 586 -2092
rect -507 -2440 215 -2439
rect -507 -3160 -506 -2440
rect 214 -3160 215 -2440
rect -507 -3161 215 -3160
rect -198 -3559 -94 -3161
rect 482 -3212 502 -2388
rect 566 -3212 586 -2388
rect 482 -3508 586 -3212
rect -507 -3560 215 -3559
rect -507 -4280 -506 -3560
rect 214 -4280 215 -3560
rect -507 -4281 215 -4280
rect -198 -4679 -94 -4281
rect 482 -4332 502 -3508
rect 566 -4332 586 -3508
rect 482 -4628 586 -4332
rect -507 -4680 215 -4679
rect -507 -5400 -506 -4680
rect 214 -5400 215 -4680
rect -507 -5401 215 -5400
rect -198 -5799 -94 -5401
rect 482 -5452 502 -4628
rect 566 -5452 586 -4628
rect 482 -5748 586 -5452
rect -507 -5800 215 -5799
rect -507 -6520 -506 -5800
rect 214 -6520 215 -5800
rect -507 -6521 215 -6520
rect -198 -6919 -94 -6521
rect 482 -6572 502 -5748
rect 566 -6572 586 -5748
rect 482 -6868 586 -6572
rect -507 -6920 215 -6919
rect -507 -7640 -506 -6920
rect 214 -7640 215 -6920
rect -507 -7641 215 -7640
rect -198 -8039 -94 -7641
rect 482 -7692 502 -6868
rect 566 -7692 586 -6868
rect 482 -7988 586 -7692
rect -507 -8040 215 -8039
rect -507 -8760 -506 -8040
rect 214 -8760 215 -8040
rect -507 -8761 215 -8760
rect -198 -8960 -94 -8761
rect 482 -8812 502 -7988
rect 566 -8812 586 -7988
rect 482 -8960 586 -8812
<< properties >>
string FIXED_BBOX -586 7960 294 8840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
