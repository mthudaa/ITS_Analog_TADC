magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< metal3 >>
rect -586 4892 586 4920
rect -586 4068 502 4892
rect 566 4068 586 4892
rect -586 4040 586 4068
rect -586 3772 586 3800
rect -586 2948 502 3772
rect 566 2948 586 3772
rect -586 2920 586 2948
rect -586 2652 586 2680
rect -586 1828 502 2652
rect 566 1828 586 2652
rect -586 1800 586 1828
rect -586 1532 586 1560
rect -586 708 502 1532
rect 566 708 586 1532
rect -586 680 586 708
rect -586 412 586 440
rect -586 -412 502 412
rect 566 -412 586 412
rect -586 -440 586 -412
rect -586 -708 586 -680
rect -586 -1532 502 -708
rect 566 -1532 586 -708
rect -586 -1560 586 -1532
rect -586 -1828 586 -1800
rect -586 -2652 502 -1828
rect 566 -2652 586 -1828
rect -586 -2680 586 -2652
rect -586 -2948 586 -2920
rect -586 -3772 502 -2948
rect 566 -3772 586 -2948
rect -586 -3800 586 -3772
rect -586 -4068 586 -4040
rect -586 -4892 502 -4068
rect 566 -4892 586 -4068
rect -586 -4920 586 -4892
<< via3 >>
rect 502 4068 566 4892
rect 502 2948 566 3772
rect 502 1828 566 2652
rect 502 708 566 1532
rect 502 -412 566 412
rect 502 -1532 566 -708
rect 502 -2652 566 -1828
rect 502 -3772 566 -2948
rect 502 -4892 566 -4068
<< mimcap >>
rect -546 4840 254 4880
rect -546 4120 -506 4840
rect 214 4120 254 4840
rect -546 4080 254 4120
rect -546 3720 254 3760
rect -546 3000 -506 3720
rect 214 3000 254 3720
rect -546 2960 254 3000
rect -546 2600 254 2640
rect -546 1880 -506 2600
rect 214 1880 254 2600
rect -546 1840 254 1880
rect -546 1480 254 1520
rect -546 760 -506 1480
rect 214 760 254 1480
rect -546 720 254 760
rect -546 360 254 400
rect -546 -360 -506 360
rect 214 -360 254 360
rect -546 -400 254 -360
rect -546 -760 254 -720
rect -546 -1480 -506 -760
rect 214 -1480 254 -760
rect -546 -1520 254 -1480
rect -546 -1880 254 -1840
rect -546 -2600 -506 -1880
rect 214 -2600 254 -1880
rect -546 -2640 254 -2600
rect -546 -3000 254 -2960
rect -546 -3720 -506 -3000
rect 214 -3720 254 -3000
rect -546 -3760 254 -3720
rect -546 -4120 254 -4080
rect -546 -4840 -506 -4120
rect 214 -4840 254 -4120
rect -546 -4880 254 -4840
<< mimcapcontact >>
rect -506 4120 214 4840
rect -506 3000 214 3720
rect -506 1880 214 2600
rect -506 760 214 1480
rect -506 -360 214 360
rect -506 -1480 214 -760
rect -506 -2600 214 -1880
rect -506 -3720 214 -3000
rect -506 -4840 214 -4120
<< metal4 >>
rect -198 4841 -94 5040
rect 482 4892 586 5040
rect -507 4840 215 4841
rect -507 4120 -506 4840
rect 214 4120 215 4840
rect -507 4119 215 4120
rect -198 3721 -94 4119
rect 482 4068 502 4892
rect 566 4068 586 4892
rect 482 3772 586 4068
rect -507 3720 215 3721
rect -507 3000 -506 3720
rect 214 3000 215 3720
rect -507 2999 215 3000
rect -198 2601 -94 2999
rect 482 2948 502 3772
rect 566 2948 586 3772
rect 482 2652 586 2948
rect -507 2600 215 2601
rect -507 1880 -506 2600
rect 214 1880 215 2600
rect -507 1879 215 1880
rect -198 1481 -94 1879
rect 482 1828 502 2652
rect 566 1828 586 2652
rect 482 1532 586 1828
rect -507 1480 215 1481
rect -507 760 -506 1480
rect 214 760 215 1480
rect -507 759 215 760
rect -198 361 -94 759
rect 482 708 502 1532
rect 566 708 586 1532
rect 482 412 586 708
rect -507 360 215 361
rect -507 -360 -506 360
rect 214 -360 215 360
rect -507 -361 215 -360
rect -198 -759 -94 -361
rect 482 -412 502 412
rect 566 -412 586 412
rect 482 -708 586 -412
rect -507 -760 215 -759
rect -507 -1480 -506 -760
rect 214 -1480 215 -760
rect -507 -1481 215 -1480
rect -198 -1879 -94 -1481
rect 482 -1532 502 -708
rect 566 -1532 586 -708
rect 482 -1828 586 -1532
rect -507 -1880 215 -1879
rect -507 -2600 -506 -1880
rect 214 -2600 215 -1880
rect -507 -2601 215 -2600
rect -198 -2999 -94 -2601
rect 482 -2652 502 -1828
rect 566 -2652 586 -1828
rect 482 -2948 586 -2652
rect -507 -3000 215 -2999
rect -507 -3720 -506 -3000
rect 214 -3720 215 -3000
rect -507 -3721 215 -3720
rect -198 -4119 -94 -3721
rect 482 -3772 502 -2948
rect 566 -3772 586 -2948
rect 482 -4068 586 -3772
rect -507 -4120 215 -4119
rect -507 -4840 -506 -4120
rect 214 -4840 215 -4120
rect -507 -4841 215 -4840
rect -198 -5040 -94 -4841
rect 482 -4892 502 -4068
rect 566 -4892 586 -4068
rect 482 -5040 586 -4892
<< properties >>
string FIXED_BBOX -586 4040 294 4920
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
