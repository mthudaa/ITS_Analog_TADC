magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< pwell >>
rect -236 -355 236 355
<< nmos >>
rect -50 55 50 155
rect -50 -155 50 -55
<< ndiff >>
rect -108 122 -50 155
rect -108 88 -96 122
rect -62 88 -50 122
rect -108 55 -50 88
rect 50 122 108 155
rect 50 88 62 122
rect 96 88 108 122
rect 50 55 108 88
rect -108 -88 -50 -55
rect -108 -122 -96 -88
rect -62 -122 -50 -88
rect -108 -155 -50 -122
rect 50 -88 108 -55
rect 50 -122 62 -88
rect 96 -122 108 -88
rect 50 -155 108 -122
<< ndiffc >>
rect -96 88 -62 122
rect 62 88 96 122
rect -96 -122 -62 -88
rect 62 -122 96 -88
<< psubdiff >>
rect -210 295 -85 329
rect -51 295 -17 329
rect 17 295 51 329
rect 85 295 210 329
rect -210 221 -176 295
rect -210 153 -176 187
rect 176 221 210 295
rect -210 85 -176 119
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect 176 -119 210 -85
rect -210 -295 -176 -221
rect 176 -187 210 -153
rect 176 -295 210 -221
rect -210 -329 -85 -295
rect -51 -329 -17 -295
rect 17 -329 51 -295
rect 85 -329 210 -295
<< psubdiffcont >>
rect -85 295 -51 329
rect -17 295 17 329
rect 51 295 85 329
rect -210 187 -176 221
rect 176 187 210 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect 176 -85 210 -51
rect 176 -153 210 -119
rect -210 -221 -176 -187
rect 176 -221 210 -187
rect -85 -329 -51 -295
rect -17 -329 17 -295
rect 51 -329 85 -295
<< poly >>
rect -50 227 50 243
rect -50 193 -17 227
rect 17 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect -50 -243 50 -227
<< polycont >>
rect -17 193 17 227
rect -17 -17 17 17
rect -17 -227 17 -193
<< locali >>
rect -210 295 -85 329
rect -51 295 -17 329
rect 17 295 51 329
rect 85 295 210 329
rect -210 221 -176 295
rect -50 193 -17 227
rect 17 193 50 227
rect 176 221 210 295
rect -210 153 -176 187
rect -210 85 -176 119
rect -96 122 -62 159
rect -96 51 -62 88
rect 62 122 96 159
rect 62 51 96 88
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect 176 17 210 51
rect -50 -17 -17 17
rect 17 -17 50 17
rect -210 -51 -176 -17
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -96 -88 -62 -51
rect -96 -159 -62 -122
rect 62 -88 96 -51
rect 62 -159 96 -122
rect 176 -119 210 -85
rect 176 -187 210 -153
rect -210 -295 -176 -221
rect -50 -227 -17 -193
rect 17 -227 50 -193
rect 176 -295 210 -221
rect -210 -329 -85 -295
rect -51 -329 -17 -295
rect 17 -329 51 -295
rect 85 -329 210 -295
<< viali >>
rect -17 193 17 227
rect -96 88 -62 122
rect 62 88 96 122
rect -17 -17 17 17
rect -96 -122 -62 -88
rect 62 -122 96 -88
rect -17 -227 17 -193
<< metal1 >>
rect -46 227 46 233
rect -46 193 -17 227
rect 17 193 46 227
rect -46 187 46 193
rect -102 122 -56 155
rect -102 88 -96 122
rect -62 88 -56 122
rect -102 55 -56 88
rect 56 122 102 155
rect 56 88 62 122
rect 96 88 102 122
rect 56 55 102 88
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -88 -56 -55
rect -102 -122 -96 -88
rect -62 -122 -56 -88
rect -102 -155 -56 -122
rect 56 -88 102 -55
rect 56 -122 62 -88
rect 96 -122 102 -88
rect 56 -155 102 -122
rect -46 -193 46 -187
rect -46 -227 -17 -193
rect 17 -227 46 -193
rect -46 -233 46 -227
<< properties >>
string FIXED_BBOX -193 -312 193 312
<< end >>
