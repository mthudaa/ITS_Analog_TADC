magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal1 >>
rect -269 116208 -149 116232
rect -269 116156 -235 116208
rect -183 116156 -149 116208
rect -269 116132 -149 116156
rect -259 114192 -159 116132
rect -59 114192 41 116437
rect 4533 116008 4653 116032
rect 4533 115956 4567 116008
rect 4619 115956 4653 116008
rect 4533 115932 4653 115956
rect 4543 114192 4643 115932
rect 4743 114192 4843 116437
rect 9345 115821 9445 115832
rect 9335 115797 9455 115821
rect 9335 115745 9369 115797
rect 9421 115745 9455 115797
rect 9335 115721 9455 115745
rect 9345 114192 9445 115721
rect 9545 114192 9645 116437
rect 14147 115619 14247 115632
rect 14137 115595 14257 115619
rect 14137 115543 14171 115595
rect 14223 115543 14257 115595
rect 14137 115519 14257 115543
rect 14147 114192 14247 115519
rect 14347 114302 14447 116437
rect 18949 115427 19049 115432
rect 18939 115403 19059 115427
rect 18939 115351 18973 115403
rect 19025 115351 19059 115403
rect 18939 115327 19059 115351
rect 14346 114192 14447 114302
rect 18949 114192 19049 115327
rect 19149 114192 19249 116437
rect 23741 115208 23861 115232
rect 23741 115156 23775 115208
rect 23827 115156 23861 115208
rect 23741 115132 23861 115156
rect 23751 114192 23851 115132
rect 23951 114192 24051 116437
rect 28543 115008 28663 115032
rect 28543 114956 28577 115008
rect 28629 114956 28663 115008
rect 28543 114932 28663 114956
rect 28553 114192 28653 114932
rect 28753 114192 28853 116437
rect 33345 114808 33465 114832
rect 33345 114756 33379 114808
rect 33431 114756 33465 114808
rect 33345 114732 33465 114756
rect 33355 114192 33455 114732
rect 33555 114192 33655 116437
rect 38147 114608 38267 114632
rect 38147 114556 38181 114608
rect 38233 114556 38267 114608
rect 38147 114532 38267 114556
rect 38157 114192 38257 114532
rect 38357 114192 38457 116437
rect 42949 114408 43069 114432
rect 42949 114356 42983 114408
rect 43035 114356 43069 114408
rect 42949 114332 43069 114356
rect 42959 114192 43059 114332
rect 43159 114192 43259 116437
rect -258 -400 -158 1640
rect -268 -424 -148 -400
rect -268 -476 -234 -424
rect -182 -476 -148 -424
rect -268 -500 -148 -476
rect -58 -705 42 1440
rect 4544 -200 4644 1640
rect 4534 -224 4654 -200
rect 4534 -276 4568 -224
rect 4620 -276 4654 -224
rect 4534 -300 4654 -276
rect 4744 -705 4844 1440
rect 9346 11 9446 1640
rect 9336 -13 9456 11
rect 9336 -65 9370 -13
rect 9422 -65 9456 -13
rect 9336 -89 9456 -65
rect 9346 -100 9446 -89
rect 9546 -705 9646 1440
rect 14148 213 14248 1640
rect 14138 189 14258 213
rect 14138 137 14172 189
rect 14224 137 14258 189
rect 14138 113 14258 137
rect 14148 100 14248 113
rect 14348 -705 14448 1440
rect 18950 405 19050 1640
rect 18940 381 19060 405
rect 18940 329 18974 381
rect 19026 329 19060 381
rect 18940 305 19060 329
rect 18950 300 19050 305
rect 19150 -705 19250 1440
rect 23752 600 23852 1640
rect 23742 576 23862 600
rect 23742 524 23776 576
rect 23828 524 23862 576
rect 23742 500 23862 524
rect 23952 -705 24052 1440
rect 28554 800 28654 1640
rect 28544 776 28664 800
rect 28544 724 28578 776
rect 28630 724 28664 776
rect 28544 700 28664 724
rect 28754 -705 28854 1440
rect 33356 1000 33456 1640
rect 33346 976 33466 1000
rect 33346 924 33380 976
rect 33432 924 33466 976
rect 33346 900 33466 924
rect 33556 -705 33656 1436
rect 38158 1200 38258 1640
rect 38148 1176 38268 1200
rect 38148 1124 38182 1176
rect 38234 1124 38268 1176
rect 38148 1100 38268 1124
rect 38358 -705 38458 1440
rect 42960 1400 43060 1640
rect 42950 1376 43070 1400
rect 42950 1324 42984 1376
rect 43036 1324 43070 1376
rect 42950 1300 43070 1324
rect 43160 -705 43260 1440
<< via1 >>
rect -235 116156 -183 116208
rect 4567 115956 4619 116008
rect 9369 115745 9421 115797
rect 14171 115543 14223 115595
rect 18973 115351 19025 115403
rect 23775 115156 23827 115208
rect 28577 114956 28629 115008
rect 33379 114756 33431 114808
rect 38181 114556 38233 114608
rect 42983 114356 43035 114408
rect -234 -476 -182 -424
rect 4568 -276 4620 -224
rect 9370 -65 9422 -13
rect 14172 137 14224 189
rect 18974 329 19026 381
rect 23776 524 23828 576
rect 28578 724 28630 776
rect 33380 924 33432 976
rect 38182 1124 38234 1176
rect 42984 1324 43036 1376
<< metal2 >>
rect -259 116232 -159 116242
rect -259 116208 50471 116232
rect -259 116156 -235 116208
rect -183 116156 50471 116208
rect -259 116132 50471 116156
rect -259 116122 -159 116132
rect 4543 116032 4643 116042
rect 4543 116008 50271 116032
rect 4543 115956 4567 116008
rect 4619 115956 50271 116008
rect 4543 115932 50271 115956
rect 4543 115922 4643 115932
rect 9345 115821 9445 115831
rect 9345 115797 50071 115821
rect 9345 115745 9369 115797
rect 9421 115745 50071 115797
rect 9345 115721 50071 115745
rect 9345 115711 9445 115721
rect 14147 115619 14247 115629
rect 14147 115595 49871 115619
rect 14147 115543 14171 115595
rect 14223 115543 49871 115595
rect 14147 115520 49871 115543
rect 14147 115519 14346 115520
rect 14147 115509 14247 115519
rect 18949 115427 19049 115437
rect 18949 115403 49671 115427
rect 18949 115351 18973 115403
rect 19025 115351 49671 115403
rect 18949 115327 49671 115351
rect 18949 115317 19049 115327
rect 23751 115232 23851 115242
rect 23751 115208 49471 115232
rect 23751 115156 23775 115208
rect 23827 115156 49471 115208
rect 23751 115132 49471 115156
rect 23751 115122 23851 115132
rect 28553 115032 28653 115042
rect 28553 115008 49271 115032
rect 28553 114956 28577 115008
rect 28629 114956 49271 115008
rect 28553 114932 49271 114956
rect 28553 114922 28653 114932
rect 33355 114832 33455 114842
rect 33355 114808 49071 114832
rect 33355 114756 33379 114808
rect 33431 114756 49071 114808
rect 33355 114732 49071 114756
rect 33355 114722 33455 114732
rect 38157 114632 38257 114642
rect 38157 114608 48871 114632
rect 38157 114556 38181 114608
rect 38233 114556 48871 114608
rect 38157 114532 48871 114556
rect 38157 114522 38257 114532
rect 42959 114432 43059 114442
rect 42959 114408 48671 114432
rect 42959 114356 42983 114408
rect 43035 114356 48671 114408
rect 42959 114332 48671 114356
rect 42959 114322 43059 114332
rect -1089 58369 -949 104859
rect -1089 58239 -948 58369
rect -1088 6313 -948 58239
rect -809 57252 -669 104803
rect -529 58311 -389 99937
rect -529 58239 -388 58311
rect -809 57052 -668 57252
rect -808 18026 -668 57052
rect -528 18124 -388 58239
rect 47771 57252 47911 112692
rect 48051 57252 48191 112892
rect 48331 57252 48471 113892
rect 48571 57252 48671 114332
rect 48771 57252 48871 114532
rect 48971 57252 49071 114732
rect 49171 57252 49271 114932
rect 49371 57252 49471 115132
rect 49571 57252 49671 115327
rect 49771 57252 49871 115520
rect 49971 57252 50071 115721
rect 50171 57252 50271 115932
rect 50371 57252 50471 116132
rect 47771 57028 47912 57252
rect 48051 57041 48192 57252
rect 47772 3040 47912 57028
rect 48052 2840 48192 57041
rect 48331 57034 48472 57252
rect 48571 57090 48672 57252
rect 48771 57114 48872 57252
rect 48332 1840 48472 57034
rect 42960 1400 43060 1410
rect 48572 1400 48672 57090
rect 42960 1376 48672 1400
rect 42960 1324 42984 1376
rect 43036 1324 48672 1376
rect 42960 1300 48672 1324
rect 42960 1290 43060 1300
rect 38158 1200 38258 1210
rect 48772 1200 48872 57114
rect 48971 57067 49072 57252
rect 49171 57137 49272 57252
rect 38158 1176 48872 1200
rect 38158 1124 38182 1176
rect 38234 1124 48872 1176
rect 38158 1100 48872 1124
rect 38158 1090 38258 1100
rect 33356 1000 33456 1010
rect 48972 1000 49072 57067
rect 33356 976 49072 1000
rect 33356 924 33380 976
rect 33432 924 49072 976
rect 33356 900 49072 924
rect 33356 890 33456 900
rect 28554 800 28654 810
rect 49172 800 49272 57137
rect 49371 57054 49472 57252
rect 49571 57160 49672 57252
rect 28554 776 49272 800
rect 28554 724 28578 776
rect 28630 724 49272 776
rect 28554 700 49272 724
rect 28554 690 28654 700
rect 23752 600 23852 610
rect 49372 600 49472 57054
rect 23752 576 49472 600
rect 23752 524 23776 576
rect 23828 524 49472 576
rect 23752 500 49472 524
rect 23752 490 23852 500
rect 18950 405 19050 415
rect 49572 405 49672 57160
rect 49771 57114 49872 57252
rect 18950 381 49672 405
rect 18950 329 18974 381
rect 19026 329 49672 381
rect 18950 305 49672 329
rect 18950 295 19050 305
rect 14148 213 14248 223
rect 14148 212 14347 213
rect 49772 212 49872 57114
rect 49971 57081 50072 57252
rect 50171 57090 50272 57252
rect 50371 57107 50472 57252
rect 14148 189 49872 212
rect 14148 137 14172 189
rect 14224 137 49872 189
rect 14148 113 49872 137
rect 14148 103 14248 113
rect 9346 11 9446 21
rect 49972 11 50072 57081
rect 9346 -13 50072 11
rect 9346 -65 9370 -13
rect 9422 -65 50072 -13
rect 9346 -89 50072 -65
rect 9346 -99 9446 -89
rect 4544 -200 4644 -190
rect 50172 -200 50272 57090
rect 4544 -224 50272 -200
rect 4544 -276 4568 -224
rect 4620 -276 50272 -224
rect 4544 -300 50272 -276
rect 4544 -310 4644 -300
rect -258 -400 -158 -390
rect 50372 -400 50472 57107
rect -258 -424 50472 -400
rect -258 -476 -234 -424
rect -182 -476 50472 -424
rect -258 -500 50472 -476
rect -258 -510 -158 -500
<< metal4 >>
rect 1898 59571 45766 59667
rect 1899 56065 45767 56161
use single_10b_cdac  single_10b_cdac_0
timestamp 1750100919
transform -1 0 47387 0 1 41235
box -1094 -40255 48486 14944
use single_10b_cdac  single_10b_cdac_1
timestamp 1750100919
transform -1 0 47387 0 -1 74497
box -1094 -40255 48486 14944
<< labels >>
flabel metal1 s 43179 116361 43239 116421 0 FreeSans 500 0 0 0 SWP_IN[0]
port 1 nsew
flabel metal1 s 38377 116359 38437 116419 0 FreeSans 500 0 0 0 SWP_IN[1]
port 2 nsew
flabel metal1 s 33574 116351 33634 116411 0 FreeSans 500 0 0 0 SWP_IN[2]
port 3 nsew
flabel metal1 s 28773 116358 28833 116418 0 FreeSans 500 0 0 0 SWP_IN[3]
port 4 nsew
flabel metal1 s 23966 116343 24026 116403 0 FreeSans 500 0 0 0 SWP_IN[4]
port 5 nsew
flabel metal1 s 19169 116339 19229 116399 0 FreeSans 500 0 0 0 SWP_IN[5]
port 6 nsew
flabel metal1 s 14366 116356 14426 116416 0 FreeSans 500 0 0 0 SWP_IN[6]
port 7 nsew
flabel metal1 s 9567 116353 9627 116413 0 FreeSans 500 0 0 0 SWP_IN[7]
port 8 nsew
flabel metal1 s 4765 116358 4825 116418 0 FreeSans 500 0 0 0 SWP_IN[8]
port 9 nsew
flabel metal1 s -38 116364 22 116424 0 FreeSans 500 0 0 0 SWP_IN[9]
port 10 nsew
flabel metal1 s 43181 -683 43241 -623 0 FreeSans 500 0 0 0 SWN_IN[0]
port 11 nsew
flabel metal1 s 38375 -683 38435 -623 0 FreeSans 500 0 0 0 SWN_IN[1]
port 12 nsew
flabel metal1 s 33571 -693 33631 -633 0 FreeSans 500 0 0 0 SWN_IN[2]
port 13 nsew
flabel metal1 s 28774 -691 28834 -631 0 FreeSans 500 0 0 0 SWN_IN[3]
port 14 nsew
flabel metal1 s 23968 -689 24028 -629 0 FreeSans 500 0 0 0 SWN_IN[4]
port 15 nsew
flabel metal1 s 19166 -687 19226 -627 0 FreeSans 500 0 0 0 SWN_IN[5]
port 16 nsew
flabel metal1 s 14366 -687 14426 -627 0 FreeSans 500 0 0 0 SWN_IN[6]
port 17 nsew
flabel metal1 s 9562 -683 9622 -623 0 FreeSans 500 0 0 0 SWN_IN[7]
port 18 nsew
flabel metal1 s 4760 -683 4820 -623 0 FreeSans 500 0 0 0 SWN_IN[8]
port 19 nsew
flabel metal1 s -42 -683 18 -623 0 FreeSans 500 0 0 0 SWN_IN[9]
port 20 nsew
flabel metal2 s 48594 1567 48654 1627 0 FreeSans 500 0 0 0 CF[0]
port 21 nsew
flabel metal2 s 48796 1577 48856 1637 0 FreeSans 500 0 0 0 CF[1]
port 22 nsew
flabel metal2 s 48992 1577 49052 1637 0 FreeSans 500 0 0 0 CF[2]
port 23 nsew
flabel metal2 s 49192 1579 49252 1639 0 FreeSans 500 0 0 0 CF[3]
port 24 nsew
flabel metal2 s 49390 1577 49450 1637 0 FreeSans 500 0 0 0 CF[4]
port 25 nsew
flabel metal2 s 49590 1571 49650 1631 0 FreeSans 500 0 0 0 CF[5]
port 26 nsew
flabel metal2 s 49790 1573 49850 1633 0 FreeSans 500 0 0 0 CF[6]
port 27 nsew
flabel metal2 s 49996 1567 50056 1627 0 FreeSans 500 0 0 0 CF[7]
port 28 nsew
flabel metal2 s 50190 1561 50250 1621 0 FreeSans 500 0 0 0 CF[8]
port 29 nsew
flabel metal2 s 50390 1563 50450 1623 0 FreeSans 500 0 0 0 CF[9]
port 30 nsew
flabel metal2 s 48373 3281 48433 3341 0 FreeSans 500 0 0 0 VCM
port 31 nsew
flabel metal2 s 48092 3275 48152 3335 0 FreeSans 500 0 0 0 VDD
port 32 nsew
flabel metal2 s 47805 3284 47865 3344 0 FreeSans 500 0 0 0 VSS
port 33 nsew
flabel metal4 s 1898 59571 1994 59667 0 FreeSans 1000 0 0 0 VCP
port 34 nsew
flabel metal4 s 1899 56065 1995 56161 0 FreeSans 1000 0 0 0 VCN
port 35 nsew
<< end >>
