magic
tech sky130A
magscale 1 2
timestamp 1757810374
<< metal3 >>
rect -892 5612 -120 5640
rect -892 5188 -204 5612
rect -140 5188 -120 5612
rect -892 5160 -120 5188
rect 120 5612 892 5640
rect 120 5188 808 5612
rect 872 5188 892 5612
rect 120 5160 892 5188
rect -892 4892 -120 4920
rect -892 4468 -204 4892
rect -140 4468 -120 4892
rect -892 4440 -120 4468
rect 120 4892 892 4920
rect 120 4468 808 4892
rect 872 4468 892 4892
rect 120 4440 892 4468
rect -892 4172 -120 4200
rect -892 3748 -204 4172
rect -140 3748 -120 4172
rect -892 3720 -120 3748
rect 120 4172 892 4200
rect 120 3748 808 4172
rect 872 3748 892 4172
rect 120 3720 892 3748
rect -892 3452 -120 3480
rect -892 3028 -204 3452
rect -140 3028 -120 3452
rect -892 3000 -120 3028
rect 120 3452 892 3480
rect 120 3028 808 3452
rect 872 3028 892 3452
rect 120 3000 892 3028
rect -892 2732 -120 2760
rect -892 2308 -204 2732
rect -140 2308 -120 2732
rect -892 2280 -120 2308
rect 120 2732 892 2760
rect 120 2308 808 2732
rect 872 2308 892 2732
rect 120 2280 892 2308
rect -892 2012 -120 2040
rect -892 1588 -204 2012
rect -140 1588 -120 2012
rect -892 1560 -120 1588
rect 120 2012 892 2040
rect 120 1588 808 2012
rect 872 1588 892 2012
rect 120 1560 892 1588
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect -892 -1588 -120 -1560
rect -892 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect -892 -2040 -120 -2012
rect 120 -1588 892 -1560
rect 120 -2012 808 -1588
rect 872 -2012 892 -1588
rect 120 -2040 892 -2012
rect -892 -2308 -120 -2280
rect -892 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect -892 -2760 -120 -2732
rect 120 -2308 892 -2280
rect 120 -2732 808 -2308
rect 872 -2732 892 -2308
rect 120 -2760 892 -2732
rect -892 -3028 -120 -3000
rect -892 -3452 -204 -3028
rect -140 -3452 -120 -3028
rect -892 -3480 -120 -3452
rect 120 -3028 892 -3000
rect 120 -3452 808 -3028
rect 872 -3452 892 -3028
rect 120 -3480 892 -3452
rect -892 -3748 -120 -3720
rect -892 -4172 -204 -3748
rect -140 -4172 -120 -3748
rect -892 -4200 -120 -4172
rect 120 -3748 892 -3720
rect 120 -4172 808 -3748
rect 872 -4172 892 -3748
rect 120 -4200 892 -4172
rect -892 -4468 -120 -4440
rect -892 -4892 -204 -4468
rect -140 -4892 -120 -4468
rect -892 -4920 -120 -4892
rect 120 -4468 892 -4440
rect 120 -4892 808 -4468
rect 872 -4892 892 -4468
rect 120 -4920 892 -4892
rect -892 -5188 -120 -5160
rect -892 -5612 -204 -5188
rect -140 -5612 -120 -5188
rect -892 -5640 -120 -5612
rect 120 -5188 892 -5160
rect 120 -5612 808 -5188
rect 872 -5612 892 -5188
rect 120 -5640 892 -5612
<< via3 >>
rect -204 5188 -140 5612
rect 808 5188 872 5612
rect -204 4468 -140 4892
rect 808 4468 872 4892
rect -204 3748 -140 4172
rect 808 3748 872 4172
rect -204 3028 -140 3452
rect 808 3028 872 3452
rect -204 2308 -140 2732
rect 808 2308 872 2732
rect -204 1588 -140 2012
rect 808 1588 872 2012
rect -204 868 -140 1292
rect 808 868 872 1292
rect -204 148 -140 572
rect 808 148 872 572
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect -204 -2012 -140 -1588
rect 808 -2012 872 -1588
rect -204 -2732 -140 -2308
rect 808 -2732 872 -2308
rect -204 -3452 -140 -3028
rect 808 -3452 872 -3028
rect -204 -4172 -140 -3748
rect 808 -4172 872 -3748
rect -204 -4892 -140 -4468
rect 808 -4892 872 -4468
rect -204 -5612 -140 -5188
rect 808 -5612 872 -5188
<< mimcap >>
rect -852 5560 -452 5600
rect -852 5240 -812 5560
rect -492 5240 -452 5560
rect -852 5200 -452 5240
rect 160 5560 560 5600
rect 160 5240 200 5560
rect 520 5240 560 5560
rect 160 5200 560 5240
rect -852 4840 -452 4880
rect -852 4520 -812 4840
rect -492 4520 -452 4840
rect -852 4480 -452 4520
rect 160 4840 560 4880
rect 160 4520 200 4840
rect 520 4520 560 4840
rect 160 4480 560 4520
rect -852 4120 -452 4160
rect -852 3800 -812 4120
rect -492 3800 -452 4120
rect -852 3760 -452 3800
rect 160 4120 560 4160
rect 160 3800 200 4120
rect 520 3800 560 4120
rect 160 3760 560 3800
rect -852 3400 -452 3440
rect -852 3080 -812 3400
rect -492 3080 -452 3400
rect -852 3040 -452 3080
rect 160 3400 560 3440
rect 160 3080 200 3400
rect 520 3080 560 3400
rect 160 3040 560 3080
rect -852 2680 -452 2720
rect -852 2360 -812 2680
rect -492 2360 -452 2680
rect -852 2320 -452 2360
rect 160 2680 560 2720
rect 160 2360 200 2680
rect 520 2360 560 2680
rect 160 2320 560 2360
rect -852 1960 -452 2000
rect -852 1640 -812 1960
rect -492 1640 -452 1960
rect -852 1600 -452 1640
rect 160 1960 560 2000
rect 160 1640 200 1960
rect 520 1640 560 1960
rect 160 1600 560 1640
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect -852 -1640 -452 -1600
rect -852 -1960 -812 -1640
rect -492 -1960 -452 -1640
rect -852 -2000 -452 -1960
rect 160 -1640 560 -1600
rect 160 -1960 200 -1640
rect 520 -1960 560 -1640
rect 160 -2000 560 -1960
rect -852 -2360 -452 -2320
rect -852 -2680 -812 -2360
rect -492 -2680 -452 -2360
rect -852 -2720 -452 -2680
rect 160 -2360 560 -2320
rect 160 -2680 200 -2360
rect 520 -2680 560 -2360
rect 160 -2720 560 -2680
rect -852 -3080 -452 -3040
rect -852 -3400 -812 -3080
rect -492 -3400 -452 -3080
rect -852 -3440 -452 -3400
rect 160 -3080 560 -3040
rect 160 -3400 200 -3080
rect 520 -3400 560 -3080
rect 160 -3440 560 -3400
rect -852 -3800 -452 -3760
rect -852 -4120 -812 -3800
rect -492 -4120 -452 -3800
rect -852 -4160 -452 -4120
rect 160 -3800 560 -3760
rect 160 -4120 200 -3800
rect 520 -4120 560 -3800
rect 160 -4160 560 -4120
rect -852 -4520 -452 -4480
rect -852 -4840 -812 -4520
rect -492 -4840 -452 -4520
rect -852 -4880 -452 -4840
rect 160 -4520 560 -4480
rect 160 -4840 200 -4520
rect 520 -4840 560 -4520
rect 160 -4880 560 -4840
rect -852 -5240 -452 -5200
rect -852 -5560 -812 -5240
rect -492 -5560 -452 -5240
rect -852 -5600 -452 -5560
rect 160 -5240 560 -5200
rect 160 -5560 200 -5240
rect 520 -5560 560 -5240
rect 160 -5600 560 -5560
<< mimcapcontact >>
rect -812 5240 -492 5560
rect 200 5240 520 5560
rect -812 4520 -492 4840
rect 200 4520 520 4840
rect -812 3800 -492 4120
rect 200 3800 520 4120
rect -812 3080 -492 3400
rect 200 3080 520 3400
rect -812 2360 -492 2680
rect 200 2360 520 2680
rect -812 1640 -492 1960
rect 200 1640 520 1960
rect -812 920 -492 1240
rect 200 920 520 1240
rect -812 200 -492 520
rect 200 200 520 520
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect -812 -1960 -492 -1640
rect 200 -1960 520 -1640
rect -812 -2680 -492 -2360
rect 200 -2680 520 -2360
rect -812 -3400 -492 -3080
rect 200 -3400 520 -3080
rect -812 -4120 -492 -3800
rect 200 -4120 520 -3800
rect -812 -4840 -492 -4520
rect 200 -4840 520 -4520
rect -812 -5560 -492 -5240
rect 200 -5560 520 -5240
<< metal4 >>
rect -704 5561 -600 5760
rect -220 5612 -124 5628
rect -813 5560 -491 5561
rect -813 5240 -812 5560
rect -492 5240 -491 5560
rect -813 5239 -491 5240
rect -704 4841 -600 5239
rect -220 5188 -204 5612
rect -140 5188 -124 5612
rect 308 5561 412 5760
rect 792 5612 888 5628
rect 199 5560 521 5561
rect 199 5240 200 5560
rect 520 5240 521 5560
rect 199 5239 521 5240
rect -220 5172 -124 5188
rect -220 4892 -124 4908
rect -813 4840 -491 4841
rect -813 4520 -812 4840
rect -492 4520 -491 4840
rect -813 4519 -491 4520
rect -704 4121 -600 4519
rect -220 4468 -204 4892
rect -140 4468 -124 4892
rect 308 4841 412 5239
rect 792 5188 808 5612
rect 872 5188 888 5612
rect 792 5172 888 5188
rect 792 4892 888 4908
rect 199 4840 521 4841
rect 199 4520 200 4840
rect 520 4520 521 4840
rect 199 4519 521 4520
rect -220 4452 -124 4468
rect -220 4172 -124 4188
rect -813 4120 -491 4121
rect -813 3800 -812 4120
rect -492 3800 -491 4120
rect -813 3799 -491 3800
rect -704 3401 -600 3799
rect -220 3748 -204 4172
rect -140 3748 -124 4172
rect 308 4121 412 4519
rect 792 4468 808 4892
rect 872 4468 888 4892
rect 792 4452 888 4468
rect 792 4172 888 4188
rect 199 4120 521 4121
rect 199 3800 200 4120
rect 520 3800 521 4120
rect 199 3799 521 3800
rect -220 3732 -124 3748
rect -220 3452 -124 3468
rect -813 3400 -491 3401
rect -813 3080 -812 3400
rect -492 3080 -491 3400
rect -813 3079 -491 3080
rect -704 2681 -600 3079
rect -220 3028 -204 3452
rect -140 3028 -124 3452
rect 308 3401 412 3799
rect 792 3748 808 4172
rect 872 3748 888 4172
rect 792 3732 888 3748
rect 792 3452 888 3468
rect 199 3400 521 3401
rect 199 3080 200 3400
rect 520 3080 521 3400
rect 199 3079 521 3080
rect -220 3012 -124 3028
rect -220 2732 -124 2748
rect -813 2680 -491 2681
rect -813 2360 -812 2680
rect -492 2360 -491 2680
rect -813 2359 -491 2360
rect -704 1961 -600 2359
rect -220 2308 -204 2732
rect -140 2308 -124 2732
rect 308 2681 412 3079
rect 792 3028 808 3452
rect 872 3028 888 3452
rect 792 3012 888 3028
rect 792 2732 888 2748
rect 199 2680 521 2681
rect 199 2360 200 2680
rect 520 2360 521 2680
rect 199 2359 521 2360
rect -220 2292 -124 2308
rect -220 2012 -124 2028
rect -813 1960 -491 1961
rect -813 1640 -812 1960
rect -492 1640 -491 1960
rect -813 1639 -491 1640
rect -704 1241 -600 1639
rect -220 1588 -204 2012
rect -140 1588 -124 2012
rect 308 1961 412 2359
rect 792 2308 808 2732
rect 872 2308 888 2732
rect 792 2292 888 2308
rect 792 2012 888 2028
rect 199 1960 521 1961
rect 199 1640 200 1960
rect 520 1640 521 1960
rect 199 1639 521 1640
rect -220 1572 -124 1588
rect -220 1292 -124 1308
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -704 521 -600 919
rect -220 868 -204 1292
rect -140 868 -124 1292
rect 308 1241 412 1639
rect 792 1588 808 2012
rect 872 1588 888 2012
rect 792 1572 888 1588
rect 792 1292 888 1308
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -220 852 -124 868
rect -220 572 -124 588
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -704 -199 -600 199
rect -220 148 -204 572
rect -140 148 -124 572
rect 308 521 412 919
rect 792 868 808 1292
rect 872 868 888 1292
rect 792 852 888 868
rect 792 572 888 588
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -220 132 -124 148
rect -220 -148 -124 -132
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -704 -919 -600 -521
rect -220 -572 -204 -148
rect -140 -572 -124 -148
rect 308 -199 412 199
rect 792 148 808 572
rect 872 148 888 572
rect 792 132 888 148
rect 792 -148 888 -132
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -220 -588 -124 -572
rect -220 -868 -124 -852
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -704 -1639 -600 -1241
rect -220 -1292 -204 -868
rect -140 -1292 -124 -868
rect 308 -919 412 -521
rect 792 -572 808 -148
rect 872 -572 888 -148
rect 792 -588 888 -572
rect 792 -868 888 -852
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -220 -1308 -124 -1292
rect -220 -1588 -124 -1572
rect -813 -1640 -491 -1639
rect -813 -1960 -812 -1640
rect -492 -1960 -491 -1640
rect -813 -1961 -491 -1960
rect -704 -2359 -600 -1961
rect -220 -2012 -204 -1588
rect -140 -2012 -124 -1588
rect 308 -1639 412 -1241
rect 792 -1292 808 -868
rect 872 -1292 888 -868
rect 792 -1308 888 -1292
rect 792 -1588 888 -1572
rect 199 -1640 521 -1639
rect 199 -1960 200 -1640
rect 520 -1960 521 -1640
rect 199 -1961 521 -1960
rect -220 -2028 -124 -2012
rect -220 -2308 -124 -2292
rect -813 -2360 -491 -2359
rect -813 -2680 -812 -2360
rect -492 -2680 -491 -2360
rect -813 -2681 -491 -2680
rect -704 -3079 -600 -2681
rect -220 -2732 -204 -2308
rect -140 -2732 -124 -2308
rect 308 -2359 412 -1961
rect 792 -2012 808 -1588
rect 872 -2012 888 -1588
rect 792 -2028 888 -2012
rect 792 -2308 888 -2292
rect 199 -2360 521 -2359
rect 199 -2680 200 -2360
rect 520 -2680 521 -2360
rect 199 -2681 521 -2680
rect -220 -2748 -124 -2732
rect -220 -3028 -124 -3012
rect -813 -3080 -491 -3079
rect -813 -3400 -812 -3080
rect -492 -3400 -491 -3080
rect -813 -3401 -491 -3400
rect -704 -3799 -600 -3401
rect -220 -3452 -204 -3028
rect -140 -3452 -124 -3028
rect 308 -3079 412 -2681
rect 792 -2732 808 -2308
rect 872 -2732 888 -2308
rect 792 -2748 888 -2732
rect 792 -3028 888 -3012
rect 199 -3080 521 -3079
rect 199 -3400 200 -3080
rect 520 -3400 521 -3080
rect 199 -3401 521 -3400
rect -220 -3468 -124 -3452
rect -220 -3748 -124 -3732
rect -813 -3800 -491 -3799
rect -813 -4120 -812 -3800
rect -492 -4120 -491 -3800
rect -813 -4121 -491 -4120
rect -704 -4519 -600 -4121
rect -220 -4172 -204 -3748
rect -140 -4172 -124 -3748
rect 308 -3799 412 -3401
rect 792 -3452 808 -3028
rect 872 -3452 888 -3028
rect 792 -3468 888 -3452
rect 792 -3748 888 -3732
rect 199 -3800 521 -3799
rect 199 -4120 200 -3800
rect 520 -4120 521 -3800
rect 199 -4121 521 -4120
rect -220 -4188 -124 -4172
rect -220 -4468 -124 -4452
rect -813 -4520 -491 -4519
rect -813 -4840 -812 -4520
rect -492 -4840 -491 -4520
rect -813 -4841 -491 -4840
rect -704 -5239 -600 -4841
rect -220 -4892 -204 -4468
rect -140 -4892 -124 -4468
rect 308 -4519 412 -4121
rect 792 -4172 808 -3748
rect 872 -4172 888 -3748
rect 792 -4188 888 -4172
rect 792 -4468 888 -4452
rect 199 -4520 521 -4519
rect 199 -4840 200 -4520
rect 520 -4840 521 -4520
rect 199 -4841 521 -4840
rect -220 -4908 -124 -4892
rect -220 -5188 -124 -5172
rect -813 -5240 -491 -5239
rect -813 -5560 -812 -5240
rect -492 -5560 -491 -5240
rect -813 -5561 -491 -5560
rect -704 -5760 -600 -5561
rect -220 -5612 -204 -5188
rect -140 -5612 -124 -5188
rect 308 -5239 412 -4841
rect 792 -4892 808 -4468
rect 872 -4892 888 -4468
rect 792 -4908 888 -4892
rect 792 -5188 888 -5172
rect 199 -5240 521 -5239
rect 199 -5560 200 -5240
rect 520 -5560 521 -5240
rect 199 -5561 521 -5560
rect -220 -5628 -124 -5612
rect 308 -5760 412 -5561
rect 792 -5612 808 -5188
rect 872 -5612 888 -5188
rect 792 -5628 888 -5612
<< properties >>
string FIXED_BBOX 120 5160 600 5640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 2 ny 16 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
