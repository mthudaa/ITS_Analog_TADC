magic
tech sky130A
magscale 1 2
timestamp 1748351693
<< error_p >>
rect -29 445 29 451
rect -29 411 -17 445
rect -29 405 29 411
<< nwell >>
rect -109 -498 109 464
<< pmos >>
rect -15 -436 15 364
<< pdiff >>
rect -73 352 -15 364
rect -73 -424 -61 352
rect -27 -424 -15 352
rect -73 -436 -15 -424
rect 15 352 73 364
rect 15 -424 27 352
rect 61 -424 73 352
rect 15 -436 73 -424
<< pdiffc >>
rect -61 -424 -27 352
rect 27 -424 61 352
<< poly >>
rect -33 445 33 461
rect -33 411 -17 445
rect 17 411 33 445
rect -33 395 33 411
rect -15 364 15 395
rect -15 -462 15 -436
<< polycont >>
rect -17 411 17 445
<< locali >>
rect -33 411 -17 445
rect 17 411 33 445
rect -61 352 -27 368
rect -61 -440 -27 -424
rect 27 352 61 368
rect 27 -440 61 -424
<< viali >>
rect -17 411 17 445
rect -61 -424 -27 352
rect 27 -424 61 352
<< metal1 >>
rect -29 445 29 451
rect -29 411 -17 445
rect 17 411 29 445
rect -29 405 29 411
rect -67 352 -21 364
rect -67 -424 -61 352
rect -27 -424 -21 352
rect -67 -436 -21 -424
rect 21 352 67 364
rect 21 -424 27 352
rect 61 -424 67 352
rect 21 -436 67 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
