magic
tech sky130A
magscale 1 2
timestamp 1748279908
<< metal3 >>
rect -17084 11732 -16312 11760
rect -17084 11308 -16396 11732
rect -16332 11308 -16312 11732
rect -17084 11280 -16312 11308
rect -16072 11732 -15300 11760
rect -16072 11308 -15384 11732
rect -15320 11308 -15300 11732
rect -16072 11280 -15300 11308
rect -15060 11732 -14288 11760
rect -15060 11308 -14372 11732
rect -14308 11308 -14288 11732
rect -15060 11280 -14288 11308
rect -14048 11732 -13276 11760
rect -14048 11308 -13360 11732
rect -13296 11308 -13276 11732
rect -14048 11280 -13276 11308
rect -13036 11732 -12264 11760
rect -13036 11308 -12348 11732
rect -12284 11308 -12264 11732
rect -13036 11280 -12264 11308
rect -12024 11732 -11252 11760
rect -12024 11308 -11336 11732
rect -11272 11308 -11252 11732
rect -12024 11280 -11252 11308
rect -11012 11732 -10240 11760
rect -11012 11308 -10324 11732
rect -10260 11308 -10240 11732
rect -11012 11280 -10240 11308
rect -10000 11732 -9228 11760
rect -10000 11308 -9312 11732
rect -9248 11308 -9228 11732
rect -10000 11280 -9228 11308
rect -8988 11732 -8216 11760
rect -8988 11308 -8300 11732
rect -8236 11308 -8216 11732
rect -8988 11280 -8216 11308
rect -7976 11732 -7204 11760
rect -7976 11308 -7288 11732
rect -7224 11308 -7204 11732
rect -7976 11280 -7204 11308
rect -6964 11732 -6192 11760
rect -6964 11308 -6276 11732
rect -6212 11308 -6192 11732
rect -6964 11280 -6192 11308
rect -5952 11732 -5180 11760
rect -5952 11308 -5264 11732
rect -5200 11308 -5180 11732
rect -5952 11280 -5180 11308
rect -4940 11732 -4168 11760
rect -4940 11308 -4252 11732
rect -4188 11308 -4168 11732
rect -4940 11280 -4168 11308
rect -3928 11732 -3156 11760
rect -3928 11308 -3240 11732
rect -3176 11308 -3156 11732
rect -3928 11280 -3156 11308
rect -2916 11732 -2144 11760
rect -2916 11308 -2228 11732
rect -2164 11308 -2144 11732
rect -2916 11280 -2144 11308
rect -1904 11732 -1132 11760
rect -1904 11308 -1216 11732
rect -1152 11308 -1132 11732
rect -1904 11280 -1132 11308
rect -892 11732 -120 11760
rect -892 11308 -204 11732
rect -140 11308 -120 11732
rect -892 11280 -120 11308
rect 120 11732 892 11760
rect 120 11308 808 11732
rect 872 11308 892 11732
rect 120 11280 892 11308
rect 1132 11732 1904 11760
rect 1132 11308 1820 11732
rect 1884 11308 1904 11732
rect 1132 11280 1904 11308
rect 2144 11732 2916 11760
rect 2144 11308 2832 11732
rect 2896 11308 2916 11732
rect 2144 11280 2916 11308
rect 3156 11732 3928 11760
rect 3156 11308 3844 11732
rect 3908 11308 3928 11732
rect 3156 11280 3928 11308
rect 4168 11732 4940 11760
rect 4168 11308 4856 11732
rect 4920 11308 4940 11732
rect 4168 11280 4940 11308
rect 5180 11732 5952 11760
rect 5180 11308 5868 11732
rect 5932 11308 5952 11732
rect 5180 11280 5952 11308
rect 6192 11732 6964 11760
rect 6192 11308 6880 11732
rect 6944 11308 6964 11732
rect 6192 11280 6964 11308
rect 7204 11732 7976 11760
rect 7204 11308 7892 11732
rect 7956 11308 7976 11732
rect 7204 11280 7976 11308
rect 8216 11732 8988 11760
rect 8216 11308 8904 11732
rect 8968 11308 8988 11732
rect 8216 11280 8988 11308
rect 9228 11732 10000 11760
rect 9228 11308 9916 11732
rect 9980 11308 10000 11732
rect 9228 11280 10000 11308
rect 10240 11732 11012 11760
rect 10240 11308 10928 11732
rect 10992 11308 11012 11732
rect 10240 11280 11012 11308
rect 11252 11732 12024 11760
rect 11252 11308 11940 11732
rect 12004 11308 12024 11732
rect 11252 11280 12024 11308
rect 12264 11732 13036 11760
rect 12264 11308 12952 11732
rect 13016 11308 13036 11732
rect 12264 11280 13036 11308
rect 13276 11732 14048 11760
rect 13276 11308 13964 11732
rect 14028 11308 14048 11732
rect 13276 11280 14048 11308
rect 14288 11732 15060 11760
rect 14288 11308 14976 11732
rect 15040 11308 15060 11732
rect 14288 11280 15060 11308
rect 15300 11732 16072 11760
rect 15300 11308 15988 11732
rect 16052 11308 16072 11732
rect 15300 11280 16072 11308
rect 16312 11732 17084 11760
rect 16312 11308 17000 11732
rect 17064 11308 17084 11732
rect 16312 11280 17084 11308
rect -17084 11012 -16312 11040
rect -17084 10588 -16396 11012
rect -16332 10588 -16312 11012
rect -17084 10560 -16312 10588
rect -16072 11012 -15300 11040
rect -16072 10588 -15384 11012
rect -15320 10588 -15300 11012
rect -16072 10560 -15300 10588
rect -15060 11012 -14288 11040
rect -15060 10588 -14372 11012
rect -14308 10588 -14288 11012
rect -15060 10560 -14288 10588
rect -14048 11012 -13276 11040
rect -14048 10588 -13360 11012
rect -13296 10588 -13276 11012
rect -14048 10560 -13276 10588
rect -13036 11012 -12264 11040
rect -13036 10588 -12348 11012
rect -12284 10588 -12264 11012
rect -13036 10560 -12264 10588
rect -12024 11012 -11252 11040
rect -12024 10588 -11336 11012
rect -11272 10588 -11252 11012
rect -12024 10560 -11252 10588
rect -11012 11012 -10240 11040
rect -11012 10588 -10324 11012
rect -10260 10588 -10240 11012
rect -11012 10560 -10240 10588
rect -10000 11012 -9228 11040
rect -10000 10588 -9312 11012
rect -9248 10588 -9228 11012
rect -10000 10560 -9228 10588
rect -8988 11012 -8216 11040
rect -8988 10588 -8300 11012
rect -8236 10588 -8216 11012
rect -8988 10560 -8216 10588
rect -7976 11012 -7204 11040
rect -7976 10588 -7288 11012
rect -7224 10588 -7204 11012
rect -7976 10560 -7204 10588
rect -6964 11012 -6192 11040
rect -6964 10588 -6276 11012
rect -6212 10588 -6192 11012
rect -6964 10560 -6192 10588
rect -5952 11012 -5180 11040
rect -5952 10588 -5264 11012
rect -5200 10588 -5180 11012
rect -5952 10560 -5180 10588
rect -4940 11012 -4168 11040
rect -4940 10588 -4252 11012
rect -4188 10588 -4168 11012
rect -4940 10560 -4168 10588
rect -3928 11012 -3156 11040
rect -3928 10588 -3240 11012
rect -3176 10588 -3156 11012
rect -3928 10560 -3156 10588
rect -2916 11012 -2144 11040
rect -2916 10588 -2228 11012
rect -2164 10588 -2144 11012
rect -2916 10560 -2144 10588
rect -1904 11012 -1132 11040
rect -1904 10588 -1216 11012
rect -1152 10588 -1132 11012
rect -1904 10560 -1132 10588
rect -892 11012 -120 11040
rect -892 10588 -204 11012
rect -140 10588 -120 11012
rect -892 10560 -120 10588
rect 120 11012 892 11040
rect 120 10588 808 11012
rect 872 10588 892 11012
rect 120 10560 892 10588
rect 1132 11012 1904 11040
rect 1132 10588 1820 11012
rect 1884 10588 1904 11012
rect 1132 10560 1904 10588
rect 2144 11012 2916 11040
rect 2144 10588 2832 11012
rect 2896 10588 2916 11012
rect 2144 10560 2916 10588
rect 3156 11012 3928 11040
rect 3156 10588 3844 11012
rect 3908 10588 3928 11012
rect 3156 10560 3928 10588
rect 4168 11012 4940 11040
rect 4168 10588 4856 11012
rect 4920 10588 4940 11012
rect 4168 10560 4940 10588
rect 5180 11012 5952 11040
rect 5180 10588 5868 11012
rect 5932 10588 5952 11012
rect 5180 10560 5952 10588
rect 6192 11012 6964 11040
rect 6192 10588 6880 11012
rect 6944 10588 6964 11012
rect 6192 10560 6964 10588
rect 7204 11012 7976 11040
rect 7204 10588 7892 11012
rect 7956 10588 7976 11012
rect 7204 10560 7976 10588
rect 8216 11012 8988 11040
rect 8216 10588 8904 11012
rect 8968 10588 8988 11012
rect 8216 10560 8988 10588
rect 9228 11012 10000 11040
rect 9228 10588 9916 11012
rect 9980 10588 10000 11012
rect 9228 10560 10000 10588
rect 10240 11012 11012 11040
rect 10240 10588 10928 11012
rect 10992 10588 11012 11012
rect 10240 10560 11012 10588
rect 11252 11012 12024 11040
rect 11252 10588 11940 11012
rect 12004 10588 12024 11012
rect 11252 10560 12024 10588
rect 12264 11012 13036 11040
rect 12264 10588 12952 11012
rect 13016 10588 13036 11012
rect 12264 10560 13036 10588
rect 13276 11012 14048 11040
rect 13276 10588 13964 11012
rect 14028 10588 14048 11012
rect 13276 10560 14048 10588
rect 14288 11012 15060 11040
rect 14288 10588 14976 11012
rect 15040 10588 15060 11012
rect 14288 10560 15060 10588
rect 15300 11012 16072 11040
rect 15300 10588 15988 11012
rect 16052 10588 16072 11012
rect 15300 10560 16072 10588
rect 16312 11012 17084 11040
rect 16312 10588 17000 11012
rect 17064 10588 17084 11012
rect 16312 10560 17084 10588
rect -17084 10292 -16312 10320
rect -17084 9868 -16396 10292
rect -16332 9868 -16312 10292
rect -17084 9840 -16312 9868
rect -16072 10292 -15300 10320
rect -16072 9868 -15384 10292
rect -15320 9868 -15300 10292
rect -16072 9840 -15300 9868
rect -15060 10292 -14288 10320
rect -15060 9868 -14372 10292
rect -14308 9868 -14288 10292
rect -15060 9840 -14288 9868
rect -14048 10292 -13276 10320
rect -14048 9868 -13360 10292
rect -13296 9868 -13276 10292
rect -14048 9840 -13276 9868
rect -13036 10292 -12264 10320
rect -13036 9868 -12348 10292
rect -12284 9868 -12264 10292
rect -13036 9840 -12264 9868
rect -12024 10292 -11252 10320
rect -12024 9868 -11336 10292
rect -11272 9868 -11252 10292
rect -12024 9840 -11252 9868
rect -11012 10292 -10240 10320
rect -11012 9868 -10324 10292
rect -10260 9868 -10240 10292
rect -11012 9840 -10240 9868
rect -10000 10292 -9228 10320
rect -10000 9868 -9312 10292
rect -9248 9868 -9228 10292
rect -10000 9840 -9228 9868
rect -8988 10292 -8216 10320
rect -8988 9868 -8300 10292
rect -8236 9868 -8216 10292
rect -8988 9840 -8216 9868
rect -7976 10292 -7204 10320
rect -7976 9868 -7288 10292
rect -7224 9868 -7204 10292
rect -7976 9840 -7204 9868
rect -6964 10292 -6192 10320
rect -6964 9868 -6276 10292
rect -6212 9868 -6192 10292
rect -6964 9840 -6192 9868
rect -5952 10292 -5180 10320
rect -5952 9868 -5264 10292
rect -5200 9868 -5180 10292
rect -5952 9840 -5180 9868
rect -4940 10292 -4168 10320
rect -4940 9868 -4252 10292
rect -4188 9868 -4168 10292
rect -4940 9840 -4168 9868
rect -3928 10292 -3156 10320
rect -3928 9868 -3240 10292
rect -3176 9868 -3156 10292
rect -3928 9840 -3156 9868
rect -2916 10292 -2144 10320
rect -2916 9868 -2228 10292
rect -2164 9868 -2144 10292
rect -2916 9840 -2144 9868
rect -1904 10292 -1132 10320
rect -1904 9868 -1216 10292
rect -1152 9868 -1132 10292
rect -1904 9840 -1132 9868
rect -892 10292 -120 10320
rect -892 9868 -204 10292
rect -140 9868 -120 10292
rect -892 9840 -120 9868
rect 120 10292 892 10320
rect 120 9868 808 10292
rect 872 9868 892 10292
rect 120 9840 892 9868
rect 1132 10292 1904 10320
rect 1132 9868 1820 10292
rect 1884 9868 1904 10292
rect 1132 9840 1904 9868
rect 2144 10292 2916 10320
rect 2144 9868 2832 10292
rect 2896 9868 2916 10292
rect 2144 9840 2916 9868
rect 3156 10292 3928 10320
rect 3156 9868 3844 10292
rect 3908 9868 3928 10292
rect 3156 9840 3928 9868
rect 4168 10292 4940 10320
rect 4168 9868 4856 10292
rect 4920 9868 4940 10292
rect 4168 9840 4940 9868
rect 5180 10292 5952 10320
rect 5180 9868 5868 10292
rect 5932 9868 5952 10292
rect 5180 9840 5952 9868
rect 6192 10292 6964 10320
rect 6192 9868 6880 10292
rect 6944 9868 6964 10292
rect 6192 9840 6964 9868
rect 7204 10292 7976 10320
rect 7204 9868 7892 10292
rect 7956 9868 7976 10292
rect 7204 9840 7976 9868
rect 8216 10292 8988 10320
rect 8216 9868 8904 10292
rect 8968 9868 8988 10292
rect 8216 9840 8988 9868
rect 9228 10292 10000 10320
rect 9228 9868 9916 10292
rect 9980 9868 10000 10292
rect 9228 9840 10000 9868
rect 10240 10292 11012 10320
rect 10240 9868 10928 10292
rect 10992 9868 11012 10292
rect 10240 9840 11012 9868
rect 11252 10292 12024 10320
rect 11252 9868 11940 10292
rect 12004 9868 12024 10292
rect 11252 9840 12024 9868
rect 12264 10292 13036 10320
rect 12264 9868 12952 10292
rect 13016 9868 13036 10292
rect 12264 9840 13036 9868
rect 13276 10292 14048 10320
rect 13276 9868 13964 10292
rect 14028 9868 14048 10292
rect 13276 9840 14048 9868
rect 14288 10292 15060 10320
rect 14288 9868 14976 10292
rect 15040 9868 15060 10292
rect 14288 9840 15060 9868
rect 15300 10292 16072 10320
rect 15300 9868 15988 10292
rect 16052 9868 16072 10292
rect 15300 9840 16072 9868
rect 16312 10292 17084 10320
rect 16312 9868 17000 10292
rect 17064 9868 17084 10292
rect 16312 9840 17084 9868
rect -17084 9572 -16312 9600
rect -17084 9148 -16396 9572
rect -16332 9148 -16312 9572
rect -17084 9120 -16312 9148
rect -16072 9572 -15300 9600
rect -16072 9148 -15384 9572
rect -15320 9148 -15300 9572
rect -16072 9120 -15300 9148
rect -15060 9572 -14288 9600
rect -15060 9148 -14372 9572
rect -14308 9148 -14288 9572
rect -15060 9120 -14288 9148
rect -14048 9572 -13276 9600
rect -14048 9148 -13360 9572
rect -13296 9148 -13276 9572
rect -14048 9120 -13276 9148
rect -13036 9572 -12264 9600
rect -13036 9148 -12348 9572
rect -12284 9148 -12264 9572
rect -13036 9120 -12264 9148
rect -12024 9572 -11252 9600
rect -12024 9148 -11336 9572
rect -11272 9148 -11252 9572
rect -12024 9120 -11252 9148
rect -11012 9572 -10240 9600
rect -11012 9148 -10324 9572
rect -10260 9148 -10240 9572
rect -11012 9120 -10240 9148
rect -10000 9572 -9228 9600
rect -10000 9148 -9312 9572
rect -9248 9148 -9228 9572
rect -10000 9120 -9228 9148
rect -8988 9572 -8216 9600
rect -8988 9148 -8300 9572
rect -8236 9148 -8216 9572
rect -8988 9120 -8216 9148
rect -7976 9572 -7204 9600
rect -7976 9148 -7288 9572
rect -7224 9148 -7204 9572
rect -7976 9120 -7204 9148
rect -6964 9572 -6192 9600
rect -6964 9148 -6276 9572
rect -6212 9148 -6192 9572
rect -6964 9120 -6192 9148
rect -5952 9572 -5180 9600
rect -5952 9148 -5264 9572
rect -5200 9148 -5180 9572
rect -5952 9120 -5180 9148
rect -4940 9572 -4168 9600
rect -4940 9148 -4252 9572
rect -4188 9148 -4168 9572
rect -4940 9120 -4168 9148
rect -3928 9572 -3156 9600
rect -3928 9148 -3240 9572
rect -3176 9148 -3156 9572
rect -3928 9120 -3156 9148
rect -2916 9572 -2144 9600
rect -2916 9148 -2228 9572
rect -2164 9148 -2144 9572
rect -2916 9120 -2144 9148
rect -1904 9572 -1132 9600
rect -1904 9148 -1216 9572
rect -1152 9148 -1132 9572
rect -1904 9120 -1132 9148
rect -892 9572 -120 9600
rect -892 9148 -204 9572
rect -140 9148 -120 9572
rect -892 9120 -120 9148
rect 120 9572 892 9600
rect 120 9148 808 9572
rect 872 9148 892 9572
rect 120 9120 892 9148
rect 1132 9572 1904 9600
rect 1132 9148 1820 9572
rect 1884 9148 1904 9572
rect 1132 9120 1904 9148
rect 2144 9572 2916 9600
rect 2144 9148 2832 9572
rect 2896 9148 2916 9572
rect 2144 9120 2916 9148
rect 3156 9572 3928 9600
rect 3156 9148 3844 9572
rect 3908 9148 3928 9572
rect 3156 9120 3928 9148
rect 4168 9572 4940 9600
rect 4168 9148 4856 9572
rect 4920 9148 4940 9572
rect 4168 9120 4940 9148
rect 5180 9572 5952 9600
rect 5180 9148 5868 9572
rect 5932 9148 5952 9572
rect 5180 9120 5952 9148
rect 6192 9572 6964 9600
rect 6192 9148 6880 9572
rect 6944 9148 6964 9572
rect 6192 9120 6964 9148
rect 7204 9572 7976 9600
rect 7204 9148 7892 9572
rect 7956 9148 7976 9572
rect 7204 9120 7976 9148
rect 8216 9572 8988 9600
rect 8216 9148 8904 9572
rect 8968 9148 8988 9572
rect 8216 9120 8988 9148
rect 9228 9572 10000 9600
rect 9228 9148 9916 9572
rect 9980 9148 10000 9572
rect 9228 9120 10000 9148
rect 10240 9572 11012 9600
rect 10240 9148 10928 9572
rect 10992 9148 11012 9572
rect 10240 9120 11012 9148
rect 11252 9572 12024 9600
rect 11252 9148 11940 9572
rect 12004 9148 12024 9572
rect 11252 9120 12024 9148
rect 12264 9572 13036 9600
rect 12264 9148 12952 9572
rect 13016 9148 13036 9572
rect 12264 9120 13036 9148
rect 13276 9572 14048 9600
rect 13276 9148 13964 9572
rect 14028 9148 14048 9572
rect 13276 9120 14048 9148
rect 14288 9572 15060 9600
rect 14288 9148 14976 9572
rect 15040 9148 15060 9572
rect 14288 9120 15060 9148
rect 15300 9572 16072 9600
rect 15300 9148 15988 9572
rect 16052 9148 16072 9572
rect 15300 9120 16072 9148
rect 16312 9572 17084 9600
rect 16312 9148 17000 9572
rect 17064 9148 17084 9572
rect 16312 9120 17084 9148
rect -17084 8852 -16312 8880
rect -17084 8428 -16396 8852
rect -16332 8428 -16312 8852
rect -17084 8400 -16312 8428
rect -16072 8852 -15300 8880
rect -16072 8428 -15384 8852
rect -15320 8428 -15300 8852
rect -16072 8400 -15300 8428
rect -15060 8852 -14288 8880
rect -15060 8428 -14372 8852
rect -14308 8428 -14288 8852
rect -15060 8400 -14288 8428
rect -14048 8852 -13276 8880
rect -14048 8428 -13360 8852
rect -13296 8428 -13276 8852
rect -14048 8400 -13276 8428
rect -13036 8852 -12264 8880
rect -13036 8428 -12348 8852
rect -12284 8428 -12264 8852
rect -13036 8400 -12264 8428
rect -12024 8852 -11252 8880
rect -12024 8428 -11336 8852
rect -11272 8428 -11252 8852
rect -12024 8400 -11252 8428
rect -11012 8852 -10240 8880
rect -11012 8428 -10324 8852
rect -10260 8428 -10240 8852
rect -11012 8400 -10240 8428
rect -10000 8852 -9228 8880
rect -10000 8428 -9312 8852
rect -9248 8428 -9228 8852
rect -10000 8400 -9228 8428
rect -8988 8852 -8216 8880
rect -8988 8428 -8300 8852
rect -8236 8428 -8216 8852
rect -8988 8400 -8216 8428
rect -7976 8852 -7204 8880
rect -7976 8428 -7288 8852
rect -7224 8428 -7204 8852
rect -7976 8400 -7204 8428
rect -6964 8852 -6192 8880
rect -6964 8428 -6276 8852
rect -6212 8428 -6192 8852
rect -6964 8400 -6192 8428
rect -5952 8852 -5180 8880
rect -5952 8428 -5264 8852
rect -5200 8428 -5180 8852
rect -5952 8400 -5180 8428
rect -4940 8852 -4168 8880
rect -4940 8428 -4252 8852
rect -4188 8428 -4168 8852
rect -4940 8400 -4168 8428
rect -3928 8852 -3156 8880
rect -3928 8428 -3240 8852
rect -3176 8428 -3156 8852
rect -3928 8400 -3156 8428
rect -2916 8852 -2144 8880
rect -2916 8428 -2228 8852
rect -2164 8428 -2144 8852
rect -2916 8400 -2144 8428
rect -1904 8852 -1132 8880
rect -1904 8428 -1216 8852
rect -1152 8428 -1132 8852
rect -1904 8400 -1132 8428
rect -892 8852 -120 8880
rect -892 8428 -204 8852
rect -140 8428 -120 8852
rect -892 8400 -120 8428
rect 120 8852 892 8880
rect 120 8428 808 8852
rect 872 8428 892 8852
rect 120 8400 892 8428
rect 1132 8852 1904 8880
rect 1132 8428 1820 8852
rect 1884 8428 1904 8852
rect 1132 8400 1904 8428
rect 2144 8852 2916 8880
rect 2144 8428 2832 8852
rect 2896 8428 2916 8852
rect 2144 8400 2916 8428
rect 3156 8852 3928 8880
rect 3156 8428 3844 8852
rect 3908 8428 3928 8852
rect 3156 8400 3928 8428
rect 4168 8852 4940 8880
rect 4168 8428 4856 8852
rect 4920 8428 4940 8852
rect 4168 8400 4940 8428
rect 5180 8852 5952 8880
rect 5180 8428 5868 8852
rect 5932 8428 5952 8852
rect 5180 8400 5952 8428
rect 6192 8852 6964 8880
rect 6192 8428 6880 8852
rect 6944 8428 6964 8852
rect 6192 8400 6964 8428
rect 7204 8852 7976 8880
rect 7204 8428 7892 8852
rect 7956 8428 7976 8852
rect 7204 8400 7976 8428
rect 8216 8852 8988 8880
rect 8216 8428 8904 8852
rect 8968 8428 8988 8852
rect 8216 8400 8988 8428
rect 9228 8852 10000 8880
rect 9228 8428 9916 8852
rect 9980 8428 10000 8852
rect 9228 8400 10000 8428
rect 10240 8852 11012 8880
rect 10240 8428 10928 8852
rect 10992 8428 11012 8852
rect 10240 8400 11012 8428
rect 11252 8852 12024 8880
rect 11252 8428 11940 8852
rect 12004 8428 12024 8852
rect 11252 8400 12024 8428
rect 12264 8852 13036 8880
rect 12264 8428 12952 8852
rect 13016 8428 13036 8852
rect 12264 8400 13036 8428
rect 13276 8852 14048 8880
rect 13276 8428 13964 8852
rect 14028 8428 14048 8852
rect 13276 8400 14048 8428
rect 14288 8852 15060 8880
rect 14288 8428 14976 8852
rect 15040 8428 15060 8852
rect 14288 8400 15060 8428
rect 15300 8852 16072 8880
rect 15300 8428 15988 8852
rect 16052 8428 16072 8852
rect 15300 8400 16072 8428
rect 16312 8852 17084 8880
rect 16312 8428 17000 8852
rect 17064 8428 17084 8852
rect 16312 8400 17084 8428
rect -17084 8132 -16312 8160
rect -17084 7708 -16396 8132
rect -16332 7708 -16312 8132
rect -17084 7680 -16312 7708
rect -16072 8132 -15300 8160
rect -16072 7708 -15384 8132
rect -15320 7708 -15300 8132
rect -16072 7680 -15300 7708
rect -15060 8132 -14288 8160
rect -15060 7708 -14372 8132
rect -14308 7708 -14288 8132
rect -15060 7680 -14288 7708
rect -14048 8132 -13276 8160
rect -14048 7708 -13360 8132
rect -13296 7708 -13276 8132
rect -14048 7680 -13276 7708
rect -13036 8132 -12264 8160
rect -13036 7708 -12348 8132
rect -12284 7708 -12264 8132
rect -13036 7680 -12264 7708
rect -12024 8132 -11252 8160
rect -12024 7708 -11336 8132
rect -11272 7708 -11252 8132
rect -12024 7680 -11252 7708
rect -11012 8132 -10240 8160
rect -11012 7708 -10324 8132
rect -10260 7708 -10240 8132
rect -11012 7680 -10240 7708
rect -10000 8132 -9228 8160
rect -10000 7708 -9312 8132
rect -9248 7708 -9228 8132
rect -10000 7680 -9228 7708
rect -8988 8132 -8216 8160
rect -8988 7708 -8300 8132
rect -8236 7708 -8216 8132
rect -8988 7680 -8216 7708
rect -7976 8132 -7204 8160
rect -7976 7708 -7288 8132
rect -7224 7708 -7204 8132
rect -7976 7680 -7204 7708
rect -6964 8132 -6192 8160
rect -6964 7708 -6276 8132
rect -6212 7708 -6192 8132
rect -6964 7680 -6192 7708
rect -5952 8132 -5180 8160
rect -5952 7708 -5264 8132
rect -5200 7708 -5180 8132
rect -5952 7680 -5180 7708
rect -4940 8132 -4168 8160
rect -4940 7708 -4252 8132
rect -4188 7708 -4168 8132
rect -4940 7680 -4168 7708
rect -3928 8132 -3156 8160
rect -3928 7708 -3240 8132
rect -3176 7708 -3156 8132
rect -3928 7680 -3156 7708
rect -2916 8132 -2144 8160
rect -2916 7708 -2228 8132
rect -2164 7708 -2144 8132
rect -2916 7680 -2144 7708
rect -1904 8132 -1132 8160
rect -1904 7708 -1216 8132
rect -1152 7708 -1132 8132
rect -1904 7680 -1132 7708
rect -892 8132 -120 8160
rect -892 7708 -204 8132
rect -140 7708 -120 8132
rect -892 7680 -120 7708
rect 120 8132 892 8160
rect 120 7708 808 8132
rect 872 7708 892 8132
rect 120 7680 892 7708
rect 1132 8132 1904 8160
rect 1132 7708 1820 8132
rect 1884 7708 1904 8132
rect 1132 7680 1904 7708
rect 2144 8132 2916 8160
rect 2144 7708 2832 8132
rect 2896 7708 2916 8132
rect 2144 7680 2916 7708
rect 3156 8132 3928 8160
rect 3156 7708 3844 8132
rect 3908 7708 3928 8132
rect 3156 7680 3928 7708
rect 4168 8132 4940 8160
rect 4168 7708 4856 8132
rect 4920 7708 4940 8132
rect 4168 7680 4940 7708
rect 5180 8132 5952 8160
rect 5180 7708 5868 8132
rect 5932 7708 5952 8132
rect 5180 7680 5952 7708
rect 6192 8132 6964 8160
rect 6192 7708 6880 8132
rect 6944 7708 6964 8132
rect 6192 7680 6964 7708
rect 7204 8132 7976 8160
rect 7204 7708 7892 8132
rect 7956 7708 7976 8132
rect 7204 7680 7976 7708
rect 8216 8132 8988 8160
rect 8216 7708 8904 8132
rect 8968 7708 8988 8132
rect 8216 7680 8988 7708
rect 9228 8132 10000 8160
rect 9228 7708 9916 8132
rect 9980 7708 10000 8132
rect 9228 7680 10000 7708
rect 10240 8132 11012 8160
rect 10240 7708 10928 8132
rect 10992 7708 11012 8132
rect 10240 7680 11012 7708
rect 11252 8132 12024 8160
rect 11252 7708 11940 8132
rect 12004 7708 12024 8132
rect 11252 7680 12024 7708
rect 12264 8132 13036 8160
rect 12264 7708 12952 8132
rect 13016 7708 13036 8132
rect 12264 7680 13036 7708
rect 13276 8132 14048 8160
rect 13276 7708 13964 8132
rect 14028 7708 14048 8132
rect 13276 7680 14048 7708
rect 14288 8132 15060 8160
rect 14288 7708 14976 8132
rect 15040 7708 15060 8132
rect 14288 7680 15060 7708
rect 15300 8132 16072 8160
rect 15300 7708 15988 8132
rect 16052 7708 16072 8132
rect 15300 7680 16072 7708
rect 16312 8132 17084 8160
rect 16312 7708 17000 8132
rect 17064 7708 17084 8132
rect 16312 7680 17084 7708
rect -17084 7412 -16312 7440
rect -17084 6988 -16396 7412
rect -16332 6988 -16312 7412
rect -17084 6960 -16312 6988
rect -16072 7412 -15300 7440
rect -16072 6988 -15384 7412
rect -15320 6988 -15300 7412
rect -16072 6960 -15300 6988
rect -15060 7412 -14288 7440
rect -15060 6988 -14372 7412
rect -14308 6988 -14288 7412
rect -15060 6960 -14288 6988
rect -14048 7412 -13276 7440
rect -14048 6988 -13360 7412
rect -13296 6988 -13276 7412
rect -14048 6960 -13276 6988
rect -13036 7412 -12264 7440
rect -13036 6988 -12348 7412
rect -12284 6988 -12264 7412
rect -13036 6960 -12264 6988
rect -12024 7412 -11252 7440
rect -12024 6988 -11336 7412
rect -11272 6988 -11252 7412
rect -12024 6960 -11252 6988
rect -11012 7412 -10240 7440
rect -11012 6988 -10324 7412
rect -10260 6988 -10240 7412
rect -11012 6960 -10240 6988
rect -10000 7412 -9228 7440
rect -10000 6988 -9312 7412
rect -9248 6988 -9228 7412
rect -10000 6960 -9228 6988
rect -8988 7412 -8216 7440
rect -8988 6988 -8300 7412
rect -8236 6988 -8216 7412
rect -8988 6960 -8216 6988
rect -7976 7412 -7204 7440
rect -7976 6988 -7288 7412
rect -7224 6988 -7204 7412
rect -7976 6960 -7204 6988
rect -6964 7412 -6192 7440
rect -6964 6988 -6276 7412
rect -6212 6988 -6192 7412
rect -6964 6960 -6192 6988
rect -5952 7412 -5180 7440
rect -5952 6988 -5264 7412
rect -5200 6988 -5180 7412
rect -5952 6960 -5180 6988
rect -4940 7412 -4168 7440
rect -4940 6988 -4252 7412
rect -4188 6988 -4168 7412
rect -4940 6960 -4168 6988
rect -3928 7412 -3156 7440
rect -3928 6988 -3240 7412
rect -3176 6988 -3156 7412
rect -3928 6960 -3156 6988
rect -2916 7412 -2144 7440
rect -2916 6988 -2228 7412
rect -2164 6988 -2144 7412
rect -2916 6960 -2144 6988
rect -1904 7412 -1132 7440
rect -1904 6988 -1216 7412
rect -1152 6988 -1132 7412
rect -1904 6960 -1132 6988
rect -892 7412 -120 7440
rect -892 6988 -204 7412
rect -140 6988 -120 7412
rect -892 6960 -120 6988
rect 120 7412 892 7440
rect 120 6988 808 7412
rect 872 6988 892 7412
rect 120 6960 892 6988
rect 1132 7412 1904 7440
rect 1132 6988 1820 7412
rect 1884 6988 1904 7412
rect 1132 6960 1904 6988
rect 2144 7412 2916 7440
rect 2144 6988 2832 7412
rect 2896 6988 2916 7412
rect 2144 6960 2916 6988
rect 3156 7412 3928 7440
rect 3156 6988 3844 7412
rect 3908 6988 3928 7412
rect 3156 6960 3928 6988
rect 4168 7412 4940 7440
rect 4168 6988 4856 7412
rect 4920 6988 4940 7412
rect 4168 6960 4940 6988
rect 5180 7412 5952 7440
rect 5180 6988 5868 7412
rect 5932 6988 5952 7412
rect 5180 6960 5952 6988
rect 6192 7412 6964 7440
rect 6192 6988 6880 7412
rect 6944 6988 6964 7412
rect 6192 6960 6964 6988
rect 7204 7412 7976 7440
rect 7204 6988 7892 7412
rect 7956 6988 7976 7412
rect 7204 6960 7976 6988
rect 8216 7412 8988 7440
rect 8216 6988 8904 7412
rect 8968 6988 8988 7412
rect 8216 6960 8988 6988
rect 9228 7412 10000 7440
rect 9228 6988 9916 7412
rect 9980 6988 10000 7412
rect 9228 6960 10000 6988
rect 10240 7412 11012 7440
rect 10240 6988 10928 7412
rect 10992 6988 11012 7412
rect 10240 6960 11012 6988
rect 11252 7412 12024 7440
rect 11252 6988 11940 7412
rect 12004 6988 12024 7412
rect 11252 6960 12024 6988
rect 12264 7412 13036 7440
rect 12264 6988 12952 7412
rect 13016 6988 13036 7412
rect 12264 6960 13036 6988
rect 13276 7412 14048 7440
rect 13276 6988 13964 7412
rect 14028 6988 14048 7412
rect 13276 6960 14048 6988
rect 14288 7412 15060 7440
rect 14288 6988 14976 7412
rect 15040 6988 15060 7412
rect 14288 6960 15060 6988
rect 15300 7412 16072 7440
rect 15300 6988 15988 7412
rect 16052 6988 16072 7412
rect 15300 6960 16072 6988
rect 16312 7412 17084 7440
rect 16312 6988 17000 7412
rect 17064 6988 17084 7412
rect 16312 6960 17084 6988
rect -17084 6692 -16312 6720
rect -17084 6268 -16396 6692
rect -16332 6268 -16312 6692
rect -17084 6240 -16312 6268
rect -16072 6692 -15300 6720
rect -16072 6268 -15384 6692
rect -15320 6268 -15300 6692
rect -16072 6240 -15300 6268
rect -15060 6692 -14288 6720
rect -15060 6268 -14372 6692
rect -14308 6268 -14288 6692
rect -15060 6240 -14288 6268
rect -14048 6692 -13276 6720
rect -14048 6268 -13360 6692
rect -13296 6268 -13276 6692
rect -14048 6240 -13276 6268
rect -13036 6692 -12264 6720
rect -13036 6268 -12348 6692
rect -12284 6268 -12264 6692
rect -13036 6240 -12264 6268
rect -12024 6692 -11252 6720
rect -12024 6268 -11336 6692
rect -11272 6268 -11252 6692
rect -12024 6240 -11252 6268
rect -11012 6692 -10240 6720
rect -11012 6268 -10324 6692
rect -10260 6268 -10240 6692
rect -11012 6240 -10240 6268
rect -10000 6692 -9228 6720
rect -10000 6268 -9312 6692
rect -9248 6268 -9228 6692
rect -10000 6240 -9228 6268
rect -8988 6692 -8216 6720
rect -8988 6268 -8300 6692
rect -8236 6268 -8216 6692
rect -8988 6240 -8216 6268
rect -7976 6692 -7204 6720
rect -7976 6268 -7288 6692
rect -7224 6268 -7204 6692
rect -7976 6240 -7204 6268
rect -6964 6692 -6192 6720
rect -6964 6268 -6276 6692
rect -6212 6268 -6192 6692
rect -6964 6240 -6192 6268
rect -5952 6692 -5180 6720
rect -5952 6268 -5264 6692
rect -5200 6268 -5180 6692
rect -5952 6240 -5180 6268
rect -4940 6692 -4168 6720
rect -4940 6268 -4252 6692
rect -4188 6268 -4168 6692
rect -4940 6240 -4168 6268
rect -3928 6692 -3156 6720
rect -3928 6268 -3240 6692
rect -3176 6268 -3156 6692
rect -3928 6240 -3156 6268
rect -2916 6692 -2144 6720
rect -2916 6268 -2228 6692
rect -2164 6268 -2144 6692
rect -2916 6240 -2144 6268
rect -1904 6692 -1132 6720
rect -1904 6268 -1216 6692
rect -1152 6268 -1132 6692
rect -1904 6240 -1132 6268
rect -892 6692 -120 6720
rect -892 6268 -204 6692
rect -140 6268 -120 6692
rect -892 6240 -120 6268
rect 120 6692 892 6720
rect 120 6268 808 6692
rect 872 6268 892 6692
rect 120 6240 892 6268
rect 1132 6692 1904 6720
rect 1132 6268 1820 6692
rect 1884 6268 1904 6692
rect 1132 6240 1904 6268
rect 2144 6692 2916 6720
rect 2144 6268 2832 6692
rect 2896 6268 2916 6692
rect 2144 6240 2916 6268
rect 3156 6692 3928 6720
rect 3156 6268 3844 6692
rect 3908 6268 3928 6692
rect 3156 6240 3928 6268
rect 4168 6692 4940 6720
rect 4168 6268 4856 6692
rect 4920 6268 4940 6692
rect 4168 6240 4940 6268
rect 5180 6692 5952 6720
rect 5180 6268 5868 6692
rect 5932 6268 5952 6692
rect 5180 6240 5952 6268
rect 6192 6692 6964 6720
rect 6192 6268 6880 6692
rect 6944 6268 6964 6692
rect 6192 6240 6964 6268
rect 7204 6692 7976 6720
rect 7204 6268 7892 6692
rect 7956 6268 7976 6692
rect 7204 6240 7976 6268
rect 8216 6692 8988 6720
rect 8216 6268 8904 6692
rect 8968 6268 8988 6692
rect 8216 6240 8988 6268
rect 9228 6692 10000 6720
rect 9228 6268 9916 6692
rect 9980 6268 10000 6692
rect 9228 6240 10000 6268
rect 10240 6692 11012 6720
rect 10240 6268 10928 6692
rect 10992 6268 11012 6692
rect 10240 6240 11012 6268
rect 11252 6692 12024 6720
rect 11252 6268 11940 6692
rect 12004 6268 12024 6692
rect 11252 6240 12024 6268
rect 12264 6692 13036 6720
rect 12264 6268 12952 6692
rect 13016 6268 13036 6692
rect 12264 6240 13036 6268
rect 13276 6692 14048 6720
rect 13276 6268 13964 6692
rect 14028 6268 14048 6692
rect 13276 6240 14048 6268
rect 14288 6692 15060 6720
rect 14288 6268 14976 6692
rect 15040 6268 15060 6692
rect 14288 6240 15060 6268
rect 15300 6692 16072 6720
rect 15300 6268 15988 6692
rect 16052 6268 16072 6692
rect 15300 6240 16072 6268
rect 16312 6692 17084 6720
rect 16312 6268 17000 6692
rect 17064 6268 17084 6692
rect 16312 6240 17084 6268
rect -17084 5972 -16312 6000
rect -17084 5548 -16396 5972
rect -16332 5548 -16312 5972
rect -17084 5520 -16312 5548
rect -16072 5972 -15300 6000
rect -16072 5548 -15384 5972
rect -15320 5548 -15300 5972
rect -16072 5520 -15300 5548
rect -15060 5972 -14288 6000
rect -15060 5548 -14372 5972
rect -14308 5548 -14288 5972
rect -15060 5520 -14288 5548
rect -14048 5972 -13276 6000
rect -14048 5548 -13360 5972
rect -13296 5548 -13276 5972
rect -14048 5520 -13276 5548
rect -13036 5972 -12264 6000
rect -13036 5548 -12348 5972
rect -12284 5548 -12264 5972
rect -13036 5520 -12264 5548
rect -12024 5972 -11252 6000
rect -12024 5548 -11336 5972
rect -11272 5548 -11252 5972
rect -12024 5520 -11252 5548
rect -11012 5972 -10240 6000
rect -11012 5548 -10324 5972
rect -10260 5548 -10240 5972
rect -11012 5520 -10240 5548
rect -10000 5972 -9228 6000
rect -10000 5548 -9312 5972
rect -9248 5548 -9228 5972
rect -10000 5520 -9228 5548
rect -8988 5972 -8216 6000
rect -8988 5548 -8300 5972
rect -8236 5548 -8216 5972
rect -8988 5520 -8216 5548
rect -7976 5972 -7204 6000
rect -7976 5548 -7288 5972
rect -7224 5548 -7204 5972
rect -7976 5520 -7204 5548
rect -6964 5972 -6192 6000
rect -6964 5548 -6276 5972
rect -6212 5548 -6192 5972
rect -6964 5520 -6192 5548
rect -5952 5972 -5180 6000
rect -5952 5548 -5264 5972
rect -5200 5548 -5180 5972
rect -5952 5520 -5180 5548
rect -4940 5972 -4168 6000
rect -4940 5548 -4252 5972
rect -4188 5548 -4168 5972
rect -4940 5520 -4168 5548
rect -3928 5972 -3156 6000
rect -3928 5548 -3240 5972
rect -3176 5548 -3156 5972
rect -3928 5520 -3156 5548
rect -2916 5972 -2144 6000
rect -2916 5548 -2228 5972
rect -2164 5548 -2144 5972
rect -2916 5520 -2144 5548
rect -1904 5972 -1132 6000
rect -1904 5548 -1216 5972
rect -1152 5548 -1132 5972
rect -1904 5520 -1132 5548
rect -892 5972 -120 6000
rect -892 5548 -204 5972
rect -140 5548 -120 5972
rect -892 5520 -120 5548
rect 120 5972 892 6000
rect 120 5548 808 5972
rect 872 5548 892 5972
rect 120 5520 892 5548
rect 1132 5972 1904 6000
rect 1132 5548 1820 5972
rect 1884 5548 1904 5972
rect 1132 5520 1904 5548
rect 2144 5972 2916 6000
rect 2144 5548 2832 5972
rect 2896 5548 2916 5972
rect 2144 5520 2916 5548
rect 3156 5972 3928 6000
rect 3156 5548 3844 5972
rect 3908 5548 3928 5972
rect 3156 5520 3928 5548
rect 4168 5972 4940 6000
rect 4168 5548 4856 5972
rect 4920 5548 4940 5972
rect 4168 5520 4940 5548
rect 5180 5972 5952 6000
rect 5180 5548 5868 5972
rect 5932 5548 5952 5972
rect 5180 5520 5952 5548
rect 6192 5972 6964 6000
rect 6192 5548 6880 5972
rect 6944 5548 6964 5972
rect 6192 5520 6964 5548
rect 7204 5972 7976 6000
rect 7204 5548 7892 5972
rect 7956 5548 7976 5972
rect 7204 5520 7976 5548
rect 8216 5972 8988 6000
rect 8216 5548 8904 5972
rect 8968 5548 8988 5972
rect 8216 5520 8988 5548
rect 9228 5972 10000 6000
rect 9228 5548 9916 5972
rect 9980 5548 10000 5972
rect 9228 5520 10000 5548
rect 10240 5972 11012 6000
rect 10240 5548 10928 5972
rect 10992 5548 11012 5972
rect 10240 5520 11012 5548
rect 11252 5972 12024 6000
rect 11252 5548 11940 5972
rect 12004 5548 12024 5972
rect 11252 5520 12024 5548
rect 12264 5972 13036 6000
rect 12264 5548 12952 5972
rect 13016 5548 13036 5972
rect 12264 5520 13036 5548
rect 13276 5972 14048 6000
rect 13276 5548 13964 5972
rect 14028 5548 14048 5972
rect 13276 5520 14048 5548
rect 14288 5972 15060 6000
rect 14288 5548 14976 5972
rect 15040 5548 15060 5972
rect 14288 5520 15060 5548
rect 15300 5972 16072 6000
rect 15300 5548 15988 5972
rect 16052 5548 16072 5972
rect 15300 5520 16072 5548
rect 16312 5972 17084 6000
rect 16312 5548 17000 5972
rect 17064 5548 17084 5972
rect 16312 5520 17084 5548
rect -17084 5252 -16312 5280
rect -17084 4828 -16396 5252
rect -16332 4828 -16312 5252
rect -17084 4800 -16312 4828
rect -16072 5252 -15300 5280
rect -16072 4828 -15384 5252
rect -15320 4828 -15300 5252
rect -16072 4800 -15300 4828
rect -15060 5252 -14288 5280
rect -15060 4828 -14372 5252
rect -14308 4828 -14288 5252
rect -15060 4800 -14288 4828
rect -14048 5252 -13276 5280
rect -14048 4828 -13360 5252
rect -13296 4828 -13276 5252
rect -14048 4800 -13276 4828
rect -13036 5252 -12264 5280
rect -13036 4828 -12348 5252
rect -12284 4828 -12264 5252
rect -13036 4800 -12264 4828
rect -12024 5252 -11252 5280
rect -12024 4828 -11336 5252
rect -11272 4828 -11252 5252
rect -12024 4800 -11252 4828
rect -11012 5252 -10240 5280
rect -11012 4828 -10324 5252
rect -10260 4828 -10240 5252
rect -11012 4800 -10240 4828
rect -10000 5252 -9228 5280
rect -10000 4828 -9312 5252
rect -9248 4828 -9228 5252
rect -10000 4800 -9228 4828
rect -8988 5252 -8216 5280
rect -8988 4828 -8300 5252
rect -8236 4828 -8216 5252
rect -8988 4800 -8216 4828
rect -7976 5252 -7204 5280
rect -7976 4828 -7288 5252
rect -7224 4828 -7204 5252
rect -7976 4800 -7204 4828
rect -6964 5252 -6192 5280
rect -6964 4828 -6276 5252
rect -6212 4828 -6192 5252
rect -6964 4800 -6192 4828
rect -5952 5252 -5180 5280
rect -5952 4828 -5264 5252
rect -5200 4828 -5180 5252
rect -5952 4800 -5180 4828
rect -4940 5252 -4168 5280
rect -4940 4828 -4252 5252
rect -4188 4828 -4168 5252
rect -4940 4800 -4168 4828
rect -3928 5252 -3156 5280
rect -3928 4828 -3240 5252
rect -3176 4828 -3156 5252
rect -3928 4800 -3156 4828
rect -2916 5252 -2144 5280
rect -2916 4828 -2228 5252
rect -2164 4828 -2144 5252
rect -2916 4800 -2144 4828
rect -1904 5252 -1132 5280
rect -1904 4828 -1216 5252
rect -1152 4828 -1132 5252
rect -1904 4800 -1132 4828
rect -892 5252 -120 5280
rect -892 4828 -204 5252
rect -140 4828 -120 5252
rect -892 4800 -120 4828
rect 120 5252 892 5280
rect 120 4828 808 5252
rect 872 4828 892 5252
rect 120 4800 892 4828
rect 1132 5252 1904 5280
rect 1132 4828 1820 5252
rect 1884 4828 1904 5252
rect 1132 4800 1904 4828
rect 2144 5252 2916 5280
rect 2144 4828 2832 5252
rect 2896 4828 2916 5252
rect 2144 4800 2916 4828
rect 3156 5252 3928 5280
rect 3156 4828 3844 5252
rect 3908 4828 3928 5252
rect 3156 4800 3928 4828
rect 4168 5252 4940 5280
rect 4168 4828 4856 5252
rect 4920 4828 4940 5252
rect 4168 4800 4940 4828
rect 5180 5252 5952 5280
rect 5180 4828 5868 5252
rect 5932 4828 5952 5252
rect 5180 4800 5952 4828
rect 6192 5252 6964 5280
rect 6192 4828 6880 5252
rect 6944 4828 6964 5252
rect 6192 4800 6964 4828
rect 7204 5252 7976 5280
rect 7204 4828 7892 5252
rect 7956 4828 7976 5252
rect 7204 4800 7976 4828
rect 8216 5252 8988 5280
rect 8216 4828 8904 5252
rect 8968 4828 8988 5252
rect 8216 4800 8988 4828
rect 9228 5252 10000 5280
rect 9228 4828 9916 5252
rect 9980 4828 10000 5252
rect 9228 4800 10000 4828
rect 10240 5252 11012 5280
rect 10240 4828 10928 5252
rect 10992 4828 11012 5252
rect 10240 4800 11012 4828
rect 11252 5252 12024 5280
rect 11252 4828 11940 5252
rect 12004 4828 12024 5252
rect 11252 4800 12024 4828
rect 12264 5252 13036 5280
rect 12264 4828 12952 5252
rect 13016 4828 13036 5252
rect 12264 4800 13036 4828
rect 13276 5252 14048 5280
rect 13276 4828 13964 5252
rect 14028 4828 14048 5252
rect 13276 4800 14048 4828
rect 14288 5252 15060 5280
rect 14288 4828 14976 5252
rect 15040 4828 15060 5252
rect 14288 4800 15060 4828
rect 15300 5252 16072 5280
rect 15300 4828 15988 5252
rect 16052 4828 16072 5252
rect 15300 4800 16072 4828
rect 16312 5252 17084 5280
rect 16312 4828 17000 5252
rect 17064 4828 17084 5252
rect 16312 4800 17084 4828
rect -17084 4532 -16312 4560
rect -17084 4108 -16396 4532
rect -16332 4108 -16312 4532
rect -17084 4080 -16312 4108
rect -16072 4532 -15300 4560
rect -16072 4108 -15384 4532
rect -15320 4108 -15300 4532
rect -16072 4080 -15300 4108
rect -15060 4532 -14288 4560
rect -15060 4108 -14372 4532
rect -14308 4108 -14288 4532
rect -15060 4080 -14288 4108
rect -14048 4532 -13276 4560
rect -14048 4108 -13360 4532
rect -13296 4108 -13276 4532
rect -14048 4080 -13276 4108
rect -13036 4532 -12264 4560
rect -13036 4108 -12348 4532
rect -12284 4108 -12264 4532
rect -13036 4080 -12264 4108
rect -12024 4532 -11252 4560
rect -12024 4108 -11336 4532
rect -11272 4108 -11252 4532
rect -12024 4080 -11252 4108
rect -11012 4532 -10240 4560
rect -11012 4108 -10324 4532
rect -10260 4108 -10240 4532
rect -11012 4080 -10240 4108
rect -10000 4532 -9228 4560
rect -10000 4108 -9312 4532
rect -9248 4108 -9228 4532
rect -10000 4080 -9228 4108
rect -8988 4532 -8216 4560
rect -8988 4108 -8300 4532
rect -8236 4108 -8216 4532
rect -8988 4080 -8216 4108
rect -7976 4532 -7204 4560
rect -7976 4108 -7288 4532
rect -7224 4108 -7204 4532
rect -7976 4080 -7204 4108
rect -6964 4532 -6192 4560
rect -6964 4108 -6276 4532
rect -6212 4108 -6192 4532
rect -6964 4080 -6192 4108
rect -5952 4532 -5180 4560
rect -5952 4108 -5264 4532
rect -5200 4108 -5180 4532
rect -5952 4080 -5180 4108
rect -4940 4532 -4168 4560
rect -4940 4108 -4252 4532
rect -4188 4108 -4168 4532
rect -4940 4080 -4168 4108
rect -3928 4532 -3156 4560
rect -3928 4108 -3240 4532
rect -3176 4108 -3156 4532
rect -3928 4080 -3156 4108
rect -2916 4532 -2144 4560
rect -2916 4108 -2228 4532
rect -2164 4108 -2144 4532
rect -2916 4080 -2144 4108
rect -1904 4532 -1132 4560
rect -1904 4108 -1216 4532
rect -1152 4108 -1132 4532
rect -1904 4080 -1132 4108
rect -892 4532 -120 4560
rect -892 4108 -204 4532
rect -140 4108 -120 4532
rect -892 4080 -120 4108
rect 120 4532 892 4560
rect 120 4108 808 4532
rect 872 4108 892 4532
rect 120 4080 892 4108
rect 1132 4532 1904 4560
rect 1132 4108 1820 4532
rect 1884 4108 1904 4532
rect 1132 4080 1904 4108
rect 2144 4532 2916 4560
rect 2144 4108 2832 4532
rect 2896 4108 2916 4532
rect 2144 4080 2916 4108
rect 3156 4532 3928 4560
rect 3156 4108 3844 4532
rect 3908 4108 3928 4532
rect 3156 4080 3928 4108
rect 4168 4532 4940 4560
rect 4168 4108 4856 4532
rect 4920 4108 4940 4532
rect 4168 4080 4940 4108
rect 5180 4532 5952 4560
rect 5180 4108 5868 4532
rect 5932 4108 5952 4532
rect 5180 4080 5952 4108
rect 6192 4532 6964 4560
rect 6192 4108 6880 4532
rect 6944 4108 6964 4532
rect 6192 4080 6964 4108
rect 7204 4532 7976 4560
rect 7204 4108 7892 4532
rect 7956 4108 7976 4532
rect 7204 4080 7976 4108
rect 8216 4532 8988 4560
rect 8216 4108 8904 4532
rect 8968 4108 8988 4532
rect 8216 4080 8988 4108
rect 9228 4532 10000 4560
rect 9228 4108 9916 4532
rect 9980 4108 10000 4532
rect 9228 4080 10000 4108
rect 10240 4532 11012 4560
rect 10240 4108 10928 4532
rect 10992 4108 11012 4532
rect 10240 4080 11012 4108
rect 11252 4532 12024 4560
rect 11252 4108 11940 4532
rect 12004 4108 12024 4532
rect 11252 4080 12024 4108
rect 12264 4532 13036 4560
rect 12264 4108 12952 4532
rect 13016 4108 13036 4532
rect 12264 4080 13036 4108
rect 13276 4532 14048 4560
rect 13276 4108 13964 4532
rect 14028 4108 14048 4532
rect 13276 4080 14048 4108
rect 14288 4532 15060 4560
rect 14288 4108 14976 4532
rect 15040 4108 15060 4532
rect 14288 4080 15060 4108
rect 15300 4532 16072 4560
rect 15300 4108 15988 4532
rect 16052 4108 16072 4532
rect 15300 4080 16072 4108
rect 16312 4532 17084 4560
rect 16312 4108 17000 4532
rect 17064 4108 17084 4532
rect 16312 4080 17084 4108
rect -17084 3812 -16312 3840
rect -17084 3388 -16396 3812
rect -16332 3388 -16312 3812
rect -17084 3360 -16312 3388
rect -16072 3812 -15300 3840
rect -16072 3388 -15384 3812
rect -15320 3388 -15300 3812
rect -16072 3360 -15300 3388
rect -15060 3812 -14288 3840
rect -15060 3388 -14372 3812
rect -14308 3388 -14288 3812
rect -15060 3360 -14288 3388
rect -14048 3812 -13276 3840
rect -14048 3388 -13360 3812
rect -13296 3388 -13276 3812
rect -14048 3360 -13276 3388
rect -13036 3812 -12264 3840
rect -13036 3388 -12348 3812
rect -12284 3388 -12264 3812
rect -13036 3360 -12264 3388
rect -12024 3812 -11252 3840
rect -12024 3388 -11336 3812
rect -11272 3388 -11252 3812
rect -12024 3360 -11252 3388
rect -11012 3812 -10240 3840
rect -11012 3388 -10324 3812
rect -10260 3388 -10240 3812
rect -11012 3360 -10240 3388
rect -10000 3812 -9228 3840
rect -10000 3388 -9312 3812
rect -9248 3388 -9228 3812
rect -10000 3360 -9228 3388
rect -8988 3812 -8216 3840
rect -8988 3388 -8300 3812
rect -8236 3388 -8216 3812
rect -8988 3360 -8216 3388
rect -7976 3812 -7204 3840
rect -7976 3388 -7288 3812
rect -7224 3388 -7204 3812
rect -7976 3360 -7204 3388
rect -6964 3812 -6192 3840
rect -6964 3388 -6276 3812
rect -6212 3388 -6192 3812
rect -6964 3360 -6192 3388
rect -5952 3812 -5180 3840
rect -5952 3388 -5264 3812
rect -5200 3388 -5180 3812
rect -5952 3360 -5180 3388
rect -4940 3812 -4168 3840
rect -4940 3388 -4252 3812
rect -4188 3388 -4168 3812
rect -4940 3360 -4168 3388
rect -3928 3812 -3156 3840
rect -3928 3388 -3240 3812
rect -3176 3388 -3156 3812
rect -3928 3360 -3156 3388
rect -2916 3812 -2144 3840
rect -2916 3388 -2228 3812
rect -2164 3388 -2144 3812
rect -2916 3360 -2144 3388
rect -1904 3812 -1132 3840
rect -1904 3388 -1216 3812
rect -1152 3388 -1132 3812
rect -1904 3360 -1132 3388
rect -892 3812 -120 3840
rect -892 3388 -204 3812
rect -140 3388 -120 3812
rect -892 3360 -120 3388
rect 120 3812 892 3840
rect 120 3388 808 3812
rect 872 3388 892 3812
rect 120 3360 892 3388
rect 1132 3812 1904 3840
rect 1132 3388 1820 3812
rect 1884 3388 1904 3812
rect 1132 3360 1904 3388
rect 2144 3812 2916 3840
rect 2144 3388 2832 3812
rect 2896 3388 2916 3812
rect 2144 3360 2916 3388
rect 3156 3812 3928 3840
rect 3156 3388 3844 3812
rect 3908 3388 3928 3812
rect 3156 3360 3928 3388
rect 4168 3812 4940 3840
rect 4168 3388 4856 3812
rect 4920 3388 4940 3812
rect 4168 3360 4940 3388
rect 5180 3812 5952 3840
rect 5180 3388 5868 3812
rect 5932 3388 5952 3812
rect 5180 3360 5952 3388
rect 6192 3812 6964 3840
rect 6192 3388 6880 3812
rect 6944 3388 6964 3812
rect 6192 3360 6964 3388
rect 7204 3812 7976 3840
rect 7204 3388 7892 3812
rect 7956 3388 7976 3812
rect 7204 3360 7976 3388
rect 8216 3812 8988 3840
rect 8216 3388 8904 3812
rect 8968 3388 8988 3812
rect 8216 3360 8988 3388
rect 9228 3812 10000 3840
rect 9228 3388 9916 3812
rect 9980 3388 10000 3812
rect 9228 3360 10000 3388
rect 10240 3812 11012 3840
rect 10240 3388 10928 3812
rect 10992 3388 11012 3812
rect 10240 3360 11012 3388
rect 11252 3812 12024 3840
rect 11252 3388 11940 3812
rect 12004 3388 12024 3812
rect 11252 3360 12024 3388
rect 12264 3812 13036 3840
rect 12264 3388 12952 3812
rect 13016 3388 13036 3812
rect 12264 3360 13036 3388
rect 13276 3812 14048 3840
rect 13276 3388 13964 3812
rect 14028 3388 14048 3812
rect 13276 3360 14048 3388
rect 14288 3812 15060 3840
rect 14288 3388 14976 3812
rect 15040 3388 15060 3812
rect 14288 3360 15060 3388
rect 15300 3812 16072 3840
rect 15300 3388 15988 3812
rect 16052 3388 16072 3812
rect 15300 3360 16072 3388
rect 16312 3812 17084 3840
rect 16312 3388 17000 3812
rect 17064 3388 17084 3812
rect 16312 3360 17084 3388
rect -17084 3092 -16312 3120
rect -17084 2668 -16396 3092
rect -16332 2668 -16312 3092
rect -17084 2640 -16312 2668
rect -16072 3092 -15300 3120
rect -16072 2668 -15384 3092
rect -15320 2668 -15300 3092
rect -16072 2640 -15300 2668
rect -15060 3092 -14288 3120
rect -15060 2668 -14372 3092
rect -14308 2668 -14288 3092
rect -15060 2640 -14288 2668
rect -14048 3092 -13276 3120
rect -14048 2668 -13360 3092
rect -13296 2668 -13276 3092
rect -14048 2640 -13276 2668
rect -13036 3092 -12264 3120
rect -13036 2668 -12348 3092
rect -12284 2668 -12264 3092
rect -13036 2640 -12264 2668
rect -12024 3092 -11252 3120
rect -12024 2668 -11336 3092
rect -11272 2668 -11252 3092
rect -12024 2640 -11252 2668
rect -11012 3092 -10240 3120
rect -11012 2668 -10324 3092
rect -10260 2668 -10240 3092
rect -11012 2640 -10240 2668
rect -10000 3092 -9228 3120
rect -10000 2668 -9312 3092
rect -9248 2668 -9228 3092
rect -10000 2640 -9228 2668
rect -8988 3092 -8216 3120
rect -8988 2668 -8300 3092
rect -8236 2668 -8216 3092
rect -8988 2640 -8216 2668
rect -7976 3092 -7204 3120
rect -7976 2668 -7288 3092
rect -7224 2668 -7204 3092
rect -7976 2640 -7204 2668
rect -6964 3092 -6192 3120
rect -6964 2668 -6276 3092
rect -6212 2668 -6192 3092
rect -6964 2640 -6192 2668
rect -5952 3092 -5180 3120
rect -5952 2668 -5264 3092
rect -5200 2668 -5180 3092
rect -5952 2640 -5180 2668
rect -4940 3092 -4168 3120
rect -4940 2668 -4252 3092
rect -4188 2668 -4168 3092
rect -4940 2640 -4168 2668
rect -3928 3092 -3156 3120
rect -3928 2668 -3240 3092
rect -3176 2668 -3156 3092
rect -3928 2640 -3156 2668
rect -2916 3092 -2144 3120
rect -2916 2668 -2228 3092
rect -2164 2668 -2144 3092
rect -2916 2640 -2144 2668
rect -1904 3092 -1132 3120
rect -1904 2668 -1216 3092
rect -1152 2668 -1132 3092
rect -1904 2640 -1132 2668
rect -892 3092 -120 3120
rect -892 2668 -204 3092
rect -140 2668 -120 3092
rect -892 2640 -120 2668
rect 120 3092 892 3120
rect 120 2668 808 3092
rect 872 2668 892 3092
rect 120 2640 892 2668
rect 1132 3092 1904 3120
rect 1132 2668 1820 3092
rect 1884 2668 1904 3092
rect 1132 2640 1904 2668
rect 2144 3092 2916 3120
rect 2144 2668 2832 3092
rect 2896 2668 2916 3092
rect 2144 2640 2916 2668
rect 3156 3092 3928 3120
rect 3156 2668 3844 3092
rect 3908 2668 3928 3092
rect 3156 2640 3928 2668
rect 4168 3092 4940 3120
rect 4168 2668 4856 3092
rect 4920 2668 4940 3092
rect 4168 2640 4940 2668
rect 5180 3092 5952 3120
rect 5180 2668 5868 3092
rect 5932 2668 5952 3092
rect 5180 2640 5952 2668
rect 6192 3092 6964 3120
rect 6192 2668 6880 3092
rect 6944 2668 6964 3092
rect 6192 2640 6964 2668
rect 7204 3092 7976 3120
rect 7204 2668 7892 3092
rect 7956 2668 7976 3092
rect 7204 2640 7976 2668
rect 8216 3092 8988 3120
rect 8216 2668 8904 3092
rect 8968 2668 8988 3092
rect 8216 2640 8988 2668
rect 9228 3092 10000 3120
rect 9228 2668 9916 3092
rect 9980 2668 10000 3092
rect 9228 2640 10000 2668
rect 10240 3092 11012 3120
rect 10240 2668 10928 3092
rect 10992 2668 11012 3092
rect 10240 2640 11012 2668
rect 11252 3092 12024 3120
rect 11252 2668 11940 3092
rect 12004 2668 12024 3092
rect 11252 2640 12024 2668
rect 12264 3092 13036 3120
rect 12264 2668 12952 3092
rect 13016 2668 13036 3092
rect 12264 2640 13036 2668
rect 13276 3092 14048 3120
rect 13276 2668 13964 3092
rect 14028 2668 14048 3092
rect 13276 2640 14048 2668
rect 14288 3092 15060 3120
rect 14288 2668 14976 3092
rect 15040 2668 15060 3092
rect 14288 2640 15060 2668
rect 15300 3092 16072 3120
rect 15300 2668 15988 3092
rect 16052 2668 16072 3092
rect 15300 2640 16072 2668
rect 16312 3092 17084 3120
rect 16312 2668 17000 3092
rect 17064 2668 17084 3092
rect 16312 2640 17084 2668
rect -17084 2372 -16312 2400
rect -17084 1948 -16396 2372
rect -16332 1948 -16312 2372
rect -17084 1920 -16312 1948
rect -16072 2372 -15300 2400
rect -16072 1948 -15384 2372
rect -15320 1948 -15300 2372
rect -16072 1920 -15300 1948
rect -15060 2372 -14288 2400
rect -15060 1948 -14372 2372
rect -14308 1948 -14288 2372
rect -15060 1920 -14288 1948
rect -14048 2372 -13276 2400
rect -14048 1948 -13360 2372
rect -13296 1948 -13276 2372
rect -14048 1920 -13276 1948
rect -13036 2372 -12264 2400
rect -13036 1948 -12348 2372
rect -12284 1948 -12264 2372
rect -13036 1920 -12264 1948
rect -12024 2372 -11252 2400
rect -12024 1948 -11336 2372
rect -11272 1948 -11252 2372
rect -12024 1920 -11252 1948
rect -11012 2372 -10240 2400
rect -11012 1948 -10324 2372
rect -10260 1948 -10240 2372
rect -11012 1920 -10240 1948
rect -10000 2372 -9228 2400
rect -10000 1948 -9312 2372
rect -9248 1948 -9228 2372
rect -10000 1920 -9228 1948
rect -8988 2372 -8216 2400
rect -8988 1948 -8300 2372
rect -8236 1948 -8216 2372
rect -8988 1920 -8216 1948
rect -7976 2372 -7204 2400
rect -7976 1948 -7288 2372
rect -7224 1948 -7204 2372
rect -7976 1920 -7204 1948
rect -6964 2372 -6192 2400
rect -6964 1948 -6276 2372
rect -6212 1948 -6192 2372
rect -6964 1920 -6192 1948
rect -5952 2372 -5180 2400
rect -5952 1948 -5264 2372
rect -5200 1948 -5180 2372
rect -5952 1920 -5180 1948
rect -4940 2372 -4168 2400
rect -4940 1948 -4252 2372
rect -4188 1948 -4168 2372
rect -4940 1920 -4168 1948
rect -3928 2372 -3156 2400
rect -3928 1948 -3240 2372
rect -3176 1948 -3156 2372
rect -3928 1920 -3156 1948
rect -2916 2372 -2144 2400
rect -2916 1948 -2228 2372
rect -2164 1948 -2144 2372
rect -2916 1920 -2144 1948
rect -1904 2372 -1132 2400
rect -1904 1948 -1216 2372
rect -1152 1948 -1132 2372
rect -1904 1920 -1132 1948
rect -892 2372 -120 2400
rect -892 1948 -204 2372
rect -140 1948 -120 2372
rect -892 1920 -120 1948
rect 120 2372 892 2400
rect 120 1948 808 2372
rect 872 1948 892 2372
rect 120 1920 892 1948
rect 1132 2372 1904 2400
rect 1132 1948 1820 2372
rect 1884 1948 1904 2372
rect 1132 1920 1904 1948
rect 2144 2372 2916 2400
rect 2144 1948 2832 2372
rect 2896 1948 2916 2372
rect 2144 1920 2916 1948
rect 3156 2372 3928 2400
rect 3156 1948 3844 2372
rect 3908 1948 3928 2372
rect 3156 1920 3928 1948
rect 4168 2372 4940 2400
rect 4168 1948 4856 2372
rect 4920 1948 4940 2372
rect 4168 1920 4940 1948
rect 5180 2372 5952 2400
rect 5180 1948 5868 2372
rect 5932 1948 5952 2372
rect 5180 1920 5952 1948
rect 6192 2372 6964 2400
rect 6192 1948 6880 2372
rect 6944 1948 6964 2372
rect 6192 1920 6964 1948
rect 7204 2372 7976 2400
rect 7204 1948 7892 2372
rect 7956 1948 7976 2372
rect 7204 1920 7976 1948
rect 8216 2372 8988 2400
rect 8216 1948 8904 2372
rect 8968 1948 8988 2372
rect 8216 1920 8988 1948
rect 9228 2372 10000 2400
rect 9228 1948 9916 2372
rect 9980 1948 10000 2372
rect 9228 1920 10000 1948
rect 10240 2372 11012 2400
rect 10240 1948 10928 2372
rect 10992 1948 11012 2372
rect 10240 1920 11012 1948
rect 11252 2372 12024 2400
rect 11252 1948 11940 2372
rect 12004 1948 12024 2372
rect 11252 1920 12024 1948
rect 12264 2372 13036 2400
rect 12264 1948 12952 2372
rect 13016 1948 13036 2372
rect 12264 1920 13036 1948
rect 13276 2372 14048 2400
rect 13276 1948 13964 2372
rect 14028 1948 14048 2372
rect 13276 1920 14048 1948
rect 14288 2372 15060 2400
rect 14288 1948 14976 2372
rect 15040 1948 15060 2372
rect 14288 1920 15060 1948
rect 15300 2372 16072 2400
rect 15300 1948 15988 2372
rect 16052 1948 16072 2372
rect 15300 1920 16072 1948
rect 16312 2372 17084 2400
rect 16312 1948 17000 2372
rect 17064 1948 17084 2372
rect 16312 1920 17084 1948
rect -17084 1652 -16312 1680
rect -17084 1228 -16396 1652
rect -16332 1228 -16312 1652
rect -17084 1200 -16312 1228
rect -16072 1652 -15300 1680
rect -16072 1228 -15384 1652
rect -15320 1228 -15300 1652
rect -16072 1200 -15300 1228
rect -15060 1652 -14288 1680
rect -15060 1228 -14372 1652
rect -14308 1228 -14288 1652
rect -15060 1200 -14288 1228
rect -14048 1652 -13276 1680
rect -14048 1228 -13360 1652
rect -13296 1228 -13276 1652
rect -14048 1200 -13276 1228
rect -13036 1652 -12264 1680
rect -13036 1228 -12348 1652
rect -12284 1228 -12264 1652
rect -13036 1200 -12264 1228
rect -12024 1652 -11252 1680
rect -12024 1228 -11336 1652
rect -11272 1228 -11252 1652
rect -12024 1200 -11252 1228
rect -11012 1652 -10240 1680
rect -11012 1228 -10324 1652
rect -10260 1228 -10240 1652
rect -11012 1200 -10240 1228
rect -10000 1652 -9228 1680
rect -10000 1228 -9312 1652
rect -9248 1228 -9228 1652
rect -10000 1200 -9228 1228
rect -8988 1652 -8216 1680
rect -8988 1228 -8300 1652
rect -8236 1228 -8216 1652
rect -8988 1200 -8216 1228
rect -7976 1652 -7204 1680
rect -7976 1228 -7288 1652
rect -7224 1228 -7204 1652
rect -7976 1200 -7204 1228
rect -6964 1652 -6192 1680
rect -6964 1228 -6276 1652
rect -6212 1228 -6192 1652
rect -6964 1200 -6192 1228
rect -5952 1652 -5180 1680
rect -5952 1228 -5264 1652
rect -5200 1228 -5180 1652
rect -5952 1200 -5180 1228
rect -4940 1652 -4168 1680
rect -4940 1228 -4252 1652
rect -4188 1228 -4168 1652
rect -4940 1200 -4168 1228
rect -3928 1652 -3156 1680
rect -3928 1228 -3240 1652
rect -3176 1228 -3156 1652
rect -3928 1200 -3156 1228
rect -2916 1652 -2144 1680
rect -2916 1228 -2228 1652
rect -2164 1228 -2144 1652
rect -2916 1200 -2144 1228
rect -1904 1652 -1132 1680
rect -1904 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -1904 1200 -1132 1228
rect -892 1652 -120 1680
rect -892 1228 -204 1652
rect -140 1228 -120 1652
rect -892 1200 -120 1228
rect 120 1652 892 1680
rect 120 1228 808 1652
rect 872 1228 892 1652
rect 120 1200 892 1228
rect 1132 1652 1904 1680
rect 1132 1228 1820 1652
rect 1884 1228 1904 1652
rect 1132 1200 1904 1228
rect 2144 1652 2916 1680
rect 2144 1228 2832 1652
rect 2896 1228 2916 1652
rect 2144 1200 2916 1228
rect 3156 1652 3928 1680
rect 3156 1228 3844 1652
rect 3908 1228 3928 1652
rect 3156 1200 3928 1228
rect 4168 1652 4940 1680
rect 4168 1228 4856 1652
rect 4920 1228 4940 1652
rect 4168 1200 4940 1228
rect 5180 1652 5952 1680
rect 5180 1228 5868 1652
rect 5932 1228 5952 1652
rect 5180 1200 5952 1228
rect 6192 1652 6964 1680
rect 6192 1228 6880 1652
rect 6944 1228 6964 1652
rect 6192 1200 6964 1228
rect 7204 1652 7976 1680
rect 7204 1228 7892 1652
rect 7956 1228 7976 1652
rect 7204 1200 7976 1228
rect 8216 1652 8988 1680
rect 8216 1228 8904 1652
rect 8968 1228 8988 1652
rect 8216 1200 8988 1228
rect 9228 1652 10000 1680
rect 9228 1228 9916 1652
rect 9980 1228 10000 1652
rect 9228 1200 10000 1228
rect 10240 1652 11012 1680
rect 10240 1228 10928 1652
rect 10992 1228 11012 1652
rect 10240 1200 11012 1228
rect 11252 1652 12024 1680
rect 11252 1228 11940 1652
rect 12004 1228 12024 1652
rect 11252 1200 12024 1228
rect 12264 1652 13036 1680
rect 12264 1228 12952 1652
rect 13016 1228 13036 1652
rect 12264 1200 13036 1228
rect 13276 1652 14048 1680
rect 13276 1228 13964 1652
rect 14028 1228 14048 1652
rect 13276 1200 14048 1228
rect 14288 1652 15060 1680
rect 14288 1228 14976 1652
rect 15040 1228 15060 1652
rect 14288 1200 15060 1228
rect 15300 1652 16072 1680
rect 15300 1228 15988 1652
rect 16052 1228 16072 1652
rect 15300 1200 16072 1228
rect 16312 1652 17084 1680
rect 16312 1228 17000 1652
rect 17064 1228 17084 1652
rect 16312 1200 17084 1228
rect -17084 932 -16312 960
rect -17084 508 -16396 932
rect -16332 508 -16312 932
rect -17084 480 -16312 508
rect -16072 932 -15300 960
rect -16072 508 -15384 932
rect -15320 508 -15300 932
rect -16072 480 -15300 508
rect -15060 932 -14288 960
rect -15060 508 -14372 932
rect -14308 508 -14288 932
rect -15060 480 -14288 508
rect -14048 932 -13276 960
rect -14048 508 -13360 932
rect -13296 508 -13276 932
rect -14048 480 -13276 508
rect -13036 932 -12264 960
rect -13036 508 -12348 932
rect -12284 508 -12264 932
rect -13036 480 -12264 508
rect -12024 932 -11252 960
rect -12024 508 -11336 932
rect -11272 508 -11252 932
rect -12024 480 -11252 508
rect -11012 932 -10240 960
rect -11012 508 -10324 932
rect -10260 508 -10240 932
rect -11012 480 -10240 508
rect -10000 932 -9228 960
rect -10000 508 -9312 932
rect -9248 508 -9228 932
rect -10000 480 -9228 508
rect -8988 932 -8216 960
rect -8988 508 -8300 932
rect -8236 508 -8216 932
rect -8988 480 -8216 508
rect -7976 932 -7204 960
rect -7976 508 -7288 932
rect -7224 508 -7204 932
rect -7976 480 -7204 508
rect -6964 932 -6192 960
rect -6964 508 -6276 932
rect -6212 508 -6192 932
rect -6964 480 -6192 508
rect -5952 932 -5180 960
rect -5952 508 -5264 932
rect -5200 508 -5180 932
rect -5952 480 -5180 508
rect -4940 932 -4168 960
rect -4940 508 -4252 932
rect -4188 508 -4168 932
rect -4940 480 -4168 508
rect -3928 932 -3156 960
rect -3928 508 -3240 932
rect -3176 508 -3156 932
rect -3928 480 -3156 508
rect -2916 932 -2144 960
rect -2916 508 -2228 932
rect -2164 508 -2144 932
rect -2916 480 -2144 508
rect -1904 932 -1132 960
rect -1904 508 -1216 932
rect -1152 508 -1132 932
rect -1904 480 -1132 508
rect -892 932 -120 960
rect -892 508 -204 932
rect -140 508 -120 932
rect -892 480 -120 508
rect 120 932 892 960
rect 120 508 808 932
rect 872 508 892 932
rect 120 480 892 508
rect 1132 932 1904 960
rect 1132 508 1820 932
rect 1884 508 1904 932
rect 1132 480 1904 508
rect 2144 932 2916 960
rect 2144 508 2832 932
rect 2896 508 2916 932
rect 2144 480 2916 508
rect 3156 932 3928 960
rect 3156 508 3844 932
rect 3908 508 3928 932
rect 3156 480 3928 508
rect 4168 932 4940 960
rect 4168 508 4856 932
rect 4920 508 4940 932
rect 4168 480 4940 508
rect 5180 932 5952 960
rect 5180 508 5868 932
rect 5932 508 5952 932
rect 5180 480 5952 508
rect 6192 932 6964 960
rect 6192 508 6880 932
rect 6944 508 6964 932
rect 6192 480 6964 508
rect 7204 932 7976 960
rect 7204 508 7892 932
rect 7956 508 7976 932
rect 7204 480 7976 508
rect 8216 932 8988 960
rect 8216 508 8904 932
rect 8968 508 8988 932
rect 8216 480 8988 508
rect 9228 932 10000 960
rect 9228 508 9916 932
rect 9980 508 10000 932
rect 9228 480 10000 508
rect 10240 932 11012 960
rect 10240 508 10928 932
rect 10992 508 11012 932
rect 10240 480 11012 508
rect 11252 932 12024 960
rect 11252 508 11940 932
rect 12004 508 12024 932
rect 11252 480 12024 508
rect 12264 932 13036 960
rect 12264 508 12952 932
rect 13016 508 13036 932
rect 12264 480 13036 508
rect 13276 932 14048 960
rect 13276 508 13964 932
rect 14028 508 14048 932
rect 13276 480 14048 508
rect 14288 932 15060 960
rect 14288 508 14976 932
rect 15040 508 15060 932
rect 14288 480 15060 508
rect 15300 932 16072 960
rect 15300 508 15988 932
rect 16052 508 16072 932
rect 15300 480 16072 508
rect 16312 932 17084 960
rect 16312 508 17000 932
rect 17064 508 17084 932
rect 16312 480 17084 508
rect -17084 212 -16312 240
rect -17084 -212 -16396 212
rect -16332 -212 -16312 212
rect -17084 -240 -16312 -212
rect -16072 212 -15300 240
rect -16072 -212 -15384 212
rect -15320 -212 -15300 212
rect -16072 -240 -15300 -212
rect -15060 212 -14288 240
rect -15060 -212 -14372 212
rect -14308 -212 -14288 212
rect -15060 -240 -14288 -212
rect -14048 212 -13276 240
rect -14048 -212 -13360 212
rect -13296 -212 -13276 212
rect -14048 -240 -13276 -212
rect -13036 212 -12264 240
rect -13036 -212 -12348 212
rect -12284 -212 -12264 212
rect -13036 -240 -12264 -212
rect -12024 212 -11252 240
rect -12024 -212 -11336 212
rect -11272 -212 -11252 212
rect -12024 -240 -11252 -212
rect -11012 212 -10240 240
rect -11012 -212 -10324 212
rect -10260 -212 -10240 212
rect -11012 -240 -10240 -212
rect -10000 212 -9228 240
rect -10000 -212 -9312 212
rect -9248 -212 -9228 212
rect -10000 -240 -9228 -212
rect -8988 212 -8216 240
rect -8988 -212 -8300 212
rect -8236 -212 -8216 212
rect -8988 -240 -8216 -212
rect -7976 212 -7204 240
rect -7976 -212 -7288 212
rect -7224 -212 -7204 212
rect -7976 -240 -7204 -212
rect -6964 212 -6192 240
rect -6964 -212 -6276 212
rect -6212 -212 -6192 212
rect -6964 -240 -6192 -212
rect -5952 212 -5180 240
rect -5952 -212 -5264 212
rect -5200 -212 -5180 212
rect -5952 -240 -5180 -212
rect -4940 212 -4168 240
rect -4940 -212 -4252 212
rect -4188 -212 -4168 212
rect -4940 -240 -4168 -212
rect -3928 212 -3156 240
rect -3928 -212 -3240 212
rect -3176 -212 -3156 212
rect -3928 -240 -3156 -212
rect -2916 212 -2144 240
rect -2916 -212 -2228 212
rect -2164 -212 -2144 212
rect -2916 -240 -2144 -212
rect -1904 212 -1132 240
rect -1904 -212 -1216 212
rect -1152 -212 -1132 212
rect -1904 -240 -1132 -212
rect -892 212 -120 240
rect -892 -212 -204 212
rect -140 -212 -120 212
rect -892 -240 -120 -212
rect 120 212 892 240
rect 120 -212 808 212
rect 872 -212 892 212
rect 120 -240 892 -212
rect 1132 212 1904 240
rect 1132 -212 1820 212
rect 1884 -212 1904 212
rect 1132 -240 1904 -212
rect 2144 212 2916 240
rect 2144 -212 2832 212
rect 2896 -212 2916 212
rect 2144 -240 2916 -212
rect 3156 212 3928 240
rect 3156 -212 3844 212
rect 3908 -212 3928 212
rect 3156 -240 3928 -212
rect 4168 212 4940 240
rect 4168 -212 4856 212
rect 4920 -212 4940 212
rect 4168 -240 4940 -212
rect 5180 212 5952 240
rect 5180 -212 5868 212
rect 5932 -212 5952 212
rect 5180 -240 5952 -212
rect 6192 212 6964 240
rect 6192 -212 6880 212
rect 6944 -212 6964 212
rect 6192 -240 6964 -212
rect 7204 212 7976 240
rect 7204 -212 7892 212
rect 7956 -212 7976 212
rect 7204 -240 7976 -212
rect 8216 212 8988 240
rect 8216 -212 8904 212
rect 8968 -212 8988 212
rect 8216 -240 8988 -212
rect 9228 212 10000 240
rect 9228 -212 9916 212
rect 9980 -212 10000 212
rect 9228 -240 10000 -212
rect 10240 212 11012 240
rect 10240 -212 10928 212
rect 10992 -212 11012 212
rect 10240 -240 11012 -212
rect 11252 212 12024 240
rect 11252 -212 11940 212
rect 12004 -212 12024 212
rect 11252 -240 12024 -212
rect 12264 212 13036 240
rect 12264 -212 12952 212
rect 13016 -212 13036 212
rect 12264 -240 13036 -212
rect 13276 212 14048 240
rect 13276 -212 13964 212
rect 14028 -212 14048 212
rect 13276 -240 14048 -212
rect 14288 212 15060 240
rect 14288 -212 14976 212
rect 15040 -212 15060 212
rect 14288 -240 15060 -212
rect 15300 212 16072 240
rect 15300 -212 15988 212
rect 16052 -212 16072 212
rect 15300 -240 16072 -212
rect 16312 212 17084 240
rect 16312 -212 17000 212
rect 17064 -212 17084 212
rect 16312 -240 17084 -212
rect -17084 -508 -16312 -480
rect -17084 -932 -16396 -508
rect -16332 -932 -16312 -508
rect -17084 -960 -16312 -932
rect -16072 -508 -15300 -480
rect -16072 -932 -15384 -508
rect -15320 -932 -15300 -508
rect -16072 -960 -15300 -932
rect -15060 -508 -14288 -480
rect -15060 -932 -14372 -508
rect -14308 -932 -14288 -508
rect -15060 -960 -14288 -932
rect -14048 -508 -13276 -480
rect -14048 -932 -13360 -508
rect -13296 -932 -13276 -508
rect -14048 -960 -13276 -932
rect -13036 -508 -12264 -480
rect -13036 -932 -12348 -508
rect -12284 -932 -12264 -508
rect -13036 -960 -12264 -932
rect -12024 -508 -11252 -480
rect -12024 -932 -11336 -508
rect -11272 -932 -11252 -508
rect -12024 -960 -11252 -932
rect -11012 -508 -10240 -480
rect -11012 -932 -10324 -508
rect -10260 -932 -10240 -508
rect -11012 -960 -10240 -932
rect -10000 -508 -9228 -480
rect -10000 -932 -9312 -508
rect -9248 -932 -9228 -508
rect -10000 -960 -9228 -932
rect -8988 -508 -8216 -480
rect -8988 -932 -8300 -508
rect -8236 -932 -8216 -508
rect -8988 -960 -8216 -932
rect -7976 -508 -7204 -480
rect -7976 -932 -7288 -508
rect -7224 -932 -7204 -508
rect -7976 -960 -7204 -932
rect -6964 -508 -6192 -480
rect -6964 -932 -6276 -508
rect -6212 -932 -6192 -508
rect -6964 -960 -6192 -932
rect -5952 -508 -5180 -480
rect -5952 -932 -5264 -508
rect -5200 -932 -5180 -508
rect -5952 -960 -5180 -932
rect -4940 -508 -4168 -480
rect -4940 -932 -4252 -508
rect -4188 -932 -4168 -508
rect -4940 -960 -4168 -932
rect -3928 -508 -3156 -480
rect -3928 -932 -3240 -508
rect -3176 -932 -3156 -508
rect -3928 -960 -3156 -932
rect -2916 -508 -2144 -480
rect -2916 -932 -2228 -508
rect -2164 -932 -2144 -508
rect -2916 -960 -2144 -932
rect -1904 -508 -1132 -480
rect -1904 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -1904 -960 -1132 -932
rect -892 -508 -120 -480
rect -892 -932 -204 -508
rect -140 -932 -120 -508
rect -892 -960 -120 -932
rect 120 -508 892 -480
rect 120 -932 808 -508
rect 872 -932 892 -508
rect 120 -960 892 -932
rect 1132 -508 1904 -480
rect 1132 -932 1820 -508
rect 1884 -932 1904 -508
rect 1132 -960 1904 -932
rect 2144 -508 2916 -480
rect 2144 -932 2832 -508
rect 2896 -932 2916 -508
rect 2144 -960 2916 -932
rect 3156 -508 3928 -480
rect 3156 -932 3844 -508
rect 3908 -932 3928 -508
rect 3156 -960 3928 -932
rect 4168 -508 4940 -480
rect 4168 -932 4856 -508
rect 4920 -932 4940 -508
rect 4168 -960 4940 -932
rect 5180 -508 5952 -480
rect 5180 -932 5868 -508
rect 5932 -932 5952 -508
rect 5180 -960 5952 -932
rect 6192 -508 6964 -480
rect 6192 -932 6880 -508
rect 6944 -932 6964 -508
rect 6192 -960 6964 -932
rect 7204 -508 7976 -480
rect 7204 -932 7892 -508
rect 7956 -932 7976 -508
rect 7204 -960 7976 -932
rect 8216 -508 8988 -480
rect 8216 -932 8904 -508
rect 8968 -932 8988 -508
rect 8216 -960 8988 -932
rect 9228 -508 10000 -480
rect 9228 -932 9916 -508
rect 9980 -932 10000 -508
rect 9228 -960 10000 -932
rect 10240 -508 11012 -480
rect 10240 -932 10928 -508
rect 10992 -932 11012 -508
rect 10240 -960 11012 -932
rect 11252 -508 12024 -480
rect 11252 -932 11940 -508
rect 12004 -932 12024 -508
rect 11252 -960 12024 -932
rect 12264 -508 13036 -480
rect 12264 -932 12952 -508
rect 13016 -932 13036 -508
rect 12264 -960 13036 -932
rect 13276 -508 14048 -480
rect 13276 -932 13964 -508
rect 14028 -932 14048 -508
rect 13276 -960 14048 -932
rect 14288 -508 15060 -480
rect 14288 -932 14976 -508
rect 15040 -932 15060 -508
rect 14288 -960 15060 -932
rect 15300 -508 16072 -480
rect 15300 -932 15988 -508
rect 16052 -932 16072 -508
rect 15300 -960 16072 -932
rect 16312 -508 17084 -480
rect 16312 -932 17000 -508
rect 17064 -932 17084 -508
rect 16312 -960 17084 -932
rect -17084 -1228 -16312 -1200
rect -17084 -1652 -16396 -1228
rect -16332 -1652 -16312 -1228
rect -17084 -1680 -16312 -1652
rect -16072 -1228 -15300 -1200
rect -16072 -1652 -15384 -1228
rect -15320 -1652 -15300 -1228
rect -16072 -1680 -15300 -1652
rect -15060 -1228 -14288 -1200
rect -15060 -1652 -14372 -1228
rect -14308 -1652 -14288 -1228
rect -15060 -1680 -14288 -1652
rect -14048 -1228 -13276 -1200
rect -14048 -1652 -13360 -1228
rect -13296 -1652 -13276 -1228
rect -14048 -1680 -13276 -1652
rect -13036 -1228 -12264 -1200
rect -13036 -1652 -12348 -1228
rect -12284 -1652 -12264 -1228
rect -13036 -1680 -12264 -1652
rect -12024 -1228 -11252 -1200
rect -12024 -1652 -11336 -1228
rect -11272 -1652 -11252 -1228
rect -12024 -1680 -11252 -1652
rect -11012 -1228 -10240 -1200
rect -11012 -1652 -10324 -1228
rect -10260 -1652 -10240 -1228
rect -11012 -1680 -10240 -1652
rect -10000 -1228 -9228 -1200
rect -10000 -1652 -9312 -1228
rect -9248 -1652 -9228 -1228
rect -10000 -1680 -9228 -1652
rect -8988 -1228 -8216 -1200
rect -8988 -1652 -8300 -1228
rect -8236 -1652 -8216 -1228
rect -8988 -1680 -8216 -1652
rect -7976 -1228 -7204 -1200
rect -7976 -1652 -7288 -1228
rect -7224 -1652 -7204 -1228
rect -7976 -1680 -7204 -1652
rect -6964 -1228 -6192 -1200
rect -6964 -1652 -6276 -1228
rect -6212 -1652 -6192 -1228
rect -6964 -1680 -6192 -1652
rect -5952 -1228 -5180 -1200
rect -5952 -1652 -5264 -1228
rect -5200 -1652 -5180 -1228
rect -5952 -1680 -5180 -1652
rect -4940 -1228 -4168 -1200
rect -4940 -1652 -4252 -1228
rect -4188 -1652 -4168 -1228
rect -4940 -1680 -4168 -1652
rect -3928 -1228 -3156 -1200
rect -3928 -1652 -3240 -1228
rect -3176 -1652 -3156 -1228
rect -3928 -1680 -3156 -1652
rect -2916 -1228 -2144 -1200
rect -2916 -1652 -2228 -1228
rect -2164 -1652 -2144 -1228
rect -2916 -1680 -2144 -1652
rect -1904 -1228 -1132 -1200
rect -1904 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -1904 -1680 -1132 -1652
rect -892 -1228 -120 -1200
rect -892 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect -892 -1680 -120 -1652
rect 120 -1228 892 -1200
rect 120 -1652 808 -1228
rect 872 -1652 892 -1228
rect 120 -1680 892 -1652
rect 1132 -1228 1904 -1200
rect 1132 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 1132 -1680 1904 -1652
rect 2144 -1228 2916 -1200
rect 2144 -1652 2832 -1228
rect 2896 -1652 2916 -1228
rect 2144 -1680 2916 -1652
rect 3156 -1228 3928 -1200
rect 3156 -1652 3844 -1228
rect 3908 -1652 3928 -1228
rect 3156 -1680 3928 -1652
rect 4168 -1228 4940 -1200
rect 4168 -1652 4856 -1228
rect 4920 -1652 4940 -1228
rect 4168 -1680 4940 -1652
rect 5180 -1228 5952 -1200
rect 5180 -1652 5868 -1228
rect 5932 -1652 5952 -1228
rect 5180 -1680 5952 -1652
rect 6192 -1228 6964 -1200
rect 6192 -1652 6880 -1228
rect 6944 -1652 6964 -1228
rect 6192 -1680 6964 -1652
rect 7204 -1228 7976 -1200
rect 7204 -1652 7892 -1228
rect 7956 -1652 7976 -1228
rect 7204 -1680 7976 -1652
rect 8216 -1228 8988 -1200
rect 8216 -1652 8904 -1228
rect 8968 -1652 8988 -1228
rect 8216 -1680 8988 -1652
rect 9228 -1228 10000 -1200
rect 9228 -1652 9916 -1228
rect 9980 -1652 10000 -1228
rect 9228 -1680 10000 -1652
rect 10240 -1228 11012 -1200
rect 10240 -1652 10928 -1228
rect 10992 -1652 11012 -1228
rect 10240 -1680 11012 -1652
rect 11252 -1228 12024 -1200
rect 11252 -1652 11940 -1228
rect 12004 -1652 12024 -1228
rect 11252 -1680 12024 -1652
rect 12264 -1228 13036 -1200
rect 12264 -1652 12952 -1228
rect 13016 -1652 13036 -1228
rect 12264 -1680 13036 -1652
rect 13276 -1228 14048 -1200
rect 13276 -1652 13964 -1228
rect 14028 -1652 14048 -1228
rect 13276 -1680 14048 -1652
rect 14288 -1228 15060 -1200
rect 14288 -1652 14976 -1228
rect 15040 -1652 15060 -1228
rect 14288 -1680 15060 -1652
rect 15300 -1228 16072 -1200
rect 15300 -1652 15988 -1228
rect 16052 -1652 16072 -1228
rect 15300 -1680 16072 -1652
rect 16312 -1228 17084 -1200
rect 16312 -1652 17000 -1228
rect 17064 -1652 17084 -1228
rect 16312 -1680 17084 -1652
rect -17084 -1948 -16312 -1920
rect -17084 -2372 -16396 -1948
rect -16332 -2372 -16312 -1948
rect -17084 -2400 -16312 -2372
rect -16072 -1948 -15300 -1920
rect -16072 -2372 -15384 -1948
rect -15320 -2372 -15300 -1948
rect -16072 -2400 -15300 -2372
rect -15060 -1948 -14288 -1920
rect -15060 -2372 -14372 -1948
rect -14308 -2372 -14288 -1948
rect -15060 -2400 -14288 -2372
rect -14048 -1948 -13276 -1920
rect -14048 -2372 -13360 -1948
rect -13296 -2372 -13276 -1948
rect -14048 -2400 -13276 -2372
rect -13036 -1948 -12264 -1920
rect -13036 -2372 -12348 -1948
rect -12284 -2372 -12264 -1948
rect -13036 -2400 -12264 -2372
rect -12024 -1948 -11252 -1920
rect -12024 -2372 -11336 -1948
rect -11272 -2372 -11252 -1948
rect -12024 -2400 -11252 -2372
rect -11012 -1948 -10240 -1920
rect -11012 -2372 -10324 -1948
rect -10260 -2372 -10240 -1948
rect -11012 -2400 -10240 -2372
rect -10000 -1948 -9228 -1920
rect -10000 -2372 -9312 -1948
rect -9248 -2372 -9228 -1948
rect -10000 -2400 -9228 -2372
rect -8988 -1948 -8216 -1920
rect -8988 -2372 -8300 -1948
rect -8236 -2372 -8216 -1948
rect -8988 -2400 -8216 -2372
rect -7976 -1948 -7204 -1920
rect -7976 -2372 -7288 -1948
rect -7224 -2372 -7204 -1948
rect -7976 -2400 -7204 -2372
rect -6964 -1948 -6192 -1920
rect -6964 -2372 -6276 -1948
rect -6212 -2372 -6192 -1948
rect -6964 -2400 -6192 -2372
rect -5952 -1948 -5180 -1920
rect -5952 -2372 -5264 -1948
rect -5200 -2372 -5180 -1948
rect -5952 -2400 -5180 -2372
rect -4940 -1948 -4168 -1920
rect -4940 -2372 -4252 -1948
rect -4188 -2372 -4168 -1948
rect -4940 -2400 -4168 -2372
rect -3928 -1948 -3156 -1920
rect -3928 -2372 -3240 -1948
rect -3176 -2372 -3156 -1948
rect -3928 -2400 -3156 -2372
rect -2916 -1948 -2144 -1920
rect -2916 -2372 -2228 -1948
rect -2164 -2372 -2144 -1948
rect -2916 -2400 -2144 -2372
rect -1904 -1948 -1132 -1920
rect -1904 -2372 -1216 -1948
rect -1152 -2372 -1132 -1948
rect -1904 -2400 -1132 -2372
rect -892 -1948 -120 -1920
rect -892 -2372 -204 -1948
rect -140 -2372 -120 -1948
rect -892 -2400 -120 -2372
rect 120 -1948 892 -1920
rect 120 -2372 808 -1948
rect 872 -2372 892 -1948
rect 120 -2400 892 -2372
rect 1132 -1948 1904 -1920
rect 1132 -2372 1820 -1948
rect 1884 -2372 1904 -1948
rect 1132 -2400 1904 -2372
rect 2144 -1948 2916 -1920
rect 2144 -2372 2832 -1948
rect 2896 -2372 2916 -1948
rect 2144 -2400 2916 -2372
rect 3156 -1948 3928 -1920
rect 3156 -2372 3844 -1948
rect 3908 -2372 3928 -1948
rect 3156 -2400 3928 -2372
rect 4168 -1948 4940 -1920
rect 4168 -2372 4856 -1948
rect 4920 -2372 4940 -1948
rect 4168 -2400 4940 -2372
rect 5180 -1948 5952 -1920
rect 5180 -2372 5868 -1948
rect 5932 -2372 5952 -1948
rect 5180 -2400 5952 -2372
rect 6192 -1948 6964 -1920
rect 6192 -2372 6880 -1948
rect 6944 -2372 6964 -1948
rect 6192 -2400 6964 -2372
rect 7204 -1948 7976 -1920
rect 7204 -2372 7892 -1948
rect 7956 -2372 7976 -1948
rect 7204 -2400 7976 -2372
rect 8216 -1948 8988 -1920
rect 8216 -2372 8904 -1948
rect 8968 -2372 8988 -1948
rect 8216 -2400 8988 -2372
rect 9228 -1948 10000 -1920
rect 9228 -2372 9916 -1948
rect 9980 -2372 10000 -1948
rect 9228 -2400 10000 -2372
rect 10240 -1948 11012 -1920
rect 10240 -2372 10928 -1948
rect 10992 -2372 11012 -1948
rect 10240 -2400 11012 -2372
rect 11252 -1948 12024 -1920
rect 11252 -2372 11940 -1948
rect 12004 -2372 12024 -1948
rect 11252 -2400 12024 -2372
rect 12264 -1948 13036 -1920
rect 12264 -2372 12952 -1948
rect 13016 -2372 13036 -1948
rect 12264 -2400 13036 -2372
rect 13276 -1948 14048 -1920
rect 13276 -2372 13964 -1948
rect 14028 -2372 14048 -1948
rect 13276 -2400 14048 -2372
rect 14288 -1948 15060 -1920
rect 14288 -2372 14976 -1948
rect 15040 -2372 15060 -1948
rect 14288 -2400 15060 -2372
rect 15300 -1948 16072 -1920
rect 15300 -2372 15988 -1948
rect 16052 -2372 16072 -1948
rect 15300 -2400 16072 -2372
rect 16312 -1948 17084 -1920
rect 16312 -2372 17000 -1948
rect 17064 -2372 17084 -1948
rect 16312 -2400 17084 -2372
rect -17084 -2668 -16312 -2640
rect -17084 -3092 -16396 -2668
rect -16332 -3092 -16312 -2668
rect -17084 -3120 -16312 -3092
rect -16072 -2668 -15300 -2640
rect -16072 -3092 -15384 -2668
rect -15320 -3092 -15300 -2668
rect -16072 -3120 -15300 -3092
rect -15060 -2668 -14288 -2640
rect -15060 -3092 -14372 -2668
rect -14308 -3092 -14288 -2668
rect -15060 -3120 -14288 -3092
rect -14048 -2668 -13276 -2640
rect -14048 -3092 -13360 -2668
rect -13296 -3092 -13276 -2668
rect -14048 -3120 -13276 -3092
rect -13036 -2668 -12264 -2640
rect -13036 -3092 -12348 -2668
rect -12284 -3092 -12264 -2668
rect -13036 -3120 -12264 -3092
rect -12024 -2668 -11252 -2640
rect -12024 -3092 -11336 -2668
rect -11272 -3092 -11252 -2668
rect -12024 -3120 -11252 -3092
rect -11012 -2668 -10240 -2640
rect -11012 -3092 -10324 -2668
rect -10260 -3092 -10240 -2668
rect -11012 -3120 -10240 -3092
rect -10000 -2668 -9228 -2640
rect -10000 -3092 -9312 -2668
rect -9248 -3092 -9228 -2668
rect -10000 -3120 -9228 -3092
rect -8988 -2668 -8216 -2640
rect -8988 -3092 -8300 -2668
rect -8236 -3092 -8216 -2668
rect -8988 -3120 -8216 -3092
rect -7976 -2668 -7204 -2640
rect -7976 -3092 -7288 -2668
rect -7224 -3092 -7204 -2668
rect -7976 -3120 -7204 -3092
rect -6964 -2668 -6192 -2640
rect -6964 -3092 -6276 -2668
rect -6212 -3092 -6192 -2668
rect -6964 -3120 -6192 -3092
rect -5952 -2668 -5180 -2640
rect -5952 -3092 -5264 -2668
rect -5200 -3092 -5180 -2668
rect -5952 -3120 -5180 -3092
rect -4940 -2668 -4168 -2640
rect -4940 -3092 -4252 -2668
rect -4188 -3092 -4168 -2668
rect -4940 -3120 -4168 -3092
rect -3928 -2668 -3156 -2640
rect -3928 -3092 -3240 -2668
rect -3176 -3092 -3156 -2668
rect -3928 -3120 -3156 -3092
rect -2916 -2668 -2144 -2640
rect -2916 -3092 -2228 -2668
rect -2164 -3092 -2144 -2668
rect -2916 -3120 -2144 -3092
rect -1904 -2668 -1132 -2640
rect -1904 -3092 -1216 -2668
rect -1152 -3092 -1132 -2668
rect -1904 -3120 -1132 -3092
rect -892 -2668 -120 -2640
rect -892 -3092 -204 -2668
rect -140 -3092 -120 -2668
rect -892 -3120 -120 -3092
rect 120 -2668 892 -2640
rect 120 -3092 808 -2668
rect 872 -3092 892 -2668
rect 120 -3120 892 -3092
rect 1132 -2668 1904 -2640
rect 1132 -3092 1820 -2668
rect 1884 -3092 1904 -2668
rect 1132 -3120 1904 -3092
rect 2144 -2668 2916 -2640
rect 2144 -3092 2832 -2668
rect 2896 -3092 2916 -2668
rect 2144 -3120 2916 -3092
rect 3156 -2668 3928 -2640
rect 3156 -3092 3844 -2668
rect 3908 -3092 3928 -2668
rect 3156 -3120 3928 -3092
rect 4168 -2668 4940 -2640
rect 4168 -3092 4856 -2668
rect 4920 -3092 4940 -2668
rect 4168 -3120 4940 -3092
rect 5180 -2668 5952 -2640
rect 5180 -3092 5868 -2668
rect 5932 -3092 5952 -2668
rect 5180 -3120 5952 -3092
rect 6192 -2668 6964 -2640
rect 6192 -3092 6880 -2668
rect 6944 -3092 6964 -2668
rect 6192 -3120 6964 -3092
rect 7204 -2668 7976 -2640
rect 7204 -3092 7892 -2668
rect 7956 -3092 7976 -2668
rect 7204 -3120 7976 -3092
rect 8216 -2668 8988 -2640
rect 8216 -3092 8904 -2668
rect 8968 -3092 8988 -2668
rect 8216 -3120 8988 -3092
rect 9228 -2668 10000 -2640
rect 9228 -3092 9916 -2668
rect 9980 -3092 10000 -2668
rect 9228 -3120 10000 -3092
rect 10240 -2668 11012 -2640
rect 10240 -3092 10928 -2668
rect 10992 -3092 11012 -2668
rect 10240 -3120 11012 -3092
rect 11252 -2668 12024 -2640
rect 11252 -3092 11940 -2668
rect 12004 -3092 12024 -2668
rect 11252 -3120 12024 -3092
rect 12264 -2668 13036 -2640
rect 12264 -3092 12952 -2668
rect 13016 -3092 13036 -2668
rect 12264 -3120 13036 -3092
rect 13276 -2668 14048 -2640
rect 13276 -3092 13964 -2668
rect 14028 -3092 14048 -2668
rect 13276 -3120 14048 -3092
rect 14288 -2668 15060 -2640
rect 14288 -3092 14976 -2668
rect 15040 -3092 15060 -2668
rect 14288 -3120 15060 -3092
rect 15300 -2668 16072 -2640
rect 15300 -3092 15988 -2668
rect 16052 -3092 16072 -2668
rect 15300 -3120 16072 -3092
rect 16312 -2668 17084 -2640
rect 16312 -3092 17000 -2668
rect 17064 -3092 17084 -2668
rect 16312 -3120 17084 -3092
rect -17084 -3388 -16312 -3360
rect -17084 -3812 -16396 -3388
rect -16332 -3812 -16312 -3388
rect -17084 -3840 -16312 -3812
rect -16072 -3388 -15300 -3360
rect -16072 -3812 -15384 -3388
rect -15320 -3812 -15300 -3388
rect -16072 -3840 -15300 -3812
rect -15060 -3388 -14288 -3360
rect -15060 -3812 -14372 -3388
rect -14308 -3812 -14288 -3388
rect -15060 -3840 -14288 -3812
rect -14048 -3388 -13276 -3360
rect -14048 -3812 -13360 -3388
rect -13296 -3812 -13276 -3388
rect -14048 -3840 -13276 -3812
rect -13036 -3388 -12264 -3360
rect -13036 -3812 -12348 -3388
rect -12284 -3812 -12264 -3388
rect -13036 -3840 -12264 -3812
rect -12024 -3388 -11252 -3360
rect -12024 -3812 -11336 -3388
rect -11272 -3812 -11252 -3388
rect -12024 -3840 -11252 -3812
rect -11012 -3388 -10240 -3360
rect -11012 -3812 -10324 -3388
rect -10260 -3812 -10240 -3388
rect -11012 -3840 -10240 -3812
rect -10000 -3388 -9228 -3360
rect -10000 -3812 -9312 -3388
rect -9248 -3812 -9228 -3388
rect -10000 -3840 -9228 -3812
rect -8988 -3388 -8216 -3360
rect -8988 -3812 -8300 -3388
rect -8236 -3812 -8216 -3388
rect -8988 -3840 -8216 -3812
rect -7976 -3388 -7204 -3360
rect -7976 -3812 -7288 -3388
rect -7224 -3812 -7204 -3388
rect -7976 -3840 -7204 -3812
rect -6964 -3388 -6192 -3360
rect -6964 -3812 -6276 -3388
rect -6212 -3812 -6192 -3388
rect -6964 -3840 -6192 -3812
rect -5952 -3388 -5180 -3360
rect -5952 -3812 -5264 -3388
rect -5200 -3812 -5180 -3388
rect -5952 -3840 -5180 -3812
rect -4940 -3388 -4168 -3360
rect -4940 -3812 -4252 -3388
rect -4188 -3812 -4168 -3388
rect -4940 -3840 -4168 -3812
rect -3928 -3388 -3156 -3360
rect -3928 -3812 -3240 -3388
rect -3176 -3812 -3156 -3388
rect -3928 -3840 -3156 -3812
rect -2916 -3388 -2144 -3360
rect -2916 -3812 -2228 -3388
rect -2164 -3812 -2144 -3388
rect -2916 -3840 -2144 -3812
rect -1904 -3388 -1132 -3360
rect -1904 -3812 -1216 -3388
rect -1152 -3812 -1132 -3388
rect -1904 -3840 -1132 -3812
rect -892 -3388 -120 -3360
rect -892 -3812 -204 -3388
rect -140 -3812 -120 -3388
rect -892 -3840 -120 -3812
rect 120 -3388 892 -3360
rect 120 -3812 808 -3388
rect 872 -3812 892 -3388
rect 120 -3840 892 -3812
rect 1132 -3388 1904 -3360
rect 1132 -3812 1820 -3388
rect 1884 -3812 1904 -3388
rect 1132 -3840 1904 -3812
rect 2144 -3388 2916 -3360
rect 2144 -3812 2832 -3388
rect 2896 -3812 2916 -3388
rect 2144 -3840 2916 -3812
rect 3156 -3388 3928 -3360
rect 3156 -3812 3844 -3388
rect 3908 -3812 3928 -3388
rect 3156 -3840 3928 -3812
rect 4168 -3388 4940 -3360
rect 4168 -3812 4856 -3388
rect 4920 -3812 4940 -3388
rect 4168 -3840 4940 -3812
rect 5180 -3388 5952 -3360
rect 5180 -3812 5868 -3388
rect 5932 -3812 5952 -3388
rect 5180 -3840 5952 -3812
rect 6192 -3388 6964 -3360
rect 6192 -3812 6880 -3388
rect 6944 -3812 6964 -3388
rect 6192 -3840 6964 -3812
rect 7204 -3388 7976 -3360
rect 7204 -3812 7892 -3388
rect 7956 -3812 7976 -3388
rect 7204 -3840 7976 -3812
rect 8216 -3388 8988 -3360
rect 8216 -3812 8904 -3388
rect 8968 -3812 8988 -3388
rect 8216 -3840 8988 -3812
rect 9228 -3388 10000 -3360
rect 9228 -3812 9916 -3388
rect 9980 -3812 10000 -3388
rect 9228 -3840 10000 -3812
rect 10240 -3388 11012 -3360
rect 10240 -3812 10928 -3388
rect 10992 -3812 11012 -3388
rect 10240 -3840 11012 -3812
rect 11252 -3388 12024 -3360
rect 11252 -3812 11940 -3388
rect 12004 -3812 12024 -3388
rect 11252 -3840 12024 -3812
rect 12264 -3388 13036 -3360
rect 12264 -3812 12952 -3388
rect 13016 -3812 13036 -3388
rect 12264 -3840 13036 -3812
rect 13276 -3388 14048 -3360
rect 13276 -3812 13964 -3388
rect 14028 -3812 14048 -3388
rect 13276 -3840 14048 -3812
rect 14288 -3388 15060 -3360
rect 14288 -3812 14976 -3388
rect 15040 -3812 15060 -3388
rect 14288 -3840 15060 -3812
rect 15300 -3388 16072 -3360
rect 15300 -3812 15988 -3388
rect 16052 -3812 16072 -3388
rect 15300 -3840 16072 -3812
rect 16312 -3388 17084 -3360
rect 16312 -3812 17000 -3388
rect 17064 -3812 17084 -3388
rect 16312 -3840 17084 -3812
rect -17084 -4108 -16312 -4080
rect -17084 -4532 -16396 -4108
rect -16332 -4532 -16312 -4108
rect -17084 -4560 -16312 -4532
rect -16072 -4108 -15300 -4080
rect -16072 -4532 -15384 -4108
rect -15320 -4532 -15300 -4108
rect -16072 -4560 -15300 -4532
rect -15060 -4108 -14288 -4080
rect -15060 -4532 -14372 -4108
rect -14308 -4532 -14288 -4108
rect -15060 -4560 -14288 -4532
rect -14048 -4108 -13276 -4080
rect -14048 -4532 -13360 -4108
rect -13296 -4532 -13276 -4108
rect -14048 -4560 -13276 -4532
rect -13036 -4108 -12264 -4080
rect -13036 -4532 -12348 -4108
rect -12284 -4532 -12264 -4108
rect -13036 -4560 -12264 -4532
rect -12024 -4108 -11252 -4080
rect -12024 -4532 -11336 -4108
rect -11272 -4532 -11252 -4108
rect -12024 -4560 -11252 -4532
rect -11012 -4108 -10240 -4080
rect -11012 -4532 -10324 -4108
rect -10260 -4532 -10240 -4108
rect -11012 -4560 -10240 -4532
rect -10000 -4108 -9228 -4080
rect -10000 -4532 -9312 -4108
rect -9248 -4532 -9228 -4108
rect -10000 -4560 -9228 -4532
rect -8988 -4108 -8216 -4080
rect -8988 -4532 -8300 -4108
rect -8236 -4532 -8216 -4108
rect -8988 -4560 -8216 -4532
rect -7976 -4108 -7204 -4080
rect -7976 -4532 -7288 -4108
rect -7224 -4532 -7204 -4108
rect -7976 -4560 -7204 -4532
rect -6964 -4108 -6192 -4080
rect -6964 -4532 -6276 -4108
rect -6212 -4532 -6192 -4108
rect -6964 -4560 -6192 -4532
rect -5952 -4108 -5180 -4080
rect -5952 -4532 -5264 -4108
rect -5200 -4532 -5180 -4108
rect -5952 -4560 -5180 -4532
rect -4940 -4108 -4168 -4080
rect -4940 -4532 -4252 -4108
rect -4188 -4532 -4168 -4108
rect -4940 -4560 -4168 -4532
rect -3928 -4108 -3156 -4080
rect -3928 -4532 -3240 -4108
rect -3176 -4532 -3156 -4108
rect -3928 -4560 -3156 -4532
rect -2916 -4108 -2144 -4080
rect -2916 -4532 -2228 -4108
rect -2164 -4532 -2144 -4108
rect -2916 -4560 -2144 -4532
rect -1904 -4108 -1132 -4080
rect -1904 -4532 -1216 -4108
rect -1152 -4532 -1132 -4108
rect -1904 -4560 -1132 -4532
rect -892 -4108 -120 -4080
rect -892 -4532 -204 -4108
rect -140 -4532 -120 -4108
rect -892 -4560 -120 -4532
rect 120 -4108 892 -4080
rect 120 -4532 808 -4108
rect 872 -4532 892 -4108
rect 120 -4560 892 -4532
rect 1132 -4108 1904 -4080
rect 1132 -4532 1820 -4108
rect 1884 -4532 1904 -4108
rect 1132 -4560 1904 -4532
rect 2144 -4108 2916 -4080
rect 2144 -4532 2832 -4108
rect 2896 -4532 2916 -4108
rect 2144 -4560 2916 -4532
rect 3156 -4108 3928 -4080
rect 3156 -4532 3844 -4108
rect 3908 -4532 3928 -4108
rect 3156 -4560 3928 -4532
rect 4168 -4108 4940 -4080
rect 4168 -4532 4856 -4108
rect 4920 -4532 4940 -4108
rect 4168 -4560 4940 -4532
rect 5180 -4108 5952 -4080
rect 5180 -4532 5868 -4108
rect 5932 -4532 5952 -4108
rect 5180 -4560 5952 -4532
rect 6192 -4108 6964 -4080
rect 6192 -4532 6880 -4108
rect 6944 -4532 6964 -4108
rect 6192 -4560 6964 -4532
rect 7204 -4108 7976 -4080
rect 7204 -4532 7892 -4108
rect 7956 -4532 7976 -4108
rect 7204 -4560 7976 -4532
rect 8216 -4108 8988 -4080
rect 8216 -4532 8904 -4108
rect 8968 -4532 8988 -4108
rect 8216 -4560 8988 -4532
rect 9228 -4108 10000 -4080
rect 9228 -4532 9916 -4108
rect 9980 -4532 10000 -4108
rect 9228 -4560 10000 -4532
rect 10240 -4108 11012 -4080
rect 10240 -4532 10928 -4108
rect 10992 -4532 11012 -4108
rect 10240 -4560 11012 -4532
rect 11252 -4108 12024 -4080
rect 11252 -4532 11940 -4108
rect 12004 -4532 12024 -4108
rect 11252 -4560 12024 -4532
rect 12264 -4108 13036 -4080
rect 12264 -4532 12952 -4108
rect 13016 -4532 13036 -4108
rect 12264 -4560 13036 -4532
rect 13276 -4108 14048 -4080
rect 13276 -4532 13964 -4108
rect 14028 -4532 14048 -4108
rect 13276 -4560 14048 -4532
rect 14288 -4108 15060 -4080
rect 14288 -4532 14976 -4108
rect 15040 -4532 15060 -4108
rect 14288 -4560 15060 -4532
rect 15300 -4108 16072 -4080
rect 15300 -4532 15988 -4108
rect 16052 -4532 16072 -4108
rect 15300 -4560 16072 -4532
rect 16312 -4108 17084 -4080
rect 16312 -4532 17000 -4108
rect 17064 -4532 17084 -4108
rect 16312 -4560 17084 -4532
rect -17084 -4828 -16312 -4800
rect -17084 -5252 -16396 -4828
rect -16332 -5252 -16312 -4828
rect -17084 -5280 -16312 -5252
rect -16072 -4828 -15300 -4800
rect -16072 -5252 -15384 -4828
rect -15320 -5252 -15300 -4828
rect -16072 -5280 -15300 -5252
rect -15060 -4828 -14288 -4800
rect -15060 -5252 -14372 -4828
rect -14308 -5252 -14288 -4828
rect -15060 -5280 -14288 -5252
rect -14048 -4828 -13276 -4800
rect -14048 -5252 -13360 -4828
rect -13296 -5252 -13276 -4828
rect -14048 -5280 -13276 -5252
rect -13036 -4828 -12264 -4800
rect -13036 -5252 -12348 -4828
rect -12284 -5252 -12264 -4828
rect -13036 -5280 -12264 -5252
rect -12024 -4828 -11252 -4800
rect -12024 -5252 -11336 -4828
rect -11272 -5252 -11252 -4828
rect -12024 -5280 -11252 -5252
rect -11012 -4828 -10240 -4800
rect -11012 -5252 -10324 -4828
rect -10260 -5252 -10240 -4828
rect -11012 -5280 -10240 -5252
rect -10000 -4828 -9228 -4800
rect -10000 -5252 -9312 -4828
rect -9248 -5252 -9228 -4828
rect -10000 -5280 -9228 -5252
rect -8988 -4828 -8216 -4800
rect -8988 -5252 -8300 -4828
rect -8236 -5252 -8216 -4828
rect -8988 -5280 -8216 -5252
rect -7976 -4828 -7204 -4800
rect -7976 -5252 -7288 -4828
rect -7224 -5252 -7204 -4828
rect -7976 -5280 -7204 -5252
rect -6964 -4828 -6192 -4800
rect -6964 -5252 -6276 -4828
rect -6212 -5252 -6192 -4828
rect -6964 -5280 -6192 -5252
rect -5952 -4828 -5180 -4800
rect -5952 -5252 -5264 -4828
rect -5200 -5252 -5180 -4828
rect -5952 -5280 -5180 -5252
rect -4940 -4828 -4168 -4800
rect -4940 -5252 -4252 -4828
rect -4188 -5252 -4168 -4828
rect -4940 -5280 -4168 -5252
rect -3928 -4828 -3156 -4800
rect -3928 -5252 -3240 -4828
rect -3176 -5252 -3156 -4828
rect -3928 -5280 -3156 -5252
rect -2916 -4828 -2144 -4800
rect -2916 -5252 -2228 -4828
rect -2164 -5252 -2144 -4828
rect -2916 -5280 -2144 -5252
rect -1904 -4828 -1132 -4800
rect -1904 -5252 -1216 -4828
rect -1152 -5252 -1132 -4828
rect -1904 -5280 -1132 -5252
rect -892 -4828 -120 -4800
rect -892 -5252 -204 -4828
rect -140 -5252 -120 -4828
rect -892 -5280 -120 -5252
rect 120 -4828 892 -4800
rect 120 -5252 808 -4828
rect 872 -5252 892 -4828
rect 120 -5280 892 -5252
rect 1132 -4828 1904 -4800
rect 1132 -5252 1820 -4828
rect 1884 -5252 1904 -4828
rect 1132 -5280 1904 -5252
rect 2144 -4828 2916 -4800
rect 2144 -5252 2832 -4828
rect 2896 -5252 2916 -4828
rect 2144 -5280 2916 -5252
rect 3156 -4828 3928 -4800
rect 3156 -5252 3844 -4828
rect 3908 -5252 3928 -4828
rect 3156 -5280 3928 -5252
rect 4168 -4828 4940 -4800
rect 4168 -5252 4856 -4828
rect 4920 -5252 4940 -4828
rect 4168 -5280 4940 -5252
rect 5180 -4828 5952 -4800
rect 5180 -5252 5868 -4828
rect 5932 -5252 5952 -4828
rect 5180 -5280 5952 -5252
rect 6192 -4828 6964 -4800
rect 6192 -5252 6880 -4828
rect 6944 -5252 6964 -4828
rect 6192 -5280 6964 -5252
rect 7204 -4828 7976 -4800
rect 7204 -5252 7892 -4828
rect 7956 -5252 7976 -4828
rect 7204 -5280 7976 -5252
rect 8216 -4828 8988 -4800
rect 8216 -5252 8904 -4828
rect 8968 -5252 8988 -4828
rect 8216 -5280 8988 -5252
rect 9228 -4828 10000 -4800
rect 9228 -5252 9916 -4828
rect 9980 -5252 10000 -4828
rect 9228 -5280 10000 -5252
rect 10240 -4828 11012 -4800
rect 10240 -5252 10928 -4828
rect 10992 -5252 11012 -4828
rect 10240 -5280 11012 -5252
rect 11252 -4828 12024 -4800
rect 11252 -5252 11940 -4828
rect 12004 -5252 12024 -4828
rect 11252 -5280 12024 -5252
rect 12264 -4828 13036 -4800
rect 12264 -5252 12952 -4828
rect 13016 -5252 13036 -4828
rect 12264 -5280 13036 -5252
rect 13276 -4828 14048 -4800
rect 13276 -5252 13964 -4828
rect 14028 -5252 14048 -4828
rect 13276 -5280 14048 -5252
rect 14288 -4828 15060 -4800
rect 14288 -5252 14976 -4828
rect 15040 -5252 15060 -4828
rect 14288 -5280 15060 -5252
rect 15300 -4828 16072 -4800
rect 15300 -5252 15988 -4828
rect 16052 -5252 16072 -4828
rect 15300 -5280 16072 -5252
rect 16312 -4828 17084 -4800
rect 16312 -5252 17000 -4828
rect 17064 -5252 17084 -4828
rect 16312 -5280 17084 -5252
rect -17084 -5548 -16312 -5520
rect -17084 -5972 -16396 -5548
rect -16332 -5972 -16312 -5548
rect -17084 -6000 -16312 -5972
rect -16072 -5548 -15300 -5520
rect -16072 -5972 -15384 -5548
rect -15320 -5972 -15300 -5548
rect -16072 -6000 -15300 -5972
rect -15060 -5548 -14288 -5520
rect -15060 -5972 -14372 -5548
rect -14308 -5972 -14288 -5548
rect -15060 -6000 -14288 -5972
rect -14048 -5548 -13276 -5520
rect -14048 -5972 -13360 -5548
rect -13296 -5972 -13276 -5548
rect -14048 -6000 -13276 -5972
rect -13036 -5548 -12264 -5520
rect -13036 -5972 -12348 -5548
rect -12284 -5972 -12264 -5548
rect -13036 -6000 -12264 -5972
rect -12024 -5548 -11252 -5520
rect -12024 -5972 -11336 -5548
rect -11272 -5972 -11252 -5548
rect -12024 -6000 -11252 -5972
rect -11012 -5548 -10240 -5520
rect -11012 -5972 -10324 -5548
rect -10260 -5972 -10240 -5548
rect -11012 -6000 -10240 -5972
rect -10000 -5548 -9228 -5520
rect -10000 -5972 -9312 -5548
rect -9248 -5972 -9228 -5548
rect -10000 -6000 -9228 -5972
rect -8988 -5548 -8216 -5520
rect -8988 -5972 -8300 -5548
rect -8236 -5972 -8216 -5548
rect -8988 -6000 -8216 -5972
rect -7976 -5548 -7204 -5520
rect -7976 -5972 -7288 -5548
rect -7224 -5972 -7204 -5548
rect -7976 -6000 -7204 -5972
rect -6964 -5548 -6192 -5520
rect -6964 -5972 -6276 -5548
rect -6212 -5972 -6192 -5548
rect -6964 -6000 -6192 -5972
rect -5952 -5548 -5180 -5520
rect -5952 -5972 -5264 -5548
rect -5200 -5972 -5180 -5548
rect -5952 -6000 -5180 -5972
rect -4940 -5548 -4168 -5520
rect -4940 -5972 -4252 -5548
rect -4188 -5972 -4168 -5548
rect -4940 -6000 -4168 -5972
rect -3928 -5548 -3156 -5520
rect -3928 -5972 -3240 -5548
rect -3176 -5972 -3156 -5548
rect -3928 -6000 -3156 -5972
rect -2916 -5548 -2144 -5520
rect -2916 -5972 -2228 -5548
rect -2164 -5972 -2144 -5548
rect -2916 -6000 -2144 -5972
rect -1904 -5548 -1132 -5520
rect -1904 -5972 -1216 -5548
rect -1152 -5972 -1132 -5548
rect -1904 -6000 -1132 -5972
rect -892 -5548 -120 -5520
rect -892 -5972 -204 -5548
rect -140 -5972 -120 -5548
rect -892 -6000 -120 -5972
rect 120 -5548 892 -5520
rect 120 -5972 808 -5548
rect 872 -5972 892 -5548
rect 120 -6000 892 -5972
rect 1132 -5548 1904 -5520
rect 1132 -5972 1820 -5548
rect 1884 -5972 1904 -5548
rect 1132 -6000 1904 -5972
rect 2144 -5548 2916 -5520
rect 2144 -5972 2832 -5548
rect 2896 -5972 2916 -5548
rect 2144 -6000 2916 -5972
rect 3156 -5548 3928 -5520
rect 3156 -5972 3844 -5548
rect 3908 -5972 3928 -5548
rect 3156 -6000 3928 -5972
rect 4168 -5548 4940 -5520
rect 4168 -5972 4856 -5548
rect 4920 -5972 4940 -5548
rect 4168 -6000 4940 -5972
rect 5180 -5548 5952 -5520
rect 5180 -5972 5868 -5548
rect 5932 -5972 5952 -5548
rect 5180 -6000 5952 -5972
rect 6192 -5548 6964 -5520
rect 6192 -5972 6880 -5548
rect 6944 -5972 6964 -5548
rect 6192 -6000 6964 -5972
rect 7204 -5548 7976 -5520
rect 7204 -5972 7892 -5548
rect 7956 -5972 7976 -5548
rect 7204 -6000 7976 -5972
rect 8216 -5548 8988 -5520
rect 8216 -5972 8904 -5548
rect 8968 -5972 8988 -5548
rect 8216 -6000 8988 -5972
rect 9228 -5548 10000 -5520
rect 9228 -5972 9916 -5548
rect 9980 -5972 10000 -5548
rect 9228 -6000 10000 -5972
rect 10240 -5548 11012 -5520
rect 10240 -5972 10928 -5548
rect 10992 -5972 11012 -5548
rect 10240 -6000 11012 -5972
rect 11252 -5548 12024 -5520
rect 11252 -5972 11940 -5548
rect 12004 -5972 12024 -5548
rect 11252 -6000 12024 -5972
rect 12264 -5548 13036 -5520
rect 12264 -5972 12952 -5548
rect 13016 -5972 13036 -5548
rect 12264 -6000 13036 -5972
rect 13276 -5548 14048 -5520
rect 13276 -5972 13964 -5548
rect 14028 -5972 14048 -5548
rect 13276 -6000 14048 -5972
rect 14288 -5548 15060 -5520
rect 14288 -5972 14976 -5548
rect 15040 -5972 15060 -5548
rect 14288 -6000 15060 -5972
rect 15300 -5548 16072 -5520
rect 15300 -5972 15988 -5548
rect 16052 -5972 16072 -5548
rect 15300 -6000 16072 -5972
rect 16312 -5548 17084 -5520
rect 16312 -5972 17000 -5548
rect 17064 -5972 17084 -5548
rect 16312 -6000 17084 -5972
rect -17084 -6268 -16312 -6240
rect -17084 -6692 -16396 -6268
rect -16332 -6692 -16312 -6268
rect -17084 -6720 -16312 -6692
rect -16072 -6268 -15300 -6240
rect -16072 -6692 -15384 -6268
rect -15320 -6692 -15300 -6268
rect -16072 -6720 -15300 -6692
rect -15060 -6268 -14288 -6240
rect -15060 -6692 -14372 -6268
rect -14308 -6692 -14288 -6268
rect -15060 -6720 -14288 -6692
rect -14048 -6268 -13276 -6240
rect -14048 -6692 -13360 -6268
rect -13296 -6692 -13276 -6268
rect -14048 -6720 -13276 -6692
rect -13036 -6268 -12264 -6240
rect -13036 -6692 -12348 -6268
rect -12284 -6692 -12264 -6268
rect -13036 -6720 -12264 -6692
rect -12024 -6268 -11252 -6240
rect -12024 -6692 -11336 -6268
rect -11272 -6692 -11252 -6268
rect -12024 -6720 -11252 -6692
rect -11012 -6268 -10240 -6240
rect -11012 -6692 -10324 -6268
rect -10260 -6692 -10240 -6268
rect -11012 -6720 -10240 -6692
rect -10000 -6268 -9228 -6240
rect -10000 -6692 -9312 -6268
rect -9248 -6692 -9228 -6268
rect -10000 -6720 -9228 -6692
rect -8988 -6268 -8216 -6240
rect -8988 -6692 -8300 -6268
rect -8236 -6692 -8216 -6268
rect -8988 -6720 -8216 -6692
rect -7976 -6268 -7204 -6240
rect -7976 -6692 -7288 -6268
rect -7224 -6692 -7204 -6268
rect -7976 -6720 -7204 -6692
rect -6964 -6268 -6192 -6240
rect -6964 -6692 -6276 -6268
rect -6212 -6692 -6192 -6268
rect -6964 -6720 -6192 -6692
rect -5952 -6268 -5180 -6240
rect -5952 -6692 -5264 -6268
rect -5200 -6692 -5180 -6268
rect -5952 -6720 -5180 -6692
rect -4940 -6268 -4168 -6240
rect -4940 -6692 -4252 -6268
rect -4188 -6692 -4168 -6268
rect -4940 -6720 -4168 -6692
rect -3928 -6268 -3156 -6240
rect -3928 -6692 -3240 -6268
rect -3176 -6692 -3156 -6268
rect -3928 -6720 -3156 -6692
rect -2916 -6268 -2144 -6240
rect -2916 -6692 -2228 -6268
rect -2164 -6692 -2144 -6268
rect -2916 -6720 -2144 -6692
rect -1904 -6268 -1132 -6240
rect -1904 -6692 -1216 -6268
rect -1152 -6692 -1132 -6268
rect -1904 -6720 -1132 -6692
rect -892 -6268 -120 -6240
rect -892 -6692 -204 -6268
rect -140 -6692 -120 -6268
rect -892 -6720 -120 -6692
rect 120 -6268 892 -6240
rect 120 -6692 808 -6268
rect 872 -6692 892 -6268
rect 120 -6720 892 -6692
rect 1132 -6268 1904 -6240
rect 1132 -6692 1820 -6268
rect 1884 -6692 1904 -6268
rect 1132 -6720 1904 -6692
rect 2144 -6268 2916 -6240
rect 2144 -6692 2832 -6268
rect 2896 -6692 2916 -6268
rect 2144 -6720 2916 -6692
rect 3156 -6268 3928 -6240
rect 3156 -6692 3844 -6268
rect 3908 -6692 3928 -6268
rect 3156 -6720 3928 -6692
rect 4168 -6268 4940 -6240
rect 4168 -6692 4856 -6268
rect 4920 -6692 4940 -6268
rect 4168 -6720 4940 -6692
rect 5180 -6268 5952 -6240
rect 5180 -6692 5868 -6268
rect 5932 -6692 5952 -6268
rect 5180 -6720 5952 -6692
rect 6192 -6268 6964 -6240
rect 6192 -6692 6880 -6268
rect 6944 -6692 6964 -6268
rect 6192 -6720 6964 -6692
rect 7204 -6268 7976 -6240
rect 7204 -6692 7892 -6268
rect 7956 -6692 7976 -6268
rect 7204 -6720 7976 -6692
rect 8216 -6268 8988 -6240
rect 8216 -6692 8904 -6268
rect 8968 -6692 8988 -6268
rect 8216 -6720 8988 -6692
rect 9228 -6268 10000 -6240
rect 9228 -6692 9916 -6268
rect 9980 -6692 10000 -6268
rect 9228 -6720 10000 -6692
rect 10240 -6268 11012 -6240
rect 10240 -6692 10928 -6268
rect 10992 -6692 11012 -6268
rect 10240 -6720 11012 -6692
rect 11252 -6268 12024 -6240
rect 11252 -6692 11940 -6268
rect 12004 -6692 12024 -6268
rect 11252 -6720 12024 -6692
rect 12264 -6268 13036 -6240
rect 12264 -6692 12952 -6268
rect 13016 -6692 13036 -6268
rect 12264 -6720 13036 -6692
rect 13276 -6268 14048 -6240
rect 13276 -6692 13964 -6268
rect 14028 -6692 14048 -6268
rect 13276 -6720 14048 -6692
rect 14288 -6268 15060 -6240
rect 14288 -6692 14976 -6268
rect 15040 -6692 15060 -6268
rect 14288 -6720 15060 -6692
rect 15300 -6268 16072 -6240
rect 15300 -6692 15988 -6268
rect 16052 -6692 16072 -6268
rect 15300 -6720 16072 -6692
rect 16312 -6268 17084 -6240
rect 16312 -6692 17000 -6268
rect 17064 -6692 17084 -6268
rect 16312 -6720 17084 -6692
rect -17084 -6988 -16312 -6960
rect -17084 -7412 -16396 -6988
rect -16332 -7412 -16312 -6988
rect -17084 -7440 -16312 -7412
rect -16072 -6988 -15300 -6960
rect -16072 -7412 -15384 -6988
rect -15320 -7412 -15300 -6988
rect -16072 -7440 -15300 -7412
rect -15060 -6988 -14288 -6960
rect -15060 -7412 -14372 -6988
rect -14308 -7412 -14288 -6988
rect -15060 -7440 -14288 -7412
rect -14048 -6988 -13276 -6960
rect -14048 -7412 -13360 -6988
rect -13296 -7412 -13276 -6988
rect -14048 -7440 -13276 -7412
rect -13036 -6988 -12264 -6960
rect -13036 -7412 -12348 -6988
rect -12284 -7412 -12264 -6988
rect -13036 -7440 -12264 -7412
rect -12024 -6988 -11252 -6960
rect -12024 -7412 -11336 -6988
rect -11272 -7412 -11252 -6988
rect -12024 -7440 -11252 -7412
rect -11012 -6988 -10240 -6960
rect -11012 -7412 -10324 -6988
rect -10260 -7412 -10240 -6988
rect -11012 -7440 -10240 -7412
rect -10000 -6988 -9228 -6960
rect -10000 -7412 -9312 -6988
rect -9248 -7412 -9228 -6988
rect -10000 -7440 -9228 -7412
rect -8988 -6988 -8216 -6960
rect -8988 -7412 -8300 -6988
rect -8236 -7412 -8216 -6988
rect -8988 -7440 -8216 -7412
rect -7976 -6988 -7204 -6960
rect -7976 -7412 -7288 -6988
rect -7224 -7412 -7204 -6988
rect -7976 -7440 -7204 -7412
rect -6964 -6988 -6192 -6960
rect -6964 -7412 -6276 -6988
rect -6212 -7412 -6192 -6988
rect -6964 -7440 -6192 -7412
rect -5952 -6988 -5180 -6960
rect -5952 -7412 -5264 -6988
rect -5200 -7412 -5180 -6988
rect -5952 -7440 -5180 -7412
rect -4940 -6988 -4168 -6960
rect -4940 -7412 -4252 -6988
rect -4188 -7412 -4168 -6988
rect -4940 -7440 -4168 -7412
rect -3928 -6988 -3156 -6960
rect -3928 -7412 -3240 -6988
rect -3176 -7412 -3156 -6988
rect -3928 -7440 -3156 -7412
rect -2916 -6988 -2144 -6960
rect -2916 -7412 -2228 -6988
rect -2164 -7412 -2144 -6988
rect -2916 -7440 -2144 -7412
rect -1904 -6988 -1132 -6960
rect -1904 -7412 -1216 -6988
rect -1152 -7412 -1132 -6988
rect -1904 -7440 -1132 -7412
rect -892 -6988 -120 -6960
rect -892 -7412 -204 -6988
rect -140 -7412 -120 -6988
rect -892 -7440 -120 -7412
rect 120 -6988 892 -6960
rect 120 -7412 808 -6988
rect 872 -7412 892 -6988
rect 120 -7440 892 -7412
rect 1132 -6988 1904 -6960
rect 1132 -7412 1820 -6988
rect 1884 -7412 1904 -6988
rect 1132 -7440 1904 -7412
rect 2144 -6988 2916 -6960
rect 2144 -7412 2832 -6988
rect 2896 -7412 2916 -6988
rect 2144 -7440 2916 -7412
rect 3156 -6988 3928 -6960
rect 3156 -7412 3844 -6988
rect 3908 -7412 3928 -6988
rect 3156 -7440 3928 -7412
rect 4168 -6988 4940 -6960
rect 4168 -7412 4856 -6988
rect 4920 -7412 4940 -6988
rect 4168 -7440 4940 -7412
rect 5180 -6988 5952 -6960
rect 5180 -7412 5868 -6988
rect 5932 -7412 5952 -6988
rect 5180 -7440 5952 -7412
rect 6192 -6988 6964 -6960
rect 6192 -7412 6880 -6988
rect 6944 -7412 6964 -6988
rect 6192 -7440 6964 -7412
rect 7204 -6988 7976 -6960
rect 7204 -7412 7892 -6988
rect 7956 -7412 7976 -6988
rect 7204 -7440 7976 -7412
rect 8216 -6988 8988 -6960
rect 8216 -7412 8904 -6988
rect 8968 -7412 8988 -6988
rect 8216 -7440 8988 -7412
rect 9228 -6988 10000 -6960
rect 9228 -7412 9916 -6988
rect 9980 -7412 10000 -6988
rect 9228 -7440 10000 -7412
rect 10240 -6988 11012 -6960
rect 10240 -7412 10928 -6988
rect 10992 -7412 11012 -6988
rect 10240 -7440 11012 -7412
rect 11252 -6988 12024 -6960
rect 11252 -7412 11940 -6988
rect 12004 -7412 12024 -6988
rect 11252 -7440 12024 -7412
rect 12264 -6988 13036 -6960
rect 12264 -7412 12952 -6988
rect 13016 -7412 13036 -6988
rect 12264 -7440 13036 -7412
rect 13276 -6988 14048 -6960
rect 13276 -7412 13964 -6988
rect 14028 -7412 14048 -6988
rect 13276 -7440 14048 -7412
rect 14288 -6988 15060 -6960
rect 14288 -7412 14976 -6988
rect 15040 -7412 15060 -6988
rect 14288 -7440 15060 -7412
rect 15300 -6988 16072 -6960
rect 15300 -7412 15988 -6988
rect 16052 -7412 16072 -6988
rect 15300 -7440 16072 -7412
rect 16312 -6988 17084 -6960
rect 16312 -7412 17000 -6988
rect 17064 -7412 17084 -6988
rect 16312 -7440 17084 -7412
rect -17084 -7708 -16312 -7680
rect -17084 -8132 -16396 -7708
rect -16332 -8132 -16312 -7708
rect -17084 -8160 -16312 -8132
rect -16072 -7708 -15300 -7680
rect -16072 -8132 -15384 -7708
rect -15320 -8132 -15300 -7708
rect -16072 -8160 -15300 -8132
rect -15060 -7708 -14288 -7680
rect -15060 -8132 -14372 -7708
rect -14308 -8132 -14288 -7708
rect -15060 -8160 -14288 -8132
rect -14048 -7708 -13276 -7680
rect -14048 -8132 -13360 -7708
rect -13296 -8132 -13276 -7708
rect -14048 -8160 -13276 -8132
rect -13036 -7708 -12264 -7680
rect -13036 -8132 -12348 -7708
rect -12284 -8132 -12264 -7708
rect -13036 -8160 -12264 -8132
rect -12024 -7708 -11252 -7680
rect -12024 -8132 -11336 -7708
rect -11272 -8132 -11252 -7708
rect -12024 -8160 -11252 -8132
rect -11012 -7708 -10240 -7680
rect -11012 -8132 -10324 -7708
rect -10260 -8132 -10240 -7708
rect -11012 -8160 -10240 -8132
rect -10000 -7708 -9228 -7680
rect -10000 -8132 -9312 -7708
rect -9248 -8132 -9228 -7708
rect -10000 -8160 -9228 -8132
rect -8988 -7708 -8216 -7680
rect -8988 -8132 -8300 -7708
rect -8236 -8132 -8216 -7708
rect -8988 -8160 -8216 -8132
rect -7976 -7708 -7204 -7680
rect -7976 -8132 -7288 -7708
rect -7224 -8132 -7204 -7708
rect -7976 -8160 -7204 -8132
rect -6964 -7708 -6192 -7680
rect -6964 -8132 -6276 -7708
rect -6212 -8132 -6192 -7708
rect -6964 -8160 -6192 -8132
rect -5952 -7708 -5180 -7680
rect -5952 -8132 -5264 -7708
rect -5200 -8132 -5180 -7708
rect -5952 -8160 -5180 -8132
rect -4940 -7708 -4168 -7680
rect -4940 -8132 -4252 -7708
rect -4188 -8132 -4168 -7708
rect -4940 -8160 -4168 -8132
rect -3928 -7708 -3156 -7680
rect -3928 -8132 -3240 -7708
rect -3176 -8132 -3156 -7708
rect -3928 -8160 -3156 -8132
rect -2916 -7708 -2144 -7680
rect -2916 -8132 -2228 -7708
rect -2164 -8132 -2144 -7708
rect -2916 -8160 -2144 -8132
rect -1904 -7708 -1132 -7680
rect -1904 -8132 -1216 -7708
rect -1152 -8132 -1132 -7708
rect -1904 -8160 -1132 -8132
rect -892 -7708 -120 -7680
rect -892 -8132 -204 -7708
rect -140 -8132 -120 -7708
rect -892 -8160 -120 -8132
rect 120 -7708 892 -7680
rect 120 -8132 808 -7708
rect 872 -8132 892 -7708
rect 120 -8160 892 -8132
rect 1132 -7708 1904 -7680
rect 1132 -8132 1820 -7708
rect 1884 -8132 1904 -7708
rect 1132 -8160 1904 -8132
rect 2144 -7708 2916 -7680
rect 2144 -8132 2832 -7708
rect 2896 -8132 2916 -7708
rect 2144 -8160 2916 -8132
rect 3156 -7708 3928 -7680
rect 3156 -8132 3844 -7708
rect 3908 -8132 3928 -7708
rect 3156 -8160 3928 -8132
rect 4168 -7708 4940 -7680
rect 4168 -8132 4856 -7708
rect 4920 -8132 4940 -7708
rect 4168 -8160 4940 -8132
rect 5180 -7708 5952 -7680
rect 5180 -8132 5868 -7708
rect 5932 -8132 5952 -7708
rect 5180 -8160 5952 -8132
rect 6192 -7708 6964 -7680
rect 6192 -8132 6880 -7708
rect 6944 -8132 6964 -7708
rect 6192 -8160 6964 -8132
rect 7204 -7708 7976 -7680
rect 7204 -8132 7892 -7708
rect 7956 -8132 7976 -7708
rect 7204 -8160 7976 -8132
rect 8216 -7708 8988 -7680
rect 8216 -8132 8904 -7708
rect 8968 -8132 8988 -7708
rect 8216 -8160 8988 -8132
rect 9228 -7708 10000 -7680
rect 9228 -8132 9916 -7708
rect 9980 -8132 10000 -7708
rect 9228 -8160 10000 -8132
rect 10240 -7708 11012 -7680
rect 10240 -8132 10928 -7708
rect 10992 -8132 11012 -7708
rect 10240 -8160 11012 -8132
rect 11252 -7708 12024 -7680
rect 11252 -8132 11940 -7708
rect 12004 -8132 12024 -7708
rect 11252 -8160 12024 -8132
rect 12264 -7708 13036 -7680
rect 12264 -8132 12952 -7708
rect 13016 -8132 13036 -7708
rect 12264 -8160 13036 -8132
rect 13276 -7708 14048 -7680
rect 13276 -8132 13964 -7708
rect 14028 -8132 14048 -7708
rect 13276 -8160 14048 -8132
rect 14288 -7708 15060 -7680
rect 14288 -8132 14976 -7708
rect 15040 -8132 15060 -7708
rect 14288 -8160 15060 -8132
rect 15300 -7708 16072 -7680
rect 15300 -8132 15988 -7708
rect 16052 -8132 16072 -7708
rect 15300 -8160 16072 -8132
rect 16312 -7708 17084 -7680
rect 16312 -8132 17000 -7708
rect 17064 -8132 17084 -7708
rect 16312 -8160 17084 -8132
rect -17084 -8428 -16312 -8400
rect -17084 -8852 -16396 -8428
rect -16332 -8852 -16312 -8428
rect -17084 -8880 -16312 -8852
rect -16072 -8428 -15300 -8400
rect -16072 -8852 -15384 -8428
rect -15320 -8852 -15300 -8428
rect -16072 -8880 -15300 -8852
rect -15060 -8428 -14288 -8400
rect -15060 -8852 -14372 -8428
rect -14308 -8852 -14288 -8428
rect -15060 -8880 -14288 -8852
rect -14048 -8428 -13276 -8400
rect -14048 -8852 -13360 -8428
rect -13296 -8852 -13276 -8428
rect -14048 -8880 -13276 -8852
rect -13036 -8428 -12264 -8400
rect -13036 -8852 -12348 -8428
rect -12284 -8852 -12264 -8428
rect -13036 -8880 -12264 -8852
rect -12024 -8428 -11252 -8400
rect -12024 -8852 -11336 -8428
rect -11272 -8852 -11252 -8428
rect -12024 -8880 -11252 -8852
rect -11012 -8428 -10240 -8400
rect -11012 -8852 -10324 -8428
rect -10260 -8852 -10240 -8428
rect -11012 -8880 -10240 -8852
rect -10000 -8428 -9228 -8400
rect -10000 -8852 -9312 -8428
rect -9248 -8852 -9228 -8428
rect -10000 -8880 -9228 -8852
rect -8988 -8428 -8216 -8400
rect -8988 -8852 -8300 -8428
rect -8236 -8852 -8216 -8428
rect -8988 -8880 -8216 -8852
rect -7976 -8428 -7204 -8400
rect -7976 -8852 -7288 -8428
rect -7224 -8852 -7204 -8428
rect -7976 -8880 -7204 -8852
rect -6964 -8428 -6192 -8400
rect -6964 -8852 -6276 -8428
rect -6212 -8852 -6192 -8428
rect -6964 -8880 -6192 -8852
rect -5952 -8428 -5180 -8400
rect -5952 -8852 -5264 -8428
rect -5200 -8852 -5180 -8428
rect -5952 -8880 -5180 -8852
rect -4940 -8428 -4168 -8400
rect -4940 -8852 -4252 -8428
rect -4188 -8852 -4168 -8428
rect -4940 -8880 -4168 -8852
rect -3928 -8428 -3156 -8400
rect -3928 -8852 -3240 -8428
rect -3176 -8852 -3156 -8428
rect -3928 -8880 -3156 -8852
rect -2916 -8428 -2144 -8400
rect -2916 -8852 -2228 -8428
rect -2164 -8852 -2144 -8428
rect -2916 -8880 -2144 -8852
rect -1904 -8428 -1132 -8400
rect -1904 -8852 -1216 -8428
rect -1152 -8852 -1132 -8428
rect -1904 -8880 -1132 -8852
rect -892 -8428 -120 -8400
rect -892 -8852 -204 -8428
rect -140 -8852 -120 -8428
rect -892 -8880 -120 -8852
rect 120 -8428 892 -8400
rect 120 -8852 808 -8428
rect 872 -8852 892 -8428
rect 120 -8880 892 -8852
rect 1132 -8428 1904 -8400
rect 1132 -8852 1820 -8428
rect 1884 -8852 1904 -8428
rect 1132 -8880 1904 -8852
rect 2144 -8428 2916 -8400
rect 2144 -8852 2832 -8428
rect 2896 -8852 2916 -8428
rect 2144 -8880 2916 -8852
rect 3156 -8428 3928 -8400
rect 3156 -8852 3844 -8428
rect 3908 -8852 3928 -8428
rect 3156 -8880 3928 -8852
rect 4168 -8428 4940 -8400
rect 4168 -8852 4856 -8428
rect 4920 -8852 4940 -8428
rect 4168 -8880 4940 -8852
rect 5180 -8428 5952 -8400
rect 5180 -8852 5868 -8428
rect 5932 -8852 5952 -8428
rect 5180 -8880 5952 -8852
rect 6192 -8428 6964 -8400
rect 6192 -8852 6880 -8428
rect 6944 -8852 6964 -8428
rect 6192 -8880 6964 -8852
rect 7204 -8428 7976 -8400
rect 7204 -8852 7892 -8428
rect 7956 -8852 7976 -8428
rect 7204 -8880 7976 -8852
rect 8216 -8428 8988 -8400
rect 8216 -8852 8904 -8428
rect 8968 -8852 8988 -8428
rect 8216 -8880 8988 -8852
rect 9228 -8428 10000 -8400
rect 9228 -8852 9916 -8428
rect 9980 -8852 10000 -8428
rect 9228 -8880 10000 -8852
rect 10240 -8428 11012 -8400
rect 10240 -8852 10928 -8428
rect 10992 -8852 11012 -8428
rect 10240 -8880 11012 -8852
rect 11252 -8428 12024 -8400
rect 11252 -8852 11940 -8428
rect 12004 -8852 12024 -8428
rect 11252 -8880 12024 -8852
rect 12264 -8428 13036 -8400
rect 12264 -8852 12952 -8428
rect 13016 -8852 13036 -8428
rect 12264 -8880 13036 -8852
rect 13276 -8428 14048 -8400
rect 13276 -8852 13964 -8428
rect 14028 -8852 14048 -8428
rect 13276 -8880 14048 -8852
rect 14288 -8428 15060 -8400
rect 14288 -8852 14976 -8428
rect 15040 -8852 15060 -8428
rect 14288 -8880 15060 -8852
rect 15300 -8428 16072 -8400
rect 15300 -8852 15988 -8428
rect 16052 -8852 16072 -8428
rect 15300 -8880 16072 -8852
rect 16312 -8428 17084 -8400
rect 16312 -8852 17000 -8428
rect 17064 -8852 17084 -8428
rect 16312 -8880 17084 -8852
rect -17084 -9148 -16312 -9120
rect -17084 -9572 -16396 -9148
rect -16332 -9572 -16312 -9148
rect -17084 -9600 -16312 -9572
rect -16072 -9148 -15300 -9120
rect -16072 -9572 -15384 -9148
rect -15320 -9572 -15300 -9148
rect -16072 -9600 -15300 -9572
rect -15060 -9148 -14288 -9120
rect -15060 -9572 -14372 -9148
rect -14308 -9572 -14288 -9148
rect -15060 -9600 -14288 -9572
rect -14048 -9148 -13276 -9120
rect -14048 -9572 -13360 -9148
rect -13296 -9572 -13276 -9148
rect -14048 -9600 -13276 -9572
rect -13036 -9148 -12264 -9120
rect -13036 -9572 -12348 -9148
rect -12284 -9572 -12264 -9148
rect -13036 -9600 -12264 -9572
rect -12024 -9148 -11252 -9120
rect -12024 -9572 -11336 -9148
rect -11272 -9572 -11252 -9148
rect -12024 -9600 -11252 -9572
rect -11012 -9148 -10240 -9120
rect -11012 -9572 -10324 -9148
rect -10260 -9572 -10240 -9148
rect -11012 -9600 -10240 -9572
rect -10000 -9148 -9228 -9120
rect -10000 -9572 -9312 -9148
rect -9248 -9572 -9228 -9148
rect -10000 -9600 -9228 -9572
rect -8988 -9148 -8216 -9120
rect -8988 -9572 -8300 -9148
rect -8236 -9572 -8216 -9148
rect -8988 -9600 -8216 -9572
rect -7976 -9148 -7204 -9120
rect -7976 -9572 -7288 -9148
rect -7224 -9572 -7204 -9148
rect -7976 -9600 -7204 -9572
rect -6964 -9148 -6192 -9120
rect -6964 -9572 -6276 -9148
rect -6212 -9572 -6192 -9148
rect -6964 -9600 -6192 -9572
rect -5952 -9148 -5180 -9120
rect -5952 -9572 -5264 -9148
rect -5200 -9572 -5180 -9148
rect -5952 -9600 -5180 -9572
rect -4940 -9148 -4168 -9120
rect -4940 -9572 -4252 -9148
rect -4188 -9572 -4168 -9148
rect -4940 -9600 -4168 -9572
rect -3928 -9148 -3156 -9120
rect -3928 -9572 -3240 -9148
rect -3176 -9572 -3156 -9148
rect -3928 -9600 -3156 -9572
rect -2916 -9148 -2144 -9120
rect -2916 -9572 -2228 -9148
rect -2164 -9572 -2144 -9148
rect -2916 -9600 -2144 -9572
rect -1904 -9148 -1132 -9120
rect -1904 -9572 -1216 -9148
rect -1152 -9572 -1132 -9148
rect -1904 -9600 -1132 -9572
rect -892 -9148 -120 -9120
rect -892 -9572 -204 -9148
rect -140 -9572 -120 -9148
rect -892 -9600 -120 -9572
rect 120 -9148 892 -9120
rect 120 -9572 808 -9148
rect 872 -9572 892 -9148
rect 120 -9600 892 -9572
rect 1132 -9148 1904 -9120
rect 1132 -9572 1820 -9148
rect 1884 -9572 1904 -9148
rect 1132 -9600 1904 -9572
rect 2144 -9148 2916 -9120
rect 2144 -9572 2832 -9148
rect 2896 -9572 2916 -9148
rect 2144 -9600 2916 -9572
rect 3156 -9148 3928 -9120
rect 3156 -9572 3844 -9148
rect 3908 -9572 3928 -9148
rect 3156 -9600 3928 -9572
rect 4168 -9148 4940 -9120
rect 4168 -9572 4856 -9148
rect 4920 -9572 4940 -9148
rect 4168 -9600 4940 -9572
rect 5180 -9148 5952 -9120
rect 5180 -9572 5868 -9148
rect 5932 -9572 5952 -9148
rect 5180 -9600 5952 -9572
rect 6192 -9148 6964 -9120
rect 6192 -9572 6880 -9148
rect 6944 -9572 6964 -9148
rect 6192 -9600 6964 -9572
rect 7204 -9148 7976 -9120
rect 7204 -9572 7892 -9148
rect 7956 -9572 7976 -9148
rect 7204 -9600 7976 -9572
rect 8216 -9148 8988 -9120
rect 8216 -9572 8904 -9148
rect 8968 -9572 8988 -9148
rect 8216 -9600 8988 -9572
rect 9228 -9148 10000 -9120
rect 9228 -9572 9916 -9148
rect 9980 -9572 10000 -9148
rect 9228 -9600 10000 -9572
rect 10240 -9148 11012 -9120
rect 10240 -9572 10928 -9148
rect 10992 -9572 11012 -9148
rect 10240 -9600 11012 -9572
rect 11252 -9148 12024 -9120
rect 11252 -9572 11940 -9148
rect 12004 -9572 12024 -9148
rect 11252 -9600 12024 -9572
rect 12264 -9148 13036 -9120
rect 12264 -9572 12952 -9148
rect 13016 -9572 13036 -9148
rect 12264 -9600 13036 -9572
rect 13276 -9148 14048 -9120
rect 13276 -9572 13964 -9148
rect 14028 -9572 14048 -9148
rect 13276 -9600 14048 -9572
rect 14288 -9148 15060 -9120
rect 14288 -9572 14976 -9148
rect 15040 -9572 15060 -9148
rect 14288 -9600 15060 -9572
rect 15300 -9148 16072 -9120
rect 15300 -9572 15988 -9148
rect 16052 -9572 16072 -9148
rect 15300 -9600 16072 -9572
rect 16312 -9148 17084 -9120
rect 16312 -9572 17000 -9148
rect 17064 -9572 17084 -9148
rect 16312 -9600 17084 -9572
rect -17084 -9868 -16312 -9840
rect -17084 -10292 -16396 -9868
rect -16332 -10292 -16312 -9868
rect -17084 -10320 -16312 -10292
rect -16072 -9868 -15300 -9840
rect -16072 -10292 -15384 -9868
rect -15320 -10292 -15300 -9868
rect -16072 -10320 -15300 -10292
rect -15060 -9868 -14288 -9840
rect -15060 -10292 -14372 -9868
rect -14308 -10292 -14288 -9868
rect -15060 -10320 -14288 -10292
rect -14048 -9868 -13276 -9840
rect -14048 -10292 -13360 -9868
rect -13296 -10292 -13276 -9868
rect -14048 -10320 -13276 -10292
rect -13036 -9868 -12264 -9840
rect -13036 -10292 -12348 -9868
rect -12284 -10292 -12264 -9868
rect -13036 -10320 -12264 -10292
rect -12024 -9868 -11252 -9840
rect -12024 -10292 -11336 -9868
rect -11272 -10292 -11252 -9868
rect -12024 -10320 -11252 -10292
rect -11012 -9868 -10240 -9840
rect -11012 -10292 -10324 -9868
rect -10260 -10292 -10240 -9868
rect -11012 -10320 -10240 -10292
rect -10000 -9868 -9228 -9840
rect -10000 -10292 -9312 -9868
rect -9248 -10292 -9228 -9868
rect -10000 -10320 -9228 -10292
rect -8988 -9868 -8216 -9840
rect -8988 -10292 -8300 -9868
rect -8236 -10292 -8216 -9868
rect -8988 -10320 -8216 -10292
rect -7976 -9868 -7204 -9840
rect -7976 -10292 -7288 -9868
rect -7224 -10292 -7204 -9868
rect -7976 -10320 -7204 -10292
rect -6964 -9868 -6192 -9840
rect -6964 -10292 -6276 -9868
rect -6212 -10292 -6192 -9868
rect -6964 -10320 -6192 -10292
rect -5952 -9868 -5180 -9840
rect -5952 -10292 -5264 -9868
rect -5200 -10292 -5180 -9868
rect -5952 -10320 -5180 -10292
rect -4940 -9868 -4168 -9840
rect -4940 -10292 -4252 -9868
rect -4188 -10292 -4168 -9868
rect -4940 -10320 -4168 -10292
rect -3928 -9868 -3156 -9840
rect -3928 -10292 -3240 -9868
rect -3176 -10292 -3156 -9868
rect -3928 -10320 -3156 -10292
rect -2916 -9868 -2144 -9840
rect -2916 -10292 -2228 -9868
rect -2164 -10292 -2144 -9868
rect -2916 -10320 -2144 -10292
rect -1904 -9868 -1132 -9840
rect -1904 -10292 -1216 -9868
rect -1152 -10292 -1132 -9868
rect -1904 -10320 -1132 -10292
rect -892 -9868 -120 -9840
rect -892 -10292 -204 -9868
rect -140 -10292 -120 -9868
rect -892 -10320 -120 -10292
rect 120 -9868 892 -9840
rect 120 -10292 808 -9868
rect 872 -10292 892 -9868
rect 120 -10320 892 -10292
rect 1132 -9868 1904 -9840
rect 1132 -10292 1820 -9868
rect 1884 -10292 1904 -9868
rect 1132 -10320 1904 -10292
rect 2144 -9868 2916 -9840
rect 2144 -10292 2832 -9868
rect 2896 -10292 2916 -9868
rect 2144 -10320 2916 -10292
rect 3156 -9868 3928 -9840
rect 3156 -10292 3844 -9868
rect 3908 -10292 3928 -9868
rect 3156 -10320 3928 -10292
rect 4168 -9868 4940 -9840
rect 4168 -10292 4856 -9868
rect 4920 -10292 4940 -9868
rect 4168 -10320 4940 -10292
rect 5180 -9868 5952 -9840
rect 5180 -10292 5868 -9868
rect 5932 -10292 5952 -9868
rect 5180 -10320 5952 -10292
rect 6192 -9868 6964 -9840
rect 6192 -10292 6880 -9868
rect 6944 -10292 6964 -9868
rect 6192 -10320 6964 -10292
rect 7204 -9868 7976 -9840
rect 7204 -10292 7892 -9868
rect 7956 -10292 7976 -9868
rect 7204 -10320 7976 -10292
rect 8216 -9868 8988 -9840
rect 8216 -10292 8904 -9868
rect 8968 -10292 8988 -9868
rect 8216 -10320 8988 -10292
rect 9228 -9868 10000 -9840
rect 9228 -10292 9916 -9868
rect 9980 -10292 10000 -9868
rect 9228 -10320 10000 -10292
rect 10240 -9868 11012 -9840
rect 10240 -10292 10928 -9868
rect 10992 -10292 11012 -9868
rect 10240 -10320 11012 -10292
rect 11252 -9868 12024 -9840
rect 11252 -10292 11940 -9868
rect 12004 -10292 12024 -9868
rect 11252 -10320 12024 -10292
rect 12264 -9868 13036 -9840
rect 12264 -10292 12952 -9868
rect 13016 -10292 13036 -9868
rect 12264 -10320 13036 -10292
rect 13276 -9868 14048 -9840
rect 13276 -10292 13964 -9868
rect 14028 -10292 14048 -9868
rect 13276 -10320 14048 -10292
rect 14288 -9868 15060 -9840
rect 14288 -10292 14976 -9868
rect 15040 -10292 15060 -9868
rect 14288 -10320 15060 -10292
rect 15300 -9868 16072 -9840
rect 15300 -10292 15988 -9868
rect 16052 -10292 16072 -9868
rect 15300 -10320 16072 -10292
rect 16312 -9868 17084 -9840
rect 16312 -10292 17000 -9868
rect 17064 -10292 17084 -9868
rect 16312 -10320 17084 -10292
rect -17084 -10588 -16312 -10560
rect -17084 -11012 -16396 -10588
rect -16332 -11012 -16312 -10588
rect -17084 -11040 -16312 -11012
rect -16072 -10588 -15300 -10560
rect -16072 -11012 -15384 -10588
rect -15320 -11012 -15300 -10588
rect -16072 -11040 -15300 -11012
rect -15060 -10588 -14288 -10560
rect -15060 -11012 -14372 -10588
rect -14308 -11012 -14288 -10588
rect -15060 -11040 -14288 -11012
rect -14048 -10588 -13276 -10560
rect -14048 -11012 -13360 -10588
rect -13296 -11012 -13276 -10588
rect -14048 -11040 -13276 -11012
rect -13036 -10588 -12264 -10560
rect -13036 -11012 -12348 -10588
rect -12284 -11012 -12264 -10588
rect -13036 -11040 -12264 -11012
rect -12024 -10588 -11252 -10560
rect -12024 -11012 -11336 -10588
rect -11272 -11012 -11252 -10588
rect -12024 -11040 -11252 -11012
rect -11012 -10588 -10240 -10560
rect -11012 -11012 -10324 -10588
rect -10260 -11012 -10240 -10588
rect -11012 -11040 -10240 -11012
rect -10000 -10588 -9228 -10560
rect -10000 -11012 -9312 -10588
rect -9248 -11012 -9228 -10588
rect -10000 -11040 -9228 -11012
rect -8988 -10588 -8216 -10560
rect -8988 -11012 -8300 -10588
rect -8236 -11012 -8216 -10588
rect -8988 -11040 -8216 -11012
rect -7976 -10588 -7204 -10560
rect -7976 -11012 -7288 -10588
rect -7224 -11012 -7204 -10588
rect -7976 -11040 -7204 -11012
rect -6964 -10588 -6192 -10560
rect -6964 -11012 -6276 -10588
rect -6212 -11012 -6192 -10588
rect -6964 -11040 -6192 -11012
rect -5952 -10588 -5180 -10560
rect -5952 -11012 -5264 -10588
rect -5200 -11012 -5180 -10588
rect -5952 -11040 -5180 -11012
rect -4940 -10588 -4168 -10560
rect -4940 -11012 -4252 -10588
rect -4188 -11012 -4168 -10588
rect -4940 -11040 -4168 -11012
rect -3928 -10588 -3156 -10560
rect -3928 -11012 -3240 -10588
rect -3176 -11012 -3156 -10588
rect -3928 -11040 -3156 -11012
rect -2916 -10588 -2144 -10560
rect -2916 -11012 -2228 -10588
rect -2164 -11012 -2144 -10588
rect -2916 -11040 -2144 -11012
rect -1904 -10588 -1132 -10560
rect -1904 -11012 -1216 -10588
rect -1152 -11012 -1132 -10588
rect -1904 -11040 -1132 -11012
rect -892 -10588 -120 -10560
rect -892 -11012 -204 -10588
rect -140 -11012 -120 -10588
rect -892 -11040 -120 -11012
rect 120 -10588 892 -10560
rect 120 -11012 808 -10588
rect 872 -11012 892 -10588
rect 120 -11040 892 -11012
rect 1132 -10588 1904 -10560
rect 1132 -11012 1820 -10588
rect 1884 -11012 1904 -10588
rect 1132 -11040 1904 -11012
rect 2144 -10588 2916 -10560
rect 2144 -11012 2832 -10588
rect 2896 -11012 2916 -10588
rect 2144 -11040 2916 -11012
rect 3156 -10588 3928 -10560
rect 3156 -11012 3844 -10588
rect 3908 -11012 3928 -10588
rect 3156 -11040 3928 -11012
rect 4168 -10588 4940 -10560
rect 4168 -11012 4856 -10588
rect 4920 -11012 4940 -10588
rect 4168 -11040 4940 -11012
rect 5180 -10588 5952 -10560
rect 5180 -11012 5868 -10588
rect 5932 -11012 5952 -10588
rect 5180 -11040 5952 -11012
rect 6192 -10588 6964 -10560
rect 6192 -11012 6880 -10588
rect 6944 -11012 6964 -10588
rect 6192 -11040 6964 -11012
rect 7204 -10588 7976 -10560
rect 7204 -11012 7892 -10588
rect 7956 -11012 7976 -10588
rect 7204 -11040 7976 -11012
rect 8216 -10588 8988 -10560
rect 8216 -11012 8904 -10588
rect 8968 -11012 8988 -10588
rect 8216 -11040 8988 -11012
rect 9228 -10588 10000 -10560
rect 9228 -11012 9916 -10588
rect 9980 -11012 10000 -10588
rect 9228 -11040 10000 -11012
rect 10240 -10588 11012 -10560
rect 10240 -11012 10928 -10588
rect 10992 -11012 11012 -10588
rect 10240 -11040 11012 -11012
rect 11252 -10588 12024 -10560
rect 11252 -11012 11940 -10588
rect 12004 -11012 12024 -10588
rect 11252 -11040 12024 -11012
rect 12264 -10588 13036 -10560
rect 12264 -11012 12952 -10588
rect 13016 -11012 13036 -10588
rect 12264 -11040 13036 -11012
rect 13276 -10588 14048 -10560
rect 13276 -11012 13964 -10588
rect 14028 -11012 14048 -10588
rect 13276 -11040 14048 -11012
rect 14288 -10588 15060 -10560
rect 14288 -11012 14976 -10588
rect 15040 -11012 15060 -10588
rect 14288 -11040 15060 -11012
rect 15300 -10588 16072 -10560
rect 15300 -11012 15988 -10588
rect 16052 -11012 16072 -10588
rect 15300 -11040 16072 -11012
rect 16312 -10588 17084 -10560
rect 16312 -11012 17000 -10588
rect 17064 -11012 17084 -10588
rect 16312 -11040 17084 -11012
rect -17084 -11308 -16312 -11280
rect -17084 -11732 -16396 -11308
rect -16332 -11732 -16312 -11308
rect -17084 -11760 -16312 -11732
rect -16072 -11308 -15300 -11280
rect -16072 -11732 -15384 -11308
rect -15320 -11732 -15300 -11308
rect -16072 -11760 -15300 -11732
rect -15060 -11308 -14288 -11280
rect -15060 -11732 -14372 -11308
rect -14308 -11732 -14288 -11308
rect -15060 -11760 -14288 -11732
rect -14048 -11308 -13276 -11280
rect -14048 -11732 -13360 -11308
rect -13296 -11732 -13276 -11308
rect -14048 -11760 -13276 -11732
rect -13036 -11308 -12264 -11280
rect -13036 -11732 -12348 -11308
rect -12284 -11732 -12264 -11308
rect -13036 -11760 -12264 -11732
rect -12024 -11308 -11252 -11280
rect -12024 -11732 -11336 -11308
rect -11272 -11732 -11252 -11308
rect -12024 -11760 -11252 -11732
rect -11012 -11308 -10240 -11280
rect -11012 -11732 -10324 -11308
rect -10260 -11732 -10240 -11308
rect -11012 -11760 -10240 -11732
rect -10000 -11308 -9228 -11280
rect -10000 -11732 -9312 -11308
rect -9248 -11732 -9228 -11308
rect -10000 -11760 -9228 -11732
rect -8988 -11308 -8216 -11280
rect -8988 -11732 -8300 -11308
rect -8236 -11732 -8216 -11308
rect -8988 -11760 -8216 -11732
rect -7976 -11308 -7204 -11280
rect -7976 -11732 -7288 -11308
rect -7224 -11732 -7204 -11308
rect -7976 -11760 -7204 -11732
rect -6964 -11308 -6192 -11280
rect -6964 -11732 -6276 -11308
rect -6212 -11732 -6192 -11308
rect -6964 -11760 -6192 -11732
rect -5952 -11308 -5180 -11280
rect -5952 -11732 -5264 -11308
rect -5200 -11732 -5180 -11308
rect -5952 -11760 -5180 -11732
rect -4940 -11308 -4168 -11280
rect -4940 -11732 -4252 -11308
rect -4188 -11732 -4168 -11308
rect -4940 -11760 -4168 -11732
rect -3928 -11308 -3156 -11280
rect -3928 -11732 -3240 -11308
rect -3176 -11732 -3156 -11308
rect -3928 -11760 -3156 -11732
rect -2916 -11308 -2144 -11280
rect -2916 -11732 -2228 -11308
rect -2164 -11732 -2144 -11308
rect -2916 -11760 -2144 -11732
rect -1904 -11308 -1132 -11280
rect -1904 -11732 -1216 -11308
rect -1152 -11732 -1132 -11308
rect -1904 -11760 -1132 -11732
rect -892 -11308 -120 -11280
rect -892 -11732 -204 -11308
rect -140 -11732 -120 -11308
rect -892 -11760 -120 -11732
rect 120 -11308 892 -11280
rect 120 -11732 808 -11308
rect 872 -11732 892 -11308
rect 120 -11760 892 -11732
rect 1132 -11308 1904 -11280
rect 1132 -11732 1820 -11308
rect 1884 -11732 1904 -11308
rect 1132 -11760 1904 -11732
rect 2144 -11308 2916 -11280
rect 2144 -11732 2832 -11308
rect 2896 -11732 2916 -11308
rect 2144 -11760 2916 -11732
rect 3156 -11308 3928 -11280
rect 3156 -11732 3844 -11308
rect 3908 -11732 3928 -11308
rect 3156 -11760 3928 -11732
rect 4168 -11308 4940 -11280
rect 4168 -11732 4856 -11308
rect 4920 -11732 4940 -11308
rect 4168 -11760 4940 -11732
rect 5180 -11308 5952 -11280
rect 5180 -11732 5868 -11308
rect 5932 -11732 5952 -11308
rect 5180 -11760 5952 -11732
rect 6192 -11308 6964 -11280
rect 6192 -11732 6880 -11308
rect 6944 -11732 6964 -11308
rect 6192 -11760 6964 -11732
rect 7204 -11308 7976 -11280
rect 7204 -11732 7892 -11308
rect 7956 -11732 7976 -11308
rect 7204 -11760 7976 -11732
rect 8216 -11308 8988 -11280
rect 8216 -11732 8904 -11308
rect 8968 -11732 8988 -11308
rect 8216 -11760 8988 -11732
rect 9228 -11308 10000 -11280
rect 9228 -11732 9916 -11308
rect 9980 -11732 10000 -11308
rect 9228 -11760 10000 -11732
rect 10240 -11308 11012 -11280
rect 10240 -11732 10928 -11308
rect 10992 -11732 11012 -11308
rect 10240 -11760 11012 -11732
rect 11252 -11308 12024 -11280
rect 11252 -11732 11940 -11308
rect 12004 -11732 12024 -11308
rect 11252 -11760 12024 -11732
rect 12264 -11308 13036 -11280
rect 12264 -11732 12952 -11308
rect 13016 -11732 13036 -11308
rect 12264 -11760 13036 -11732
rect 13276 -11308 14048 -11280
rect 13276 -11732 13964 -11308
rect 14028 -11732 14048 -11308
rect 13276 -11760 14048 -11732
rect 14288 -11308 15060 -11280
rect 14288 -11732 14976 -11308
rect 15040 -11732 15060 -11308
rect 14288 -11760 15060 -11732
rect 15300 -11308 16072 -11280
rect 15300 -11732 15988 -11308
rect 16052 -11732 16072 -11308
rect 15300 -11760 16072 -11732
rect 16312 -11308 17084 -11280
rect 16312 -11732 17000 -11308
rect 17064 -11732 17084 -11308
rect 16312 -11760 17084 -11732
<< via3 >>
rect -16396 11308 -16332 11732
rect -15384 11308 -15320 11732
rect -14372 11308 -14308 11732
rect -13360 11308 -13296 11732
rect -12348 11308 -12284 11732
rect -11336 11308 -11272 11732
rect -10324 11308 -10260 11732
rect -9312 11308 -9248 11732
rect -8300 11308 -8236 11732
rect -7288 11308 -7224 11732
rect -6276 11308 -6212 11732
rect -5264 11308 -5200 11732
rect -4252 11308 -4188 11732
rect -3240 11308 -3176 11732
rect -2228 11308 -2164 11732
rect -1216 11308 -1152 11732
rect -204 11308 -140 11732
rect 808 11308 872 11732
rect 1820 11308 1884 11732
rect 2832 11308 2896 11732
rect 3844 11308 3908 11732
rect 4856 11308 4920 11732
rect 5868 11308 5932 11732
rect 6880 11308 6944 11732
rect 7892 11308 7956 11732
rect 8904 11308 8968 11732
rect 9916 11308 9980 11732
rect 10928 11308 10992 11732
rect 11940 11308 12004 11732
rect 12952 11308 13016 11732
rect 13964 11308 14028 11732
rect 14976 11308 15040 11732
rect 15988 11308 16052 11732
rect 17000 11308 17064 11732
rect -16396 10588 -16332 11012
rect -15384 10588 -15320 11012
rect -14372 10588 -14308 11012
rect -13360 10588 -13296 11012
rect -12348 10588 -12284 11012
rect -11336 10588 -11272 11012
rect -10324 10588 -10260 11012
rect -9312 10588 -9248 11012
rect -8300 10588 -8236 11012
rect -7288 10588 -7224 11012
rect -6276 10588 -6212 11012
rect -5264 10588 -5200 11012
rect -4252 10588 -4188 11012
rect -3240 10588 -3176 11012
rect -2228 10588 -2164 11012
rect -1216 10588 -1152 11012
rect -204 10588 -140 11012
rect 808 10588 872 11012
rect 1820 10588 1884 11012
rect 2832 10588 2896 11012
rect 3844 10588 3908 11012
rect 4856 10588 4920 11012
rect 5868 10588 5932 11012
rect 6880 10588 6944 11012
rect 7892 10588 7956 11012
rect 8904 10588 8968 11012
rect 9916 10588 9980 11012
rect 10928 10588 10992 11012
rect 11940 10588 12004 11012
rect 12952 10588 13016 11012
rect 13964 10588 14028 11012
rect 14976 10588 15040 11012
rect 15988 10588 16052 11012
rect 17000 10588 17064 11012
rect -16396 9868 -16332 10292
rect -15384 9868 -15320 10292
rect -14372 9868 -14308 10292
rect -13360 9868 -13296 10292
rect -12348 9868 -12284 10292
rect -11336 9868 -11272 10292
rect -10324 9868 -10260 10292
rect -9312 9868 -9248 10292
rect -8300 9868 -8236 10292
rect -7288 9868 -7224 10292
rect -6276 9868 -6212 10292
rect -5264 9868 -5200 10292
rect -4252 9868 -4188 10292
rect -3240 9868 -3176 10292
rect -2228 9868 -2164 10292
rect -1216 9868 -1152 10292
rect -204 9868 -140 10292
rect 808 9868 872 10292
rect 1820 9868 1884 10292
rect 2832 9868 2896 10292
rect 3844 9868 3908 10292
rect 4856 9868 4920 10292
rect 5868 9868 5932 10292
rect 6880 9868 6944 10292
rect 7892 9868 7956 10292
rect 8904 9868 8968 10292
rect 9916 9868 9980 10292
rect 10928 9868 10992 10292
rect 11940 9868 12004 10292
rect 12952 9868 13016 10292
rect 13964 9868 14028 10292
rect 14976 9868 15040 10292
rect 15988 9868 16052 10292
rect 17000 9868 17064 10292
rect -16396 9148 -16332 9572
rect -15384 9148 -15320 9572
rect -14372 9148 -14308 9572
rect -13360 9148 -13296 9572
rect -12348 9148 -12284 9572
rect -11336 9148 -11272 9572
rect -10324 9148 -10260 9572
rect -9312 9148 -9248 9572
rect -8300 9148 -8236 9572
rect -7288 9148 -7224 9572
rect -6276 9148 -6212 9572
rect -5264 9148 -5200 9572
rect -4252 9148 -4188 9572
rect -3240 9148 -3176 9572
rect -2228 9148 -2164 9572
rect -1216 9148 -1152 9572
rect -204 9148 -140 9572
rect 808 9148 872 9572
rect 1820 9148 1884 9572
rect 2832 9148 2896 9572
rect 3844 9148 3908 9572
rect 4856 9148 4920 9572
rect 5868 9148 5932 9572
rect 6880 9148 6944 9572
rect 7892 9148 7956 9572
rect 8904 9148 8968 9572
rect 9916 9148 9980 9572
rect 10928 9148 10992 9572
rect 11940 9148 12004 9572
rect 12952 9148 13016 9572
rect 13964 9148 14028 9572
rect 14976 9148 15040 9572
rect 15988 9148 16052 9572
rect 17000 9148 17064 9572
rect -16396 8428 -16332 8852
rect -15384 8428 -15320 8852
rect -14372 8428 -14308 8852
rect -13360 8428 -13296 8852
rect -12348 8428 -12284 8852
rect -11336 8428 -11272 8852
rect -10324 8428 -10260 8852
rect -9312 8428 -9248 8852
rect -8300 8428 -8236 8852
rect -7288 8428 -7224 8852
rect -6276 8428 -6212 8852
rect -5264 8428 -5200 8852
rect -4252 8428 -4188 8852
rect -3240 8428 -3176 8852
rect -2228 8428 -2164 8852
rect -1216 8428 -1152 8852
rect -204 8428 -140 8852
rect 808 8428 872 8852
rect 1820 8428 1884 8852
rect 2832 8428 2896 8852
rect 3844 8428 3908 8852
rect 4856 8428 4920 8852
rect 5868 8428 5932 8852
rect 6880 8428 6944 8852
rect 7892 8428 7956 8852
rect 8904 8428 8968 8852
rect 9916 8428 9980 8852
rect 10928 8428 10992 8852
rect 11940 8428 12004 8852
rect 12952 8428 13016 8852
rect 13964 8428 14028 8852
rect 14976 8428 15040 8852
rect 15988 8428 16052 8852
rect 17000 8428 17064 8852
rect -16396 7708 -16332 8132
rect -15384 7708 -15320 8132
rect -14372 7708 -14308 8132
rect -13360 7708 -13296 8132
rect -12348 7708 -12284 8132
rect -11336 7708 -11272 8132
rect -10324 7708 -10260 8132
rect -9312 7708 -9248 8132
rect -8300 7708 -8236 8132
rect -7288 7708 -7224 8132
rect -6276 7708 -6212 8132
rect -5264 7708 -5200 8132
rect -4252 7708 -4188 8132
rect -3240 7708 -3176 8132
rect -2228 7708 -2164 8132
rect -1216 7708 -1152 8132
rect -204 7708 -140 8132
rect 808 7708 872 8132
rect 1820 7708 1884 8132
rect 2832 7708 2896 8132
rect 3844 7708 3908 8132
rect 4856 7708 4920 8132
rect 5868 7708 5932 8132
rect 6880 7708 6944 8132
rect 7892 7708 7956 8132
rect 8904 7708 8968 8132
rect 9916 7708 9980 8132
rect 10928 7708 10992 8132
rect 11940 7708 12004 8132
rect 12952 7708 13016 8132
rect 13964 7708 14028 8132
rect 14976 7708 15040 8132
rect 15988 7708 16052 8132
rect 17000 7708 17064 8132
rect -16396 6988 -16332 7412
rect -15384 6988 -15320 7412
rect -14372 6988 -14308 7412
rect -13360 6988 -13296 7412
rect -12348 6988 -12284 7412
rect -11336 6988 -11272 7412
rect -10324 6988 -10260 7412
rect -9312 6988 -9248 7412
rect -8300 6988 -8236 7412
rect -7288 6988 -7224 7412
rect -6276 6988 -6212 7412
rect -5264 6988 -5200 7412
rect -4252 6988 -4188 7412
rect -3240 6988 -3176 7412
rect -2228 6988 -2164 7412
rect -1216 6988 -1152 7412
rect -204 6988 -140 7412
rect 808 6988 872 7412
rect 1820 6988 1884 7412
rect 2832 6988 2896 7412
rect 3844 6988 3908 7412
rect 4856 6988 4920 7412
rect 5868 6988 5932 7412
rect 6880 6988 6944 7412
rect 7892 6988 7956 7412
rect 8904 6988 8968 7412
rect 9916 6988 9980 7412
rect 10928 6988 10992 7412
rect 11940 6988 12004 7412
rect 12952 6988 13016 7412
rect 13964 6988 14028 7412
rect 14976 6988 15040 7412
rect 15988 6988 16052 7412
rect 17000 6988 17064 7412
rect -16396 6268 -16332 6692
rect -15384 6268 -15320 6692
rect -14372 6268 -14308 6692
rect -13360 6268 -13296 6692
rect -12348 6268 -12284 6692
rect -11336 6268 -11272 6692
rect -10324 6268 -10260 6692
rect -9312 6268 -9248 6692
rect -8300 6268 -8236 6692
rect -7288 6268 -7224 6692
rect -6276 6268 -6212 6692
rect -5264 6268 -5200 6692
rect -4252 6268 -4188 6692
rect -3240 6268 -3176 6692
rect -2228 6268 -2164 6692
rect -1216 6268 -1152 6692
rect -204 6268 -140 6692
rect 808 6268 872 6692
rect 1820 6268 1884 6692
rect 2832 6268 2896 6692
rect 3844 6268 3908 6692
rect 4856 6268 4920 6692
rect 5868 6268 5932 6692
rect 6880 6268 6944 6692
rect 7892 6268 7956 6692
rect 8904 6268 8968 6692
rect 9916 6268 9980 6692
rect 10928 6268 10992 6692
rect 11940 6268 12004 6692
rect 12952 6268 13016 6692
rect 13964 6268 14028 6692
rect 14976 6268 15040 6692
rect 15988 6268 16052 6692
rect 17000 6268 17064 6692
rect -16396 5548 -16332 5972
rect -15384 5548 -15320 5972
rect -14372 5548 -14308 5972
rect -13360 5548 -13296 5972
rect -12348 5548 -12284 5972
rect -11336 5548 -11272 5972
rect -10324 5548 -10260 5972
rect -9312 5548 -9248 5972
rect -8300 5548 -8236 5972
rect -7288 5548 -7224 5972
rect -6276 5548 -6212 5972
rect -5264 5548 -5200 5972
rect -4252 5548 -4188 5972
rect -3240 5548 -3176 5972
rect -2228 5548 -2164 5972
rect -1216 5548 -1152 5972
rect -204 5548 -140 5972
rect 808 5548 872 5972
rect 1820 5548 1884 5972
rect 2832 5548 2896 5972
rect 3844 5548 3908 5972
rect 4856 5548 4920 5972
rect 5868 5548 5932 5972
rect 6880 5548 6944 5972
rect 7892 5548 7956 5972
rect 8904 5548 8968 5972
rect 9916 5548 9980 5972
rect 10928 5548 10992 5972
rect 11940 5548 12004 5972
rect 12952 5548 13016 5972
rect 13964 5548 14028 5972
rect 14976 5548 15040 5972
rect 15988 5548 16052 5972
rect 17000 5548 17064 5972
rect -16396 4828 -16332 5252
rect -15384 4828 -15320 5252
rect -14372 4828 -14308 5252
rect -13360 4828 -13296 5252
rect -12348 4828 -12284 5252
rect -11336 4828 -11272 5252
rect -10324 4828 -10260 5252
rect -9312 4828 -9248 5252
rect -8300 4828 -8236 5252
rect -7288 4828 -7224 5252
rect -6276 4828 -6212 5252
rect -5264 4828 -5200 5252
rect -4252 4828 -4188 5252
rect -3240 4828 -3176 5252
rect -2228 4828 -2164 5252
rect -1216 4828 -1152 5252
rect -204 4828 -140 5252
rect 808 4828 872 5252
rect 1820 4828 1884 5252
rect 2832 4828 2896 5252
rect 3844 4828 3908 5252
rect 4856 4828 4920 5252
rect 5868 4828 5932 5252
rect 6880 4828 6944 5252
rect 7892 4828 7956 5252
rect 8904 4828 8968 5252
rect 9916 4828 9980 5252
rect 10928 4828 10992 5252
rect 11940 4828 12004 5252
rect 12952 4828 13016 5252
rect 13964 4828 14028 5252
rect 14976 4828 15040 5252
rect 15988 4828 16052 5252
rect 17000 4828 17064 5252
rect -16396 4108 -16332 4532
rect -15384 4108 -15320 4532
rect -14372 4108 -14308 4532
rect -13360 4108 -13296 4532
rect -12348 4108 -12284 4532
rect -11336 4108 -11272 4532
rect -10324 4108 -10260 4532
rect -9312 4108 -9248 4532
rect -8300 4108 -8236 4532
rect -7288 4108 -7224 4532
rect -6276 4108 -6212 4532
rect -5264 4108 -5200 4532
rect -4252 4108 -4188 4532
rect -3240 4108 -3176 4532
rect -2228 4108 -2164 4532
rect -1216 4108 -1152 4532
rect -204 4108 -140 4532
rect 808 4108 872 4532
rect 1820 4108 1884 4532
rect 2832 4108 2896 4532
rect 3844 4108 3908 4532
rect 4856 4108 4920 4532
rect 5868 4108 5932 4532
rect 6880 4108 6944 4532
rect 7892 4108 7956 4532
rect 8904 4108 8968 4532
rect 9916 4108 9980 4532
rect 10928 4108 10992 4532
rect 11940 4108 12004 4532
rect 12952 4108 13016 4532
rect 13964 4108 14028 4532
rect 14976 4108 15040 4532
rect 15988 4108 16052 4532
rect 17000 4108 17064 4532
rect -16396 3388 -16332 3812
rect -15384 3388 -15320 3812
rect -14372 3388 -14308 3812
rect -13360 3388 -13296 3812
rect -12348 3388 -12284 3812
rect -11336 3388 -11272 3812
rect -10324 3388 -10260 3812
rect -9312 3388 -9248 3812
rect -8300 3388 -8236 3812
rect -7288 3388 -7224 3812
rect -6276 3388 -6212 3812
rect -5264 3388 -5200 3812
rect -4252 3388 -4188 3812
rect -3240 3388 -3176 3812
rect -2228 3388 -2164 3812
rect -1216 3388 -1152 3812
rect -204 3388 -140 3812
rect 808 3388 872 3812
rect 1820 3388 1884 3812
rect 2832 3388 2896 3812
rect 3844 3388 3908 3812
rect 4856 3388 4920 3812
rect 5868 3388 5932 3812
rect 6880 3388 6944 3812
rect 7892 3388 7956 3812
rect 8904 3388 8968 3812
rect 9916 3388 9980 3812
rect 10928 3388 10992 3812
rect 11940 3388 12004 3812
rect 12952 3388 13016 3812
rect 13964 3388 14028 3812
rect 14976 3388 15040 3812
rect 15988 3388 16052 3812
rect 17000 3388 17064 3812
rect -16396 2668 -16332 3092
rect -15384 2668 -15320 3092
rect -14372 2668 -14308 3092
rect -13360 2668 -13296 3092
rect -12348 2668 -12284 3092
rect -11336 2668 -11272 3092
rect -10324 2668 -10260 3092
rect -9312 2668 -9248 3092
rect -8300 2668 -8236 3092
rect -7288 2668 -7224 3092
rect -6276 2668 -6212 3092
rect -5264 2668 -5200 3092
rect -4252 2668 -4188 3092
rect -3240 2668 -3176 3092
rect -2228 2668 -2164 3092
rect -1216 2668 -1152 3092
rect -204 2668 -140 3092
rect 808 2668 872 3092
rect 1820 2668 1884 3092
rect 2832 2668 2896 3092
rect 3844 2668 3908 3092
rect 4856 2668 4920 3092
rect 5868 2668 5932 3092
rect 6880 2668 6944 3092
rect 7892 2668 7956 3092
rect 8904 2668 8968 3092
rect 9916 2668 9980 3092
rect 10928 2668 10992 3092
rect 11940 2668 12004 3092
rect 12952 2668 13016 3092
rect 13964 2668 14028 3092
rect 14976 2668 15040 3092
rect 15988 2668 16052 3092
rect 17000 2668 17064 3092
rect -16396 1948 -16332 2372
rect -15384 1948 -15320 2372
rect -14372 1948 -14308 2372
rect -13360 1948 -13296 2372
rect -12348 1948 -12284 2372
rect -11336 1948 -11272 2372
rect -10324 1948 -10260 2372
rect -9312 1948 -9248 2372
rect -8300 1948 -8236 2372
rect -7288 1948 -7224 2372
rect -6276 1948 -6212 2372
rect -5264 1948 -5200 2372
rect -4252 1948 -4188 2372
rect -3240 1948 -3176 2372
rect -2228 1948 -2164 2372
rect -1216 1948 -1152 2372
rect -204 1948 -140 2372
rect 808 1948 872 2372
rect 1820 1948 1884 2372
rect 2832 1948 2896 2372
rect 3844 1948 3908 2372
rect 4856 1948 4920 2372
rect 5868 1948 5932 2372
rect 6880 1948 6944 2372
rect 7892 1948 7956 2372
rect 8904 1948 8968 2372
rect 9916 1948 9980 2372
rect 10928 1948 10992 2372
rect 11940 1948 12004 2372
rect 12952 1948 13016 2372
rect 13964 1948 14028 2372
rect 14976 1948 15040 2372
rect 15988 1948 16052 2372
rect 17000 1948 17064 2372
rect -16396 1228 -16332 1652
rect -15384 1228 -15320 1652
rect -14372 1228 -14308 1652
rect -13360 1228 -13296 1652
rect -12348 1228 -12284 1652
rect -11336 1228 -11272 1652
rect -10324 1228 -10260 1652
rect -9312 1228 -9248 1652
rect -8300 1228 -8236 1652
rect -7288 1228 -7224 1652
rect -6276 1228 -6212 1652
rect -5264 1228 -5200 1652
rect -4252 1228 -4188 1652
rect -3240 1228 -3176 1652
rect -2228 1228 -2164 1652
rect -1216 1228 -1152 1652
rect -204 1228 -140 1652
rect 808 1228 872 1652
rect 1820 1228 1884 1652
rect 2832 1228 2896 1652
rect 3844 1228 3908 1652
rect 4856 1228 4920 1652
rect 5868 1228 5932 1652
rect 6880 1228 6944 1652
rect 7892 1228 7956 1652
rect 8904 1228 8968 1652
rect 9916 1228 9980 1652
rect 10928 1228 10992 1652
rect 11940 1228 12004 1652
rect 12952 1228 13016 1652
rect 13964 1228 14028 1652
rect 14976 1228 15040 1652
rect 15988 1228 16052 1652
rect 17000 1228 17064 1652
rect -16396 508 -16332 932
rect -15384 508 -15320 932
rect -14372 508 -14308 932
rect -13360 508 -13296 932
rect -12348 508 -12284 932
rect -11336 508 -11272 932
rect -10324 508 -10260 932
rect -9312 508 -9248 932
rect -8300 508 -8236 932
rect -7288 508 -7224 932
rect -6276 508 -6212 932
rect -5264 508 -5200 932
rect -4252 508 -4188 932
rect -3240 508 -3176 932
rect -2228 508 -2164 932
rect -1216 508 -1152 932
rect -204 508 -140 932
rect 808 508 872 932
rect 1820 508 1884 932
rect 2832 508 2896 932
rect 3844 508 3908 932
rect 4856 508 4920 932
rect 5868 508 5932 932
rect 6880 508 6944 932
rect 7892 508 7956 932
rect 8904 508 8968 932
rect 9916 508 9980 932
rect 10928 508 10992 932
rect 11940 508 12004 932
rect 12952 508 13016 932
rect 13964 508 14028 932
rect 14976 508 15040 932
rect 15988 508 16052 932
rect 17000 508 17064 932
rect -16396 -212 -16332 212
rect -15384 -212 -15320 212
rect -14372 -212 -14308 212
rect -13360 -212 -13296 212
rect -12348 -212 -12284 212
rect -11336 -212 -11272 212
rect -10324 -212 -10260 212
rect -9312 -212 -9248 212
rect -8300 -212 -8236 212
rect -7288 -212 -7224 212
rect -6276 -212 -6212 212
rect -5264 -212 -5200 212
rect -4252 -212 -4188 212
rect -3240 -212 -3176 212
rect -2228 -212 -2164 212
rect -1216 -212 -1152 212
rect -204 -212 -140 212
rect 808 -212 872 212
rect 1820 -212 1884 212
rect 2832 -212 2896 212
rect 3844 -212 3908 212
rect 4856 -212 4920 212
rect 5868 -212 5932 212
rect 6880 -212 6944 212
rect 7892 -212 7956 212
rect 8904 -212 8968 212
rect 9916 -212 9980 212
rect 10928 -212 10992 212
rect 11940 -212 12004 212
rect 12952 -212 13016 212
rect 13964 -212 14028 212
rect 14976 -212 15040 212
rect 15988 -212 16052 212
rect 17000 -212 17064 212
rect -16396 -932 -16332 -508
rect -15384 -932 -15320 -508
rect -14372 -932 -14308 -508
rect -13360 -932 -13296 -508
rect -12348 -932 -12284 -508
rect -11336 -932 -11272 -508
rect -10324 -932 -10260 -508
rect -9312 -932 -9248 -508
rect -8300 -932 -8236 -508
rect -7288 -932 -7224 -508
rect -6276 -932 -6212 -508
rect -5264 -932 -5200 -508
rect -4252 -932 -4188 -508
rect -3240 -932 -3176 -508
rect -2228 -932 -2164 -508
rect -1216 -932 -1152 -508
rect -204 -932 -140 -508
rect 808 -932 872 -508
rect 1820 -932 1884 -508
rect 2832 -932 2896 -508
rect 3844 -932 3908 -508
rect 4856 -932 4920 -508
rect 5868 -932 5932 -508
rect 6880 -932 6944 -508
rect 7892 -932 7956 -508
rect 8904 -932 8968 -508
rect 9916 -932 9980 -508
rect 10928 -932 10992 -508
rect 11940 -932 12004 -508
rect 12952 -932 13016 -508
rect 13964 -932 14028 -508
rect 14976 -932 15040 -508
rect 15988 -932 16052 -508
rect 17000 -932 17064 -508
rect -16396 -1652 -16332 -1228
rect -15384 -1652 -15320 -1228
rect -14372 -1652 -14308 -1228
rect -13360 -1652 -13296 -1228
rect -12348 -1652 -12284 -1228
rect -11336 -1652 -11272 -1228
rect -10324 -1652 -10260 -1228
rect -9312 -1652 -9248 -1228
rect -8300 -1652 -8236 -1228
rect -7288 -1652 -7224 -1228
rect -6276 -1652 -6212 -1228
rect -5264 -1652 -5200 -1228
rect -4252 -1652 -4188 -1228
rect -3240 -1652 -3176 -1228
rect -2228 -1652 -2164 -1228
rect -1216 -1652 -1152 -1228
rect -204 -1652 -140 -1228
rect 808 -1652 872 -1228
rect 1820 -1652 1884 -1228
rect 2832 -1652 2896 -1228
rect 3844 -1652 3908 -1228
rect 4856 -1652 4920 -1228
rect 5868 -1652 5932 -1228
rect 6880 -1652 6944 -1228
rect 7892 -1652 7956 -1228
rect 8904 -1652 8968 -1228
rect 9916 -1652 9980 -1228
rect 10928 -1652 10992 -1228
rect 11940 -1652 12004 -1228
rect 12952 -1652 13016 -1228
rect 13964 -1652 14028 -1228
rect 14976 -1652 15040 -1228
rect 15988 -1652 16052 -1228
rect 17000 -1652 17064 -1228
rect -16396 -2372 -16332 -1948
rect -15384 -2372 -15320 -1948
rect -14372 -2372 -14308 -1948
rect -13360 -2372 -13296 -1948
rect -12348 -2372 -12284 -1948
rect -11336 -2372 -11272 -1948
rect -10324 -2372 -10260 -1948
rect -9312 -2372 -9248 -1948
rect -8300 -2372 -8236 -1948
rect -7288 -2372 -7224 -1948
rect -6276 -2372 -6212 -1948
rect -5264 -2372 -5200 -1948
rect -4252 -2372 -4188 -1948
rect -3240 -2372 -3176 -1948
rect -2228 -2372 -2164 -1948
rect -1216 -2372 -1152 -1948
rect -204 -2372 -140 -1948
rect 808 -2372 872 -1948
rect 1820 -2372 1884 -1948
rect 2832 -2372 2896 -1948
rect 3844 -2372 3908 -1948
rect 4856 -2372 4920 -1948
rect 5868 -2372 5932 -1948
rect 6880 -2372 6944 -1948
rect 7892 -2372 7956 -1948
rect 8904 -2372 8968 -1948
rect 9916 -2372 9980 -1948
rect 10928 -2372 10992 -1948
rect 11940 -2372 12004 -1948
rect 12952 -2372 13016 -1948
rect 13964 -2372 14028 -1948
rect 14976 -2372 15040 -1948
rect 15988 -2372 16052 -1948
rect 17000 -2372 17064 -1948
rect -16396 -3092 -16332 -2668
rect -15384 -3092 -15320 -2668
rect -14372 -3092 -14308 -2668
rect -13360 -3092 -13296 -2668
rect -12348 -3092 -12284 -2668
rect -11336 -3092 -11272 -2668
rect -10324 -3092 -10260 -2668
rect -9312 -3092 -9248 -2668
rect -8300 -3092 -8236 -2668
rect -7288 -3092 -7224 -2668
rect -6276 -3092 -6212 -2668
rect -5264 -3092 -5200 -2668
rect -4252 -3092 -4188 -2668
rect -3240 -3092 -3176 -2668
rect -2228 -3092 -2164 -2668
rect -1216 -3092 -1152 -2668
rect -204 -3092 -140 -2668
rect 808 -3092 872 -2668
rect 1820 -3092 1884 -2668
rect 2832 -3092 2896 -2668
rect 3844 -3092 3908 -2668
rect 4856 -3092 4920 -2668
rect 5868 -3092 5932 -2668
rect 6880 -3092 6944 -2668
rect 7892 -3092 7956 -2668
rect 8904 -3092 8968 -2668
rect 9916 -3092 9980 -2668
rect 10928 -3092 10992 -2668
rect 11940 -3092 12004 -2668
rect 12952 -3092 13016 -2668
rect 13964 -3092 14028 -2668
rect 14976 -3092 15040 -2668
rect 15988 -3092 16052 -2668
rect 17000 -3092 17064 -2668
rect -16396 -3812 -16332 -3388
rect -15384 -3812 -15320 -3388
rect -14372 -3812 -14308 -3388
rect -13360 -3812 -13296 -3388
rect -12348 -3812 -12284 -3388
rect -11336 -3812 -11272 -3388
rect -10324 -3812 -10260 -3388
rect -9312 -3812 -9248 -3388
rect -8300 -3812 -8236 -3388
rect -7288 -3812 -7224 -3388
rect -6276 -3812 -6212 -3388
rect -5264 -3812 -5200 -3388
rect -4252 -3812 -4188 -3388
rect -3240 -3812 -3176 -3388
rect -2228 -3812 -2164 -3388
rect -1216 -3812 -1152 -3388
rect -204 -3812 -140 -3388
rect 808 -3812 872 -3388
rect 1820 -3812 1884 -3388
rect 2832 -3812 2896 -3388
rect 3844 -3812 3908 -3388
rect 4856 -3812 4920 -3388
rect 5868 -3812 5932 -3388
rect 6880 -3812 6944 -3388
rect 7892 -3812 7956 -3388
rect 8904 -3812 8968 -3388
rect 9916 -3812 9980 -3388
rect 10928 -3812 10992 -3388
rect 11940 -3812 12004 -3388
rect 12952 -3812 13016 -3388
rect 13964 -3812 14028 -3388
rect 14976 -3812 15040 -3388
rect 15988 -3812 16052 -3388
rect 17000 -3812 17064 -3388
rect -16396 -4532 -16332 -4108
rect -15384 -4532 -15320 -4108
rect -14372 -4532 -14308 -4108
rect -13360 -4532 -13296 -4108
rect -12348 -4532 -12284 -4108
rect -11336 -4532 -11272 -4108
rect -10324 -4532 -10260 -4108
rect -9312 -4532 -9248 -4108
rect -8300 -4532 -8236 -4108
rect -7288 -4532 -7224 -4108
rect -6276 -4532 -6212 -4108
rect -5264 -4532 -5200 -4108
rect -4252 -4532 -4188 -4108
rect -3240 -4532 -3176 -4108
rect -2228 -4532 -2164 -4108
rect -1216 -4532 -1152 -4108
rect -204 -4532 -140 -4108
rect 808 -4532 872 -4108
rect 1820 -4532 1884 -4108
rect 2832 -4532 2896 -4108
rect 3844 -4532 3908 -4108
rect 4856 -4532 4920 -4108
rect 5868 -4532 5932 -4108
rect 6880 -4532 6944 -4108
rect 7892 -4532 7956 -4108
rect 8904 -4532 8968 -4108
rect 9916 -4532 9980 -4108
rect 10928 -4532 10992 -4108
rect 11940 -4532 12004 -4108
rect 12952 -4532 13016 -4108
rect 13964 -4532 14028 -4108
rect 14976 -4532 15040 -4108
rect 15988 -4532 16052 -4108
rect 17000 -4532 17064 -4108
rect -16396 -5252 -16332 -4828
rect -15384 -5252 -15320 -4828
rect -14372 -5252 -14308 -4828
rect -13360 -5252 -13296 -4828
rect -12348 -5252 -12284 -4828
rect -11336 -5252 -11272 -4828
rect -10324 -5252 -10260 -4828
rect -9312 -5252 -9248 -4828
rect -8300 -5252 -8236 -4828
rect -7288 -5252 -7224 -4828
rect -6276 -5252 -6212 -4828
rect -5264 -5252 -5200 -4828
rect -4252 -5252 -4188 -4828
rect -3240 -5252 -3176 -4828
rect -2228 -5252 -2164 -4828
rect -1216 -5252 -1152 -4828
rect -204 -5252 -140 -4828
rect 808 -5252 872 -4828
rect 1820 -5252 1884 -4828
rect 2832 -5252 2896 -4828
rect 3844 -5252 3908 -4828
rect 4856 -5252 4920 -4828
rect 5868 -5252 5932 -4828
rect 6880 -5252 6944 -4828
rect 7892 -5252 7956 -4828
rect 8904 -5252 8968 -4828
rect 9916 -5252 9980 -4828
rect 10928 -5252 10992 -4828
rect 11940 -5252 12004 -4828
rect 12952 -5252 13016 -4828
rect 13964 -5252 14028 -4828
rect 14976 -5252 15040 -4828
rect 15988 -5252 16052 -4828
rect 17000 -5252 17064 -4828
rect -16396 -5972 -16332 -5548
rect -15384 -5972 -15320 -5548
rect -14372 -5972 -14308 -5548
rect -13360 -5972 -13296 -5548
rect -12348 -5972 -12284 -5548
rect -11336 -5972 -11272 -5548
rect -10324 -5972 -10260 -5548
rect -9312 -5972 -9248 -5548
rect -8300 -5972 -8236 -5548
rect -7288 -5972 -7224 -5548
rect -6276 -5972 -6212 -5548
rect -5264 -5972 -5200 -5548
rect -4252 -5972 -4188 -5548
rect -3240 -5972 -3176 -5548
rect -2228 -5972 -2164 -5548
rect -1216 -5972 -1152 -5548
rect -204 -5972 -140 -5548
rect 808 -5972 872 -5548
rect 1820 -5972 1884 -5548
rect 2832 -5972 2896 -5548
rect 3844 -5972 3908 -5548
rect 4856 -5972 4920 -5548
rect 5868 -5972 5932 -5548
rect 6880 -5972 6944 -5548
rect 7892 -5972 7956 -5548
rect 8904 -5972 8968 -5548
rect 9916 -5972 9980 -5548
rect 10928 -5972 10992 -5548
rect 11940 -5972 12004 -5548
rect 12952 -5972 13016 -5548
rect 13964 -5972 14028 -5548
rect 14976 -5972 15040 -5548
rect 15988 -5972 16052 -5548
rect 17000 -5972 17064 -5548
rect -16396 -6692 -16332 -6268
rect -15384 -6692 -15320 -6268
rect -14372 -6692 -14308 -6268
rect -13360 -6692 -13296 -6268
rect -12348 -6692 -12284 -6268
rect -11336 -6692 -11272 -6268
rect -10324 -6692 -10260 -6268
rect -9312 -6692 -9248 -6268
rect -8300 -6692 -8236 -6268
rect -7288 -6692 -7224 -6268
rect -6276 -6692 -6212 -6268
rect -5264 -6692 -5200 -6268
rect -4252 -6692 -4188 -6268
rect -3240 -6692 -3176 -6268
rect -2228 -6692 -2164 -6268
rect -1216 -6692 -1152 -6268
rect -204 -6692 -140 -6268
rect 808 -6692 872 -6268
rect 1820 -6692 1884 -6268
rect 2832 -6692 2896 -6268
rect 3844 -6692 3908 -6268
rect 4856 -6692 4920 -6268
rect 5868 -6692 5932 -6268
rect 6880 -6692 6944 -6268
rect 7892 -6692 7956 -6268
rect 8904 -6692 8968 -6268
rect 9916 -6692 9980 -6268
rect 10928 -6692 10992 -6268
rect 11940 -6692 12004 -6268
rect 12952 -6692 13016 -6268
rect 13964 -6692 14028 -6268
rect 14976 -6692 15040 -6268
rect 15988 -6692 16052 -6268
rect 17000 -6692 17064 -6268
rect -16396 -7412 -16332 -6988
rect -15384 -7412 -15320 -6988
rect -14372 -7412 -14308 -6988
rect -13360 -7412 -13296 -6988
rect -12348 -7412 -12284 -6988
rect -11336 -7412 -11272 -6988
rect -10324 -7412 -10260 -6988
rect -9312 -7412 -9248 -6988
rect -8300 -7412 -8236 -6988
rect -7288 -7412 -7224 -6988
rect -6276 -7412 -6212 -6988
rect -5264 -7412 -5200 -6988
rect -4252 -7412 -4188 -6988
rect -3240 -7412 -3176 -6988
rect -2228 -7412 -2164 -6988
rect -1216 -7412 -1152 -6988
rect -204 -7412 -140 -6988
rect 808 -7412 872 -6988
rect 1820 -7412 1884 -6988
rect 2832 -7412 2896 -6988
rect 3844 -7412 3908 -6988
rect 4856 -7412 4920 -6988
rect 5868 -7412 5932 -6988
rect 6880 -7412 6944 -6988
rect 7892 -7412 7956 -6988
rect 8904 -7412 8968 -6988
rect 9916 -7412 9980 -6988
rect 10928 -7412 10992 -6988
rect 11940 -7412 12004 -6988
rect 12952 -7412 13016 -6988
rect 13964 -7412 14028 -6988
rect 14976 -7412 15040 -6988
rect 15988 -7412 16052 -6988
rect 17000 -7412 17064 -6988
rect -16396 -8132 -16332 -7708
rect -15384 -8132 -15320 -7708
rect -14372 -8132 -14308 -7708
rect -13360 -8132 -13296 -7708
rect -12348 -8132 -12284 -7708
rect -11336 -8132 -11272 -7708
rect -10324 -8132 -10260 -7708
rect -9312 -8132 -9248 -7708
rect -8300 -8132 -8236 -7708
rect -7288 -8132 -7224 -7708
rect -6276 -8132 -6212 -7708
rect -5264 -8132 -5200 -7708
rect -4252 -8132 -4188 -7708
rect -3240 -8132 -3176 -7708
rect -2228 -8132 -2164 -7708
rect -1216 -8132 -1152 -7708
rect -204 -8132 -140 -7708
rect 808 -8132 872 -7708
rect 1820 -8132 1884 -7708
rect 2832 -8132 2896 -7708
rect 3844 -8132 3908 -7708
rect 4856 -8132 4920 -7708
rect 5868 -8132 5932 -7708
rect 6880 -8132 6944 -7708
rect 7892 -8132 7956 -7708
rect 8904 -8132 8968 -7708
rect 9916 -8132 9980 -7708
rect 10928 -8132 10992 -7708
rect 11940 -8132 12004 -7708
rect 12952 -8132 13016 -7708
rect 13964 -8132 14028 -7708
rect 14976 -8132 15040 -7708
rect 15988 -8132 16052 -7708
rect 17000 -8132 17064 -7708
rect -16396 -8852 -16332 -8428
rect -15384 -8852 -15320 -8428
rect -14372 -8852 -14308 -8428
rect -13360 -8852 -13296 -8428
rect -12348 -8852 -12284 -8428
rect -11336 -8852 -11272 -8428
rect -10324 -8852 -10260 -8428
rect -9312 -8852 -9248 -8428
rect -8300 -8852 -8236 -8428
rect -7288 -8852 -7224 -8428
rect -6276 -8852 -6212 -8428
rect -5264 -8852 -5200 -8428
rect -4252 -8852 -4188 -8428
rect -3240 -8852 -3176 -8428
rect -2228 -8852 -2164 -8428
rect -1216 -8852 -1152 -8428
rect -204 -8852 -140 -8428
rect 808 -8852 872 -8428
rect 1820 -8852 1884 -8428
rect 2832 -8852 2896 -8428
rect 3844 -8852 3908 -8428
rect 4856 -8852 4920 -8428
rect 5868 -8852 5932 -8428
rect 6880 -8852 6944 -8428
rect 7892 -8852 7956 -8428
rect 8904 -8852 8968 -8428
rect 9916 -8852 9980 -8428
rect 10928 -8852 10992 -8428
rect 11940 -8852 12004 -8428
rect 12952 -8852 13016 -8428
rect 13964 -8852 14028 -8428
rect 14976 -8852 15040 -8428
rect 15988 -8852 16052 -8428
rect 17000 -8852 17064 -8428
rect -16396 -9572 -16332 -9148
rect -15384 -9572 -15320 -9148
rect -14372 -9572 -14308 -9148
rect -13360 -9572 -13296 -9148
rect -12348 -9572 -12284 -9148
rect -11336 -9572 -11272 -9148
rect -10324 -9572 -10260 -9148
rect -9312 -9572 -9248 -9148
rect -8300 -9572 -8236 -9148
rect -7288 -9572 -7224 -9148
rect -6276 -9572 -6212 -9148
rect -5264 -9572 -5200 -9148
rect -4252 -9572 -4188 -9148
rect -3240 -9572 -3176 -9148
rect -2228 -9572 -2164 -9148
rect -1216 -9572 -1152 -9148
rect -204 -9572 -140 -9148
rect 808 -9572 872 -9148
rect 1820 -9572 1884 -9148
rect 2832 -9572 2896 -9148
rect 3844 -9572 3908 -9148
rect 4856 -9572 4920 -9148
rect 5868 -9572 5932 -9148
rect 6880 -9572 6944 -9148
rect 7892 -9572 7956 -9148
rect 8904 -9572 8968 -9148
rect 9916 -9572 9980 -9148
rect 10928 -9572 10992 -9148
rect 11940 -9572 12004 -9148
rect 12952 -9572 13016 -9148
rect 13964 -9572 14028 -9148
rect 14976 -9572 15040 -9148
rect 15988 -9572 16052 -9148
rect 17000 -9572 17064 -9148
rect -16396 -10292 -16332 -9868
rect -15384 -10292 -15320 -9868
rect -14372 -10292 -14308 -9868
rect -13360 -10292 -13296 -9868
rect -12348 -10292 -12284 -9868
rect -11336 -10292 -11272 -9868
rect -10324 -10292 -10260 -9868
rect -9312 -10292 -9248 -9868
rect -8300 -10292 -8236 -9868
rect -7288 -10292 -7224 -9868
rect -6276 -10292 -6212 -9868
rect -5264 -10292 -5200 -9868
rect -4252 -10292 -4188 -9868
rect -3240 -10292 -3176 -9868
rect -2228 -10292 -2164 -9868
rect -1216 -10292 -1152 -9868
rect -204 -10292 -140 -9868
rect 808 -10292 872 -9868
rect 1820 -10292 1884 -9868
rect 2832 -10292 2896 -9868
rect 3844 -10292 3908 -9868
rect 4856 -10292 4920 -9868
rect 5868 -10292 5932 -9868
rect 6880 -10292 6944 -9868
rect 7892 -10292 7956 -9868
rect 8904 -10292 8968 -9868
rect 9916 -10292 9980 -9868
rect 10928 -10292 10992 -9868
rect 11940 -10292 12004 -9868
rect 12952 -10292 13016 -9868
rect 13964 -10292 14028 -9868
rect 14976 -10292 15040 -9868
rect 15988 -10292 16052 -9868
rect 17000 -10292 17064 -9868
rect -16396 -11012 -16332 -10588
rect -15384 -11012 -15320 -10588
rect -14372 -11012 -14308 -10588
rect -13360 -11012 -13296 -10588
rect -12348 -11012 -12284 -10588
rect -11336 -11012 -11272 -10588
rect -10324 -11012 -10260 -10588
rect -9312 -11012 -9248 -10588
rect -8300 -11012 -8236 -10588
rect -7288 -11012 -7224 -10588
rect -6276 -11012 -6212 -10588
rect -5264 -11012 -5200 -10588
rect -4252 -11012 -4188 -10588
rect -3240 -11012 -3176 -10588
rect -2228 -11012 -2164 -10588
rect -1216 -11012 -1152 -10588
rect -204 -11012 -140 -10588
rect 808 -11012 872 -10588
rect 1820 -11012 1884 -10588
rect 2832 -11012 2896 -10588
rect 3844 -11012 3908 -10588
rect 4856 -11012 4920 -10588
rect 5868 -11012 5932 -10588
rect 6880 -11012 6944 -10588
rect 7892 -11012 7956 -10588
rect 8904 -11012 8968 -10588
rect 9916 -11012 9980 -10588
rect 10928 -11012 10992 -10588
rect 11940 -11012 12004 -10588
rect 12952 -11012 13016 -10588
rect 13964 -11012 14028 -10588
rect 14976 -11012 15040 -10588
rect 15988 -11012 16052 -10588
rect 17000 -11012 17064 -10588
rect -16396 -11732 -16332 -11308
rect -15384 -11732 -15320 -11308
rect -14372 -11732 -14308 -11308
rect -13360 -11732 -13296 -11308
rect -12348 -11732 -12284 -11308
rect -11336 -11732 -11272 -11308
rect -10324 -11732 -10260 -11308
rect -9312 -11732 -9248 -11308
rect -8300 -11732 -8236 -11308
rect -7288 -11732 -7224 -11308
rect -6276 -11732 -6212 -11308
rect -5264 -11732 -5200 -11308
rect -4252 -11732 -4188 -11308
rect -3240 -11732 -3176 -11308
rect -2228 -11732 -2164 -11308
rect -1216 -11732 -1152 -11308
rect -204 -11732 -140 -11308
rect 808 -11732 872 -11308
rect 1820 -11732 1884 -11308
rect 2832 -11732 2896 -11308
rect 3844 -11732 3908 -11308
rect 4856 -11732 4920 -11308
rect 5868 -11732 5932 -11308
rect 6880 -11732 6944 -11308
rect 7892 -11732 7956 -11308
rect 8904 -11732 8968 -11308
rect 9916 -11732 9980 -11308
rect 10928 -11732 10992 -11308
rect 11940 -11732 12004 -11308
rect 12952 -11732 13016 -11308
rect 13964 -11732 14028 -11308
rect 14976 -11732 15040 -11308
rect 15988 -11732 16052 -11308
rect 17000 -11732 17064 -11308
<< mimcap >>
rect -17044 11680 -16644 11720
rect -17044 11360 -17004 11680
rect -16684 11360 -16644 11680
rect -17044 11320 -16644 11360
rect -16032 11680 -15632 11720
rect -16032 11360 -15992 11680
rect -15672 11360 -15632 11680
rect -16032 11320 -15632 11360
rect -15020 11680 -14620 11720
rect -15020 11360 -14980 11680
rect -14660 11360 -14620 11680
rect -15020 11320 -14620 11360
rect -14008 11680 -13608 11720
rect -14008 11360 -13968 11680
rect -13648 11360 -13608 11680
rect -14008 11320 -13608 11360
rect -12996 11680 -12596 11720
rect -12996 11360 -12956 11680
rect -12636 11360 -12596 11680
rect -12996 11320 -12596 11360
rect -11984 11680 -11584 11720
rect -11984 11360 -11944 11680
rect -11624 11360 -11584 11680
rect -11984 11320 -11584 11360
rect -10972 11680 -10572 11720
rect -10972 11360 -10932 11680
rect -10612 11360 -10572 11680
rect -10972 11320 -10572 11360
rect -9960 11680 -9560 11720
rect -9960 11360 -9920 11680
rect -9600 11360 -9560 11680
rect -9960 11320 -9560 11360
rect -8948 11680 -8548 11720
rect -8948 11360 -8908 11680
rect -8588 11360 -8548 11680
rect -8948 11320 -8548 11360
rect -7936 11680 -7536 11720
rect -7936 11360 -7896 11680
rect -7576 11360 -7536 11680
rect -7936 11320 -7536 11360
rect -6924 11680 -6524 11720
rect -6924 11360 -6884 11680
rect -6564 11360 -6524 11680
rect -6924 11320 -6524 11360
rect -5912 11680 -5512 11720
rect -5912 11360 -5872 11680
rect -5552 11360 -5512 11680
rect -5912 11320 -5512 11360
rect -4900 11680 -4500 11720
rect -4900 11360 -4860 11680
rect -4540 11360 -4500 11680
rect -4900 11320 -4500 11360
rect -3888 11680 -3488 11720
rect -3888 11360 -3848 11680
rect -3528 11360 -3488 11680
rect -3888 11320 -3488 11360
rect -2876 11680 -2476 11720
rect -2876 11360 -2836 11680
rect -2516 11360 -2476 11680
rect -2876 11320 -2476 11360
rect -1864 11680 -1464 11720
rect -1864 11360 -1824 11680
rect -1504 11360 -1464 11680
rect -1864 11320 -1464 11360
rect -852 11680 -452 11720
rect -852 11360 -812 11680
rect -492 11360 -452 11680
rect -852 11320 -452 11360
rect 160 11680 560 11720
rect 160 11360 200 11680
rect 520 11360 560 11680
rect 160 11320 560 11360
rect 1172 11680 1572 11720
rect 1172 11360 1212 11680
rect 1532 11360 1572 11680
rect 1172 11320 1572 11360
rect 2184 11680 2584 11720
rect 2184 11360 2224 11680
rect 2544 11360 2584 11680
rect 2184 11320 2584 11360
rect 3196 11680 3596 11720
rect 3196 11360 3236 11680
rect 3556 11360 3596 11680
rect 3196 11320 3596 11360
rect 4208 11680 4608 11720
rect 4208 11360 4248 11680
rect 4568 11360 4608 11680
rect 4208 11320 4608 11360
rect 5220 11680 5620 11720
rect 5220 11360 5260 11680
rect 5580 11360 5620 11680
rect 5220 11320 5620 11360
rect 6232 11680 6632 11720
rect 6232 11360 6272 11680
rect 6592 11360 6632 11680
rect 6232 11320 6632 11360
rect 7244 11680 7644 11720
rect 7244 11360 7284 11680
rect 7604 11360 7644 11680
rect 7244 11320 7644 11360
rect 8256 11680 8656 11720
rect 8256 11360 8296 11680
rect 8616 11360 8656 11680
rect 8256 11320 8656 11360
rect 9268 11680 9668 11720
rect 9268 11360 9308 11680
rect 9628 11360 9668 11680
rect 9268 11320 9668 11360
rect 10280 11680 10680 11720
rect 10280 11360 10320 11680
rect 10640 11360 10680 11680
rect 10280 11320 10680 11360
rect 11292 11680 11692 11720
rect 11292 11360 11332 11680
rect 11652 11360 11692 11680
rect 11292 11320 11692 11360
rect 12304 11680 12704 11720
rect 12304 11360 12344 11680
rect 12664 11360 12704 11680
rect 12304 11320 12704 11360
rect 13316 11680 13716 11720
rect 13316 11360 13356 11680
rect 13676 11360 13716 11680
rect 13316 11320 13716 11360
rect 14328 11680 14728 11720
rect 14328 11360 14368 11680
rect 14688 11360 14728 11680
rect 14328 11320 14728 11360
rect 15340 11680 15740 11720
rect 15340 11360 15380 11680
rect 15700 11360 15740 11680
rect 15340 11320 15740 11360
rect 16352 11680 16752 11720
rect 16352 11360 16392 11680
rect 16712 11360 16752 11680
rect 16352 11320 16752 11360
rect -17044 10960 -16644 11000
rect -17044 10640 -17004 10960
rect -16684 10640 -16644 10960
rect -17044 10600 -16644 10640
rect -16032 10960 -15632 11000
rect -16032 10640 -15992 10960
rect -15672 10640 -15632 10960
rect -16032 10600 -15632 10640
rect -15020 10960 -14620 11000
rect -15020 10640 -14980 10960
rect -14660 10640 -14620 10960
rect -15020 10600 -14620 10640
rect -14008 10960 -13608 11000
rect -14008 10640 -13968 10960
rect -13648 10640 -13608 10960
rect -14008 10600 -13608 10640
rect -12996 10960 -12596 11000
rect -12996 10640 -12956 10960
rect -12636 10640 -12596 10960
rect -12996 10600 -12596 10640
rect -11984 10960 -11584 11000
rect -11984 10640 -11944 10960
rect -11624 10640 -11584 10960
rect -11984 10600 -11584 10640
rect -10972 10960 -10572 11000
rect -10972 10640 -10932 10960
rect -10612 10640 -10572 10960
rect -10972 10600 -10572 10640
rect -9960 10960 -9560 11000
rect -9960 10640 -9920 10960
rect -9600 10640 -9560 10960
rect -9960 10600 -9560 10640
rect -8948 10960 -8548 11000
rect -8948 10640 -8908 10960
rect -8588 10640 -8548 10960
rect -8948 10600 -8548 10640
rect -7936 10960 -7536 11000
rect -7936 10640 -7896 10960
rect -7576 10640 -7536 10960
rect -7936 10600 -7536 10640
rect -6924 10960 -6524 11000
rect -6924 10640 -6884 10960
rect -6564 10640 -6524 10960
rect -6924 10600 -6524 10640
rect -5912 10960 -5512 11000
rect -5912 10640 -5872 10960
rect -5552 10640 -5512 10960
rect -5912 10600 -5512 10640
rect -4900 10960 -4500 11000
rect -4900 10640 -4860 10960
rect -4540 10640 -4500 10960
rect -4900 10600 -4500 10640
rect -3888 10960 -3488 11000
rect -3888 10640 -3848 10960
rect -3528 10640 -3488 10960
rect -3888 10600 -3488 10640
rect -2876 10960 -2476 11000
rect -2876 10640 -2836 10960
rect -2516 10640 -2476 10960
rect -2876 10600 -2476 10640
rect -1864 10960 -1464 11000
rect -1864 10640 -1824 10960
rect -1504 10640 -1464 10960
rect -1864 10600 -1464 10640
rect -852 10960 -452 11000
rect -852 10640 -812 10960
rect -492 10640 -452 10960
rect -852 10600 -452 10640
rect 160 10960 560 11000
rect 160 10640 200 10960
rect 520 10640 560 10960
rect 160 10600 560 10640
rect 1172 10960 1572 11000
rect 1172 10640 1212 10960
rect 1532 10640 1572 10960
rect 1172 10600 1572 10640
rect 2184 10960 2584 11000
rect 2184 10640 2224 10960
rect 2544 10640 2584 10960
rect 2184 10600 2584 10640
rect 3196 10960 3596 11000
rect 3196 10640 3236 10960
rect 3556 10640 3596 10960
rect 3196 10600 3596 10640
rect 4208 10960 4608 11000
rect 4208 10640 4248 10960
rect 4568 10640 4608 10960
rect 4208 10600 4608 10640
rect 5220 10960 5620 11000
rect 5220 10640 5260 10960
rect 5580 10640 5620 10960
rect 5220 10600 5620 10640
rect 6232 10960 6632 11000
rect 6232 10640 6272 10960
rect 6592 10640 6632 10960
rect 6232 10600 6632 10640
rect 7244 10960 7644 11000
rect 7244 10640 7284 10960
rect 7604 10640 7644 10960
rect 7244 10600 7644 10640
rect 8256 10960 8656 11000
rect 8256 10640 8296 10960
rect 8616 10640 8656 10960
rect 8256 10600 8656 10640
rect 9268 10960 9668 11000
rect 9268 10640 9308 10960
rect 9628 10640 9668 10960
rect 9268 10600 9668 10640
rect 10280 10960 10680 11000
rect 10280 10640 10320 10960
rect 10640 10640 10680 10960
rect 10280 10600 10680 10640
rect 11292 10960 11692 11000
rect 11292 10640 11332 10960
rect 11652 10640 11692 10960
rect 11292 10600 11692 10640
rect 12304 10960 12704 11000
rect 12304 10640 12344 10960
rect 12664 10640 12704 10960
rect 12304 10600 12704 10640
rect 13316 10960 13716 11000
rect 13316 10640 13356 10960
rect 13676 10640 13716 10960
rect 13316 10600 13716 10640
rect 14328 10960 14728 11000
rect 14328 10640 14368 10960
rect 14688 10640 14728 10960
rect 14328 10600 14728 10640
rect 15340 10960 15740 11000
rect 15340 10640 15380 10960
rect 15700 10640 15740 10960
rect 15340 10600 15740 10640
rect 16352 10960 16752 11000
rect 16352 10640 16392 10960
rect 16712 10640 16752 10960
rect 16352 10600 16752 10640
rect -17044 10240 -16644 10280
rect -17044 9920 -17004 10240
rect -16684 9920 -16644 10240
rect -17044 9880 -16644 9920
rect -16032 10240 -15632 10280
rect -16032 9920 -15992 10240
rect -15672 9920 -15632 10240
rect -16032 9880 -15632 9920
rect -15020 10240 -14620 10280
rect -15020 9920 -14980 10240
rect -14660 9920 -14620 10240
rect -15020 9880 -14620 9920
rect -14008 10240 -13608 10280
rect -14008 9920 -13968 10240
rect -13648 9920 -13608 10240
rect -14008 9880 -13608 9920
rect -12996 10240 -12596 10280
rect -12996 9920 -12956 10240
rect -12636 9920 -12596 10240
rect -12996 9880 -12596 9920
rect -11984 10240 -11584 10280
rect -11984 9920 -11944 10240
rect -11624 9920 -11584 10240
rect -11984 9880 -11584 9920
rect -10972 10240 -10572 10280
rect -10972 9920 -10932 10240
rect -10612 9920 -10572 10240
rect -10972 9880 -10572 9920
rect -9960 10240 -9560 10280
rect -9960 9920 -9920 10240
rect -9600 9920 -9560 10240
rect -9960 9880 -9560 9920
rect -8948 10240 -8548 10280
rect -8948 9920 -8908 10240
rect -8588 9920 -8548 10240
rect -8948 9880 -8548 9920
rect -7936 10240 -7536 10280
rect -7936 9920 -7896 10240
rect -7576 9920 -7536 10240
rect -7936 9880 -7536 9920
rect -6924 10240 -6524 10280
rect -6924 9920 -6884 10240
rect -6564 9920 -6524 10240
rect -6924 9880 -6524 9920
rect -5912 10240 -5512 10280
rect -5912 9920 -5872 10240
rect -5552 9920 -5512 10240
rect -5912 9880 -5512 9920
rect -4900 10240 -4500 10280
rect -4900 9920 -4860 10240
rect -4540 9920 -4500 10240
rect -4900 9880 -4500 9920
rect -3888 10240 -3488 10280
rect -3888 9920 -3848 10240
rect -3528 9920 -3488 10240
rect -3888 9880 -3488 9920
rect -2876 10240 -2476 10280
rect -2876 9920 -2836 10240
rect -2516 9920 -2476 10240
rect -2876 9880 -2476 9920
rect -1864 10240 -1464 10280
rect -1864 9920 -1824 10240
rect -1504 9920 -1464 10240
rect -1864 9880 -1464 9920
rect -852 10240 -452 10280
rect -852 9920 -812 10240
rect -492 9920 -452 10240
rect -852 9880 -452 9920
rect 160 10240 560 10280
rect 160 9920 200 10240
rect 520 9920 560 10240
rect 160 9880 560 9920
rect 1172 10240 1572 10280
rect 1172 9920 1212 10240
rect 1532 9920 1572 10240
rect 1172 9880 1572 9920
rect 2184 10240 2584 10280
rect 2184 9920 2224 10240
rect 2544 9920 2584 10240
rect 2184 9880 2584 9920
rect 3196 10240 3596 10280
rect 3196 9920 3236 10240
rect 3556 9920 3596 10240
rect 3196 9880 3596 9920
rect 4208 10240 4608 10280
rect 4208 9920 4248 10240
rect 4568 9920 4608 10240
rect 4208 9880 4608 9920
rect 5220 10240 5620 10280
rect 5220 9920 5260 10240
rect 5580 9920 5620 10240
rect 5220 9880 5620 9920
rect 6232 10240 6632 10280
rect 6232 9920 6272 10240
rect 6592 9920 6632 10240
rect 6232 9880 6632 9920
rect 7244 10240 7644 10280
rect 7244 9920 7284 10240
rect 7604 9920 7644 10240
rect 7244 9880 7644 9920
rect 8256 10240 8656 10280
rect 8256 9920 8296 10240
rect 8616 9920 8656 10240
rect 8256 9880 8656 9920
rect 9268 10240 9668 10280
rect 9268 9920 9308 10240
rect 9628 9920 9668 10240
rect 9268 9880 9668 9920
rect 10280 10240 10680 10280
rect 10280 9920 10320 10240
rect 10640 9920 10680 10240
rect 10280 9880 10680 9920
rect 11292 10240 11692 10280
rect 11292 9920 11332 10240
rect 11652 9920 11692 10240
rect 11292 9880 11692 9920
rect 12304 10240 12704 10280
rect 12304 9920 12344 10240
rect 12664 9920 12704 10240
rect 12304 9880 12704 9920
rect 13316 10240 13716 10280
rect 13316 9920 13356 10240
rect 13676 9920 13716 10240
rect 13316 9880 13716 9920
rect 14328 10240 14728 10280
rect 14328 9920 14368 10240
rect 14688 9920 14728 10240
rect 14328 9880 14728 9920
rect 15340 10240 15740 10280
rect 15340 9920 15380 10240
rect 15700 9920 15740 10240
rect 15340 9880 15740 9920
rect 16352 10240 16752 10280
rect 16352 9920 16392 10240
rect 16712 9920 16752 10240
rect 16352 9880 16752 9920
rect -17044 9520 -16644 9560
rect -17044 9200 -17004 9520
rect -16684 9200 -16644 9520
rect -17044 9160 -16644 9200
rect -16032 9520 -15632 9560
rect -16032 9200 -15992 9520
rect -15672 9200 -15632 9520
rect -16032 9160 -15632 9200
rect -15020 9520 -14620 9560
rect -15020 9200 -14980 9520
rect -14660 9200 -14620 9520
rect -15020 9160 -14620 9200
rect -14008 9520 -13608 9560
rect -14008 9200 -13968 9520
rect -13648 9200 -13608 9520
rect -14008 9160 -13608 9200
rect -12996 9520 -12596 9560
rect -12996 9200 -12956 9520
rect -12636 9200 -12596 9520
rect -12996 9160 -12596 9200
rect -11984 9520 -11584 9560
rect -11984 9200 -11944 9520
rect -11624 9200 -11584 9520
rect -11984 9160 -11584 9200
rect -10972 9520 -10572 9560
rect -10972 9200 -10932 9520
rect -10612 9200 -10572 9520
rect -10972 9160 -10572 9200
rect -9960 9520 -9560 9560
rect -9960 9200 -9920 9520
rect -9600 9200 -9560 9520
rect -9960 9160 -9560 9200
rect -8948 9520 -8548 9560
rect -8948 9200 -8908 9520
rect -8588 9200 -8548 9520
rect -8948 9160 -8548 9200
rect -7936 9520 -7536 9560
rect -7936 9200 -7896 9520
rect -7576 9200 -7536 9520
rect -7936 9160 -7536 9200
rect -6924 9520 -6524 9560
rect -6924 9200 -6884 9520
rect -6564 9200 -6524 9520
rect -6924 9160 -6524 9200
rect -5912 9520 -5512 9560
rect -5912 9200 -5872 9520
rect -5552 9200 -5512 9520
rect -5912 9160 -5512 9200
rect -4900 9520 -4500 9560
rect -4900 9200 -4860 9520
rect -4540 9200 -4500 9520
rect -4900 9160 -4500 9200
rect -3888 9520 -3488 9560
rect -3888 9200 -3848 9520
rect -3528 9200 -3488 9520
rect -3888 9160 -3488 9200
rect -2876 9520 -2476 9560
rect -2876 9200 -2836 9520
rect -2516 9200 -2476 9520
rect -2876 9160 -2476 9200
rect -1864 9520 -1464 9560
rect -1864 9200 -1824 9520
rect -1504 9200 -1464 9520
rect -1864 9160 -1464 9200
rect -852 9520 -452 9560
rect -852 9200 -812 9520
rect -492 9200 -452 9520
rect -852 9160 -452 9200
rect 160 9520 560 9560
rect 160 9200 200 9520
rect 520 9200 560 9520
rect 160 9160 560 9200
rect 1172 9520 1572 9560
rect 1172 9200 1212 9520
rect 1532 9200 1572 9520
rect 1172 9160 1572 9200
rect 2184 9520 2584 9560
rect 2184 9200 2224 9520
rect 2544 9200 2584 9520
rect 2184 9160 2584 9200
rect 3196 9520 3596 9560
rect 3196 9200 3236 9520
rect 3556 9200 3596 9520
rect 3196 9160 3596 9200
rect 4208 9520 4608 9560
rect 4208 9200 4248 9520
rect 4568 9200 4608 9520
rect 4208 9160 4608 9200
rect 5220 9520 5620 9560
rect 5220 9200 5260 9520
rect 5580 9200 5620 9520
rect 5220 9160 5620 9200
rect 6232 9520 6632 9560
rect 6232 9200 6272 9520
rect 6592 9200 6632 9520
rect 6232 9160 6632 9200
rect 7244 9520 7644 9560
rect 7244 9200 7284 9520
rect 7604 9200 7644 9520
rect 7244 9160 7644 9200
rect 8256 9520 8656 9560
rect 8256 9200 8296 9520
rect 8616 9200 8656 9520
rect 8256 9160 8656 9200
rect 9268 9520 9668 9560
rect 9268 9200 9308 9520
rect 9628 9200 9668 9520
rect 9268 9160 9668 9200
rect 10280 9520 10680 9560
rect 10280 9200 10320 9520
rect 10640 9200 10680 9520
rect 10280 9160 10680 9200
rect 11292 9520 11692 9560
rect 11292 9200 11332 9520
rect 11652 9200 11692 9520
rect 11292 9160 11692 9200
rect 12304 9520 12704 9560
rect 12304 9200 12344 9520
rect 12664 9200 12704 9520
rect 12304 9160 12704 9200
rect 13316 9520 13716 9560
rect 13316 9200 13356 9520
rect 13676 9200 13716 9520
rect 13316 9160 13716 9200
rect 14328 9520 14728 9560
rect 14328 9200 14368 9520
rect 14688 9200 14728 9520
rect 14328 9160 14728 9200
rect 15340 9520 15740 9560
rect 15340 9200 15380 9520
rect 15700 9200 15740 9520
rect 15340 9160 15740 9200
rect 16352 9520 16752 9560
rect 16352 9200 16392 9520
rect 16712 9200 16752 9520
rect 16352 9160 16752 9200
rect -17044 8800 -16644 8840
rect -17044 8480 -17004 8800
rect -16684 8480 -16644 8800
rect -17044 8440 -16644 8480
rect -16032 8800 -15632 8840
rect -16032 8480 -15992 8800
rect -15672 8480 -15632 8800
rect -16032 8440 -15632 8480
rect -15020 8800 -14620 8840
rect -15020 8480 -14980 8800
rect -14660 8480 -14620 8800
rect -15020 8440 -14620 8480
rect -14008 8800 -13608 8840
rect -14008 8480 -13968 8800
rect -13648 8480 -13608 8800
rect -14008 8440 -13608 8480
rect -12996 8800 -12596 8840
rect -12996 8480 -12956 8800
rect -12636 8480 -12596 8800
rect -12996 8440 -12596 8480
rect -11984 8800 -11584 8840
rect -11984 8480 -11944 8800
rect -11624 8480 -11584 8800
rect -11984 8440 -11584 8480
rect -10972 8800 -10572 8840
rect -10972 8480 -10932 8800
rect -10612 8480 -10572 8800
rect -10972 8440 -10572 8480
rect -9960 8800 -9560 8840
rect -9960 8480 -9920 8800
rect -9600 8480 -9560 8800
rect -9960 8440 -9560 8480
rect -8948 8800 -8548 8840
rect -8948 8480 -8908 8800
rect -8588 8480 -8548 8800
rect -8948 8440 -8548 8480
rect -7936 8800 -7536 8840
rect -7936 8480 -7896 8800
rect -7576 8480 -7536 8800
rect -7936 8440 -7536 8480
rect -6924 8800 -6524 8840
rect -6924 8480 -6884 8800
rect -6564 8480 -6524 8800
rect -6924 8440 -6524 8480
rect -5912 8800 -5512 8840
rect -5912 8480 -5872 8800
rect -5552 8480 -5512 8800
rect -5912 8440 -5512 8480
rect -4900 8800 -4500 8840
rect -4900 8480 -4860 8800
rect -4540 8480 -4500 8800
rect -4900 8440 -4500 8480
rect -3888 8800 -3488 8840
rect -3888 8480 -3848 8800
rect -3528 8480 -3488 8800
rect -3888 8440 -3488 8480
rect -2876 8800 -2476 8840
rect -2876 8480 -2836 8800
rect -2516 8480 -2476 8800
rect -2876 8440 -2476 8480
rect -1864 8800 -1464 8840
rect -1864 8480 -1824 8800
rect -1504 8480 -1464 8800
rect -1864 8440 -1464 8480
rect -852 8800 -452 8840
rect -852 8480 -812 8800
rect -492 8480 -452 8800
rect -852 8440 -452 8480
rect 160 8800 560 8840
rect 160 8480 200 8800
rect 520 8480 560 8800
rect 160 8440 560 8480
rect 1172 8800 1572 8840
rect 1172 8480 1212 8800
rect 1532 8480 1572 8800
rect 1172 8440 1572 8480
rect 2184 8800 2584 8840
rect 2184 8480 2224 8800
rect 2544 8480 2584 8800
rect 2184 8440 2584 8480
rect 3196 8800 3596 8840
rect 3196 8480 3236 8800
rect 3556 8480 3596 8800
rect 3196 8440 3596 8480
rect 4208 8800 4608 8840
rect 4208 8480 4248 8800
rect 4568 8480 4608 8800
rect 4208 8440 4608 8480
rect 5220 8800 5620 8840
rect 5220 8480 5260 8800
rect 5580 8480 5620 8800
rect 5220 8440 5620 8480
rect 6232 8800 6632 8840
rect 6232 8480 6272 8800
rect 6592 8480 6632 8800
rect 6232 8440 6632 8480
rect 7244 8800 7644 8840
rect 7244 8480 7284 8800
rect 7604 8480 7644 8800
rect 7244 8440 7644 8480
rect 8256 8800 8656 8840
rect 8256 8480 8296 8800
rect 8616 8480 8656 8800
rect 8256 8440 8656 8480
rect 9268 8800 9668 8840
rect 9268 8480 9308 8800
rect 9628 8480 9668 8800
rect 9268 8440 9668 8480
rect 10280 8800 10680 8840
rect 10280 8480 10320 8800
rect 10640 8480 10680 8800
rect 10280 8440 10680 8480
rect 11292 8800 11692 8840
rect 11292 8480 11332 8800
rect 11652 8480 11692 8800
rect 11292 8440 11692 8480
rect 12304 8800 12704 8840
rect 12304 8480 12344 8800
rect 12664 8480 12704 8800
rect 12304 8440 12704 8480
rect 13316 8800 13716 8840
rect 13316 8480 13356 8800
rect 13676 8480 13716 8800
rect 13316 8440 13716 8480
rect 14328 8800 14728 8840
rect 14328 8480 14368 8800
rect 14688 8480 14728 8800
rect 14328 8440 14728 8480
rect 15340 8800 15740 8840
rect 15340 8480 15380 8800
rect 15700 8480 15740 8800
rect 15340 8440 15740 8480
rect 16352 8800 16752 8840
rect 16352 8480 16392 8800
rect 16712 8480 16752 8800
rect 16352 8440 16752 8480
rect -17044 8080 -16644 8120
rect -17044 7760 -17004 8080
rect -16684 7760 -16644 8080
rect -17044 7720 -16644 7760
rect -16032 8080 -15632 8120
rect -16032 7760 -15992 8080
rect -15672 7760 -15632 8080
rect -16032 7720 -15632 7760
rect -15020 8080 -14620 8120
rect -15020 7760 -14980 8080
rect -14660 7760 -14620 8080
rect -15020 7720 -14620 7760
rect -14008 8080 -13608 8120
rect -14008 7760 -13968 8080
rect -13648 7760 -13608 8080
rect -14008 7720 -13608 7760
rect -12996 8080 -12596 8120
rect -12996 7760 -12956 8080
rect -12636 7760 -12596 8080
rect -12996 7720 -12596 7760
rect -11984 8080 -11584 8120
rect -11984 7760 -11944 8080
rect -11624 7760 -11584 8080
rect -11984 7720 -11584 7760
rect -10972 8080 -10572 8120
rect -10972 7760 -10932 8080
rect -10612 7760 -10572 8080
rect -10972 7720 -10572 7760
rect -9960 8080 -9560 8120
rect -9960 7760 -9920 8080
rect -9600 7760 -9560 8080
rect -9960 7720 -9560 7760
rect -8948 8080 -8548 8120
rect -8948 7760 -8908 8080
rect -8588 7760 -8548 8080
rect -8948 7720 -8548 7760
rect -7936 8080 -7536 8120
rect -7936 7760 -7896 8080
rect -7576 7760 -7536 8080
rect -7936 7720 -7536 7760
rect -6924 8080 -6524 8120
rect -6924 7760 -6884 8080
rect -6564 7760 -6524 8080
rect -6924 7720 -6524 7760
rect -5912 8080 -5512 8120
rect -5912 7760 -5872 8080
rect -5552 7760 -5512 8080
rect -5912 7720 -5512 7760
rect -4900 8080 -4500 8120
rect -4900 7760 -4860 8080
rect -4540 7760 -4500 8080
rect -4900 7720 -4500 7760
rect -3888 8080 -3488 8120
rect -3888 7760 -3848 8080
rect -3528 7760 -3488 8080
rect -3888 7720 -3488 7760
rect -2876 8080 -2476 8120
rect -2876 7760 -2836 8080
rect -2516 7760 -2476 8080
rect -2876 7720 -2476 7760
rect -1864 8080 -1464 8120
rect -1864 7760 -1824 8080
rect -1504 7760 -1464 8080
rect -1864 7720 -1464 7760
rect -852 8080 -452 8120
rect -852 7760 -812 8080
rect -492 7760 -452 8080
rect -852 7720 -452 7760
rect 160 8080 560 8120
rect 160 7760 200 8080
rect 520 7760 560 8080
rect 160 7720 560 7760
rect 1172 8080 1572 8120
rect 1172 7760 1212 8080
rect 1532 7760 1572 8080
rect 1172 7720 1572 7760
rect 2184 8080 2584 8120
rect 2184 7760 2224 8080
rect 2544 7760 2584 8080
rect 2184 7720 2584 7760
rect 3196 8080 3596 8120
rect 3196 7760 3236 8080
rect 3556 7760 3596 8080
rect 3196 7720 3596 7760
rect 4208 8080 4608 8120
rect 4208 7760 4248 8080
rect 4568 7760 4608 8080
rect 4208 7720 4608 7760
rect 5220 8080 5620 8120
rect 5220 7760 5260 8080
rect 5580 7760 5620 8080
rect 5220 7720 5620 7760
rect 6232 8080 6632 8120
rect 6232 7760 6272 8080
rect 6592 7760 6632 8080
rect 6232 7720 6632 7760
rect 7244 8080 7644 8120
rect 7244 7760 7284 8080
rect 7604 7760 7644 8080
rect 7244 7720 7644 7760
rect 8256 8080 8656 8120
rect 8256 7760 8296 8080
rect 8616 7760 8656 8080
rect 8256 7720 8656 7760
rect 9268 8080 9668 8120
rect 9268 7760 9308 8080
rect 9628 7760 9668 8080
rect 9268 7720 9668 7760
rect 10280 8080 10680 8120
rect 10280 7760 10320 8080
rect 10640 7760 10680 8080
rect 10280 7720 10680 7760
rect 11292 8080 11692 8120
rect 11292 7760 11332 8080
rect 11652 7760 11692 8080
rect 11292 7720 11692 7760
rect 12304 8080 12704 8120
rect 12304 7760 12344 8080
rect 12664 7760 12704 8080
rect 12304 7720 12704 7760
rect 13316 8080 13716 8120
rect 13316 7760 13356 8080
rect 13676 7760 13716 8080
rect 13316 7720 13716 7760
rect 14328 8080 14728 8120
rect 14328 7760 14368 8080
rect 14688 7760 14728 8080
rect 14328 7720 14728 7760
rect 15340 8080 15740 8120
rect 15340 7760 15380 8080
rect 15700 7760 15740 8080
rect 15340 7720 15740 7760
rect 16352 8080 16752 8120
rect 16352 7760 16392 8080
rect 16712 7760 16752 8080
rect 16352 7720 16752 7760
rect -17044 7360 -16644 7400
rect -17044 7040 -17004 7360
rect -16684 7040 -16644 7360
rect -17044 7000 -16644 7040
rect -16032 7360 -15632 7400
rect -16032 7040 -15992 7360
rect -15672 7040 -15632 7360
rect -16032 7000 -15632 7040
rect -15020 7360 -14620 7400
rect -15020 7040 -14980 7360
rect -14660 7040 -14620 7360
rect -15020 7000 -14620 7040
rect -14008 7360 -13608 7400
rect -14008 7040 -13968 7360
rect -13648 7040 -13608 7360
rect -14008 7000 -13608 7040
rect -12996 7360 -12596 7400
rect -12996 7040 -12956 7360
rect -12636 7040 -12596 7360
rect -12996 7000 -12596 7040
rect -11984 7360 -11584 7400
rect -11984 7040 -11944 7360
rect -11624 7040 -11584 7360
rect -11984 7000 -11584 7040
rect -10972 7360 -10572 7400
rect -10972 7040 -10932 7360
rect -10612 7040 -10572 7360
rect -10972 7000 -10572 7040
rect -9960 7360 -9560 7400
rect -9960 7040 -9920 7360
rect -9600 7040 -9560 7360
rect -9960 7000 -9560 7040
rect -8948 7360 -8548 7400
rect -8948 7040 -8908 7360
rect -8588 7040 -8548 7360
rect -8948 7000 -8548 7040
rect -7936 7360 -7536 7400
rect -7936 7040 -7896 7360
rect -7576 7040 -7536 7360
rect -7936 7000 -7536 7040
rect -6924 7360 -6524 7400
rect -6924 7040 -6884 7360
rect -6564 7040 -6524 7360
rect -6924 7000 -6524 7040
rect -5912 7360 -5512 7400
rect -5912 7040 -5872 7360
rect -5552 7040 -5512 7360
rect -5912 7000 -5512 7040
rect -4900 7360 -4500 7400
rect -4900 7040 -4860 7360
rect -4540 7040 -4500 7360
rect -4900 7000 -4500 7040
rect -3888 7360 -3488 7400
rect -3888 7040 -3848 7360
rect -3528 7040 -3488 7360
rect -3888 7000 -3488 7040
rect -2876 7360 -2476 7400
rect -2876 7040 -2836 7360
rect -2516 7040 -2476 7360
rect -2876 7000 -2476 7040
rect -1864 7360 -1464 7400
rect -1864 7040 -1824 7360
rect -1504 7040 -1464 7360
rect -1864 7000 -1464 7040
rect -852 7360 -452 7400
rect -852 7040 -812 7360
rect -492 7040 -452 7360
rect -852 7000 -452 7040
rect 160 7360 560 7400
rect 160 7040 200 7360
rect 520 7040 560 7360
rect 160 7000 560 7040
rect 1172 7360 1572 7400
rect 1172 7040 1212 7360
rect 1532 7040 1572 7360
rect 1172 7000 1572 7040
rect 2184 7360 2584 7400
rect 2184 7040 2224 7360
rect 2544 7040 2584 7360
rect 2184 7000 2584 7040
rect 3196 7360 3596 7400
rect 3196 7040 3236 7360
rect 3556 7040 3596 7360
rect 3196 7000 3596 7040
rect 4208 7360 4608 7400
rect 4208 7040 4248 7360
rect 4568 7040 4608 7360
rect 4208 7000 4608 7040
rect 5220 7360 5620 7400
rect 5220 7040 5260 7360
rect 5580 7040 5620 7360
rect 5220 7000 5620 7040
rect 6232 7360 6632 7400
rect 6232 7040 6272 7360
rect 6592 7040 6632 7360
rect 6232 7000 6632 7040
rect 7244 7360 7644 7400
rect 7244 7040 7284 7360
rect 7604 7040 7644 7360
rect 7244 7000 7644 7040
rect 8256 7360 8656 7400
rect 8256 7040 8296 7360
rect 8616 7040 8656 7360
rect 8256 7000 8656 7040
rect 9268 7360 9668 7400
rect 9268 7040 9308 7360
rect 9628 7040 9668 7360
rect 9268 7000 9668 7040
rect 10280 7360 10680 7400
rect 10280 7040 10320 7360
rect 10640 7040 10680 7360
rect 10280 7000 10680 7040
rect 11292 7360 11692 7400
rect 11292 7040 11332 7360
rect 11652 7040 11692 7360
rect 11292 7000 11692 7040
rect 12304 7360 12704 7400
rect 12304 7040 12344 7360
rect 12664 7040 12704 7360
rect 12304 7000 12704 7040
rect 13316 7360 13716 7400
rect 13316 7040 13356 7360
rect 13676 7040 13716 7360
rect 13316 7000 13716 7040
rect 14328 7360 14728 7400
rect 14328 7040 14368 7360
rect 14688 7040 14728 7360
rect 14328 7000 14728 7040
rect 15340 7360 15740 7400
rect 15340 7040 15380 7360
rect 15700 7040 15740 7360
rect 15340 7000 15740 7040
rect 16352 7360 16752 7400
rect 16352 7040 16392 7360
rect 16712 7040 16752 7360
rect 16352 7000 16752 7040
rect -17044 6640 -16644 6680
rect -17044 6320 -17004 6640
rect -16684 6320 -16644 6640
rect -17044 6280 -16644 6320
rect -16032 6640 -15632 6680
rect -16032 6320 -15992 6640
rect -15672 6320 -15632 6640
rect -16032 6280 -15632 6320
rect -15020 6640 -14620 6680
rect -15020 6320 -14980 6640
rect -14660 6320 -14620 6640
rect -15020 6280 -14620 6320
rect -14008 6640 -13608 6680
rect -14008 6320 -13968 6640
rect -13648 6320 -13608 6640
rect -14008 6280 -13608 6320
rect -12996 6640 -12596 6680
rect -12996 6320 -12956 6640
rect -12636 6320 -12596 6640
rect -12996 6280 -12596 6320
rect -11984 6640 -11584 6680
rect -11984 6320 -11944 6640
rect -11624 6320 -11584 6640
rect -11984 6280 -11584 6320
rect -10972 6640 -10572 6680
rect -10972 6320 -10932 6640
rect -10612 6320 -10572 6640
rect -10972 6280 -10572 6320
rect -9960 6640 -9560 6680
rect -9960 6320 -9920 6640
rect -9600 6320 -9560 6640
rect -9960 6280 -9560 6320
rect -8948 6640 -8548 6680
rect -8948 6320 -8908 6640
rect -8588 6320 -8548 6640
rect -8948 6280 -8548 6320
rect -7936 6640 -7536 6680
rect -7936 6320 -7896 6640
rect -7576 6320 -7536 6640
rect -7936 6280 -7536 6320
rect -6924 6640 -6524 6680
rect -6924 6320 -6884 6640
rect -6564 6320 -6524 6640
rect -6924 6280 -6524 6320
rect -5912 6640 -5512 6680
rect -5912 6320 -5872 6640
rect -5552 6320 -5512 6640
rect -5912 6280 -5512 6320
rect -4900 6640 -4500 6680
rect -4900 6320 -4860 6640
rect -4540 6320 -4500 6640
rect -4900 6280 -4500 6320
rect -3888 6640 -3488 6680
rect -3888 6320 -3848 6640
rect -3528 6320 -3488 6640
rect -3888 6280 -3488 6320
rect -2876 6640 -2476 6680
rect -2876 6320 -2836 6640
rect -2516 6320 -2476 6640
rect -2876 6280 -2476 6320
rect -1864 6640 -1464 6680
rect -1864 6320 -1824 6640
rect -1504 6320 -1464 6640
rect -1864 6280 -1464 6320
rect -852 6640 -452 6680
rect -852 6320 -812 6640
rect -492 6320 -452 6640
rect -852 6280 -452 6320
rect 160 6640 560 6680
rect 160 6320 200 6640
rect 520 6320 560 6640
rect 160 6280 560 6320
rect 1172 6640 1572 6680
rect 1172 6320 1212 6640
rect 1532 6320 1572 6640
rect 1172 6280 1572 6320
rect 2184 6640 2584 6680
rect 2184 6320 2224 6640
rect 2544 6320 2584 6640
rect 2184 6280 2584 6320
rect 3196 6640 3596 6680
rect 3196 6320 3236 6640
rect 3556 6320 3596 6640
rect 3196 6280 3596 6320
rect 4208 6640 4608 6680
rect 4208 6320 4248 6640
rect 4568 6320 4608 6640
rect 4208 6280 4608 6320
rect 5220 6640 5620 6680
rect 5220 6320 5260 6640
rect 5580 6320 5620 6640
rect 5220 6280 5620 6320
rect 6232 6640 6632 6680
rect 6232 6320 6272 6640
rect 6592 6320 6632 6640
rect 6232 6280 6632 6320
rect 7244 6640 7644 6680
rect 7244 6320 7284 6640
rect 7604 6320 7644 6640
rect 7244 6280 7644 6320
rect 8256 6640 8656 6680
rect 8256 6320 8296 6640
rect 8616 6320 8656 6640
rect 8256 6280 8656 6320
rect 9268 6640 9668 6680
rect 9268 6320 9308 6640
rect 9628 6320 9668 6640
rect 9268 6280 9668 6320
rect 10280 6640 10680 6680
rect 10280 6320 10320 6640
rect 10640 6320 10680 6640
rect 10280 6280 10680 6320
rect 11292 6640 11692 6680
rect 11292 6320 11332 6640
rect 11652 6320 11692 6640
rect 11292 6280 11692 6320
rect 12304 6640 12704 6680
rect 12304 6320 12344 6640
rect 12664 6320 12704 6640
rect 12304 6280 12704 6320
rect 13316 6640 13716 6680
rect 13316 6320 13356 6640
rect 13676 6320 13716 6640
rect 13316 6280 13716 6320
rect 14328 6640 14728 6680
rect 14328 6320 14368 6640
rect 14688 6320 14728 6640
rect 14328 6280 14728 6320
rect 15340 6640 15740 6680
rect 15340 6320 15380 6640
rect 15700 6320 15740 6640
rect 15340 6280 15740 6320
rect 16352 6640 16752 6680
rect 16352 6320 16392 6640
rect 16712 6320 16752 6640
rect 16352 6280 16752 6320
rect -17044 5920 -16644 5960
rect -17044 5600 -17004 5920
rect -16684 5600 -16644 5920
rect -17044 5560 -16644 5600
rect -16032 5920 -15632 5960
rect -16032 5600 -15992 5920
rect -15672 5600 -15632 5920
rect -16032 5560 -15632 5600
rect -15020 5920 -14620 5960
rect -15020 5600 -14980 5920
rect -14660 5600 -14620 5920
rect -15020 5560 -14620 5600
rect -14008 5920 -13608 5960
rect -14008 5600 -13968 5920
rect -13648 5600 -13608 5920
rect -14008 5560 -13608 5600
rect -12996 5920 -12596 5960
rect -12996 5600 -12956 5920
rect -12636 5600 -12596 5920
rect -12996 5560 -12596 5600
rect -11984 5920 -11584 5960
rect -11984 5600 -11944 5920
rect -11624 5600 -11584 5920
rect -11984 5560 -11584 5600
rect -10972 5920 -10572 5960
rect -10972 5600 -10932 5920
rect -10612 5600 -10572 5920
rect -10972 5560 -10572 5600
rect -9960 5920 -9560 5960
rect -9960 5600 -9920 5920
rect -9600 5600 -9560 5920
rect -9960 5560 -9560 5600
rect -8948 5920 -8548 5960
rect -8948 5600 -8908 5920
rect -8588 5600 -8548 5920
rect -8948 5560 -8548 5600
rect -7936 5920 -7536 5960
rect -7936 5600 -7896 5920
rect -7576 5600 -7536 5920
rect -7936 5560 -7536 5600
rect -6924 5920 -6524 5960
rect -6924 5600 -6884 5920
rect -6564 5600 -6524 5920
rect -6924 5560 -6524 5600
rect -5912 5920 -5512 5960
rect -5912 5600 -5872 5920
rect -5552 5600 -5512 5920
rect -5912 5560 -5512 5600
rect -4900 5920 -4500 5960
rect -4900 5600 -4860 5920
rect -4540 5600 -4500 5920
rect -4900 5560 -4500 5600
rect -3888 5920 -3488 5960
rect -3888 5600 -3848 5920
rect -3528 5600 -3488 5920
rect -3888 5560 -3488 5600
rect -2876 5920 -2476 5960
rect -2876 5600 -2836 5920
rect -2516 5600 -2476 5920
rect -2876 5560 -2476 5600
rect -1864 5920 -1464 5960
rect -1864 5600 -1824 5920
rect -1504 5600 -1464 5920
rect -1864 5560 -1464 5600
rect -852 5920 -452 5960
rect -852 5600 -812 5920
rect -492 5600 -452 5920
rect -852 5560 -452 5600
rect 160 5920 560 5960
rect 160 5600 200 5920
rect 520 5600 560 5920
rect 160 5560 560 5600
rect 1172 5920 1572 5960
rect 1172 5600 1212 5920
rect 1532 5600 1572 5920
rect 1172 5560 1572 5600
rect 2184 5920 2584 5960
rect 2184 5600 2224 5920
rect 2544 5600 2584 5920
rect 2184 5560 2584 5600
rect 3196 5920 3596 5960
rect 3196 5600 3236 5920
rect 3556 5600 3596 5920
rect 3196 5560 3596 5600
rect 4208 5920 4608 5960
rect 4208 5600 4248 5920
rect 4568 5600 4608 5920
rect 4208 5560 4608 5600
rect 5220 5920 5620 5960
rect 5220 5600 5260 5920
rect 5580 5600 5620 5920
rect 5220 5560 5620 5600
rect 6232 5920 6632 5960
rect 6232 5600 6272 5920
rect 6592 5600 6632 5920
rect 6232 5560 6632 5600
rect 7244 5920 7644 5960
rect 7244 5600 7284 5920
rect 7604 5600 7644 5920
rect 7244 5560 7644 5600
rect 8256 5920 8656 5960
rect 8256 5600 8296 5920
rect 8616 5600 8656 5920
rect 8256 5560 8656 5600
rect 9268 5920 9668 5960
rect 9268 5600 9308 5920
rect 9628 5600 9668 5920
rect 9268 5560 9668 5600
rect 10280 5920 10680 5960
rect 10280 5600 10320 5920
rect 10640 5600 10680 5920
rect 10280 5560 10680 5600
rect 11292 5920 11692 5960
rect 11292 5600 11332 5920
rect 11652 5600 11692 5920
rect 11292 5560 11692 5600
rect 12304 5920 12704 5960
rect 12304 5600 12344 5920
rect 12664 5600 12704 5920
rect 12304 5560 12704 5600
rect 13316 5920 13716 5960
rect 13316 5600 13356 5920
rect 13676 5600 13716 5920
rect 13316 5560 13716 5600
rect 14328 5920 14728 5960
rect 14328 5600 14368 5920
rect 14688 5600 14728 5920
rect 14328 5560 14728 5600
rect 15340 5920 15740 5960
rect 15340 5600 15380 5920
rect 15700 5600 15740 5920
rect 15340 5560 15740 5600
rect 16352 5920 16752 5960
rect 16352 5600 16392 5920
rect 16712 5600 16752 5920
rect 16352 5560 16752 5600
rect -17044 5200 -16644 5240
rect -17044 4880 -17004 5200
rect -16684 4880 -16644 5200
rect -17044 4840 -16644 4880
rect -16032 5200 -15632 5240
rect -16032 4880 -15992 5200
rect -15672 4880 -15632 5200
rect -16032 4840 -15632 4880
rect -15020 5200 -14620 5240
rect -15020 4880 -14980 5200
rect -14660 4880 -14620 5200
rect -15020 4840 -14620 4880
rect -14008 5200 -13608 5240
rect -14008 4880 -13968 5200
rect -13648 4880 -13608 5200
rect -14008 4840 -13608 4880
rect -12996 5200 -12596 5240
rect -12996 4880 -12956 5200
rect -12636 4880 -12596 5200
rect -12996 4840 -12596 4880
rect -11984 5200 -11584 5240
rect -11984 4880 -11944 5200
rect -11624 4880 -11584 5200
rect -11984 4840 -11584 4880
rect -10972 5200 -10572 5240
rect -10972 4880 -10932 5200
rect -10612 4880 -10572 5200
rect -10972 4840 -10572 4880
rect -9960 5200 -9560 5240
rect -9960 4880 -9920 5200
rect -9600 4880 -9560 5200
rect -9960 4840 -9560 4880
rect -8948 5200 -8548 5240
rect -8948 4880 -8908 5200
rect -8588 4880 -8548 5200
rect -8948 4840 -8548 4880
rect -7936 5200 -7536 5240
rect -7936 4880 -7896 5200
rect -7576 4880 -7536 5200
rect -7936 4840 -7536 4880
rect -6924 5200 -6524 5240
rect -6924 4880 -6884 5200
rect -6564 4880 -6524 5200
rect -6924 4840 -6524 4880
rect -5912 5200 -5512 5240
rect -5912 4880 -5872 5200
rect -5552 4880 -5512 5200
rect -5912 4840 -5512 4880
rect -4900 5200 -4500 5240
rect -4900 4880 -4860 5200
rect -4540 4880 -4500 5200
rect -4900 4840 -4500 4880
rect -3888 5200 -3488 5240
rect -3888 4880 -3848 5200
rect -3528 4880 -3488 5200
rect -3888 4840 -3488 4880
rect -2876 5200 -2476 5240
rect -2876 4880 -2836 5200
rect -2516 4880 -2476 5200
rect -2876 4840 -2476 4880
rect -1864 5200 -1464 5240
rect -1864 4880 -1824 5200
rect -1504 4880 -1464 5200
rect -1864 4840 -1464 4880
rect -852 5200 -452 5240
rect -852 4880 -812 5200
rect -492 4880 -452 5200
rect -852 4840 -452 4880
rect 160 5200 560 5240
rect 160 4880 200 5200
rect 520 4880 560 5200
rect 160 4840 560 4880
rect 1172 5200 1572 5240
rect 1172 4880 1212 5200
rect 1532 4880 1572 5200
rect 1172 4840 1572 4880
rect 2184 5200 2584 5240
rect 2184 4880 2224 5200
rect 2544 4880 2584 5200
rect 2184 4840 2584 4880
rect 3196 5200 3596 5240
rect 3196 4880 3236 5200
rect 3556 4880 3596 5200
rect 3196 4840 3596 4880
rect 4208 5200 4608 5240
rect 4208 4880 4248 5200
rect 4568 4880 4608 5200
rect 4208 4840 4608 4880
rect 5220 5200 5620 5240
rect 5220 4880 5260 5200
rect 5580 4880 5620 5200
rect 5220 4840 5620 4880
rect 6232 5200 6632 5240
rect 6232 4880 6272 5200
rect 6592 4880 6632 5200
rect 6232 4840 6632 4880
rect 7244 5200 7644 5240
rect 7244 4880 7284 5200
rect 7604 4880 7644 5200
rect 7244 4840 7644 4880
rect 8256 5200 8656 5240
rect 8256 4880 8296 5200
rect 8616 4880 8656 5200
rect 8256 4840 8656 4880
rect 9268 5200 9668 5240
rect 9268 4880 9308 5200
rect 9628 4880 9668 5200
rect 9268 4840 9668 4880
rect 10280 5200 10680 5240
rect 10280 4880 10320 5200
rect 10640 4880 10680 5200
rect 10280 4840 10680 4880
rect 11292 5200 11692 5240
rect 11292 4880 11332 5200
rect 11652 4880 11692 5200
rect 11292 4840 11692 4880
rect 12304 5200 12704 5240
rect 12304 4880 12344 5200
rect 12664 4880 12704 5200
rect 12304 4840 12704 4880
rect 13316 5200 13716 5240
rect 13316 4880 13356 5200
rect 13676 4880 13716 5200
rect 13316 4840 13716 4880
rect 14328 5200 14728 5240
rect 14328 4880 14368 5200
rect 14688 4880 14728 5200
rect 14328 4840 14728 4880
rect 15340 5200 15740 5240
rect 15340 4880 15380 5200
rect 15700 4880 15740 5200
rect 15340 4840 15740 4880
rect 16352 5200 16752 5240
rect 16352 4880 16392 5200
rect 16712 4880 16752 5200
rect 16352 4840 16752 4880
rect -17044 4480 -16644 4520
rect -17044 4160 -17004 4480
rect -16684 4160 -16644 4480
rect -17044 4120 -16644 4160
rect -16032 4480 -15632 4520
rect -16032 4160 -15992 4480
rect -15672 4160 -15632 4480
rect -16032 4120 -15632 4160
rect -15020 4480 -14620 4520
rect -15020 4160 -14980 4480
rect -14660 4160 -14620 4480
rect -15020 4120 -14620 4160
rect -14008 4480 -13608 4520
rect -14008 4160 -13968 4480
rect -13648 4160 -13608 4480
rect -14008 4120 -13608 4160
rect -12996 4480 -12596 4520
rect -12996 4160 -12956 4480
rect -12636 4160 -12596 4480
rect -12996 4120 -12596 4160
rect -11984 4480 -11584 4520
rect -11984 4160 -11944 4480
rect -11624 4160 -11584 4480
rect -11984 4120 -11584 4160
rect -10972 4480 -10572 4520
rect -10972 4160 -10932 4480
rect -10612 4160 -10572 4480
rect -10972 4120 -10572 4160
rect -9960 4480 -9560 4520
rect -9960 4160 -9920 4480
rect -9600 4160 -9560 4480
rect -9960 4120 -9560 4160
rect -8948 4480 -8548 4520
rect -8948 4160 -8908 4480
rect -8588 4160 -8548 4480
rect -8948 4120 -8548 4160
rect -7936 4480 -7536 4520
rect -7936 4160 -7896 4480
rect -7576 4160 -7536 4480
rect -7936 4120 -7536 4160
rect -6924 4480 -6524 4520
rect -6924 4160 -6884 4480
rect -6564 4160 -6524 4480
rect -6924 4120 -6524 4160
rect -5912 4480 -5512 4520
rect -5912 4160 -5872 4480
rect -5552 4160 -5512 4480
rect -5912 4120 -5512 4160
rect -4900 4480 -4500 4520
rect -4900 4160 -4860 4480
rect -4540 4160 -4500 4480
rect -4900 4120 -4500 4160
rect -3888 4480 -3488 4520
rect -3888 4160 -3848 4480
rect -3528 4160 -3488 4480
rect -3888 4120 -3488 4160
rect -2876 4480 -2476 4520
rect -2876 4160 -2836 4480
rect -2516 4160 -2476 4480
rect -2876 4120 -2476 4160
rect -1864 4480 -1464 4520
rect -1864 4160 -1824 4480
rect -1504 4160 -1464 4480
rect -1864 4120 -1464 4160
rect -852 4480 -452 4520
rect -852 4160 -812 4480
rect -492 4160 -452 4480
rect -852 4120 -452 4160
rect 160 4480 560 4520
rect 160 4160 200 4480
rect 520 4160 560 4480
rect 160 4120 560 4160
rect 1172 4480 1572 4520
rect 1172 4160 1212 4480
rect 1532 4160 1572 4480
rect 1172 4120 1572 4160
rect 2184 4480 2584 4520
rect 2184 4160 2224 4480
rect 2544 4160 2584 4480
rect 2184 4120 2584 4160
rect 3196 4480 3596 4520
rect 3196 4160 3236 4480
rect 3556 4160 3596 4480
rect 3196 4120 3596 4160
rect 4208 4480 4608 4520
rect 4208 4160 4248 4480
rect 4568 4160 4608 4480
rect 4208 4120 4608 4160
rect 5220 4480 5620 4520
rect 5220 4160 5260 4480
rect 5580 4160 5620 4480
rect 5220 4120 5620 4160
rect 6232 4480 6632 4520
rect 6232 4160 6272 4480
rect 6592 4160 6632 4480
rect 6232 4120 6632 4160
rect 7244 4480 7644 4520
rect 7244 4160 7284 4480
rect 7604 4160 7644 4480
rect 7244 4120 7644 4160
rect 8256 4480 8656 4520
rect 8256 4160 8296 4480
rect 8616 4160 8656 4480
rect 8256 4120 8656 4160
rect 9268 4480 9668 4520
rect 9268 4160 9308 4480
rect 9628 4160 9668 4480
rect 9268 4120 9668 4160
rect 10280 4480 10680 4520
rect 10280 4160 10320 4480
rect 10640 4160 10680 4480
rect 10280 4120 10680 4160
rect 11292 4480 11692 4520
rect 11292 4160 11332 4480
rect 11652 4160 11692 4480
rect 11292 4120 11692 4160
rect 12304 4480 12704 4520
rect 12304 4160 12344 4480
rect 12664 4160 12704 4480
rect 12304 4120 12704 4160
rect 13316 4480 13716 4520
rect 13316 4160 13356 4480
rect 13676 4160 13716 4480
rect 13316 4120 13716 4160
rect 14328 4480 14728 4520
rect 14328 4160 14368 4480
rect 14688 4160 14728 4480
rect 14328 4120 14728 4160
rect 15340 4480 15740 4520
rect 15340 4160 15380 4480
rect 15700 4160 15740 4480
rect 15340 4120 15740 4160
rect 16352 4480 16752 4520
rect 16352 4160 16392 4480
rect 16712 4160 16752 4480
rect 16352 4120 16752 4160
rect -17044 3760 -16644 3800
rect -17044 3440 -17004 3760
rect -16684 3440 -16644 3760
rect -17044 3400 -16644 3440
rect -16032 3760 -15632 3800
rect -16032 3440 -15992 3760
rect -15672 3440 -15632 3760
rect -16032 3400 -15632 3440
rect -15020 3760 -14620 3800
rect -15020 3440 -14980 3760
rect -14660 3440 -14620 3760
rect -15020 3400 -14620 3440
rect -14008 3760 -13608 3800
rect -14008 3440 -13968 3760
rect -13648 3440 -13608 3760
rect -14008 3400 -13608 3440
rect -12996 3760 -12596 3800
rect -12996 3440 -12956 3760
rect -12636 3440 -12596 3760
rect -12996 3400 -12596 3440
rect -11984 3760 -11584 3800
rect -11984 3440 -11944 3760
rect -11624 3440 -11584 3760
rect -11984 3400 -11584 3440
rect -10972 3760 -10572 3800
rect -10972 3440 -10932 3760
rect -10612 3440 -10572 3760
rect -10972 3400 -10572 3440
rect -9960 3760 -9560 3800
rect -9960 3440 -9920 3760
rect -9600 3440 -9560 3760
rect -9960 3400 -9560 3440
rect -8948 3760 -8548 3800
rect -8948 3440 -8908 3760
rect -8588 3440 -8548 3760
rect -8948 3400 -8548 3440
rect -7936 3760 -7536 3800
rect -7936 3440 -7896 3760
rect -7576 3440 -7536 3760
rect -7936 3400 -7536 3440
rect -6924 3760 -6524 3800
rect -6924 3440 -6884 3760
rect -6564 3440 -6524 3760
rect -6924 3400 -6524 3440
rect -5912 3760 -5512 3800
rect -5912 3440 -5872 3760
rect -5552 3440 -5512 3760
rect -5912 3400 -5512 3440
rect -4900 3760 -4500 3800
rect -4900 3440 -4860 3760
rect -4540 3440 -4500 3760
rect -4900 3400 -4500 3440
rect -3888 3760 -3488 3800
rect -3888 3440 -3848 3760
rect -3528 3440 -3488 3760
rect -3888 3400 -3488 3440
rect -2876 3760 -2476 3800
rect -2876 3440 -2836 3760
rect -2516 3440 -2476 3760
rect -2876 3400 -2476 3440
rect -1864 3760 -1464 3800
rect -1864 3440 -1824 3760
rect -1504 3440 -1464 3760
rect -1864 3400 -1464 3440
rect -852 3760 -452 3800
rect -852 3440 -812 3760
rect -492 3440 -452 3760
rect -852 3400 -452 3440
rect 160 3760 560 3800
rect 160 3440 200 3760
rect 520 3440 560 3760
rect 160 3400 560 3440
rect 1172 3760 1572 3800
rect 1172 3440 1212 3760
rect 1532 3440 1572 3760
rect 1172 3400 1572 3440
rect 2184 3760 2584 3800
rect 2184 3440 2224 3760
rect 2544 3440 2584 3760
rect 2184 3400 2584 3440
rect 3196 3760 3596 3800
rect 3196 3440 3236 3760
rect 3556 3440 3596 3760
rect 3196 3400 3596 3440
rect 4208 3760 4608 3800
rect 4208 3440 4248 3760
rect 4568 3440 4608 3760
rect 4208 3400 4608 3440
rect 5220 3760 5620 3800
rect 5220 3440 5260 3760
rect 5580 3440 5620 3760
rect 5220 3400 5620 3440
rect 6232 3760 6632 3800
rect 6232 3440 6272 3760
rect 6592 3440 6632 3760
rect 6232 3400 6632 3440
rect 7244 3760 7644 3800
rect 7244 3440 7284 3760
rect 7604 3440 7644 3760
rect 7244 3400 7644 3440
rect 8256 3760 8656 3800
rect 8256 3440 8296 3760
rect 8616 3440 8656 3760
rect 8256 3400 8656 3440
rect 9268 3760 9668 3800
rect 9268 3440 9308 3760
rect 9628 3440 9668 3760
rect 9268 3400 9668 3440
rect 10280 3760 10680 3800
rect 10280 3440 10320 3760
rect 10640 3440 10680 3760
rect 10280 3400 10680 3440
rect 11292 3760 11692 3800
rect 11292 3440 11332 3760
rect 11652 3440 11692 3760
rect 11292 3400 11692 3440
rect 12304 3760 12704 3800
rect 12304 3440 12344 3760
rect 12664 3440 12704 3760
rect 12304 3400 12704 3440
rect 13316 3760 13716 3800
rect 13316 3440 13356 3760
rect 13676 3440 13716 3760
rect 13316 3400 13716 3440
rect 14328 3760 14728 3800
rect 14328 3440 14368 3760
rect 14688 3440 14728 3760
rect 14328 3400 14728 3440
rect 15340 3760 15740 3800
rect 15340 3440 15380 3760
rect 15700 3440 15740 3760
rect 15340 3400 15740 3440
rect 16352 3760 16752 3800
rect 16352 3440 16392 3760
rect 16712 3440 16752 3760
rect 16352 3400 16752 3440
rect -17044 3040 -16644 3080
rect -17044 2720 -17004 3040
rect -16684 2720 -16644 3040
rect -17044 2680 -16644 2720
rect -16032 3040 -15632 3080
rect -16032 2720 -15992 3040
rect -15672 2720 -15632 3040
rect -16032 2680 -15632 2720
rect -15020 3040 -14620 3080
rect -15020 2720 -14980 3040
rect -14660 2720 -14620 3040
rect -15020 2680 -14620 2720
rect -14008 3040 -13608 3080
rect -14008 2720 -13968 3040
rect -13648 2720 -13608 3040
rect -14008 2680 -13608 2720
rect -12996 3040 -12596 3080
rect -12996 2720 -12956 3040
rect -12636 2720 -12596 3040
rect -12996 2680 -12596 2720
rect -11984 3040 -11584 3080
rect -11984 2720 -11944 3040
rect -11624 2720 -11584 3040
rect -11984 2680 -11584 2720
rect -10972 3040 -10572 3080
rect -10972 2720 -10932 3040
rect -10612 2720 -10572 3040
rect -10972 2680 -10572 2720
rect -9960 3040 -9560 3080
rect -9960 2720 -9920 3040
rect -9600 2720 -9560 3040
rect -9960 2680 -9560 2720
rect -8948 3040 -8548 3080
rect -8948 2720 -8908 3040
rect -8588 2720 -8548 3040
rect -8948 2680 -8548 2720
rect -7936 3040 -7536 3080
rect -7936 2720 -7896 3040
rect -7576 2720 -7536 3040
rect -7936 2680 -7536 2720
rect -6924 3040 -6524 3080
rect -6924 2720 -6884 3040
rect -6564 2720 -6524 3040
rect -6924 2680 -6524 2720
rect -5912 3040 -5512 3080
rect -5912 2720 -5872 3040
rect -5552 2720 -5512 3040
rect -5912 2680 -5512 2720
rect -4900 3040 -4500 3080
rect -4900 2720 -4860 3040
rect -4540 2720 -4500 3040
rect -4900 2680 -4500 2720
rect -3888 3040 -3488 3080
rect -3888 2720 -3848 3040
rect -3528 2720 -3488 3040
rect -3888 2680 -3488 2720
rect -2876 3040 -2476 3080
rect -2876 2720 -2836 3040
rect -2516 2720 -2476 3040
rect -2876 2680 -2476 2720
rect -1864 3040 -1464 3080
rect -1864 2720 -1824 3040
rect -1504 2720 -1464 3040
rect -1864 2680 -1464 2720
rect -852 3040 -452 3080
rect -852 2720 -812 3040
rect -492 2720 -452 3040
rect -852 2680 -452 2720
rect 160 3040 560 3080
rect 160 2720 200 3040
rect 520 2720 560 3040
rect 160 2680 560 2720
rect 1172 3040 1572 3080
rect 1172 2720 1212 3040
rect 1532 2720 1572 3040
rect 1172 2680 1572 2720
rect 2184 3040 2584 3080
rect 2184 2720 2224 3040
rect 2544 2720 2584 3040
rect 2184 2680 2584 2720
rect 3196 3040 3596 3080
rect 3196 2720 3236 3040
rect 3556 2720 3596 3040
rect 3196 2680 3596 2720
rect 4208 3040 4608 3080
rect 4208 2720 4248 3040
rect 4568 2720 4608 3040
rect 4208 2680 4608 2720
rect 5220 3040 5620 3080
rect 5220 2720 5260 3040
rect 5580 2720 5620 3040
rect 5220 2680 5620 2720
rect 6232 3040 6632 3080
rect 6232 2720 6272 3040
rect 6592 2720 6632 3040
rect 6232 2680 6632 2720
rect 7244 3040 7644 3080
rect 7244 2720 7284 3040
rect 7604 2720 7644 3040
rect 7244 2680 7644 2720
rect 8256 3040 8656 3080
rect 8256 2720 8296 3040
rect 8616 2720 8656 3040
rect 8256 2680 8656 2720
rect 9268 3040 9668 3080
rect 9268 2720 9308 3040
rect 9628 2720 9668 3040
rect 9268 2680 9668 2720
rect 10280 3040 10680 3080
rect 10280 2720 10320 3040
rect 10640 2720 10680 3040
rect 10280 2680 10680 2720
rect 11292 3040 11692 3080
rect 11292 2720 11332 3040
rect 11652 2720 11692 3040
rect 11292 2680 11692 2720
rect 12304 3040 12704 3080
rect 12304 2720 12344 3040
rect 12664 2720 12704 3040
rect 12304 2680 12704 2720
rect 13316 3040 13716 3080
rect 13316 2720 13356 3040
rect 13676 2720 13716 3040
rect 13316 2680 13716 2720
rect 14328 3040 14728 3080
rect 14328 2720 14368 3040
rect 14688 2720 14728 3040
rect 14328 2680 14728 2720
rect 15340 3040 15740 3080
rect 15340 2720 15380 3040
rect 15700 2720 15740 3040
rect 15340 2680 15740 2720
rect 16352 3040 16752 3080
rect 16352 2720 16392 3040
rect 16712 2720 16752 3040
rect 16352 2680 16752 2720
rect -17044 2320 -16644 2360
rect -17044 2000 -17004 2320
rect -16684 2000 -16644 2320
rect -17044 1960 -16644 2000
rect -16032 2320 -15632 2360
rect -16032 2000 -15992 2320
rect -15672 2000 -15632 2320
rect -16032 1960 -15632 2000
rect -15020 2320 -14620 2360
rect -15020 2000 -14980 2320
rect -14660 2000 -14620 2320
rect -15020 1960 -14620 2000
rect -14008 2320 -13608 2360
rect -14008 2000 -13968 2320
rect -13648 2000 -13608 2320
rect -14008 1960 -13608 2000
rect -12996 2320 -12596 2360
rect -12996 2000 -12956 2320
rect -12636 2000 -12596 2320
rect -12996 1960 -12596 2000
rect -11984 2320 -11584 2360
rect -11984 2000 -11944 2320
rect -11624 2000 -11584 2320
rect -11984 1960 -11584 2000
rect -10972 2320 -10572 2360
rect -10972 2000 -10932 2320
rect -10612 2000 -10572 2320
rect -10972 1960 -10572 2000
rect -9960 2320 -9560 2360
rect -9960 2000 -9920 2320
rect -9600 2000 -9560 2320
rect -9960 1960 -9560 2000
rect -8948 2320 -8548 2360
rect -8948 2000 -8908 2320
rect -8588 2000 -8548 2320
rect -8948 1960 -8548 2000
rect -7936 2320 -7536 2360
rect -7936 2000 -7896 2320
rect -7576 2000 -7536 2320
rect -7936 1960 -7536 2000
rect -6924 2320 -6524 2360
rect -6924 2000 -6884 2320
rect -6564 2000 -6524 2320
rect -6924 1960 -6524 2000
rect -5912 2320 -5512 2360
rect -5912 2000 -5872 2320
rect -5552 2000 -5512 2320
rect -5912 1960 -5512 2000
rect -4900 2320 -4500 2360
rect -4900 2000 -4860 2320
rect -4540 2000 -4500 2320
rect -4900 1960 -4500 2000
rect -3888 2320 -3488 2360
rect -3888 2000 -3848 2320
rect -3528 2000 -3488 2320
rect -3888 1960 -3488 2000
rect -2876 2320 -2476 2360
rect -2876 2000 -2836 2320
rect -2516 2000 -2476 2320
rect -2876 1960 -2476 2000
rect -1864 2320 -1464 2360
rect -1864 2000 -1824 2320
rect -1504 2000 -1464 2320
rect -1864 1960 -1464 2000
rect -852 2320 -452 2360
rect -852 2000 -812 2320
rect -492 2000 -452 2320
rect -852 1960 -452 2000
rect 160 2320 560 2360
rect 160 2000 200 2320
rect 520 2000 560 2320
rect 160 1960 560 2000
rect 1172 2320 1572 2360
rect 1172 2000 1212 2320
rect 1532 2000 1572 2320
rect 1172 1960 1572 2000
rect 2184 2320 2584 2360
rect 2184 2000 2224 2320
rect 2544 2000 2584 2320
rect 2184 1960 2584 2000
rect 3196 2320 3596 2360
rect 3196 2000 3236 2320
rect 3556 2000 3596 2320
rect 3196 1960 3596 2000
rect 4208 2320 4608 2360
rect 4208 2000 4248 2320
rect 4568 2000 4608 2320
rect 4208 1960 4608 2000
rect 5220 2320 5620 2360
rect 5220 2000 5260 2320
rect 5580 2000 5620 2320
rect 5220 1960 5620 2000
rect 6232 2320 6632 2360
rect 6232 2000 6272 2320
rect 6592 2000 6632 2320
rect 6232 1960 6632 2000
rect 7244 2320 7644 2360
rect 7244 2000 7284 2320
rect 7604 2000 7644 2320
rect 7244 1960 7644 2000
rect 8256 2320 8656 2360
rect 8256 2000 8296 2320
rect 8616 2000 8656 2320
rect 8256 1960 8656 2000
rect 9268 2320 9668 2360
rect 9268 2000 9308 2320
rect 9628 2000 9668 2320
rect 9268 1960 9668 2000
rect 10280 2320 10680 2360
rect 10280 2000 10320 2320
rect 10640 2000 10680 2320
rect 10280 1960 10680 2000
rect 11292 2320 11692 2360
rect 11292 2000 11332 2320
rect 11652 2000 11692 2320
rect 11292 1960 11692 2000
rect 12304 2320 12704 2360
rect 12304 2000 12344 2320
rect 12664 2000 12704 2320
rect 12304 1960 12704 2000
rect 13316 2320 13716 2360
rect 13316 2000 13356 2320
rect 13676 2000 13716 2320
rect 13316 1960 13716 2000
rect 14328 2320 14728 2360
rect 14328 2000 14368 2320
rect 14688 2000 14728 2320
rect 14328 1960 14728 2000
rect 15340 2320 15740 2360
rect 15340 2000 15380 2320
rect 15700 2000 15740 2320
rect 15340 1960 15740 2000
rect 16352 2320 16752 2360
rect 16352 2000 16392 2320
rect 16712 2000 16752 2320
rect 16352 1960 16752 2000
rect -17044 1600 -16644 1640
rect -17044 1280 -17004 1600
rect -16684 1280 -16644 1600
rect -17044 1240 -16644 1280
rect -16032 1600 -15632 1640
rect -16032 1280 -15992 1600
rect -15672 1280 -15632 1600
rect -16032 1240 -15632 1280
rect -15020 1600 -14620 1640
rect -15020 1280 -14980 1600
rect -14660 1280 -14620 1600
rect -15020 1240 -14620 1280
rect -14008 1600 -13608 1640
rect -14008 1280 -13968 1600
rect -13648 1280 -13608 1600
rect -14008 1240 -13608 1280
rect -12996 1600 -12596 1640
rect -12996 1280 -12956 1600
rect -12636 1280 -12596 1600
rect -12996 1240 -12596 1280
rect -11984 1600 -11584 1640
rect -11984 1280 -11944 1600
rect -11624 1280 -11584 1600
rect -11984 1240 -11584 1280
rect -10972 1600 -10572 1640
rect -10972 1280 -10932 1600
rect -10612 1280 -10572 1600
rect -10972 1240 -10572 1280
rect -9960 1600 -9560 1640
rect -9960 1280 -9920 1600
rect -9600 1280 -9560 1600
rect -9960 1240 -9560 1280
rect -8948 1600 -8548 1640
rect -8948 1280 -8908 1600
rect -8588 1280 -8548 1600
rect -8948 1240 -8548 1280
rect -7936 1600 -7536 1640
rect -7936 1280 -7896 1600
rect -7576 1280 -7536 1600
rect -7936 1240 -7536 1280
rect -6924 1600 -6524 1640
rect -6924 1280 -6884 1600
rect -6564 1280 -6524 1600
rect -6924 1240 -6524 1280
rect -5912 1600 -5512 1640
rect -5912 1280 -5872 1600
rect -5552 1280 -5512 1600
rect -5912 1240 -5512 1280
rect -4900 1600 -4500 1640
rect -4900 1280 -4860 1600
rect -4540 1280 -4500 1600
rect -4900 1240 -4500 1280
rect -3888 1600 -3488 1640
rect -3888 1280 -3848 1600
rect -3528 1280 -3488 1600
rect -3888 1240 -3488 1280
rect -2876 1600 -2476 1640
rect -2876 1280 -2836 1600
rect -2516 1280 -2476 1600
rect -2876 1240 -2476 1280
rect -1864 1600 -1464 1640
rect -1864 1280 -1824 1600
rect -1504 1280 -1464 1600
rect -1864 1240 -1464 1280
rect -852 1600 -452 1640
rect -852 1280 -812 1600
rect -492 1280 -452 1600
rect -852 1240 -452 1280
rect 160 1600 560 1640
rect 160 1280 200 1600
rect 520 1280 560 1600
rect 160 1240 560 1280
rect 1172 1600 1572 1640
rect 1172 1280 1212 1600
rect 1532 1280 1572 1600
rect 1172 1240 1572 1280
rect 2184 1600 2584 1640
rect 2184 1280 2224 1600
rect 2544 1280 2584 1600
rect 2184 1240 2584 1280
rect 3196 1600 3596 1640
rect 3196 1280 3236 1600
rect 3556 1280 3596 1600
rect 3196 1240 3596 1280
rect 4208 1600 4608 1640
rect 4208 1280 4248 1600
rect 4568 1280 4608 1600
rect 4208 1240 4608 1280
rect 5220 1600 5620 1640
rect 5220 1280 5260 1600
rect 5580 1280 5620 1600
rect 5220 1240 5620 1280
rect 6232 1600 6632 1640
rect 6232 1280 6272 1600
rect 6592 1280 6632 1600
rect 6232 1240 6632 1280
rect 7244 1600 7644 1640
rect 7244 1280 7284 1600
rect 7604 1280 7644 1600
rect 7244 1240 7644 1280
rect 8256 1600 8656 1640
rect 8256 1280 8296 1600
rect 8616 1280 8656 1600
rect 8256 1240 8656 1280
rect 9268 1600 9668 1640
rect 9268 1280 9308 1600
rect 9628 1280 9668 1600
rect 9268 1240 9668 1280
rect 10280 1600 10680 1640
rect 10280 1280 10320 1600
rect 10640 1280 10680 1600
rect 10280 1240 10680 1280
rect 11292 1600 11692 1640
rect 11292 1280 11332 1600
rect 11652 1280 11692 1600
rect 11292 1240 11692 1280
rect 12304 1600 12704 1640
rect 12304 1280 12344 1600
rect 12664 1280 12704 1600
rect 12304 1240 12704 1280
rect 13316 1600 13716 1640
rect 13316 1280 13356 1600
rect 13676 1280 13716 1600
rect 13316 1240 13716 1280
rect 14328 1600 14728 1640
rect 14328 1280 14368 1600
rect 14688 1280 14728 1600
rect 14328 1240 14728 1280
rect 15340 1600 15740 1640
rect 15340 1280 15380 1600
rect 15700 1280 15740 1600
rect 15340 1240 15740 1280
rect 16352 1600 16752 1640
rect 16352 1280 16392 1600
rect 16712 1280 16752 1600
rect 16352 1240 16752 1280
rect -17044 880 -16644 920
rect -17044 560 -17004 880
rect -16684 560 -16644 880
rect -17044 520 -16644 560
rect -16032 880 -15632 920
rect -16032 560 -15992 880
rect -15672 560 -15632 880
rect -16032 520 -15632 560
rect -15020 880 -14620 920
rect -15020 560 -14980 880
rect -14660 560 -14620 880
rect -15020 520 -14620 560
rect -14008 880 -13608 920
rect -14008 560 -13968 880
rect -13648 560 -13608 880
rect -14008 520 -13608 560
rect -12996 880 -12596 920
rect -12996 560 -12956 880
rect -12636 560 -12596 880
rect -12996 520 -12596 560
rect -11984 880 -11584 920
rect -11984 560 -11944 880
rect -11624 560 -11584 880
rect -11984 520 -11584 560
rect -10972 880 -10572 920
rect -10972 560 -10932 880
rect -10612 560 -10572 880
rect -10972 520 -10572 560
rect -9960 880 -9560 920
rect -9960 560 -9920 880
rect -9600 560 -9560 880
rect -9960 520 -9560 560
rect -8948 880 -8548 920
rect -8948 560 -8908 880
rect -8588 560 -8548 880
rect -8948 520 -8548 560
rect -7936 880 -7536 920
rect -7936 560 -7896 880
rect -7576 560 -7536 880
rect -7936 520 -7536 560
rect -6924 880 -6524 920
rect -6924 560 -6884 880
rect -6564 560 -6524 880
rect -6924 520 -6524 560
rect -5912 880 -5512 920
rect -5912 560 -5872 880
rect -5552 560 -5512 880
rect -5912 520 -5512 560
rect -4900 880 -4500 920
rect -4900 560 -4860 880
rect -4540 560 -4500 880
rect -4900 520 -4500 560
rect -3888 880 -3488 920
rect -3888 560 -3848 880
rect -3528 560 -3488 880
rect -3888 520 -3488 560
rect -2876 880 -2476 920
rect -2876 560 -2836 880
rect -2516 560 -2476 880
rect -2876 520 -2476 560
rect -1864 880 -1464 920
rect -1864 560 -1824 880
rect -1504 560 -1464 880
rect -1864 520 -1464 560
rect -852 880 -452 920
rect -852 560 -812 880
rect -492 560 -452 880
rect -852 520 -452 560
rect 160 880 560 920
rect 160 560 200 880
rect 520 560 560 880
rect 160 520 560 560
rect 1172 880 1572 920
rect 1172 560 1212 880
rect 1532 560 1572 880
rect 1172 520 1572 560
rect 2184 880 2584 920
rect 2184 560 2224 880
rect 2544 560 2584 880
rect 2184 520 2584 560
rect 3196 880 3596 920
rect 3196 560 3236 880
rect 3556 560 3596 880
rect 3196 520 3596 560
rect 4208 880 4608 920
rect 4208 560 4248 880
rect 4568 560 4608 880
rect 4208 520 4608 560
rect 5220 880 5620 920
rect 5220 560 5260 880
rect 5580 560 5620 880
rect 5220 520 5620 560
rect 6232 880 6632 920
rect 6232 560 6272 880
rect 6592 560 6632 880
rect 6232 520 6632 560
rect 7244 880 7644 920
rect 7244 560 7284 880
rect 7604 560 7644 880
rect 7244 520 7644 560
rect 8256 880 8656 920
rect 8256 560 8296 880
rect 8616 560 8656 880
rect 8256 520 8656 560
rect 9268 880 9668 920
rect 9268 560 9308 880
rect 9628 560 9668 880
rect 9268 520 9668 560
rect 10280 880 10680 920
rect 10280 560 10320 880
rect 10640 560 10680 880
rect 10280 520 10680 560
rect 11292 880 11692 920
rect 11292 560 11332 880
rect 11652 560 11692 880
rect 11292 520 11692 560
rect 12304 880 12704 920
rect 12304 560 12344 880
rect 12664 560 12704 880
rect 12304 520 12704 560
rect 13316 880 13716 920
rect 13316 560 13356 880
rect 13676 560 13716 880
rect 13316 520 13716 560
rect 14328 880 14728 920
rect 14328 560 14368 880
rect 14688 560 14728 880
rect 14328 520 14728 560
rect 15340 880 15740 920
rect 15340 560 15380 880
rect 15700 560 15740 880
rect 15340 520 15740 560
rect 16352 880 16752 920
rect 16352 560 16392 880
rect 16712 560 16752 880
rect 16352 520 16752 560
rect -17044 160 -16644 200
rect -17044 -160 -17004 160
rect -16684 -160 -16644 160
rect -17044 -200 -16644 -160
rect -16032 160 -15632 200
rect -16032 -160 -15992 160
rect -15672 -160 -15632 160
rect -16032 -200 -15632 -160
rect -15020 160 -14620 200
rect -15020 -160 -14980 160
rect -14660 -160 -14620 160
rect -15020 -200 -14620 -160
rect -14008 160 -13608 200
rect -14008 -160 -13968 160
rect -13648 -160 -13608 160
rect -14008 -200 -13608 -160
rect -12996 160 -12596 200
rect -12996 -160 -12956 160
rect -12636 -160 -12596 160
rect -12996 -200 -12596 -160
rect -11984 160 -11584 200
rect -11984 -160 -11944 160
rect -11624 -160 -11584 160
rect -11984 -200 -11584 -160
rect -10972 160 -10572 200
rect -10972 -160 -10932 160
rect -10612 -160 -10572 160
rect -10972 -200 -10572 -160
rect -9960 160 -9560 200
rect -9960 -160 -9920 160
rect -9600 -160 -9560 160
rect -9960 -200 -9560 -160
rect -8948 160 -8548 200
rect -8948 -160 -8908 160
rect -8588 -160 -8548 160
rect -8948 -200 -8548 -160
rect -7936 160 -7536 200
rect -7936 -160 -7896 160
rect -7576 -160 -7536 160
rect -7936 -200 -7536 -160
rect -6924 160 -6524 200
rect -6924 -160 -6884 160
rect -6564 -160 -6524 160
rect -6924 -200 -6524 -160
rect -5912 160 -5512 200
rect -5912 -160 -5872 160
rect -5552 -160 -5512 160
rect -5912 -200 -5512 -160
rect -4900 160 -4500 200
rect -4900 -160 -4860 160
rect -4540 -160 -4500 160
rect -4900 -200 -4500 -160
rect -3888 160 -3488 200
rect -3888 -160 -3848 160
rect -3528 -160 -3488 160
rect -3888 -200 -3488 -160
rect -2876 160 -2476 200
rect -2876 -160 -2836 160
rect -2516 -160 -2476 160
rect -2876 -200 -2476 -160
rect -1864 160 -1464 200
rect -1864 -160 -1824 160
rect -1504 -160 -1464 160
rect -1864 -200 -1464 -160
rect -852 160 -452 200
rect -852 -160 -812 160
rect -492 -160 -452 160
rect -852 -200 -452 -160
rect 160 160 560 200
rect 160 -160 200 160
rect 520 -160 560 160
rect 160 -200 560 -160
rect 1172 160 1572 200
rect 1172 -160 1212 160
rect 1532 -160 1572 160
rect 1172 -200 1572 -160
rect 2184 160 2584 200
rect 2184 -160 2224 160
rect 2544 -160 2584 160
rect 2184 -200 2584 -160
rect 3196 160 3596 200
rect 3196 -160 3236 160
rect 3556 -160 3596 160
rect 3196 -200 3596 -160
rect 4208 160 4608 200
rect 4208 -160 4248 160
rect 4568 -160 4608 160
rect 4208 -200 4608 -160
rect 5220 160 5620 200
rect 5220 -160 5260 160
rect 5580 -160 5620 160
rect 5220 -200 5620 -160
rect 6232 160 6632 200
rect 6232 -160 6272 160
rect 6592 -160 6632 160
rect 6232 -200 6632 -160
rect 7244 160 7644 200
rect 7244 -160 7284 160
rect 7604 -160 7644 160
rect 7244 -200 7644 -160
rect 8256 160 8656 200
rect 8256 -160 8296 160
rect 8616 -160 8656 160
rect 8256 -200 8656 -160
rect 9268 160 9668 200
rect 9268 -160 9308 160
rect 9628 -160 9668 160
rect 9268 -200 9668 -160
rect 10280 160 10680 200
rect 10280 -160 10320 160
rect 10640 -160 10680 160
rect 10280 -200 10680 -160
rect 11292 160 11692 200
rect 11292 -160 11332 160
rect 11652 -160 11692 160
rect 11292 -200 11692 -160
rect 12304 160 12704 200
rect 12304 -160 12344 160
rect 12664 -160 12704 160
rect 12304 -200 12704 -160
rect 13316 160 13716 200
rect 13316 -160 13356 160
rect 13676 -160 13716 160
rect 13316 -200 13716 -160
rect 14328 160 14728 200
rect 14328 -160 14368 160
rect 14688 -160 14728 160
rect 14328 -200 14728 -160
rect 15340 160 15740 200
rect 15340 -160 15380 160
rect 15700 -160 15740 160
rect 15340 -200 15740 -160
rect 16352 160 16752 200
rect 16352 -160 16392 160
rect 16712 -160 16752 160
rect 16352 -200 16752 -160
rect -17044 -560 -16644 -520
rect -17044 -880 -17004 -560
rect -16684 -880 -16644 -560
rect -17044 -920 -16644 -880
rect -16032 -560 -15632 -520
rect -16032 -880 -15992 -560
rect -15672 -880 -15632 -560
rect -16032 -920 -15632 -880
rect -15020 -560 -14620 -520
rect -15020 -880 -14980 -560
rect -14660 -880 -14620 -560
rect -15020 -920 -14620 -880
rect -14008 -560 -13608 -520
rect -14008 -880 -13968 -560
rect -13648 -880 -13608 -560
rect -14008 -920 -13608 -880
rect -12996 -560 -12596 -520
rect -12996 -880 -12956 -560
rect -12636 -880 -12596 -560
rect -12996 -920 -12596 -880
rect -11984 -560 -11584 -520
rect -11984 -880 -11944 -560
rect -11624 -880 -11584 -560
rect -11984 -920 -11584 -880
rect -10972 -560 -10572 -520
rect -10972 -880 -10932 -560
rect -10612 -880 -10572 -560
rect -10972 -920 -10572 -880
rect -9960 -560 -9560 -520
rect -9960 -880 -9920 -560
rect -9600 -880 -9560 -560
rect -9960 -920 -9560 -880
rect -8948 -560 -8548 -520
rect -8948 -880 -8908 -560
rect -8588 -880 -8548 -560
rect -8948 -920 -8548 -880
rect -7936 -560 -7536 -520
rect -7936 -880 -7896 -560
rect -7576 -880 -7536 -560
rect -7936 -920 -7536 -880
rect -6924 -560 -6524 -520
rect -6924 -880 -6884 -560
rect -6564 -880 -6524 -560
rect -6924 -920 -6524 -880
rect -5912 -560 -5512 -520
rect -5912 -880 -5872 -560
rect -5552 -880 -5512 -560
rect -5912 -920 -5512 -880
rect -4900 -560 -4500 -520
rect -4900 -880 -4860 -560
rect -4540 -880 -4500 -560
rect -4900 -920 -4500 -880
rect -3888 -560 -3488 -520
rect -3888 -880 -3848 -560
rect -3528 -880 -3488 -560
rect -3888 -920 -3488 -880
rect -2876 -560 -2476 -520
rect -2876 -880 -2836 -560
rect -2516 -880 -2476 -560
rect -2876 -920 -2476 -880
rect -1864 -560 -1464 -520
rect -1864 -880 -1824 -560
rect -1504 -880 -1464 -560
rect -1864 -920 -1464 -880
rect -852 -560 -452 -520
rect -852 -880 -812 -560
rect -492 -880 -452 -560
rect -852 -920 -452 -880
rect 160 -560 560 -520
rect 160 -880 200 -560
rect 520 -880 560 -560
rect 160 -920 560 -880
rect 1172 -560 1572 -520
rect 1172 -880 1212 -560
rect 1532 -880 1572 -560
rect 1172 -920 1572 -880
rect 2184 -560 2584 -520
rect 2184 -880 2224 -560
rect 2544 -880 2584 -560
rect 2184 -920 2584 -880
rect 3196 -560 3596 -520
rect 3196 -880 3236 -560
rect 3556 -880 3596 -560
rect 3196 -920 3596 -880
rect 4208 -560 4608 -520
rect 4208 -880 4248 -560
rect 4568 -880 4608 -560
rect 4208 -920 4608 -880
rect 5220 -560 5620 -520
rect 5220 -880 5260 -560
rect 5580 -880 5620 -560
rect 5220 -920 5620 -880
rect 6232 -560 6632 -520
rect 6232 -880 6272 -560
rect 6592 -880 6632 -560
rect 6232 -920 6632 -880
rect 7244 -560 7644 -520
rect 7244 -880 7284 -560
rect 7604 -880 7644 -560
rect 7244 -920 7644 -880
rect 8256 -560 8656 -520
rect 8256 -880 8296 -560
rect 8616 -880 8656 -560
rect 8256 -920 8656 -880
rect 9268 -560 9668 -520
rect 9268 -880 9308 -560
rect 9628 -880 9668 -560
rect 9268 -920 9668 -880
rect 10280 -560 10680 -520
rect 10280 -880 10320 -560
rect 10640 -880 10680 -560
rect 10280 -920 10680 -880
rect 11292 -560 11692 -520
rect 11292 -880 11332 -560
rect 11652 -880 11692 -560
rect 11292 -920 11692 -880
rect 12304 -560 12704 -520
rect 12304 -880 12344 -560
rect 12664 -880 12704 -560
rect 12304 -920 12704 -880
rect 13316 -560 13716 -520
rect 13316 -880 13356 -560
rect 13676 -880 13716 -560
rect 13316 -920 13716 -880
rect 14328 -560 14728 -520
rect 14328 -880 14368 -560
rect 14688 -880 14728 -560
rect 14328 -920 14728 -880
rect 15340 -560 15740 -520
rect 15340 -880 15380 -560
rect 15700 -880 15740 -560
rect 15340 -920 15740 -880
rect 16352 -560 16752 -520
rect 16352 -880 16392 -560
rect 16712 -880 16752 -560
rect 16352 -920 16752 -880
rect -17044 -1280 -16644 -1240
rect -17044 -1600 -17004 -1280
rect -16684 -1600 -16644 -1280
rect -17044 -1640 -16644 -1600
rect -16032 -1280 -15632 -1240
rect -16032 -1600 -15992 -1280
rect -15672 -1600 -15632 -1280
rect -16032 -1640 -15632 -1600
rect -15020 -1280 -14620 -1240
rect -15020 -1600 -14980 -1280
rect -14660 -1600 -14620 -1280
rect -15020 -1640 -14620 -1600
rect -14008 -1280 -13608 -1240
rect -14008 -1600 -13968 -1280
rect -13648 -1600 -13608 -1280
rect -14008 -1640 -13608 -1600
rect -12996 -1280 -12596 -1240
rect -12996 -1600 -12956 -1280
rect -12636 -1600 -12596 -1280
rect -12996 -1640 -12596 -1600
rect -11984 -1280 -11584 -1240
rect -11984 -1600 -11944 -1280
rect -11624 -1600 -11584 -1280
rect -11984 -1640 -11584 -1600
rect -10972 -1280 -10572 -1240
rect -10972 -1600 -10932 -1280
rect -10612 -1600 -10572 -1280
rect -10972 -1640 -10572 -1600
rect -9960 -1280 -9560 -1240
rect -9960 -1600 -9920 -1280
rect -9600 -1600 -9560 -1280
rect -9960 -1640 -9560 -1600
rect -8948 -1280 -8548 -1240
rect -8948 -1600 -8908 -1280
rect -8588 -1600 -8548 -1280
rect -8948 -1640 -8548 -1600
rect -7936 -1280 -7536 -1240
rect -7936 -1600 -7896 -1280
rect -7576 -1600 -7536 -1280
rect -7936 -1640 -7536 -1600
rect -6924 -1280 -6524 -1240
rect -6924 -1600 -6884 -1280
rect -6564 -1600 -6524 -1280
rect -6924 -1640 -6524 -1600
rect -5912 -1280 -5512 -1240
rect -5912 -1600 -5872 -1280
rect -5552 -1600 -5512 -1280
rect -5912 -1640 -5512 -1600
rect -4900 -1280 -4500 -1240
rect -4900 -1600 -4860 -1280
rect -4540 -1600 -4500 -1280
rect -4900 -1640 -4500 -1600
rect -3888 -1280 -3488 -1240
rect -3888 -1600 -3848 -1280
rect -3528 -1600 -3488 -1280
rect -3888 -1640 -3488 -1600
rect -2876 -1280 -2476 -1240
rect -2876 -1600 -2836 -1280
rect -2516 -1600 -2476 -1280
rect -2876 -1640 -2476 -1600
rect -1864 -1280 -1464 -1240
rect -1864 -1600 -1824 -1280
rect -1504 -1600 -1464 -1280
rect -1864 -1640 -1464 -1600
rect -852 -1280 -452 -1240
rect -852 -1600 -812 -1280
rect -492 -1600 -452 -1280
rect -852 -1640 -452 -1600
rect 160 -1280 560 -1240
rect 160 -1600 200 -1280
rect 520 -1600 560 -1280
rect 160 -1640 560 -1600
rect 1172 -1280 1572 -1240
rect 1172 -1600 1212 -1280
rect 1532 -1600 1572 -1280
rect 1172 -1640 1572 -1600
rect 2184 -1280 2584 -1240
rect 2184 -1600 2224 -1280
rect 2544 -1600 2584 -1280
rect 2184 -1640 2584 -1600
rect 3196 -1280 3596 -1240
rect 3196 -1600 3236 -1280
rect 3556 -1600 3596 -1280
rect 3196 -1640 3596 -1600
rect 4208 -1280 4608 -1240
rect 4208 -1600 4248 -1280
rect 4568 -1600 4608 -1280
rect 4208 -1640 4608 -1600
rect 5220 -1280 5620 -1240
rect 5220 -1600 5260 -1280
rect 5580 -1600 5620 -1280
rect 5220 -1640 5620 -1600
rect 6232 -1280 6632 -1240
rect 6232 -1600 6272 -1280
rect 6592 -1600 6632 -1280
rect 6232 -1640 6632 -1600
rect 7244 -1280 7644 -1240
rect 7244 -1600 7284 -1280
rect 7604 -1600 7644 -1280
rect 7244 -1640 7644 -1600
rect 8256 -1280 8656 -1240
rect 8256 -1600 8296 -1280
rect 8616 -1600 8656 -1280
rect 8256 -1640 8656 -1600
rect 9268 -1280 9668 -1240
rect 9268 -1600 9308 -1280
rect 9628 -1600 9668 -1280
rect 9268 -1640 9668 -1600
rect 10280 -1280 10680 -1240
rect 10280 -1600 10320 -1280
rect 10640 -1600 10680 -1280
rect 10280 -1640 10680 -1600
rect 11292 -1280 11692 -1240
rect 11292 -1600 11332 -1280
rect 11652 -1600 11692 -1280
rect 11292 -1640 11692 -1600
rect 12304 -1280 12704 -1240
rect 12304 -1600 12344 -1280
rect 12664 -1600 12704 -1280
rect 12304 -1640 12704 -1600
rect 13316 -1280 13716 -1240
rect 13316 -1600 13356 -1280
rect 13676 -1600 13716 -1280
rect 13316 -1640 13716 -1600
rect 14328 -1280 14728 -1240
rect 14328 -1600 14368 -1280
rect 14688 -1600 14728 -1280
rect 14328 -1640 14728 -1600
rect 15340 -1280 15740 -1240
rect 15340 -1600 15380 -1280
rect 15700 -1600 15740 -1280
rect 15340 -1640 15740 -1600
rect 16352 -1280 16752 -1240
rect 16352 -1600 16392 -1280
rect 16712 -1600 16752 -1280
rect 16352 -1640 16752 -1600
rect -17044 -2000 -16644 -1960
rect -17044 -2320 -17004 -2000
rect -16684 -2320 -16644 -2000
rect -17044 -2360 -16644 -2320
rect -16032 -2000 -15632 -1960
rect -16032 -2320 -15992 -2000
rect -15672 -2320 -15632 -2000
rect -16032 -2360 -15632 -2320
rect -15020 -2000 -14620 -1960
rect -15020 -2320 -14980 -2000
rect -14660 -2320 -14620 -2000
rect -15020 -2360 -14620 -2320
rect -14008 -2000 -13608 -1960
rect -14008 -2320 -13968 -2000
rect -13648 -2320 -13608 -2000
rect -14008 -2360 -13608 -2320
rect -12996 -2000 -12596 -1960
rect -12996 -2320 -12956 -2000
rect -12636 -2320 -12596 -2000
rect -12996 -2360 -12596 -2320
rect -11984 -2000 -11584 -1960
rect -11984 -2320 -11944 -2000
rect -11624 -2320 -11584 -2000
rect -11984 -2360 -11584 -2320
rect -10972 -2000 -10572 -1960
rect -10972 -2320 -10932 -2000
rect -10612 -2320 -10572 -2000
rect -10972 -2360 -10572 -2320
rect -9960 -2000 -9560 -1960
rect -9960 -2320 -9920 -2000
rect -9600 -2320 -9560 -2000
rect -9960 -2360 -9560 -2320
rect -8948 -2000 -8548 -1960
rect -8948 -2320 -8908 -2000
rect -8588 -2320 -8548 -2000
rect -8948 -2360 -8548 -2320
rect -7936 -2000 -7536 -1960
rect -7936 -2320 -7896 -2000
rect -7576 -2320 -7536 -2000
rect -7936 -2360 -7536 -2320
rect -6924 -2000 -6524 -1960
rect -6924 -2320 -6884 -2000
rect -6564 -2320 -6524 -2000
rect -6924 -2360 -6524 -2320
rect -5912 -2000 -5512 -1960
rect -5912 -2320 -5872 -2000
rect -5552 -2320 -5512 -2000
rect -5912 -2360 -5512 -2320
rect -4900 -2000 -4500 -1960
rect -4900 -2320 -4860 -2000
rect -4540 -2320 -4500 -2000
rect -4900 -2360 -4500 -2320
rect -3888 -2000 -3488 -1960
rect -3888 -2320 -3848 -2000
rect -3528 -2320 -3488 -2000
rect -3888 -2360 -3488 -2320
rect -2876 -2000 -2476 -1960
rect -2876 -2320 -2836 -2000
rect -2516 -2320 -2476 -2000
rect -2876 -2360 -2476 -2320
rect -1864 -2000 -1464 -1960
rect -1864 -2320 -1824 -2000
rect -1504 -2320 -1464 -2000
rect -1864 -2360 -1464 -2320
rect -852 -2000 -452 -1960
rect -852 -2320 -812 -2000
rect -492 -2320 -452 -2000
rect -852 -2360 -452 -2320
rect 160 -2000 560 -1960
rect 160 -2320 200 -2000
rect 520 -2320 560 -2000
rect 160 -2360 560 -2320
rect 1172 -2000 1572 -1960
rect 1172 -2320 1212 -2000
rect 1532 -2320 1572 -2000
rect 1172 -2360 1572 -2320
rect 2184 -2000 2584 -1960
rect 2184 -2320 2224 -2000
rect 2544 -2320 2584 -2000
rect 2184 -2360 2584 -2320
rect 3196 -2000 3596 -1960
rect 3196 -2320 3236 -2000
rect 3556 -2320 3596 -2000
rect 3196 -2360 3596 -2320
rect 4208 -2000 4608 -1960
rect 4208 -2320 4248 -2000
rect 4568 -2320 4608 -2000
rect 4208 -2360 4608 -2320
rect 5220 -2000 5620 -1960
rect 5220 -2320 5260 -2000
rect 5580 -2320 5620 -2000
rect 5220 -2360 5620 -2320
rect 6232 -2000 6632 -1960
rect 6232 -2320 6272 -2000
rect 6592 -2320 6632 -2000
rect 6232 -2360 6632 -2320
rect 7244 -2000 7644 -1960
rect 7244 -2320 7284 -2000
rect 7604 -2320 7644 -2000
rect 7244 -2360 7644 -2320
rect 8256 -2000 8656 -1960
rect 8256 -2320 8296 -2000
rect 8616 -2320 8656 -2000
rect 8256 -2360 8656 -2320
rect 9268 -2000 9668 -1960
rect 9268 -2320 9308 -2000
rect 9628 -2320 9668 -2000
rect 9268 -2360 9668 -2320
rect 10280 -2000 10680 -1960
rect 10280 -2320 10320 -2000
rect 10640 -2320 10680 -2000
rect 10280 -2360 10680 -2320
rect 11292 -2000 11692 -1960
rect 11292 -2320 11332 -2000
rect 11652 -2320 11692 -2000
rect 11292 -2360 11692 -2320
rect 12304 -2000 12704 -1960
rect 12304 -2320 12344 -2000
rect 12664 -2320 12704 -2000
rect 12304 -2360 12704 -2320
rect 13316 -2000 13716 -1960
rect 13316 -2320 13356 -2000
rect 13676 -2320 13716 -2000
rect 13316 -2360 13716 -2320
rect 14328 -2000 14728 -1960
rect 14328 -2320 14368 -2000
rect 14688 -2320 14728 -2000
rect 14328 -2360 14728 -2320
rect 15340 -2000 15740 -1960
rect 15340 -2320 15380 -2000
rect 15700 -2320 15740 -2000
rect 15340 -2360 15740 -2320
rect 16352 -2000 16752 -1960
rect 16352 -2320 16392 -2000
rect 16712 -2320 16752 -2000
rect 16352 -2360 16752 -2320
rect -17044 -2720 -16644 -2680
rect -17044 -3040 -17004 -2720
rect -16684 -3040 -16644 -2720
rect -17044 -3080 -16644 -3040
rect -16032 -2720 -15632 -2680
rect -16032 -3040 -15992 -2720
rect -15672 -3040 -15632 -2720
rect -16032 -3080 -15632 -3040
rect -15020 -2720 -14620 -2680
rect -15020 -3040 -14980 -2720
rect -14660 -3040 -14620 -2720
rect -15020 -3080 -14620 -3040
rect -14008 -2720 -13608 -2680
rect -14008 -3040 -13968 -2720
rect -13648 -3040 -13608 -2720
rect -14008 -3080 -13608 -3040
rect -12996 -2720 -12596 -2680
rect -12996 -3040 -12956 -2720
rect -12636 -3040 -12596 -2720
rect -12996 -3080 -12596 -3040
rect -11984 -2720 -11584 -2680
rect -11984 -3040 -11944 -2720
rect -11624 -3040 -11584 -2720
rect -11984 -3080 -11584 -3040
rect -10972 -2720 -10572 -2680
rect -10972 -3040 -10932 -2720
rect -10612 -3040 -10572 -2720
rect -10972 -3080 -10572 -3040
rect -9960 -2720 -9560 -2680
rect -9960 -3040 -9920 -2720
rect -9600 -3040 -9560 -2720
rect -9960 -3080 -9560 -3040
rect -8948 -2720 -8548 -2680
rect -8948 -3040 -8908 -2720
rect -8588 -3040 -8548 -2720
rect -8948 -3080 -8548 -3040
rect -7936 -2720 -7536 -2680
rect -7936 -3040 -7896 -2720
rect -7576 -3040 -7536 -2720
rect -7936 -3080 -7536 -3040
rect -6924 -2720 -6524 -2680
rect -6924 -3040 -6884 -2720
rect -6564 -3040 -6524 -2720
rect -6924 -3080 -6524 -3040
rect -5912 -2720 -5512 -2680
rect -5912 -3040 -5872 -2720
rect -5552 -3040 -5512 -2720
rect -5912 -3080 -5512 -3040
rect -4900 -2720 -4500 -2680
rect -4900 -3040 -4860 -2720
rect -4540 -3040 -4500 -2720
rect -4900 -3080 -4500 -3040
rect -3888 -2720 -3488 -2680
rect -3888 -3040 -3848 -2720
rect -3528 -3040 -3488 -2720
rect -3888 -3080 -3488 -3040
rect -2876 -2720 -2476 -2680
rect -2876 -3040 -2836 -2720
rect -2516 -3040 -2476 -2720
rect -2876 -3080 -2476 -3040
rect -1864 -2720 -1464 -2680
rect -1864 -3040 -1824 -2720
rect -1504 -3040 -1464 -2720
rect -1864 -3080 -1464 -3040
rect -852 -2720 -452 -2680
rect -852 -3040 -812 -2720
rect -492 -3040 -452 -2720
rect -852 -3080 -452 -3040
rect 160 -2720 560 -2680
rect 160 -3040 200 -2720
rect 520 -3040 560 -2720
rect 160 -3080 560 -3040
rect 1172 -2720 1572 -2680
rect 1172 -3040 1212 -2720
rect 1532 -3040 1572 -2720
rect 1172 -3080 1572 -3040
rect 2184 -2720 2584 -2680
rect 2184 -3040 2224 -2720
rect 2544 -3040 2584 -2720
rect 2184 -3080 2584 -3040
rect 3196 -2720 3596 -2680
rect 3196 -3040 3236 -2720
rect 3556 -3040 3596 -2720
rect 3196 -3080 3596 -3040
rect 4208 -2720 4608 -2680
rect 4208 -3040 4248 -2720
rect 4568 -3040 4608 -2720
rect 4208 -3080 4608 -3040
rect 5220 -2720 5620 -2680
rect 5220 -3040 5260 -2720
rect 5580 -3040 5620 -2720
rect 5220 -3080 5620 -3040
rect 6232 -2720 6632 -2680
rect 6232 -3040 6272 -2720
rect 6592 -3040 6632 -2720
rect 6232 -3080 6632 -3040
rect 7244 -2720 7644 -2680
rect 7244 -3040 7284 -2720
rect 7604 -3040 7644 -2720
rect 7244 -3080 7644 -3040
rect 8256 -2720 8656 -2680
rect 8256 -3040 8296 -2720
rect 8616 -3040 8656 -2720
rect 8256 -3080 8656 -3040
rect 9268 -2720 9668 -2680
rect 9268 -3040 9308 -2720
rect 9628 -3040 9668 -2720
rect 9268 -3080 9668 -3040
rect 10280 -2720 10680 -2680
rect 10280 -3040 10320 -2720
rect 10640 -3040 10680 -2720
rect 10280 -3080 10680 -3040
rect 11292 -2720 11692 -2680
rect 11292 -3040 11332 -2720
rect 11652 -3040 11692 -2720
rect 11292 -3080 11692 -3040
rect 12304 -2720 12704 -2680
rect 12304 -3040 12344 -2720
rect 12664 -3040 12704 -2720
rect 12304 -3080 12704 -3040
rect 13316 -2720 13716 -2680
rect 13316 -3040 13356 -2720
rect 13676 -3040 13716 -2720
rect 13316 -3080 13716 -3040
rect 14328 -2720 14728 -2680
rect 14328 -3040 14368 -2720
rect 14688 -3040 14728 -2720
rect 14328 -3080 14728 -3040
rect 15340 -2720 15740 -2680
rect 15340 -3040 15380 -2720
rect 15700 -3040 15740 -2720
rect 15340 -3080 15740 -3040
rect 16352 -2720 16752 -2680
rect 16352 -3040 16392 -2720
rect 16712 -3040 16752 -2720
rect 16352 -3080 16752 -3040
rect -17044 -3440 -16644 -3400
rect -17044 -3760 -17004 -3440
rect -16684 -3760 -16644 -3440
rect -17044 -3800 -16644 -3760
rect -16032 -3440 -15632 -3400
rect -16032 -3760 -15992 -3440
rect -15672 -3760 -15632 -3440
rect -16032 -3800 -15632 -3760
rect -15020 -3440 -14620 -3400
rect -15020 -3760 -14980 -3440
rect -14660 -3760 -14620 -3440
rect -15020 -3800 -14620 -3760
rect -14008 -3440 -13608 -3400
rect -14008 -3760 -13968 -3440
rect -13648 -3760 -13608 -3440
rect -14008 -3800 -13608 -3760
rect -12996 -3440 -12596 -3400
rect -12996 -3760 -12956 -3440
rect -12636 -3760 -12596 -3440
rect -12996 -3800 -12596 -3760
rect -11984 -3440 -11584 -3400
rect -11984 -3760 -11944 -3440
rect -11624 -3760 -11584 -3440
rect -11984 -3800 -11584 -3760
rect -10972 -3440 -10572 -3400
rect -10972 -3760 -10932 -3440
rect -10612 -3760 -10572 -3440
rect -10972 -3800 -10572 -3760
rect -9960 -3440 -9560 -3400
rect -9960 -3760 -9920 -3440
rect -9600 -3760 -9560 -3440
rect -9960 -3800 -9560 -3760
rect -8948 -3440 -8548 -3400
rect -8948 -3760 -8908 -3440
rect -8588 -3760 -8548 -3440
rect -8948 -3800 -8548 -3760
rect -7936 -3440 -7536 -3400
rect -7936 -3760 -7896 -3440
rect -7576 -3760 -7536 -3440
rect -7936 -3800 -7536 -3760
rect -6924 -3440 -6524 -3400
rect -6924 -3760 -6884 -3440
rect -6564 -3760 -6524 -3440
rect -6924 -3800 -6524 -3760
rect -5912 -3440 -5512 -3400
rect -5912 -3760 -5872 -3440
rect -5552 -3760 -5512 -3440
rect -5912 -3800 -5512 -3760
rect -4900 -3440 -4500 -3400
rect -4900 -3760 -4860 -3440
rect -4540 -3760 -4500 -3440
rect -4900 -3800 -4500 -3760
rect -3888 -3440 -3488 -3400
rect -3888 -3760 -3848 -3440
rect -3528 -3760 -3488 -3440
rect -3888 -3800 -3488 -3760
rect -2876 -3440 -2476 -3400
rect -2876 -3760 -2836 -3440
rect -2516 -3760 -2476 -3440
rect -2876 -3800 -2476 -3760
rect -1864 -3440 -1464 -3400
rect -1864 -3760 -1824 -3440
rect -1504 -3760 -1464 -3440
rect -1864 -3800 -1464 -3760
rect -852 -3440 -452 -3400
rect -852 -3760 -812 -3440
rect -492 -3760 -452 -3440
rect -852 -3800 -452 -3760
rect 160 -3440 560 -3400
rect 160 -3760 200 -3440
rect 520 -3760 560 -3440
rect 160 -3800 560 -3760
rect 1172 -3440 1572 -3400
rect 1172 -3760 1212 -3440
rect 1532 -3760 1572 -3440
rect 1172 -3800 1572 -3760
rect 2184 -3440 2584 -3400
rect 2184 -3760 2224 -3440
rect 2544 -3760 2584 -3440
rect 2184 -3800 2584 -3760
rect 3196 -3440 3596 -3400
rect 3196 -3760 3236 -3440
rect 3556 -3760 3596 -3440
rect 3196 -3800 3596 -3760
rect 4208 -3440 4608 -3400
rect 4208 -3760 4248 -3440
rect 4568 -3760 4608 -3440
rect 4208 -3800 4608 -3760
rect 5220 -3440 5620 -3400
rect 5220 -3760 5260 -3440
rect 5580 -3760 5620 -3440
rect 5220 -3800 5620 -3760
rect 6232 -3440 6632 -3400
rect 6232 -3760 6272 -3440
rect 6592 -3760 6632 -3440
rect 6232 -3800 6632 -3760
rect 7244 -3440 7644 -3400
rect 7244 -3760 7284 -3440
rect 7604 -3760 7644 -3440
rect 7244 -3800 7644 -3760
rect 8256 -3440 8656 -3400
rect 8256 -3760 8296 -3440
rect 8616 -3760 8656 -3440
rect 8256 -3800 8656 -3760
rect 9268 -3440 9668 -3400
rect 9268 -3760 9308 -3440
rect 9628 -3760 9668 -3440
rect 9268 -3800 9668 -3760
rect 10280 -3440 10680 -3400
rect 10280 -3760 10320 -3440
rect 10640 -3760 10680 -3440
rect 10280 -3800 10680 -3760
rect 11292 -3440 11692 -3400
rect 11292 -3760 11332 -3440
rect 11652 -3760 11692 -3440
rect 11292 -3800 11692 -3760
rect 12304 -3440 12704 -3400
rect 12304 -3760 12344 -3440
rect 12664 -3760 12704 -3440
rect 12304 -3800 12704 -3760
rect 13316 -3440 13716 -3400
rect 13316 -3760 13356 -3440
rect 13676 -3760 13716 -3440
rect 13316 -3800 13716 -3760
rect 14328 -3440 14728 -3400
rect 14328 -3760 14368 -3440
rect 14688 -3760 14728 -3440
rect 14328 -3800 14728 -3760
rect 15340 -3440 15740 -3400
rect 15340 -3760 15380 -3440
rect 15700 -3760 15740 -3440
rect 15340 -3800 15740 -3760
rect 16352 -3440 16752 -3400
rect 16352 -3760 16392 -3440
rect 16712 -3760 16752 -3440
rect 16352 -3800 16752 -3760
rect -17044 -4160 -16644 -4120
rect -17044 -4480 -17004 -4160
rect -16684 -4480 -16644 -4160
rect -17044 -4520 -16644 -4480
rect -16032 -4160 -15632 -4120
rect -16032 -4480 -15992 -4160
rect -15672 -4480 -15632 -4160
rect -16032 -4520 -15632 -4480
rect -15020 -4160 -14620 -4120
rect -15020 -4480 -14980 -4160
rect -14660 -4480 -14620 -4160
rect -15020 -4520 -14620 -4480
rect -14008 -4160 -13608 -4120
rect -14008 -4480 -13968 -4160
rect -13648 -4480 -13608 -4160
rect -14008 -4520 -13608 -4480
rect -12996 -4160 -12596 -4120
rect -12996 -4480 -12956 -4160
rect -12636 -4480 -12596 -4160
rect -12996 -4520 -12596 -4480
rect -11984 -4160 -11584 -4120
rect -11984 -4480 -11944 -4160
rect -11624 -4480 -11584 -4160
rect -11984 -4520 -11584 -4480
rect -10972 -4160 -10572 -4120
rect -10972 -4480 -10932 -4160
rect -10612 -4480 -10572 -4160
rect -10972 -4520 -10572 -4480
rect -9960 -4160 -9560 -4120
rect -9960 -4480 -9920 -4160
rect -9600 -4480 -9560 -4160
rect -9960 -4520 -9560 -4480
rect -8948 -4160 -8548 -4120
rect -8948 -4480 -8908 -4160
rect -8588 -4480 -8548 -4160
rect -8948 -4520 -8548 -4480
rect -7936 -4160 -7536 -4120
rect -7936 -4480 -7896 -4160
rect -7576 -4480 -7536 -4160
rect -7936 -4520 -7536 -4480
rect -6924 -4160 -6524 -4120
rect -6924 -4480 -6884 -4160
rect -6564 -4480 -6524 -4160
rect -6924 -4520 -6524 -4480
rect -5912 -4160 -5512 -4120
rect -5912 -4480 -5872 -4160
rect -5552 -4480 -5512 -4160
rect -5912 -4520 -5512 -4480
rect -4900 -4160 -4500 -4120
rect -4900 -4480 -4860 -4160
rect -4540 -4480 -4500 -4160
rect -4900 -4520 -4500 -4480
rect -3888 -4160 -3488 -4120
rect -3888 -4480 -3848 -4160
rect -3528 -4480 -3488 -4160
rect -3888 -4520 -3488 -4480
rect -2876 -4160 -2476 -4120
rect -2876 -4480 -2836 -4160
rect -2516 -4480 -2476 -4160
rect -2876 -4520 -2476 -4480
rect -1864 -4160 -1464 -4120
rect -1864 -4480 -1824 -4160
rect -1504 -4480 -1464 -4160
rect -1864 -4520 -1464 -4480
rect -852 -4160 -452 -4120
rect -852 -4480 -812 -4160
rect -492 -4480 -452 -4160
rect -852 -4520 -452 -4480
rect 160 -4160 560 -4120
rect 160 -4480 200 -4160
rect 520 -4480 560 -4160
rect 160 -4520 560 -4480
rect 1172 -4160 1572 -4120
rect 1172 -4480 1212 -4160
rect 1532 -4480 1572 -4160
rect 1172 -4520 1572 -4480
rect 2184 -4160 2584 -4120
rect 2184 -4480 2224 -4160
rect 2544 -4480 2584 -4160
rect 2184 -4520 2584 -4480
rect 3196 -4160 3596 -4120
rect 3196 -4480 3236 -4160
rect 3556 -4480 3596 -4160
rect 3196 -4520 3596 -4480
rect 4208 -4160 4608 -4120
rect 4208 -4480 4248 -4160
rect 4568 -4480 4608 -4160
rect 4208 -4520 4608 -4480
rect 5220 -4160 5620 -4120
rect 5220 -4480 5260 -4160
rect 5580 -4480 5620 -4160
rect 5220 -4520 5620 -4480
rect 6232 -4160 6632 -4120
rect 6232 -4480 6272 -4160
rect 6592 -4480 6632 -4160
rect 6232 -4520 6632 -4480
rect 7244 -4160 7644 -4120
rect 7244 -4480 7284 -4160
rect 7604 -4480 7644 -4160
rect 7244 -4520 7644 -4480
rect 8256 -4160 8656 -4120
rect 8256 -4480 8296 -4160
rect 8616 -4480 8656 -4160
rect 8256 -4520 8656 -4480
rect 9268 -4160 9668 -4120
rect 9268 -4480 9308 -4160
rect 9628 -4480 9668 -4160
rect 9268 -4520 9668 -4480
rect 10280 -4160 10680 -4120
rect 10280 -4480 10320 -4160
rect 10640 -4480 10680 -4160
rect 10280 -4520 10680 -4480
rect 11292 -4160 11692 -4120
rect 11292 -4480 11332 -4160
rect 11652 -4480 11692 -4160
rect 11292 -4520 11692 -4480
rect 12304 -4160 12704 -4120
rect 12304 -4480 12344 -4160
rect 12664 -4480 12704 -4160
rect 12304 -4520 12704 -4480
rect 13316 -4160 13716 -4120
rect 13316 -4480 13356 -4160
rect 13676 -4480 13716 -4160
rect 13316 -4520 13716 -4480
rect 14328 -4160 14728 -4120
rect 14328 -4480 14368 -4160
rect 14688 -4480 14728 -4160
rect 14328 -4520 14728 -4480
rect 15340 -4160 15740 -4120
rect 15340 -4480 15380 -4160
rect 15700 -4480 15740 -4160
rect 15340 -4520 15740 -4480
rect 16352 -4160 16752 -4120
rect 16352 -4480 16392 -4160
rect 16712 -4480 16752 -4160
rect 16352 -4520 16752 -4480
rect -17044 -4880 -16644 -4840
rect -17044 -5200 -17004 -4880
rect -16684 -5200 -16644 -4880
rect -17044 -5240 -16644 -5200
rect -16032 -4880 -15632 -4840
rect -16032 -5200 -15992 -4880
rect -15672 -5200 -15632 -4880
rect -16032 -5240 -15632 -5200
rect -15020 -4880 -14620 -4840
rect -15020 -5200 -14980 -4880
rect -14660 -5200 -14620 -4880
rect -15020 -5240 -14620 -5200
rect -14008 -4880 -13608 -4840
rect -14008 -5200 -13968 -4880
rect -13648 -5200 -13608 -4880
rect -14008 -5240 -13608 -5200
rect -12996 -4880 -12596 -4840
rect -12996 -5200 -12956 -4880
rect -12636 -5200 -12596 -4880
rect -12996 -5240 -12596 -5200
rect -11984 -4880 -11584 -4840
rect -11984 -5200 -11944 -4880
rect -11624 -5200 -11584 -4880
rect -11984 -5240 -11584 -5200
rect -10972 -4880 -10572 -4840
rect -10972 -5200 -10932 -4880
rect -10612 -5200 -10572 -4880
rect -10972 -5240 -10572 -5200
rect -9960 -4880 -9560 -4840
rect -9960 -5200 -9920 -4880
rect -9600 -5200 -9560 -4880
rect -9960 -5240 -9560 -5200
rect -8948 -4880 -8548 -4840
rect -8948 -5200 -8908 -4880
rect -8588 -5200 -8548 -4880
rect -8948 -5240 -8548 -5200
rect -7936 -4880 -7536 -4840
rect -7936 -5200 -7896 -4880
rect -7576 -5200 -7536 -4880
rect -7936 -5240 -7536 -5200
rect -6924 -4880 -6524 -4840
rect -6924 -5200 -6884 -4880
rect -6564 -5200 -6524 -4880
rect -6924 -5240 -6524 -5200
rect -5912 -4880 -5512 -4840
rect -5912 -5200 -5872 -4880
rect -5552 -5200 -5512 -4880
rect -5912 -5240 -5512 -5200
rect -4900 -4880 -4500 -4840
rect -4900 -5200 -4860 -4880
rect -4540 -5200 -4500 -4880
rect -4900 -5240 -4500 -5200
rect -3888 -4880 -3488 -4840
rect -3888 -5200 -3848 -4880
rect -3528 -5200 -3488 -4880
rect -3888 -5240 -3488 -5200
rect -2876 -4880 -2476 -4840
rect -2876 -5200 -2836 -4880
rect -2516 -5200 -2476 -4880
rect -2876 -5240 -2476 -5200
rect -1864 -4880 -1464 -4840
rect -1864 -5200 -1824 -4880
rect -1504 -5200 -1464 -4880
rect -1864 -5240 -1464 -5200
rect -852 -4880 -452 -4840
rect -852 -5200 -812 -4880
rect -492 -5200 -452 -4880
rect -852 -5240 -452 -5200
rect 160 -4880 560 -4840
rect 160 -5200 200 -4880
rect 520 -5200 560 -4880
rect 160 -5240 560 -5200
rect 1172 -4880 1572 -4840
rect 1172 -5200 1212 -4880
rect 1532 -5200 1572 -4880
rect 1172 -5240 1572 -5200
rect 2184 -4880 2584 -4840
rect 2184 -5200 2224 -4880
rect 2544 -5200 2584 -4880
rect 2184 -5240 2584 -5200
rect 3196 -4880 3596 -4840
rect 3196 -5200 3236 -4880
rect 3556 -5200 3596 -4880
rect 3196 -5240 3596 -5200
rect 4208 -4880 4608 -4840
rect 4208 -5200 4248 -4880
rect 4568 -5200 4608 -4880
rect 4208 -5240 4608 -5200
rect 5220 -4880 5620 -4840
rect 5220 -5200 5260 -4880
rect 5580 -5200 5620 -4880
rect 5220 -5240 5620 -5200
rect 6232 -4880 6632 -4840
rect 6232 -5200 6272 -4880
rect 6592 -5200 6632 -4880
rect 6232 -5240 6632 -5200
rect 7244 -4880 7644 -4840
rect 7244 -5200 7284 -4880
rect 7604 -5200 7644 -4880
rect 7244 -5240 7644 -5200
rect 8256 -4880 8656 -4840
rect 8256 -5200 8296 -4880
rect 8616 -5200 8656 -4880
rect 8256 -5240 8656 -5200
rect 9268 -4880 9668 -4840
rect 9268 -5200 9308 -4880
rect 9628 -5200 9668 -4880
rect 9268 -5240 9668 -5200
rect 10280 -4880 10680 -4840
rect 10280 -5200 10320 -4880
rect 10640 -5200 10680 -4880
rect 10280 -5240 10680 -5200
rect 11292 -4880 11692 -4840
rect 11292 -5200 11332 -4880
rect 11652 -5200 11692 -4880
rect 11292 -5240 11692 -5200
rect 12304 -4880 12704 -4840
rect 12304 -5200 12344 -4880
rect 12664 -5200 12704 -4880
rect 12304 -5240 12704 -5200
rect 13316 -4880 13716 -4840
rect 13316 -5200 13356 -4880
rect 13676 -5200 13716 -4880
rect 13316 -5240 13716 -5200
rect 14328 -4880 14728 -4840
rect 14328 -5200 14368 -4880
rect 14688 -5200 14728 -4880
rect 14328 -5240 14728 -5200
rect 15340 -4880 15740 -4840
rect 15340 -5200 15380 -4880
rect 15700 -5200 15740 -4880
rect 15340 -5240 15740 -5200
rect 16352 -4880 16752 -4840
rect 16352 -5200 16392 -4880
rect 16712 -5200 16752 -4880
rect 16352 -5240 16752 -5200
rect -17044 -5600 -16644 -5560
rect -17044 -5920 -17004 -5600
rect -16684 -5920 -16644 -5600
rect -17044 -5960 -16644 -5920
rect -16032 -5600 -15632 -5560
rect -16032 -5920 -15992 -5600
rect -15672 -5920 -15632 -5600
rect -16032 -5960 -15632 -5920
rect -15020 -5600 -14620 -5560
rect -15020 -5920 -14980 -5600
rect -14660 -5920 -14620 -5600
rect -15020 -5960 -14620 -5920
rect -14008 -5600 -13608 -5560
rect -14008 -5920 -13968 -5600
rect -13648 -5920 -13608 -5600
rect -14008 -5960 -13608 -5920
rect -12996 -5600 -12596 -5560
rect -12996 -5920 -12956 -5600
rect -12636 -5920 -12596 -5600
rect -12996 -5960 -12596 -5920
rect -11984 -5600 -11584 -5560
rect -11984 -5920 -11944 -5600
rect -11624 -5920 -11584 -5600
rect -11984 -5960 -11584 -5920
rect -10972 -5600 -10572 -5560
rect -10972 -5920 -10932 -5600
rect -10612 -5920 -10572 -5600
rect -10972 -5960 -10572 -5920
rect -9960 -5600 -9560 -5560
rect -9960 -5920 -9920 -5600
rect -9600 -5920 -9560 -5600
rect -9960 -5960 -9560 -5920
rect -8948 -5600 -8548 -5560
rect -8948 -5920 -8908 -5600
rect -8588 -5920 -8548 -5600
rect -8948 -5960 -8548 -5920
rect -7936 -5600 -7536 -5560
rect -7936 -5920 -7896 -5600
rect -7576 -5920 -7536 -5600
rect -7936 -5960 -7536 -5920
rect -6924 -5600 -6524 -5560
rect -6924 -5920 -6884 -5600
rect -6564 -5920 -6524 -5600
rect -6924 -5960 -6524 -5920
rect -5912 -5600 -5512 -5560
rect -5912 -5920 -5872 -5600
rect -5552 -5920 -5512 -5600
rect -5912 -5960 -5512 -5920
rect -4900 -5600 -4500 -5560
rect -4900 -5920 -4860 -5600
rect -4540 -5920 -4500 -5600
rect -4900 -5960 -4500 -5920
rect -3888 -5600 -3488 -5560
rect -3888 -5920 -3848 -5600
rect -3528 -5920 -3488 -5600
rect -3888 -5960 -3488 -5920
rect -2876 -5600 -2476 -5560
rect -2876 -5920 -2836 -5600
rect -2516 -5920 -2476 -5600
rect -2876 -5960 -2476 -5920
rect -1864 -5600 -1464 -5560
rect -1864 -5920 -1824 -5600
rect -1504 -5920 -1464 -5600
rect -1864 -5960 -1464 -5920
rect -852 -5600 -452 -5560
rect -852 -5920 -812 -5600
rect -492 -5920 -452 -5600
rect -852 -5960 -452 -5920
rect 160 -5600 560 -5560
rect 160 -5920 200 -5600
rect 520 -5920 560 -5600
rect 160 -5960 560 -5920
rect 1172 -5600 1572 -5560
rect 1172 -5920 1212 -5600
rect 1532 -5920 1572 -5600
rect 1172 -5960 1572 -5920
rect 2184 -5600 2584 -5560
rect 2184 -5920 2224 -5600
rect 2544 -5920 2584 -5600
rect 2184 -5960 2584 -5920
rect 3196 -5600 3596 -5560
rect 3196 -5920 3236 -5600
rect 3556 -5920 3596 -5600
rect 3196 -5960 3596 -5920
rect 4208 -5600 4608 -5560
rect 4208 -5920 4248 -5600
rect 4568 -5920 4608 -5600
rect 4208 -5960 4608 -5920
rect 5220 -5600 5620 -5560
rect 5220 -5920 5260 -5600
rect 5580 -5920 5620 -5600
rect 5220 -5960 5620 -5920
rect 6232 -5600 6632 -5560
rect 6232 -5920 6272 -5600
rect 6592 -5920 6632 -5600
rect 6232 -5960 6632 -5920
rect 7244 -5600 7644 -5560
rect 7244 -5920 7284 -5600
rect 7604 -5920 7644 -5600
rect 7244 -5960 7644 -5920
rect 8256 -5600 8656 -5560
rect 8256 -5920 8296 -5600
rect 8616 -5920 8656 -5600
rect 8256 -5960 8656 -5920
rect 9268 -5600 9668 -5560
rect 9268 -5920 9308 -5600
rect 9628 -5920 9668 -5600
rect 9268 -5960 9668 -5920
rect 10280 -5600 10680 -5560
rect 10280 -5920 10320 -5600
rect 10640 -5920 10680 -5600
rect 10280 -5960 10680 -5920
rect 11292 -5600 11692 -5560
rect 11292 -5920 11332 -5600
rect 11652 -5920 11692 -5600
rect 11292 -5960 11692 -5920
rect 12304 -5600 12704 -5560
rect 12304 -5920 12344 -5600
rect 12664 -5920 12704 -5600
rect 12304 -5960 12704 -5920
rect 13316 -5600 13716 -5560
rect 13316 -5920 13356 -5600
rect 13676 -5920 13716 -5600
rect 13316 -5960 13716 -5920
rect 14328 -5600 14728 -5560
rect 14328 -5920 14368 -5600
rect 14688 -5920 14728 -5600
rect 14328 -5960 14728 -5920
rect 15340 -5600 15740 -5560
rect 15340 -5920 15380 -5600
rect 15700 -5920 15740 -5600
rect 15340 -5960 15740 -5920
rect 16352 -5600 16752 -5560
rect 16352 -5920 16392 -5600
rect 16712 -5920 16752 -5600
rect 16352 -5960 16752 -5920
rect -17044 -6320 -16644 -6280
rect -17044 -6640 -17004 -6320
rect -16684 -6640 -16644 -6320
rect -17044 -6680 -16644 -6640
rect -16032 -6320 -15632 -6280
rect -16032 -6640 -15992 -6320
rect -15672 -6640 -15632 -6320
rect -16032 -6680 -15632 -6640
rect -15020 -6320 -14620 -6280
rect -15020 -6640 -14980 -6320
rect -14660 -6640 -14620 -6320
rect -15020 -6680 -14620 -6640
rect -14008 -6320 -13608 -6280
rect -14008 -6640 -13968 -6320
rect -13648 -6640 -13608 -6320
rect -14008 -6680 -13608 -6640
rect -12996 -6320 -12596 -6280
rect -12996 -6640 -12956 -6320
rect -12636 -6640 -12596 -6320
rect -12996 -6680 -12596 -6640
rect -11984 -6320 -11584 -6280
rect -11984 -6640 -11944 -6320
rect -11624 -6640 -11584 -6320
rect -11984 -6680 -11584 -6640
rect -10972 -6320 -10572 -6280
rect -10972 -6640 -10932 -6320
rect -10612 -6640 -10572 -6320
rect -10972 -6680 -10572 -6640
rect -9960 -6320 -9560 -6280
rect -9960 -6640 -9920 -6320
rect -9600 -6640 -9560 -6320
rect -9960 -6680 -9560 -6640
rect -8948 -6320 -8548 -6280
rect -8948 -6640 -8908 -6320
rect -8588 -6640 -8548 -6320
rect -8948 -6680 -8548 -6640
rect -7936 -6320 -7536 -6280
rect -7936 -6640 -7896 -6320
rect -7576 -6640 -7536 -6320
rect -7936 -6680 -7536 -6640
rect -6924 -6320 -6524 -6280
rect -6924 -6640 -6884 -6320
rect -6564 -6640 -6524 -6320
rect -6924 -6680 -6524 -6640
rect -5912 -6320 -5512 -6280
rect -5912 -6640 -5872 -6320
rect -5552 -6640 -5512 -6320
rect -5912 -6680 -5512 -6640
rect -4900 -6320 -4500 -6280
rect -4900 -6640 -4860 -6320
rect -4540 -6640 -4500 -6320
rect -4900 -6680 -4500 -6640
rect -3888 -6320 -3488 -6280
rect -3888 -6640 -3848 -6320
rect -3528 -6640 -3488 -6320
rect -3888 -6680 -3488 -6640
rect -2876 -6320 -2476 -6280
rect -2876 -6640 -2836 -6320
rect -2516 -6640 -2476 -6320
rect -2876 -6680 -2476 -6640
rect -1864 -6320 -1464 -6280
rect -1864 -6640 -1824 -6320
rect -1504 -6640 -1464 -6320
rect -1864 -6680 -1464 -6640
rect -852 -6320 -452 -6280
rect -852 -6640 -812 -6320
rect -492 -6640 -452 -6320
rect -852 -6680 -452 -6640
rect 160 -6320 560 -6280
rect 160 -6640 200 -6320
rect 520 -6640 560 -6320
rect 160 -6680 560 -6640
rect 1172 -6320 1572 -6280
rect 1172 -6640 1212 -6320
rect 1532 -6640 1572 -6320
rect 1172 -6680 1572 -6640
rect 2184 -6320 2584 -6280
rect 2184 -6640 2224 -6320
rect 2544 -6640 2584 -6320
rect 2184 -6680 2584 -6640
rect 3196 -6320 3596 -6280
rect 3196 -6640 3236 -6320
rect 3556 -6640 3596 -6320
rect 3196 -6680 3596 -6640
rect 4208 -6320 4608 -6280
rect 4208 -6640 4248 -6320
rect 4568 -6640 4608 -6320
rect 4208 -6680 4608 -6640
rect 5220 -6320 5620 -6280
rect 5220 -6640 5260 -6320
rect 5580 -6640 5620 -6320
rect 5220 -6680 5620 -6640
rect 6232 -6320 6632 -6280
rect 6232 -6640 6272 -6320
rect 6592 -6640 6632 -6320
rect 6232 -6680 6632 -6640
rect 7244 -6320 7644 -6280
rect 7244 -6640 7284 -6320
rect 7604 -6640 7644 -6320
rect 7244 -6680 7644 -6640
rect 8256 -6320 8656 -6280
rect 8256 -6640 8296 -6320
rect 8616 -6640 8656 -6320
rect 8256 -6680 8656 -6640
rect 9268 -6320 9668 -6280
rect 9268 -6640 9308 -6320
rect 9628 -6640 9668 -6320
rect 9268 -6680 9668 -6640
rect 10280 -6320 10680 -6280
rect 10280 -6640 10320 -6320
rect 10640 -6640 10680 -6320
rect 10280 -6680 10680 -6640
rect 11292 -6320 11692 -6280
rect 11292 -6640 11332 -6320
rect 11652 -6640 11692 -6320
rect 11292 -6680 11692 -6640
rect 12304 -6320 12704 -6280
rect 12304 -6640 12344 -6320
rect 12664 -6640 12704 -6320
rect 12304 -6680 12704 -6640
rect 13316 -6320 13716 -6280
rect 13316 -6640 13356 -6320
rect 13676 -6640 13716 -6320
rect 13316 -6680 13716 -6640
rect 14328 -6320 14728 -6280
rect 14328 -6640 14368 -6320
rect 14688 -6640 14728 -6320
rect 14328 -6680 14728 -6640
rect 15340 -6320 15740 -6280
rect 15340 -6640 15380 -6320
rect 15700 -6640 15740 -6320
rect 15340 -6680 15740 -6640
rect 16352 -6320 16752 -6280
rect 16352 -6640 16392 -6320
rect 16712 -6640 16752 -6320
rect 16352 -6680 16752 -6640
rect -17044 -7040 -16644 -7000
rect -17044 -7360 -17004 -7040
rect -16684 -7360 -16644 -7040
rect -17044 -7400 -16644 -7360
rect -16032 -7040 -15632 -7000
rect -16032 -7360 -15992 -7040
rect -15672 -7360 -15632 -7040
rect -16032 -7400 -15632 -7360
rect -15020 -7040 -14620 -7000
rect -15020 -7360 -14980 -7040
rect -14660 -7360 -14620 -7040
rect -15020 -7400 -14620 -7360
rect -14008 -7040 -13608 -7000
rect -14008 -7360 -13968 -7040
rect -13648 -7360 -13608 -7040
rect -14008 -7400 -13608 -7360
rect -12996 -7040 -12596 -7000
rect -12996 -7360 -12956 -7040
rect -12636 -7360 -12596 -7040
rect -12996 -7400 -12596 -7360
rect -11984 -7040 -11584 -7000
rect -11984 -7360 -11944 -7040
rect -11624 -7360 -11584 -7040
rect -11984 -7400 -11584 -7360
rect -10972 -7040 -10572 -7000
rect -10972 -7360 -10932 -7040
rect -10612 -7360 -10572 -7040
rect -10972 -7400 -10572 -7360
rect -9960 -7040 -9560 -7000
rect -9960 -7360 -9920 -7040
rect -9600 -7360 -9560 -7040
rect -9960 -7400 -9560 -7360
rect -8948 -7040 -8548 -7000
rect -8948 -7360 -8908 -7040
rect -8588 -7360 -8548 -7040
rect -8948 -7400 -8548 -7360
rect -7936 -7040 -7536 -7000
rect -7936 -7360 -7896 -7040
rect -7576 -7360 -7536 -7040
rect -7936 -7400 -7536 -7360
rect -6924 -7040 -6524 -7000
rect -6924 -7360 -6884 -7040
rect -6564 -7360 -6524 -7040
rect -6924 -7400 -6524 -7360
rect -5912 -7040 -5512 -7000
rect -5912 -7360 -5872 -7040
rect -5552 -7360 -5512 -7040
rect -5912 -7400 -5512 -7360
rect -4900 -7040 -4500 -7000
rect -4900 -7360 -4860 -7040
rect -4540 -7360 -4500 -7040
rect -4900 -7400 -4500 -7360
rect -3888 -7040 -3488 -7000
rect -3888 -7360 -3848 -7040
rect -3528 -7360 -3488 -7040
rect -3888 -7400 -3488 -7360
rect -2876 -7040 -2476 -7000
rect -2876 -7360 -2836 -7040
rect -2516 -7360 -2476 -7040
rect -2876 -7400 -2476 -7360
rect -1864 -7040 -1464 -7000
rect -1864 -7360 -1824 -7040
rect -1504 -7360 -1464 -7040
rect -1864 -7400 -1464 -7360
rect -852 -7040 -452 -7000
rect -852 -7360 -812 -7040
rect -492 -7360 -452 -7040
rect -852 -7400 -452 -7360
rect 160 -7040 560 -7000
rect 160 -7360 200 -7040
rect 520 -7360 560 -7040
rect 160 -7400 560 -7360
rect 1172 -7040 1572 -7000
rect 1172 -7360 1212 -7040
rect 1532 -7360 1572 -7040
rect 1172 -7400 1572 -7360
rect 2184 -7040 2584 -7000
rect 2184 -7360 2224 -7040
rect 2544 -7360 2584 -7040
rect 2184 -7400 2584 -7360
rect 3196 -7040 3596 -7000
rect 3196 -7360 3236 -7040
rect 3556 -7360 3596 -7040
rect 3196 -7400 3596 -7360
rect 4208 -7040 4608 -7000
rect 4208 -7360 4248 -7040
rect 4568 -7360 4608 -7040
rect 4208 -7400 4608 -7360
rect 5220 -7040 5620 -7000
rect 5220 -7360 5260 -7040
rect 5580 -7360 5620 -7040
rect 5220 -7400 5620 -7360
rect 6232 -7040 6632 -7000
rect 6232 -7360 6272 -7040
rect 6592 -7360 6632 -7040
rect 6232 -7400 6632 -7360
rect 7244 -7040 7644 -7000
rect 7244 -7360 7284 -7040
rect 7604 -7360 7644 -7040
rect 7244 -7400 7644 -7360
rect 8256 -7040 8656 -7000
rect 8256 -7360 8296 -7040
rect 8616 -7360 8656 -7040
rect 8256 -7400 8656 -7360
rect 9268 -7040 9668 -7000
rect 9268 -7360 9308 -7040
rect 9628 -7360 9668 -7040
rect 9268 -7400 9668 -7360
rect 10280 -7040 10680 -7000
rect 10280 -7360 10320 -7040
rect 10640 -7360 10680 -7040
rect 10280 -7400 10680 -7360
rect 11292 -7040 11692 -7000
rect 11292 -7360 11332 -7040
rect 11652 -7360 11692 -7040
rect 11292 -7400 11692 -7360
rect 12304 -7040 12704 -7000
rect 12304 -7360 12344 -7040
rect 12664 -7360 12704 -7040
rect 12304 -7400 12704 -7360
rect 13316 -7040 13716 -7000
rect 13316 -7360 13356 -7040
rect 13676 -7360 13716 -7040
rect 13316 -7400 13716 -7360
rect 14328 -7040 14728 -7000
rect 14328 -7360 14368 -7040
rect 14688 -7360 14728 -7040
rect 14328 -7400 14728 -7360
rect 15340 -7040 15740 -7000
rect 15340 -7360 15380 -7040
rect 15700 -7360 15740 -7040
rect 15340 -7400 15740 -7360
rect 16352 -7040 16752 -7000
rect 16352 -7360 16392 -7040
rect 16712 -7360 16752 -7040
rect 16352 -7400 16752 -7360
rect -17044 -7760 -16644 -7720
rect -17044 -8080 -17004 -7760
rect -16684 -8080 -16644 -7760
rect -17044 -8120 -16644 -8080
rect -16032 -7760 -15632 -7720
rect -16032 -8080 -15992 -7760
rect -15672 -8080 -15632 -7760
rect -16032 -8120 -15632 -8080
rect -15020 -7760 -14620 -7720
rect -15020 -8080 -14980 -7760
rect -14660 -8080 -14620 -7760
rect -15020 -8120 -14620 -8080
rect -14008 -7760 -13608 -7720
rect -14008 -8080 -13968 -7760
rect -13648 -8080 -13608 -7760
rect -14008 -8120 -13608 -8080
rect -12996 -7760 -12596 -7720
rect -12996 -8080 -12956 -7760
rect -12636 -8080 -12596 -7760
rect -12996 -8120 -12596 -8080
rect -11984 -7760 -11584 -7720
rect -11984 -8080 -11944 -7760
rect -11624 -8080 -11584 -7760
rect -11984 -8120 -11584 -8080
rect -10972 -7760 -10572 -7720
rect -10972 -8080 -10932 -7760
rect -10612 -8080 -10572 -7760
rect -10972 -8120 -10572 -8080
rect -9960 -7760 -9560 -7720
rect -9960 -8080 -9920 -7760
rect -9600 -8080 -9560 -7760
rect -9960 -8120 -9560 -8080
rect -8948 -7760 -8548 -7720
rect -8948 -8080 -8908 -7760
rect -8588 -8080 -8548 -7760
rect -8948 -8120 -8548 -8080
rect -7936 -7760 -7536 -7720
rect -7936 -8080 -7896 -7760
rect -7576 -8080 -7536 -7760
rect -7936 -8120 -7536 -8080
rect -6924 -7760 -6524 -7720
rect -6924 -8080 -6884 -7760
rect -6564 -8080 -6524 -7760
rect -6924 -8120 -6524 -8080
rect -5912 -7760 -5512 -7720
rect -5912 -8080 -5872 -7760
rect -5552 -8080 -5512 -7760
rect -5912 -8120 -5512 -8080
rect -4900 -7760 -4500 -7720
rect -4900 -8080 -4860 -7760
rect -4540 -8080 -4500 -7760
rect -4900 -8120 -4500 -8080
rect -3888 -7760 -3488 -7720
rect -3888 -8080 -3848 -7760
rect -3528 -8080 -3488 -7760
rect -3888 -8120 -3488 -8080
rect -2876 -7760 -2476 -7720
rect -2876 -8080 -2836 -7760
rect -2516 -8080 -2476 -7760
rect -2876 -8120 -2476 -8080
rect -1864 -7760 -1464 -7720
rect -1864 -8080 -1824 -7760
rect -1504 -8080 -1464 -7760
rect -1864 -8120 -1464 -8080
rect -852 -7760 -452 -7720
rect -852 -8080 -812 -7760
rect -492 -8080 -452 -7760
rect -852 -8120 -452 -8080
rect 160 -7760 560 -7720
rect 160 -8080 200 -7760
rect 520 -8080 560 -7760
rect 160 -8120 560 -8080
rect 1172 -7760 1572 -7720
rect 1172 -8080 1212 -7760
rect 1532 -8080 1572 -7760
rect 1172 -8120 1572 -8080
rect 2184 -7760 2584 -7720
rect 2184 -8080 2224 -7760
rect 2544 -8080 2584 -7760
rect 2184 -8120 2584 -8080
rect 3196 -7760 3596 -7720
rect 3196 -8080 3236 -7760
rect 3556 -8080 3596 -7760
rect 3196 -8120 3596 -8080
rect 4208 -7760 4608 -7720
rect 4208 -8080 4248 -7760
rect 4568 -8080 4608 -7760
rect 4208 -8120 4608 -8080
rect 5220 -7760 5620 -7720
rect 5220 -8080 5260 -7760
rect 5580 -8080 5620 -7760
rect 5220 -8120 5620 -8080
rect 6232 -7760 6632 -7720
rect 6232 -8080 6272 -7760
rect 6592 -8080 6632 -7760
rect 6232 -8120 6632 -8080
rect 7244 -7760 7644 -7720
rect 7244 -8080 7284 -7760
rect 7604 -8080 7644 -7760
rect 7244 -8120 7644 -8080
rect 8256 -7760 8656 -7720
rect 8256 -8080 8296 -7760
rect 8616 -8080 8656 -7760
rect 8256 -8120 8656 -8080
rect 9268 -7760 9668 -7720
rect 9268 -8080 9308 -7760
rect 9628 -8080 9668 -7760
rect 9268 -8120 9668 -8080
rect 10280 -7760 10680 -7720
rect 10280 -8080 10320 -7760
rect 10640 -8080 10680 -7760
rect 10280 -8120 10680 -8080
rect 11292 -7760 11692 -7720
rect 11292 -8080 11332 -7760
rect 11652 -8080 11692 -7760
rect 11292 -8120 11692 -8080
rect 12304 -7760 12704 -7720
rect 12304 -8080 12344 -7760
rect 12664 -8080 12704 -7760
rect 12304 -8120 12704 -8080
rect 13316 -7760 13716 -7720
rect 13316 -8080 13356 -7760
rect 13676 -8080 13716 -7760
rect 13316 -8120 13716 -8080
rect 14328 -7760 14728 -7720
rect 14328 -8080 14368 -7760
rect 14688 -8080 14728 -7760
rect 14328 -8120 14728 -8080
rect 15340 -7760 15740 -7720
rect 15340 -8080 15380 -7760
rect 15700 -8080 15740 -7760
rect 15340 -8120 15740 -8080
rect 16352 -7760 16752 -7720
rect 16352 -8080 16392 -7760
rect 16712 -8080 16752 -7760
rect 16352 -8120 16752 -8080
rect -17044 -8480 -16644 -8440
rect -17044 -8800 -17004 -8480
rect -16684 -8800 -16644 -8480
rect -17044 -8840 -16644 -8800
rect -16032 -8480 -15632 -8440
rect -16032 -8800 -15992 -8480
rect -15672 -8800 -15632 -8480
rect -16032 -8840 -15632 -8800
rect -15020 -8480 -14620 -8440
rect -15020 -8800 -14980 -8480
rect -14660 -8800 -14620 -8480
rect -15020 -8840 -14620 -8800
rect -14008 -8480 -13608 -8440
rect -14008 -8800 -13968 -8480
rect -13648 -8800 -13608 -8480
rect -14008 -8840 -13608 -8800
rect -12996 -8480 -12596 -8440
rect -12996 -8800 -12956 -8480
rect -12636 -8800 -12596 -8480
rect -12996 -8840 -12596 -8800
rect -11984 -8480 -11584 -8440
rect -11984 -8800 -11944 -8480
rect -11624 -8800 -11584 -8480
rect -11984 -8840 -11584 -8800
rect -10972 -8480 -10572 -8440
rect -10972 -8800 -10932 -8480
rect -10612 -8800 -10572 -8480
rect -10972 -8840 -10572 -8800
rect -9960 -8480 -9560 -8440
rect -9960 -8800 -9920 -8480
rect -9600 -8800 -9560 -8480
rect -9960 -8840 -9560 -8800
rect -8948 -8480 -8548 -8440
rect -8948 -8800 -8908 -8480
rect -8588 -8800 -8548 -8480
rect -8948 -8840 -8548 -8800
rect -7936 -8480 -7536 -8440
rect -7936 -8800 -7896 -8480
rect -7576 -8800 -7536 -8480
rect -7936 -8840 -7536 -8800
rect -6924 -8480 -6524 -8440
rect -6924 -8800 -6884 -8480
rect -6564 -8800 -6524 -8480
rect -6924 -8840 -6524 -8800
rect -5912 -8480 -5512 -8440
rect -5912 -8800 -5872 -8480
rect -5552 -8800 -5512 -8480
rect -5912 -8840 -5512 -8800
rect -4900 -8480 -4500 -8440
rect -4900 -8800 -4860 -8480
rect -4540 -8800 -4500 -8480
rect -4900 -8840 -4500 -8800
rect -3888 -8480 -3488 -8440
rect -3888 -8800 -3848 -8480
rect -3528 -8800 -3488 -8480
rect -3888 -8840 -3488 -8800
rect -2876 -8480 -2476 -8440
rect -2876 -8800 -2836 -8480
rect -2516 -8800 -2476 -8480
rect -2876 -8840 -2476 -8800
rect -1864 -8480 -1464 -8440
rect -1864 -8800 -1824 -8480
rect -1504 -8800 -1464 -8480
rect -1864 -8840 -1464 -8800
rect -852 -8480 -452 -8440
rect -852 -8800 -812 -8480
rect -492 -8800 -452 -8480
rect -852 -8840 -452 -8800
rect 160 -8480 560 -8440
rect 160 -8800 200 -8480
rect 520 -8800 560 -8480
rect 160 -8840 560 -8800
rect 1172 -8480 1572 -8440
rect 1172 -8800 1212 -8480
rect 1532 -8800 1572 -8480
rect 1172 -8840 1572 -8800
rect 2184 -8480 2584 -8440
rect 2184 -8800 2224 -8480
rect 2544 -8800 2584 -8480
rect 2184 -8840 2584 -8800
rect 3196 -8480 3596 -8440
rect 3196 -8800 3236 -8480
rect 3556 -8800 3596 -8480
rect 3196 -8840 3596 -8800
rect 4208 -8480 4608 -8440
rect 4208 -8800 4248 -8480
rect 4568 -8800 4608 -8480
rect 4208 -8840 4608 -8800
rect 5220 -8480 5620 -8440
rect 5220 -8800 5260 -8480
rect 5580 -8800 5620 -8480
rect 5220 -8840 5620 -8800
rect 6232 -8480 6632 -8440
rect 6232 -8800 6272 -8480
rect 6592 -8800 6632 -8480
rect 6232 -8840 6632 -8800
rect 7244 -8480 7644 -8440
rect 7244 -8800 7284 -8480
rect 7604 -8800 7644 -8480
rect 7244 -8840 7644 -8800
rect 8256 -8480 8656 -8440
rect 8256 -8800 8296 -8480
rect 8616 -8800 8656 -8480
rect 8256 -8840 8656 -8800
rect 9268 -8480 9668 -8440
rect 9268 -8800 9308 -8480
rect 9628 -8800 9668 -8480
rect 9268 -8840 9668 -8800
rect 10280 -8480 10680 -8440
rect 10280 -8800 10320 -8480
rect 10640 -8800 10680 -8480
rect 10280 -8840 10680 -8800
rect 11292 -8480 11692 -8440
rect 11292 -8800 11332 -8480
rect 11652 -8800 11692 -8480
rect 11292 -8840 11692 -8800
rect 12304 -8480 12704 -8440
rect 12304 -8800 12344 -8480
rect 12664 -8800 12704 -8480
rect 12304 -8840 12704 -8800
rect 13316 -8480 13716 -8440
rect 13316 -8800 13356 -8480
rect 13676 -8800 13716 -8480
rect 13316 -8840 13716 -8800
rect 14328 -8480 14728 -8440
rect 14328 -8800 14368 -8480
rect 14688 -8800 14728 -8480
rect 14328 -8840 14728 -8800
rect 15340 -8480 15740 -8440
rect 15340 -8800 15380 -8480
rect 15700 -8800 15740 -8480
rect 15340 -8840 15740 -8800
rect 16352 -8480 16752 -8440
rect 16352 -8800 16392 -8480
rect 16712 -8800 16752 -8480
rect 16352 -8840 16752 -8800
rect -17044 -9200 -16644 -9160
rect -17044 -9520 -17004 -9200
rect -16684 -9520 -16644 -9200
rect -17044 -9560 -16644 -9520
rect -16032 -9200 -15632 -9160
rect -16032 -9520 -15992 -9200
rect -15672 -9520 -15632 -9200
rect -16032 -9560 -15632 -9520
rect -15020 -9200 -14620 -9160
rect -15020 -9520 -14980 -9200
rect -14660 -9520 -14620 -9200
rect -15020 -9560 -14620 -9520
rect -14008 -9200 -13608 -9160
rect -14008 -9520 -13968 -9200
rect -13648 -9520 -13608 -9200
rect -14008 -9560 -13608 -9520
rect -12996 -9200 -12596 -9160
rect -12996 -9520 -12956 -9200
rect -12636 -9520 -12596 -9200
rect -12996 -9560 -12596 -9520
rect -11984 -9200 -11584 -9160
rect -11984 -9520 -11944 -9200
rect -11624 -9520 -11584 -9200
rect -11984 -9560 -11584 -9520
rect -10972 -9200 -10572 -9160
rect -10972 -9520 -10932 -9200
rect -10612 -9520 -10572 -9200
rect -10972 -9560 -10572 -9520
rect -9960 -9200 -9560 -9160
rect -9960 -9520 -9920 -9200
rect -9600 -9520 -9560 -9200
rect -9960 -9560 -9560 -9520
rect -8948 -9200 -8548 -9160
rect -8948 -9520 -8908 -9200
rect -8588 -9520 -8548 -9200
rect -8948 -9560 -8548 -9520
rect -7936 -9200 -7536 -9160
rect -7936 -9520 -7896 -9200
rect -7576 -9520 -7536 -9200
rect -7936 -9560 -7536 -9520
rect -6924 -9200 -6524 -9160
rect -6924 -9520 -6884 -9200
rect -6564 -9520 -6524 -9200
rect -6924 -9560 -6524 -9520
rect -5912 -9200 -5512 -9160
rect -5912 -9520 -5872 -9200
rect -5552 -9520 -5512 -9200
rect -5912 -9560 -5512 -9520
rect -4900 -9200 -4500 -9160
rect -4900 -9520 -4860 -9200
rect -4540 -9520 -4500 -9200
rect -4900 -9560 -4500 -9520
rect -3888 -9200 -3488 -9160
rect -3888 -9520 -3848 -9200
rect -3528 -9520 -3488 -9200
rect -3888 -9560 -3488 -9520
rect -2876 -9200 -2476 -9160
rect -2876 -9520 -2836 -9200
rect -2516 -9520 -2476 -9200
rect -2876 -9560 -2476 -9520
rect -1864 -9200 -1464 -9160
rect -1864 -9520 -1824 -9200
rect -1504 -9520 -1464 -9200
rect -1864 -9560 -1464 -9520
rect -852 -9200 -452 -9160
rect -852 -9520 -812 -9200
rect -492 -9520 -452 -9200
rect -852 -9560 -452 -9520
rect 160 -9200 560 -9160
rect 160 -9520 200 -9200
rect 520 -9520 560 -9200
rect 160 -9560 560 -9520
rect 1172 -9200 1572 -9160
rect 1172 -9520 1212 -9200
rect 1532 -9520 1572 -9200
rect 1172 -9560 1572 -9520
rect 2184 -9200 2584 -9160
rect 2184 -9520 2224 -9200
rect 2544 -9520 2584 -9200
rect 2184 -9560 2584 -9520
rect 3196 -9200 3596 -9160
rect 3196 -9520 3236 -9200
rect 3556 -9520 3596 -9200
rect 3196 -9560 3596 -9520
rect 4208 -9200 4608 -9160
rect 4208 -9520 4248 -9200
rect 4568 -9520 4608 -9200
rect 4208 -9560 4608 -9520
rect 5220 -9200 5620 -9160
rect 5220 -9520 5260 -9200
rect 5580 -9520 5620 -9200
rect 5220 -9560 5620 -9520
rect 6232 -9200 6632 -9160
rect 6232 -9520 6272 -9200
rect 6592 -9520 6632 -9200
rect 6232 -9560 6632 -9520
rect 7244 -9200 7644 -9160
rect 7244 -9520 7284 -9200
rect 7604 -9520 7644 -9200
rect 7244 -9560 7644 -9520
rect 8256 -9200 8656 -9160
rect 8256 -9520 8296 -9200
rect 8616 -9520 8656 -9200
rect 8256 -9560 8656 -9520
rect 9268 -9200 9668 -9160
rect 9268 -9520 9308 -9200
rect 9628 -9520 9668 -9200
rect 9268 -9560 9668 -9520
rect 10280 -9200 10680 -9160
rect 10280 -9520 10320 -9200
rect 10640 -9520 10680 -9200
rect 10280 -9560 10680 -9520
rect 11292 -9200 11692 -9160
rect 11292 -9520 11332 -9200
rect 11652 -9520 11692 -9200
rect 11292 -9560 11692 -9520
rect 12304 -9200 12704 -9160
rect 12304 -9520 12344 -9200
rect 12664 -9520 12704 -9200
rect 12304 -9560 12704 -9520
rect 13316 -9200 13716 -9160
rect 13316 -9520 13356 -9200
rect 13676 -9520 13716 -9200
rect 13316 -9560 13716 -9520
rect 14328 -9200 14728 -9160
rect 14328 -9520 14368 -9200
rect 14688 -9520 14728 -9200
rect 14328 -9560 14728 -9520
rect 15340 -9200 15740 -9160
rect 15340 -9520 15380 -9200
rect 15700 -9520 15740 -9200
rect 15340 -9560 15740 -9520
rect 16352 -9200 16752 -9160
rect 16352 -9520 16392 -9200
rect 16712 -9520 16752 -9200
rect 16352 -9560 16752 -9520
rect -17044 -9920 -16644 -9880
rect -17044 -10240 -17004 -9920
rect -16684 -10240 -16644 -9920
rect -17044 -10280 -16644 -10240
rect -16032 -9920 -15632 -9880
rect -16032 -10240 -15992 -9920
rect -15672 -10240 -15632 -9920
rect -16032 -10280 -15632 -10240
rect -15020 -9920 -14620 -9880
rect -15020 -10240 -14980 -9920
rect -14660 -10240 -14620 -9920
rect -15020 -10280 -14620 -10240
rect -14008 -9920 -13608 -9880
rect -14008 -10240 -13968 -9920
rect -13648 -10240 -13608 -9920
rect -14008 -10280 -13608 -10240
rect -12996 -9920 -12596 -9880
rect -12996 -10240 -12956 -9920
rect -12636 -10240 -12596 -9920
rect -12996 -10280 -12596 -10240
rect -11984 -9920 -11584 -9880
rect -11984 -10240 -11944 -9920
rect -11624 -10240 -11584 -9920
rect -11984 -10280 -11584 -10240
rect -10972 -9920 -10572 -9880
rect -10972 -10240 -10932 -9920
rect -10612 -10240 -10572 -9920
rect -10972 -10280 -10572 -10240
rect -9960 -9920 -9560 -9880
rect -9960 -10240 -9920 -9920
rect -9600 -10240 -9560 -9920
rect -9960 -10280 -9560 -10240
rect -8948 -9920 -8548 -9880
rect -8948 -10240 -8908 -9920
rect -8588 -10240 -8548 -9920
rect -8948 -10280 -8548 -10240
rect -7936 -9920 -7536 -9880
rect -7936 -10240 -7896 -9920
rect -7576 -10240 -7536 -9920
rect -7936 -10280 -7536 -10240
rect -6924 -9920 -6524 -9880
rect -6924 -10240 -6884 -9920
rect -6564 -10240 -6524 -9920
rect -6924 -10280 -6524 -10240
rect -5912 -9920 -5512 -9880
rect -5912 -10240 -5872 -9920
rect -5552 -10240 -5512 -9920
rect -5912 -10280 -5512 -10240
rect -4900 -9920 -4500 -9880
rect -4900 -10240 -4860 -9920
rect -4540 -10240 -4500 -9920
rect -4900 -10280 -4500 -10240
rect -3888 -9920 -3488 -9880
rect -3888 -10240 -3848 -9920
rect -3528 -10240 -3488 -9920
rect -3888 -10280 -3488 -10240
rect -2876 -9920 -2476 -9880
rect -2876 -10240 -2836 -9920
rect -2516 -10240 -2476 -9920
rect -2876 -10280 -2476 -10240
rect -1864 -9920 -1464 -9880
rect -1864 -10240 -1824 -9920
rect -1504 -10240 -1464 -9920
rect -1864 -10280 -1464 -10240
rect -852 -9920 -452 -9880
rect -852 -10240 -812 -9920
rect -492 -10240 -452 -9920
rect -852 -10280 -452 -10240
rect 160 -9920 560 -9880
rect 160 -10240 200 -9920
rect 520 -10240 560 -9920
rect 160 -10280 560 -10240
rect 1172 -9920 1572 -9880
rect 1172 -10240 1212 -9920
rect 1532 -10240 1572 -9920
rect 1172 -10280 1572 -10240
rect 2184 -9920 2584 -9880
rect 2184 -10240 2224 -9920
rect 2544 -10240 2584 -9920
rect 2184 -10280 2584 -10240
rect 3196 -9920 3596 -9880
rect 3196 -10240 3236 -9920
rect 3556 -10240 3596 -9920
rect 3196 -10280 3596 -10240
rect 4208 -9920 4608 -9880
rect 4208 -10240 4248 -9920
rect 4568 -10240 4608 -9920
rect 4208 -10280 4608 -10240
rect 5220 -9920 5620 -9880
rect 5220 -10240 5260 -9920
rect 5580 -10240 5620 -9920
rect 5220 -10280 5620 -10240
rect 6232 -9920 6632 -9880
rect 6232 -10240 6272 -9920
rect 6592 -10240 6632 -9920
rect 6232 -10280 6632 -10240
rect 7244 -9920 7644 -9880
rect 7244 -10240 7284 -9920
rect 7604 -10240 7644 -9920
rect 7244 -10280 7644 -10240
rect 8256 -9920 8656 -9880
rect 8256 -10240 8296 -9920
rect 8616 -10240 8656 -9920
rect 8256 -10280 8656 -10240
rect 9268 -9920 9668 -9880
rect 9268 -10240 9308 -9920
rect 9628 -10240 9668 -9920
rect 9268 -10280 9668 -10240
rect 10280 -9920 10680 -9880
rect 10280 -10240 10320 -9920
rect 10640 -10240 10680 -9920
rect 10280 -10280 10680 -10240
rect 11292 -9920 11692 -9880
rect 11292 -10240 11332 -9920
rect 11652 -10240 11692 -9920
rect 11292 -10280 11692 -10240
rect 12304 -9920 12704 -9880
rect 12304 -10240 12344 -9920
rect 12664 -10240 12704 -9920
rect 12304 -10280 12704 -10240
rect 13316 -9920 13716 -9880
rect 13316 -10240 13356 -9920
rect 13676 -10240 13716 -9920
rect 13316 -10280 13716 -10240
rect 14328 -9920 14728 -9880
rect 14328 -10240 14368 -9920
rect 14688 -10240 14728 -9920
rect 14328 -10280 14728 -10240
rect 15340 -9920 15740 -9880
rect 15340 -10240 15380 -9920
rect 15700 -10240 15740 -9920
rect 15340 -10280 15740 -10240
rect 16352 -9920 16752 -9880
rect 16352 -10240 16392 -9920
rect 16712 -10240 16752 -9920
rect 16352 -10280 16752 -10240
rect -17044 -10640 -16644 -10600
rect -17044 -10960 -17004 -10640
rect -16684 -10960 -16644 -10640
rect -17044 -11000 -16644 -10960
rect -16032 -10640 -15632 -10600
rect -16032 -10960 -15992 -10640
rect -15672 -10960 -15632 -10640
rect -16032 -11000 -15632 -10960
rect -15020 -10640 -14620 -10600
rect -15020 -10960 -14980 -10640
rect -14660 -10960 -14620 -10640
rect -15020 -11000 -14620 -10960
rect -14008 -10640 -13608 -10600
rect -14008 -10960 -13968 -10640
rect -13648 -10960 -13608 -10640
rect -14008 -11000 -13608 -10960
rect -12996 -10640 -12596 -10600
rect -12996 -10960 -12956 -10640
rect -12636 -10960 -12596 -10640
rect -12996 -11000 -12596 -10960
rect -11984 -10640 -11584 -10600
rect -11984 -10960 -11944 -10640
rect -11624 -10960 -11584 -10640
rect -11984 -11000 -11584 -10960
rect -10972 -10640 -10572 -10600
rect -10972 -10960 -10932 -10640
rect -10612 -10960 -10572 -10640
rect -10972 -11000 -10572 -10960
rect -9960 -10640 -9560 -10600
rect -9960 -10960 -9920 -10640
rect -9600 -10960 -9560 -10640
rect -9960 -11000 -9560 -10960
rect -8948 -10640 -8548 -10600
rect -8948 -10960 -8908 -10640
rect -8588 -10960 -8548 -10640
rect -8948 -11000 -8548 -10960
rect -7936 -10640 -7536 -10600
rect -7936 -10960 -7896 -10640
rect -7576 -10960 -7536 -10640
rect -7936 -11000 -7536 -10960
rect -6924 -10640 -6524 -10600
rect -6924 -10960 -6884 -10640
rect -6564 -10960 -6524 -10640
rect -6924 -11000 -6524 -10960
rect -5912 -10640 -5512 -10600
rect -5912 -10960 -5872 -10640
rect -5552 -10960 -5512 -10640
rect -5912 -11000 -5512 -10960
rect -4900 -10640 -4500 -10600
rect -4900 -10960 -4860 -10640
rect -4540 -10960 -4500 -10640
rect -4900 -11000 -4500 -10960
rect -3888 -10640 -3488 -10600
rect -3888 -10960 -3848 -10640
rect -3528 -10960 -3488 -10640
rect -3888 -11000 -3488 -10960
rect -2876 -10640 -2476 -10600
rect -2876 -10960 -2836 -10640
rect -2516 -10960 -2476 -10640
rect -2876 -11000 -2476 -10960
rect -1864 -10640 -1464 -10600
rect -1864 -10960 -1824 -10640
rect -1504 -10960 -1464 -10640
rect -1864 -11000 -1464 -10960
rect -852 -10640 -452 -10600
rect -852 -10960 -812 -10640
rect -492 -10960 -452 -10640
rect -852 -11000 -452 -10960
rect 160 -10640 560 -10600
rect 160 -10960 200 -10640
rect 520 -10960 560 -10640
rect 160 -11000 560 -10960
rect 1172 -10640 1572 -10600
rect 1172 -10960 1212 -10640
rect 1532 -10960 1572 -10640
rect 1172 -11000 1572 -10960
rect 2184 -10640 2584 -10600
rect 2184 -10960 2224 -10640
rect 2544 -10960 2584 -10640
rect 2184 -11000 2584 -10960
rect 3196 -10640 3596 -10600
rect 3196 -10960 3236 -10640
rect 3556 -10960 3596 -10640
rect 3196 -11000 3596 -10960
rect 4208 -10640 4608 -10600
rect 4208 -10960 4248 -10640
rect 4568 -10960 4608 -10640
rect 4208 -11000 4608 -10960
rect 5220 -10640 5620 -10600
rect 5220 -10960 5260 -10640
rect 5580 -10960 5620 -10640
rect 5220 -11000 5620 -10960
rect 6232 -10640 6632 -10600
rect 6232 -10960 6272 -10640
rect 6592 -10960 6632 -10640
rect 6232 -11000 6632 -10960
rect 7244 -10640 7644 -10600
rect 7244 -10960 7284 -10640
rect 7604 -10960 7644 -10640
rect 7244 -11000 7644 -10960
rect 8256 -10640 8656 -10600
rect 8256 -10960 8296 -10640
rect 8616 -10960 8656 -10640
rect 8256 -11000 8656 -10960
rect 9268 -10640 9668 -10600
rect 9268 -10960 9308 -10640
rect 9628 -10960 9668 -10640
rect 9268 -11000 9668 -10960
rect 10280 -10640 10680 -10600
rect 10280 -10960 10320 -10640
rect 10640 -10960 10680 -10640
rect 10280 -11000 10680 -10960
rect 11292 -10640 11692 -10600
rect 11292 -10960 11332 -10640
rect 11652 -10960 11692 -10640
rect 11292 -11000 11692 -10960
rect 12304 -10640 12704 -10600
rect 12304 -10960 12344 -10640
rect 12664 -10960 12704 -10640
rect 12304 -11000 12704 -10960
rect 13316 -10640 13716 -10600
rect 13316 -10960 13356 -10640
rect 13676 -10960 13716 -10640
rect 13316 -11000 13716 -10960
rect 14328 -10640 14728 -10600
rect 14328 -10960 14368 -10640
rect 14688 -10960 14728 -10640
rect 14328 -11000 14728 -10960
rect 15340 -10640 15740 -10600
rect 15340 -10960 15380 -10640
rect 15700 -10960 15740 -10640
rect 15340 -11000 15740 -10960
rect 16352 -10640 16752 -10600
rect 16352 -10960 16392 -10640
rect 16712 -10960 16752 -10640
rect 16352 -11000 16752 -10960
rect -17044 -11360 -16644 -11320
rect -17044 -11680 -17004 -11360
rect -16684 -11680 -16644 -11360
rect -17044 -11720 -16644 -11680
rect -16032 -11360 -15632 -11320
rect -16032 -11680 -15992 -11360
rect -15672 -11680 -15632 -11360
rect -16032 -11720 -15632 -11680
rect -15020 -11360 -14620 -11320
rect -15020 -11680 -14980 -11360
rect -14660 -11680 -14620 -11360
rect -15020 -11720 -14620 -11680
rect -14008 -11360 -13608 -11320
rect -14008 -11680 -13968 -11360
rect -13648 -11680 -13608 -11360
rect -14008 -11720 -13608 -11680
rect -12996 -11360 -12596 -11320
rect -12996 -11680 -12956 -11360
rect -12636 -11680 -12596 -11360
rect -12996 -11720 -12596 -11680
rect -11984 -11360 -11584 -11320
rect -11984 -11680 -11944 -11360
rect -11624 -11680 -11584 -11360
rect -11984 -11720 -11584 -11680
rect -10972 -11360 -10572 -11320
rect -10972 -11680 -10932 -11360
rect -10612 -11680 -10572 -11360
rect -10972 -11720 -10572 -11680
rect -9960 -11360 -9560 -11320
rect -9960 -11680 -9920 -11360
rect -9600 -11680 -9560 -11360
rect -9960 -11720 -9560 -11680
rect -8948 -11360 -8548 -11320
rect -8948 -11680 -8908 -11360
rect -8588 -11680 -8548 -11360
rect -8948 -11720 -8548 -11680
rect -7936 -11360 -7536 -11320
rect -7936 -11680 -7896 -11360
rect -7576 -11680 -7536 -11360
rect -7936 -11720 -7536 -11680
rect -6924 -11360 -6524 -11320
rect -6924 -11680 -6884 -11360
rect -6564 -11680 -6524 -11360
rect -6924 -11720 -6524 -11680
rect -5912 -11360 -5512 -11320
rect -5912 -11680 -5872 -11360
rect -5552 -11680 -5512 -11360
rect -5912 -11720 -5512 -11680
rect -4900 -11360 -4500 -11320
rect -4900 -11680 -4860 -11360
rect -4540 -11680 -4500 -11360
rect -4900 -11720 -4500 -11680
rect -3888 -11360 -3488 -11320
rect -3888 -11680 -3848 -11360
rect -3528 -11680 -3488 -11360
rect -3888 -11720 -3488 -11680
rect -2876 -11360 -2476 -11320
rect -2876 -11680 -2836 -11360
rect -2516 -11680 -2476 -11360
rect -2876 -11720 -2476 -11680
rect -1864 -11360 -1464 -11320
rect -1864 -11680 -1824 -11360
rect -1504 -11680 -1464 -11360
rect -1864 -11720 -1464 -11680
rect -852 -11360 -452 -11320
rect -852 -11680 -812 -11360
rect -492 -11680 -452 -11360
rect -852 -11720 -452 -11680
rect 160 -11360 560 -11320
rect 160 -11680 200 -11360
rect 520 -11680 560 -11360
rect 160 -11720 560 -11680
rect 1172 -11360 1572 -11320
rect 1172 -11680 1212 -11360
rect 1532 -11680 1572 -11360
rect 1172 -11720 1572 -11680
rect 2184 -11360 2584 -11320
rect 2184 -11680 2224 -11360
rect 2544 -11680 2584 -11360
rect 2184 -11720 2584 -11680
rect 3196 -11360 3596 -11320
rect 3196 -11680 3236 -11360
rect 3556 -11680 3596 -11360
rect 3196 -11720 3596 -11680
rect 4208 -11360 4608 -11320
rect 4208 -11680 4248 -11360
rect 4568 -11680 4608 -11360
rect 4208 -11720 4608 -11680
rect 5220 -11360 5620 -11320
rect 5220 -11680 5260 -11360
rect 5580 -11680 5620 -11360
rect 5220 -11720 5620 -11680
rect 6232 -11360 6632 -11320
rect 6232 -11680 6272 -11360
rect 6592 -11680 6632 -11360
rect 6232 -11720 6632 -11680
rect 7244 -11360 7644 -11320
rect 7244 -11680 7284 -11360
rect 7604 -11680 7644 -11360
rect 7244 -11720 7644 -11680
rect 8256 -11360 8656 -11320
rect 8256 -11680 8296 -11360
rect 8616 -11680 8656 -11360
rect 8256 -11720 8656 -11680
rect 9268 -11360 9668 -11320
rect 9268 -11680 9308 -11360
rect 9628 -11680 9668 -11360
rect 9268 -11720 9668 -11680
rect 10280 -11360 10680 -11320
rect 10280 -11680 10320 -11360
rect 10640 -11680 10680 -11360
rect 10280 -11720 10680 -11680
rect 11292 -11360 11692 -11320
rect 11292 -11680 11332 -11360
rect 11652 -11680 11692 -11360
rect 11292 -11720 11692 -11680
rect 12304 -11360 12704 -11320
rect 12304 -11680 12344 -11360
rect 12664 -11680 12704 -11360
rect 12304 -11720 12704 -11680
rect 13316 -11360 13716 -11320
rect 13316 -11680 13356 -11360
rect 13676 -11680 13716 -11360
rect 13316 -11720 13716 -11680
rect 14328 -11360 14728 -11320
rect 14328 -11680 14368 -11360
rect 14688 -11680 14728 -11360
rect 14328 -11720 14728 -11680
rect 15340 -11360 15740 -11320
rect 15340 -11680 15380 -11360
rect 15700 -11680 15740 -11360
rect 15340 -11720 15740 -11680
rect 16352 -11360 16752 -11320
rect 16352 -11680 16392 -11360
rect 16712 -11680 16752 -11360
rect 16352 -11720 16752 -11680
<< mimcapcontact >>
rect -17004 11360 -16684 11680
rect -15992 11360 -15672 11680
rect -14980 11360 -14660 11680
rect -13968 11360 -13648 11680
rect -12956 11360 -12636 11680
rect -11944 11360 -11624 11680
rect -10932 11360 -10612 11680
rect -9920 11360 -9600 11680
rect -8908 11360 -8588 11680
rect -7896 11360 -7576 11680
rect -6884 11360 -6564 11680
rect -5872 11360 -5552 11680
rect -4860 11360 -4540 11680
rect -3848 11360 -3528 11680
rect -2836 11360 -2516 11680
rect -1824 11360 -1504 11680
rect -812 11360 -492 11680
rect 200 11360 520 11680
rect 1212 11360 1532 11680
rect 2224 11360 2544 11680
rect 3236 11360 3556 11680
rect 4248 11360 4568 11680
rect 5260 11360 5580 11680
rect 6272 11360 6592 11680
rect 7284 11360 7604 11680
rect 8296 11360 8616 11680
rect 9308 11360 9628 11680
rect 10320 11360 10640 11680
rect 11332 11360 11652 11680
rect 12344 11360 12664 11680
rect 13356 11360 13676 11680
rect 14368 11360 14688 11680
rect 15380 11360 15700 11680
rect 16392 11360 16712 11680
rect -17004 10640 -16684 10960
rect -15992 10640 -15672 10960
rect -14980 10640 -14660 10960
rect -13968 10640 -13648 10960
rect -12956 10640 -12636 10960
rect -11944 10640 -11624 10960
rect -10932 10640 -10612 10960
rect -9920 10640 -9600 10960
rect -8908 10640 -8588 10960
rect -7896 10640 -7576 10960
rect -6884 10640 -6564 10960
rect -5872 10640 -5552 10960
rect -4860 10640 -4540 10960
rect -3848 10640 -3528 10960
rect -2836 10640 -2516 10960
rect -1824 10640 -1504 10960
rect -812 10640 -492 10960
rect 200 10640 520 10960
rect 1212 10640 1532 10960
rect 2224 10640 2544 10960
rect 3236 10640 3556 10960
rect 4248 10640 4568 10960
rect 5260 10640 5580 10960
rect 6272 10640 6592 10960
rect 7284 10640 7604 10960
rect 8296 10640 8616 10960
rect 9308 10640 9628 10960
rect 10320 10640 10640 10960
rect 11332 10640 11652 10960
rect 12344 10640 12664 10960
rect 13356 10640 13676 10960
rect 14368 10640 14688 10960
rect 15380 10640 15700 10960
rect 16392 10640 16712 10960
rect -17004 9920 -16684 10240
rect -15992 9920 -15672 10240
rect -14980 9920 -14660 10240
rect -13968 9920 -13648 10240
rect -12956 9920 -12636 10240
rect -11944 9920 -11624 10240
rect -10932 9920 -10612 10240
rect -9920 9920 -9600 10240
rect -8908 9920 -8588 10240
rect -7896 9920 -7576 10240
rect -6884 9920 -6564 10240
rect -5872 9920 -5552 10240
rect -4860 9920 -4540 10240
rect -3848 9920 -3528 10240
rect -2836 9920 -2516 10240
rect -1824 9920 -1504 10240
rect -812 9920 -492 10240
rect 200 9920 520 10240
rect 1212 9920 1532 10240
rect 2224 9920 2544 10240
rect 3236 9920 3556 10240
rect 4248 9920 4568 10240
rect 5260 9920 5580 10240
rect 6272 9920 6592 10240
rect 7284 9920 7604 10240
rect 8296 9920 8616 10240
rect 9308 9920 9628 10240
rect 10320 9920 10640 10240
rect 11332 9920 11652 10240
rect 12344 9920 12664 10240
rect 13356 9920 13676 10240
rect 14368 9920 14688 10240
rect 15380 9920 15700 10240
rect 16392 9920 16712 10240
rect -17004 9200 -16684 9520
rect -15992 9200 -15672 9520
rect -14980 9200 -14660 9520
rect -13968 9200 -13648 9520
rect -12956 9200 -12636 9520
rect -11944 9200 -11624 9520
rect -10932 9200 -10612 9520
rect -9920 9200 -9600 9520
rect -8908 9200 -8588 9520
rect -7896 9200 -7576 9520
rect -6884 9200 -6564 9520
rect -5872 9200 -5552 9520
rect -4860 9200 -4540 9520
rect -3848 9200 -3528 9520
rect -2836 9200 -2516 9520
rect -1824 9200 -1504 9520
rect -812 9200 -492 9520
rect 200 9200 520 9520
rect 1212 9200 1532 9520
rect 2224 9200 2544 9520
rect 3236 9200 3556 9520
rect 4248 9200 4568 9520
rect 5260 9200 5580 9520
rect 6272 9200 6592 9520
rect 7284 9200 7604 9520
rect 8296 9200 8616 9520
rect 9308 9200 9628 9520
rect 10320 9200 10640 9520
rect 11332 9200 11652 9520
rect 12344 9200 12664 9520
rect 13356 9200 13676 9520
rect 14368 9200 14688 9520
rect 15380 9200 15700 9520
rect 16392 9200 16712 9520
rect -17004 8480 -16684 8800
rect -15992 8480 -15672 8800
rect -14980 8480 -14660 8800
rect -13968 8480 -13648 8800
rect -12956 8480 -12636 8800
rect -11944 8480 -11624 8800
rect -10932 8480 -10612 8800
rect -9920 8480 -9600 8800
rect -8908 8480 -8588 8800
rect -7896 8480 -7576 8800
rect -6884 8480 -6564 8800
rect -5872 8480 -5552 8800
rect -4860 8480 -4540 8800
rect -3848 8480 -3528 8800
rect -2836 8480 -2516 8800
rect -1824 8480 -1504 8800
rect -812 8480 -492 8800
rect 200 8480 520 8800
rect 1212 8480 1532 8800
rect 2224 8480 2544 8800
rect 3236 8480 3556 8800
rect 4248 8480 4568 8800
rect 5260 8480 5580 8800
rect 6272 8480 6592 8800
rect 7284 8480 7604 8800
rect 8296 8480 8616 8800
rect 9308 8480 9628 8800
rect 10320 8480 10640 8800
rect 11332 8480 11652 8800
rect 12344 8480 12664 8800
rect 13356 8480 13676 8800
rect 14368 8480 14688 8800
rect 15380 8480 15700 8800
rect 16392 8480 16712 8800
rect -17004 7760 -16684 8080
rect -15992 7760 -15672 8080
rect -14980 7760 -14660 8080
rect -13968 7760 -13648 8080
rect -12956 7760 -12636 8080
rect -11944 7760 -11624 8080
rect -10932 7760 -10612 8080
rect -9920 7760 -9600 8080
rect -8908 7760 -8588 8080
rect -7896 7760 -7576 8080
rect -6884 7760 -6564 8080
rect -5872 7760 -5552 8080
rect -4860 7760 -4540 8080
rect -3848 7760 -3528 8080
rect -2836 7760 -2516 8080
rect -1824 7760 -1504 8080
rect -812 7760 -492 8080
rect 200 7760 520 8080
rect 1212 7760 1532 8080
rect 2224 7760 2544 8080
rect 3236 7760 3556 8080
rect 4248 7760 4568 8080
rect 5260 7760 5580 8080
rect 6272 7760 6592 8080
rect 7284 7760 7604 8080
rect 8296 7760 8616 8080
rect 9308 7760 9628 8080
rect 10320 7760 10640 8080
rect 11332 7760 11652 8080
rect 12344 7760 12664 8080
rect 13356 7760 13676 8080
rect 14368 7760 14688 8080
rect 15380 7760 15700 8080
rect 16392 7760 16712 8080
rect -17004 7040 -16684 7360
rect -15992 7040 -15672 7360
rect -14980 7040 -14660 7360
rect -13968 7040 -13648 7360
rect -12956 7040 -12636 7360
rect -11944 7040 -11624 7360
rect -10932 7040 -10612 7360
rect -9920 7040 -9600 7360
rect -8908 7040 -8588 7360
rect -7896 7040 -7576 7360
rect -6884 7040 -6564 7360
rect -5872 7040 -5552 7360
rect -4860 7040 -4540 7360
rect -3848 7040 -3528 7360
rect -2836 7040 -2516 7360
rect -1824 7040 -1504 7360
rect -812 7040 -492 7360
rect 200 7040 520 7360
rect 1212 7040 1532 7360
rect 2224 7040 2544 7360
rect 3236 7040 3556 7360
rect 4248 7040 4568 7360
rect 5260 7040 5580 7360
rect 6272 7040 6592 7360
rect 7284 7040 7604 7360
rect 8296 7040 8616 7360
rect 9308 7040 9628 7360
rect 10320 7040 10640 7360
rect 11332 7040 11652 7360
rect 12344 7040 12664 7360
rect 13356 7040 13676 7360
rect 14368 7040 14688 7360
rect 15380 7040 15700 7360
rect 16392 7040 16712 7360
rect -17004 6320 -16684 6640
rect -15992 6320 -15672 6640
rect -14980 6320 -14660 6640
rect -13968 6320 -13648 6640
rect -12956 6320 -12636 6640
rect -11944 6320 -11624 6640
rect -10932 6320 -10612 6640
rect -9920 6320 -9600 6640
rect -8908 6320 -8588 6640
rect -7896 6320 -7576 6640
rect -6884 6320 -6564 6640
rect -5872 6320 -5552 6640
rect -4860 6320 -4540 6640
rect -3848 6320 -3528 6640
rect -2836 6320 -2516 6640
rect -1824 6320 -1504 6640
rect -812 6320 -492 6640
rect 200 6320 520 6640
rect 1212 6320 1532 6640
rect 2224 6320 2544 6640
rect 3236 6320 3556 6640
rect 4248 6320 4568 6640
rect 5260 6320 5580 6640
rect 6272 6320 6592 6640
rect 7284 6320 7604 6640
rect 8296 6320 8616 6640
rect 9308 6320 9628 6640
rect 10320 6320 10640 6640
rect 11332 6320 11652 6640
rect 12344 6320 12664 6640
rect 13356 6320 13676 6640
rect 14368 6320 14688 6640
rect 15380 6320 15700 6640
rect 16392 6320 16712 6640
rect -17004 5600 -16684 5920
rect -15992 5600 -15672 5920
rect -14980 5600 -14660 5920
rect -13968 5600 -13648 5920
rect -12956 5600 -12636 5920
rect -11944 5600 -11624 5920
rect -10932 5600 -10612 5920
rect -9920 5600 -9600 5920
rect -8908 5600 -8588 5920
rect -7896 5600 -7576 5920
rect -6884 5600 -6564 5920
rect -5872 5600 -5552 5920
rect -4860 5600 -4540 5920
rect -3848 5600 -3528 5920
rect -2836 5600 -2516 5920
rect -1824 5600 -1504 5920
rect -812 5600 -492 5920
rect 200 5600 520 5920
rect 1212 5600 1532 5920
rect 2224 5600 2544 5920
rect 3236 5600 3556 5920
rect 4248 5600 4568 5920
rect 5260 5600 5580 5920
rect 6272 5600 6592 5920
rect 7284 5600 7604 5920
rect 8296 5600 8616 5920
rect 9308 5600 9628 5920
rect 10320 5600 10640 5920
rect 11332 5600 11652 5920
rect 12344 5600 12664 5920
rect 13356 5600 13676 5920
rect 14368 5600 14688 5920
rect 15380 5600 15700 5920
rect 16392 5600 16712 5920
rect -17004 4880 -16684 5200
rect -15992 4880 -15672 5200
rect -14980 4880 -14660 5200
rect -13968 4880 -13648 5200
rect -12956 4880 -12636 5200
rect -11944 4880 -11624 5200
rect -10932 4880 -10612 5200
rect -9920 4880 -9600 5200
rect -8908 4880 -8588 5200
rect -7896 4880 -7576 5200
rect -6884 4880 -6564 5200
rect -5872 4880 -5552 5200
rect -4860 4880 -4540 5200
rect -3848 4880 -3528 5200
rect -2836 4880 -2516 5200
rect -1824 4880 -1504 5200
rect -812 4880 -492 5200
rect 200 4880 520 5200
rect 1212 4880 1532 5200
rect 2224 4880 2544 5200
rect 3236 4880 3556 5200
rect 4248 4880 4568 5200
rect 5260 4880 5580 5200
rect 6272 4880 6592 5200
rect 7284 4880 7604 5200
rect 8296 4880 8616 5200
rect 9308 4880 9628 5200
rect 10320 4880 10640 5200
rect 11332 4880 11652 5200
rect 12344 4880 12664 5200
rect 13356 4880 13676 5200
rect 14368 4880 14688 5200
rect 15380 4880 15700 5200
rect 16392 4880 16712 5200
rect -17004 4160 -16684 4480
rect -15992 4160 -15672 4480
rect -14980 4160 -14660 4480
rect -13968 4160 -13648 4480
rect -12956 4160 -12636 4480
rect -11944 4160 -11624 4480
rect -10932 4160 -10612 4480
rect -9920 4160 -9600 4480
rect -8908 4160 -8588 4480
rect -7896 4160 -7576 4480
rect -6884 4160 -6564 4480
rect -5872 4160 -5552 4480
rect -4860 4160 -4540 4480
rect -3848 4160 -3528 4480
rect -2836 4160 -2516 4480
rect -1824 4160 -1504 4480
rect -812 4160 -492 4480
rect 200 4160 520 4480
rect 1212 4160 1532 4480
rect 2224 4160 2544 4480
rect 3236 4160 3556 4480
rect 4248 4160 4568 4480
rect 5260 4160 5580 4480
rect 6272 4160 6592 4480
rect 7284 4160 7604 4480
rect 8296 4160 8616 4480
rect 9308 4160 9628 4480
rect 10320 4160 10640 4480
rect 11332 4160 11652 4480
rect 12344 4160 12664 4480
rect 13356 4160 13676 4480
rect 14368 4160 14688 4480
rect 15380 4160 15700 4480
rect 16392 4160 16712 4480
rect -17004 3440 -16684 3760
rect -15992 3440 -15672 3760
rect -14980 3440 -14660 3760
rect -13968 3440 -13648 3760
rect -12956 3440 -12636 3760
rect -11944 3440 -11624 3760
rect -10932 3440 -10612 3760
rect -9920 3440 -9600 3760
rect -8908 3440 -8588 3760
rect -7896 3440 -7576 3760
rect -6884 3440 -6564 3760
rect -5872 3440 -5552 3760
rect -4860 3440 -4540 3760
rect -3848 3440 -3528 3760
rect -2836 3440 -2516 3760
rect -1824 3440 -1504 3760
rect -812 3440 -492 3760
rect 200 3440 520 3760
rect 1212 3440 1532 3760
rect 2224 3440 2544 3760
rect 3236 3440 3556 3760
rect 4248 3440 4568 3760
rect 5260 3440 5580 3760
rect 6272 3440 6592 3760
rect 7284 3440 7604 3760
rect 8296 3440 8616 3760
rect 9308 3440 9628 3760
rect 10320 3440 10640 3760
rect 11332 3440 11652 3760
rect 12344 3440 12664 3760
rect 13356 3440 13676 3760
rect 14368 3440 14688 3760
rect 15380 3440 15700 3760
rect 16392 3440 16712 3760
rect -17004 2720 -16684 3040
rect -15992 2720 -15672 3040
rect -14980 2720 -14660 3040
rect -13968 2720 -13648 3040
rect -12956 2720 -12636 3040
rect -11944 2720 -11624 3040
rect -10932 2720 -10612 3040
rect -9920 2720 -9600 3040
rect -8908 2720 -8588 3040
rect -7896 2720 -7576 3040
rect -6884 2720 -6564 3040
rect -5872 2720 -5552 3040
rect -4860 2720 -4540 3040
rect -3848 2720 -3528 3040
rect -2836 2720 -2516 3040
rect -1824 2720 -1504 3040
rect -812 2720 -492 3040
rect 200 2720 520 3040
rect 1212 2720 1532 3040
rect 2224 2720 2544 3040
rect 3236 2720 3556 3040
rect 4248 2720 4568 3040
rect 5260 2720 5580 3040
rect 6272 2720 6592 3040
rect 7284 2720 7604 3040
rect 8296 2720 8616 3040
rect 9308 2720 9628 3040
rect 10320 2720 10640 3040
rect 11332 2720 11652 3040
rect 12344 2720 12664 3040
rect 13356 2720 13676 3040
rect 14368 2720 14688 3040
rect 15380 2720 15700 3040
rect 16392 2720 16712 3040
rect -17004 2000 -16684 2320
rect -15992 2000 -15672 2320
rect -14980 2000 -14660 2320
rect -13968 2000 -13648 2320
rect -12956 2000 -12636 2320
rect -11944 2000 -11624 2320
rect -10932 2000 -10612 2320
rect -9920 2000 -9600 2320
rect -8908 2000 -8588 2320
rect -7896 2000 -7576 2320
rect -6884 2000 -6564 2320
rect -5872 2000 -5552 2320
rect -4860 2000 -4540 2320
rect -3848 2000 -3528 2320
rect -2836 2000 -2516 2320
rect -1824 2000 -1504 2320
rect -812 2000 -492 2320
rect 200 2000 520 2320
rect 1212 2000 1532 2320
rect 2224 2000 2544 2320
rect 3236 2000 3556 2320
rect 4248 2000 4568 2320
rect 5260 2000 5580 2320
rect 6272 2000 6592 2320
rect 7284 2000 7604 2320
rect 8296 2000 8616 2320
rect 9308 2000 9628 2320
rect 10320 2000 10640 2320
rect 11332 2000 11652 2320
rect 12344 2000 12664 2320
rect 13356 2000 13676 2320
rect 14368 2000 14688 2320
rect 15380 2000 15700 2320
rect 16392 2000 16712 2320
rect -17004 1280 -16684 1600
rect -15992 1280 -15672 1600
rect -14980 1280 -14660 1600
rect -13968 1280 -13648 1600
rect -12956 1280 -12636 1600
rect -11944 1280 -11624 1600
rect -10932 1280 -10612 1600
rect -9920 1280 -9600 1600
rect -8908 1280 -8588 1600
rect -7896 1280 -7576 1600
rect -6884 1280 -6564 1600
rect -5872 1280 -5552 1600
rect -4860 1280 -4540 1600
rect -3848 1280 -3528 1600
rect -2836 1280 -2516 1600
rect -1824 1280 -1504 1600
rect -812 1280 -492 1600
rect 200 1280 520 1600
rect 1212 1280 1532 1600
rect 2224 1280 2544 1600
rect 3236 1280 3556 1600
rect 4248 1280 4568 1600
rect 5260 1280 5580 1600
rect 6272 1280 6592 1600
rect 7284 1280 7604 1600
rect 8296 1280 8616 1600
rect 9308 1280 9628 1600
rect 10320 1280 10640 1600
rect 11332 1280 11652 1600
rect 12344 1280 12664 1600
rect 13356 1280 13676 1600
rect 14368 1280 14688 1600
rect 15380 1280 15700 1600
rect 16392 1280 16712 1600
rect -17004 560 -16684 880
rect -15992 560 -15672 880
rect -14980 560 -14660 880
rect -13968 560 -13648 880
rect -12956 560 -12636 880
rect -11944 560 -11624 880
rect -10932 560 -10612 880
rect -9920 560 -9600 880
rect -8908 560 -8588 880
rect -7896 560 -7576 880
rect -6884 560 -6564 880
rect -5872 560 -5552 880
rect -4860 560 -4540 880
rect -3848 560 -3528 880
rect -2836 560 -2516 880
rect -1824 560 -1504 880
rect -812 560 -492 880
rect 200 560 520 880
rect 1212 560 1532 880
rect 2224 560 2544 880
rect 3236 560 3556 880
rect 4248 560 4568 880
rect 5260 560 5580 880
rect 6272 560 6592 880
rect 7284 560 7604 880
rect 8296 560 8616 880
rect 9308 560 9628 880
rect 10320 560 10640 880
rect 11332 560 11652 880
rect 12344 560 12664 880
rect 13356 560 13676 880
rect 14368 560 14688 880
rect 15380 560 15700 880
rect 16392 560 16712 880
rect -17004 -160 -16684 160
rect -15992 -160 -15672 160
rect -14980 -160 -14660 160
rect -13968 -160 -13648 160
rect -12956 -160 -12636 160
rect -11944 -160 -11624 160
rect -10932 -160 -10612 160
rect -9920 -160 -9600 160
rect -8908 -160 -8588 160
rect -7896 -160 -7576 160
rect -6884 -160 -6564 160
rect -5872 -160 -5552 160
rect -4860 -160 -4540 160
rect -3848 -160 -3528 160
rect -2836 -160 -2516 160
rect -1824 -160 -1504 160
rect -812 -160 -492 160
rect 200 -160 520 160
rect 1212 -160 1532 160
rect 2224 -160 2544 160
rect 3236 -160 3556 160
rect 4248 -160 4568 160
rect 5260 -160 5580 160
rect 6272 -160 6592 160
rect 7284 -160 7604 160
rect 8296 -160 8616 160
rect 9308 -160 9628 160
rect 10320 -160 10640 160
rect 11332 -160 11652 160
rect 12344 -160 12664 160
rect 13356 -160 13676 160
rect 14368 -160 14688 160
rect 15380 -160 15700 160
rect 16392 -160 16712 160
rect -17004 -880 -16684 -560
rect -15992 -880 -15672 -560
rect -14980 -880 -14660 -560
rect -13968 -880 -13648 -560
rect -12956 -880 -12636 -560
rect -11944 -880 -11624 -560
rect -10932 -880 -10612 -560
rect -9920 -880 -9600 -560
rect -8908 -880 -8588 -560
rect -7896 -880 -7576 -560
rect -6884 -880 -6564 -560
rect -5872 -880 -5552 -560
rect -4860 -880 -4540 -560
rect -3848 -880 -3528 -560
rect -2836 -880 -2516 -560
rect -1824 -880 -1504 -560
rect -812 -880 -492 -560
rect 200 -880 520 -560
rect 1212 -880 1532 -560
rect 2224 -880 2544 -560
rect 3236 -880 3556 -560
rect 4248 -880 4568 -560
rect 5260 -880 5580 -560
rect 6272 -880 6592 -560
rect 7284 -880 7604 -560
rect 8296 -880 8616 -560
rect 9308 -880 9628 -560
rect 10320 -880 10640 -560
rect 11332 -880 11652 -560
rect 12344 -880 12664 -560
rect 13356 -880 13676 -560
rect 14368 -880 14688 -560
rect 15380 -880 15700 -560
rect 16392 -880 16712 -560
rect -17004 -1600 -16684 -1280
rect -15992 -1600 -15672 -1280
rect -14980 -1600 -14660 -1280
rect -13968 -1600 -13648 -1280
rect -12956 -1600 -12636 -1280
rect -11944 -1600 -11624 -1280
rect -10932 -1600 -10612 -1280
rect -9920 -1600 -9600 -1280
rect -8908 -1600 -8588 -1280
rect -7896 -1600 -7576 -1280
rect -6884 -1600 -6564 -1280
rect -5872 -1600 -5552 -1280
rect -4860 -1600 -4540 -1280
rect -3848 -1600 -3528 -1280
rect -2836 -1600 -2516 -1280
rect -1824 -1600 -1504 -1280
rect -812 -1600 -492 -1280
rect 200 -1600 520 -1280
rect 1212 -1600 1532 -1280
rect 2224 -1600 2544 -1280
rect 3236 -1600 3556 -1280
rect 4248 -1600 4568 -1280
rect 5260 -1600 5580 -1280
rect 6272 -1600 6592 -1280
rect 7284 -1600 7604 -1280
rect 8296 -1600 8616 -1280
rect 9308 -1600 9628 -1280
rect 10320 -1600 10640 -1280
rect 11332 -1600 11652 -1280
rect 12344 -1600 12664 -1280
rect 13356 -1600 13676 -1280
rect 14368 -1600 14688 -1280
rect 15380 -1600 15700 -1280
rect 16392 -1600 16712 -1280
rect -17004 -2320 -16684 -2000
rect -15992 -2320 -15672 -2000
rect -14980 -2320 -14660 -2000
rect -13968 -2320 -13648 -2000
rect -12956 -2320 -12636 -2000
rect -11944 -2320 -11624 -2000
rect -10932 -2320 -10612 -2000
rect -9920 -2320 -9600 -2000
rect -8908 -2320 -8588 -2000
rect -7896 -2320 -7576 -2000
rect -6884 -2320 -6564 -2000
rect -5872 -2320 -5552 -2000
rect -4860 -2320 -4540 -2000
rect -3848 -2320 -3528 -2000
rect -2836 -2320 -2516 -2000
rect -1824 -2320 -1504 -2000
rect -812 -2320 -492 -2000
rect 200 -2320 520 -2000
rect 1212 -2320 1532 -2000
rect 2224 -2320 2544 -2000
rect 3236 -2320 3556 -2000
rect 4248 -2320 4568 -2000
rect 5260 -2320 5580 -2000
rect 6272 -2320 6592 -2000
rect 7284 -2320 7604 -2000
rect 8296 -2320 8616 -2000
rect 9308 -2320 9628 -2000
rect 10320 -2320 10640 -2000
rect 11332 -2320 11652 -2000
rect 12344 -2320 12664 -2000
rect 13356 -2320 13676 -2000
rect 14368 -2320 14688 -2000
rect 15380 -2320 15700 -2000
rect 16392 -2320 16712 -2000
rect -17004 -3040 -16684 -2720
rect -15992 -3040 -15672 -2720
rect -14980 -3040 -14660 -2720
rect -13968 -3040 -13648 -2720
rect -12956 -3040 -12636 -2720
rect -11944 -3040 -11624 -2720
rect -10932 -3040 -10612 -2720
rect -9920 -3040 -9600 -2720
rect -8908 -3040 -8588 -2720
rect -7896 -3040 -7576 -2720
rect -6884 -3040 -6564 -2720
rect -5872 -3040 -5552 -2720
rect -4860 -3040 -4540 -2720
rect -3848 -3040 -3528 -2720
rect -2836 -3040 -2516 -2720
rect -1824 -3040 -1504 -2720
rect -812 -3040 -492 -2720
rect 200 -3040 520 -2720
rect 1212 -3040 1532 -2720
rect 2224 -3040 2544 -2720
rect 3236 -3040 3556 -2720
rect 4248 -3040 4568 -2720
rect 5260 -3040 5580 -2720
rect 6272 -3040 6592 -2720
rect 7284 -3040 7604 -2720
rect 8296 -3040 8616 -2720
rect 9308 -3040 9628 -2720
rect 10320 -3040 10640 -2720
rect 11332 -3040 11652 -2720
rect 12344 -3040 12664 -2720
rect 13356 -3040 13676 -2720
rect 14368 -3040 14688 -2720
rect 15380 -3040 15700 -2720
rect 16392 -3040 16712 -2720
rect -17004 -3760 -16684 -3440
rect -15992 -3760 -15672 -3440
rect -14980 -3760 -14660 -3440
rect -13968 -3760 -13648 -3440
rect -12956 -3760 -12636 -3440
rect -11944 -3760 -11624 -3440
rect -10932 -3760 -10612 -3440
rect -9920 -3760 -9600 -3440
rect -8908 -3760 -8588 -3440
rect -7896 -3760 -7576 -3440
rect -6884 -3760 -6564 -3440
rect -5872 -3760 -5552 -3440
rect -4860 -3760 -4540 -3440
rect -3848 -3760 -3528 -3440
rect -2836 -3760 -2516 -3440
rect -1824 -3760 -1504 -3440
rect -812 -3760 -492 -3440
rect 200 -3760 520 -3440
rect 1212 -3760 1532 -3440
rect 2224 -3760 2544 -3440
rect 3236 -3760 3556 -3440
rect 4248 -3760 4568 -3440
rect 5260 -3760 5580 -3440
rect 6272 -3760 6592 -3440
rect 7284 -3760 7604 -3440
rect 8296 -3760 8616 -3440
rect 9308 -3760 9628 -3440
rect 10320 -3760 10640 -3440
rect 11332 -3760 11652 -3440
rect 12344 -3760 12664 -3440
rect 13356 -3760 13676 -3440
rect 14368 -3760 14688 -3440
rect 15380 -3760 15700 -3440
rect 16392 -3760 16712 -3440
rect -17004 -4480 -16684 -4160
rect -15992 -4480 -15672 -4160
rect -14980 -4480 -14660 -4160
rect -13968 -4480 -13648 -4160
rect -12956 -4480 -12636 -4160
rect -11944 -4480 -11624 -4160
rect -10932 -4480 -10612 -4160
rect -9920 -4480 -9600 -4160
rect -8908 -4480 -8588 -4160
rect -7896 -4480 -7576 -4160
rect -6884 -4480 -6564 -4160
rect -5872 -4480 -5552 -4160
rect -4860 -4480 -4540 -4160
rect -3848 -4480 -3528 -4160
rect -2836 -4480 -2516 -4160
rect -1824 -4480 -1504 -4160
rect -812 -4480 -492 -4160
rect 200 -4480 520 -4160
rect 1212 -4480 1532 -4160
rect 2224 -4480 2544 -4160
rect 3236 -4480 3556 -4160
rect 4248 -4480 4568 -4160
rect 5260 -4480 5580 -4160
rect 6272 -4480 6592 -4160
rect 7284 -4480 7604 -4160
rect 8296 -4480 8616 -4160
rect 9308 -4480 9628 -4160
rect 10320 -4480 10640 -4160
rect 11332 -4480 11652 -4160
rect 12344 -4480 12664 -4160
rect 13356 -4480 13676 -4160
rect 14368 -4480 14688 -4160
rect 15380 -4480 15700 -4160
rect 16392 -4480 16712 -4160
rect -17004 -5200 -16684 -4880
rect -15992 -5200 -15672 -4880
rect -14980 -5200 -14660 -4880
rect -13968 -5200 -13648 -4880
rect -12956 -5200 -12636 -4880
rect -11944 -5200 -11624 -4880
rect -10932 -5200 -10612 -4880
rect -9920 -5200 -9600 -4880
rect -8908 -5200 -8588 -4880
rect -7896 -5200 -7576 -4880
rect -6884 -5200 -6564 -4880
rect -5872 -5200 -5552 -4880
rect -4860 -5200 -4540 -4880
rect -3848 -5200 -3528 -4880
rect -2836 -5200 -2516 -4880
rect -1824 -5200 -1504 -4880
rect -812 -5200 -492 -4880
rect 200 -5200 520 -4880
rect 1212 -5200 1532 -4880
rect 2224 -5200 2544 -4880
rect 3236 -5200 3556 -4880
rect 4248 -5200 4568 -4880
rect 5260 -5200 5580 -4880
rect 6272 -5200 6592 -4880
rect 7284 -5200 7604 -4880
rect 8296 -5200 8616 -4880
rect 9308 -5200 9628 -4880
rect 10320 -5200 10640 -4880
rect 11332 -5200 11652 -4880
rect 12344 -5200 12664 -4880
rect 13356 -5200 13676 -4880
rect 14368 -5200 14688 -4880
rect 15380 -5200 15700 -4880
rect 16392 -5200 16712 -4880
rect -17004 -5920 -16684 -5600
rect -15992 -5920 -15672 -5600
rect -14980 -5920 -14660 -5600
rect -13968 -5920 -13648 -5600
rect -12956 -5920 -12636 -5600
rect -11944 -5920 -11624 -5600
rect -10932 -5920 -10612 -5600
rect -9920 -5920 -9600 -5600
rect -8908 -5920 -8588 -5600
rect -7896 -5920 -7576 -5600
rect -6884 -5920 -6564 -5600
rect -5872 -5920 -5552 -5600
rect -4860 -5920 -4540 -5600
rect -3848 -5920 -3528 -5600
rect -2836 -5920 -2516 -5600
rect -1824 -5920 -1504 -5600
rect -812 -5920 -492 -5600
rect 200 -5920 520 -5600
rect 1212 -5920 1532 -5600
rect 2224 -5920 2544 -5600
rect 3236 -5920 3556 -5600
rect 4248 -5920 4568 -5600
rect 5260 -5920 5580 -5600
rect 6272 -5920 6592 -5600
rect 7284 -5920 7604 -5600
rect 8296 -5920 8616 -5600
rect 9308 -5920 9628 -5600
rect 10320 -5920 10640 -5600
rect 11332 -5920 11652 -5600
rect 12344 -5920 12664 -5600
rect 13356 -5920 13676 -5600
rect 14368 -5920 14688 -5600
rect 15380 -5920 15700 -5600
rect 16392 -5920 16712 -5600
rect -17004 -6640 -16684 -6320
rect -15992 -6640 -15672 -6320
rect -14980 -6640 -14660 -6320
rect -13968 -6640 -13648 -6320
rect -12956 -6640 -12636 -6320
rect -11944 -6640 -11624 -6320
rect -10932 -6640 -10612 -6320
rect -9920 -6640 -9600 -6320
rect -8908 -6640 -8588 -6320
rect -7896 -6640 -7576 -6320
rect -6884 -6640 -6564 -6320
rect -5872 -6640 -5552 -6320
rect -4860 -6640 -4540 -6320
rect -3848 -6640 -3528 -6320
rect -2836 -6640 -2516 -6320
rect -1824 -6640 -1504 -6320
rect -812 -6640 -492 -6320
rect 200 -6640 520 -6320
rect 1212 -6640 1532 -6320
rect 2224 -6640 2544 -6320
rect 3236 -6640 3556 -6320
rect 4248 -6640 4568 -6320
rect 5260 -6640 5580 -6320
rect 6272 -6640 6592 -6320
rect 7284 -6640 7604 -6320
rect 8296 -6640 8616 -6320
rect 9308 -6640 9628 -6320
rect 10320 -6640 10640 -6320
rect 11332 -6640 11652 -6320
rect 12344 -6640 12664 -6320
rect 13356 -6640 13676 -6320
rect 14368 -6640 14688 -6320
rect 15380 -6640 15700 -6320
rect 16392 -6640 16712 -6320
rect -17004 -7360 -16684 -7040
rect -15992 -7360 -15672 -7040
rect -14980 -7360 -14660 -7040
rect -13968 -7360 -13648 -7040
rect -12956 -7360 -12636 -7040
rect -11944 -7360 -11624 -7040
rect -10932 -7360 -10612 -7040
rect -9920 -7360 -9600 -7040
rect -8908 -7360 -8588 -7040
rect -7896 -7360 -7576 -7040
rect -6884 -7360 -6564 -7040
rect -5872 -7360 -5552 -7040
rect -4860 -7360 -4540 -7040
rect -3848 -7360 -3528 -7040
rect -2836 -7360 -2516 -7040
rect -1824 -7360 -1504 -7040
rect -812 -7360 -492 -7040
rect 200 -7360 520 -7040
rect 1212 -7360 1532 -7040
rect 2224 -7360 2544 -7040
rect 3236 -7360 3556 -7040
rect 4248 -7360 4568 -7040
rect 5260 -7360 5580 -7040
rect 6272 -7360 6592 -7040
rect 7284 -7360 7604 -7040
rect 8296 -7360 8616 -7040
rect 9308 -7360 9628 -7040
rect 10320 -7360 10640 -7040
rect 11332 -7360 11652 -7040
rect 12344 -7360 12664 -7040
rect 13356 -7360 13676 -7040
rect 14368 -7360 14688 -7040
rect 15380 -7360 15700 -7040
rect 16392 -7360 16712 -7040
rect -17004 -8080 -16684 -7760
rect -15992 -8080 -15672 -7760
rect -14980 -8080 -14660 -7760
rect -13968 -8080 -13648 -7760
rect -12956 -8080 -12636 -7760
rect -11944 -8080 -11624 -7760
rect -10932 -8080 -10612 -7760
rect -9920 -8080 -9600 -7760
rect -8908 -8080 -8588 -7760
rect -7896 -8080 -7576 -7760
rect -6884 -8080 -6564 -7760
rect -5872 -8080 -5552 -7760
rect -4860 -8080 -4540 -7760
rect -3848 -8080 -3528 -7760
rect -2836 -8080 -2516 -7760
rect -1824 -8080 -1504 -7760
rect -812 -8080 -492 -7760
rect 200 -8080 520 -7760
rect 1212 -8080 1532 -7760
rect 2224 -8080 2544 -7760
rect 3236 -8080 3556 -7760
rect 4248 -8080 4568 -7760
rect 5260 -8080 5580 -7760
rect 6272 -8080 6592 -7760
rect 7284 -8080 7604 -7760
rect 8296 -8080 8616 -7760
rect 9308 -8080 9628 -7760
rect 10320 -8080 10640 -7760
rect 11332 -8080 11652 -7760
rect 12344 -8080 12664 -7760
rect 13356 -8080 13676 -7760
rect 14368 -8080 14688 -7760
rect 15380 -8080 15700 -7760
rect 16392 -8080 16712 -7760
rect -17004 -8800 -16684 -8480
rect -15992 -8800 -15672 -8480
rect -14980 -8800 -14660 -8480
rect -13968 -8800 -13648 -8480
rect -12956 -8800 -12636 -8480
rect -11944 -8800 -11624 -8480
rect -10932 -8800 -10612 -8480
rect -9920 -8800 -9600 -8480
rect -8908 -8800 -8588 -8480
rect -7896 -8800 -7576 -8480
rect -6884 -8800 -6564 -8480
rect -5872 -8800 -5552 -8480
rect -4860 -8800 -4540 -8480
rect -3848 -8800 -3528 -8480
rect -2836 -8800 -2516 -8480
rect -1824 -8800 -1504 -8480
rect -812 -8800 -492 -8480
rect 200 -8800 520 -8480
rect 1212 -8800 1532 -8480
rect 2224 -8800 2544 -8480
rect 3236 -8800 3556 -8480
rect 4248 -8800 4568 -8480
rect 5260 -8800 5580 -8480
rect 6272 -8800 6592 -8480
rect 7284 -8800 7604 -8480
rect 8296 -8800 8616 -8480
rect 9308 -8800 9628 -8480
rect 10320 -8800 10640 -8480
rect 11332 -8800 11652 -8480
rect 12344 -8800 12664 -8480
rect 13356 -8800 13676 -8480
rect 14368 -8800 14688 -8480
rect 15380 -8800 15700 -8480
rect 16392 -8800 16712 -8480
rect -17004 -9520 -16684 -9200
rect -15992 -9520 -15672 -9200
rect -14980 -9520 -14660 -9200
rect -13968 -9520 -13648 -9200
rect -12956 -9520 -12636 -9200
rect -11944 -9520 -11624 -9200
rect -10932 -9520 -10612 -9200
rect -9920 -9520 -9600 -9200
rect -8908 -9520 -8588 -9200
rect -7896 -9520 -7576 -9200
rect -6884 -9520 -6564 -9200
rect -5872 -9520 -5552 -9200
rect -4860 -9520 -4540 -9200
rect -3848 -9520 -3528 -9200
rect -2836 -9520 -2516 -9200
rect -1824 -9520 -1504 -9200
rect -812 -9520 -492 -9200
rect 200 -9520 520 -9200
rect 1212 -9520 1532 -9200
rect 2224 -9520 2544 -9200
rect 3236 -9520 3556 -9200
rect 4248 -9520 4568 -9200
rect 5260 -9520 5580 -9200
rect 6272 -9520 6592 -9200
rect 7284 -9520 7604 -9200
rect 8296 -9520 8616 -9200
rect 9308 -9520 9628 -9200
rect 10320 -9520 10640 -9200
rect 11332 -9520 11652 -9200
rect 12344 -9520 12664 -9200
rect 13356 -9520 13676 -9200
rect 14368 -9520 14688 -9200
rect 15380 -9520 15700 -9200
rect 16392 -9520 16712 -9200
rect -17004 -10240 -16684 -9920
rect -15992 -10240 -15672 -9920
rect -14980 -10240 -14660 -9920
rect -13968 -10240 -13648 -9920
rect -12956 -10240 -12636 -9920
rect -11944 -10240 -11624 -9920
rect -10932 -10240 -10612 -9920
rect -9920 -10240 -9600 -9920
rect -8908 -10240 -8588 -9920
rect -7896 -10240 -7576 -9920
rect -6884 -10240 -6564 -9920
rect -5872 -10240 -5552 -9920
rect -4860 -10240 -4540 -9920
rect -3848 -10240 -3528 -9920
rect -2836 -10240 -2516 -9920
rect -1824 -10240 -1504 -9920
rect -812 -10240 -492 -9920
rect 200 -10240 520 -9920
rect 1212 -10240 1532 -9920
rect 2224 -10240 2544 -9920
rect 3236 -10240 3556 -9920
rect 4248 -10240 4568 -9920
rect 5260 -10240 5580 -9920
rect 6272 -10240 6592 -9920
rect 7284 -10240 7604 -9920
rect 8296 -10240 8616 -9920
rect 9308 -10240 9628 -9920
rect 10320 -10240 10640 -9920
rect 11332 -10240 11652 -9920
rect 12344 -10240 12664 -9920
rect 13356 -10240 13676 -9920
rect 14368 -10240 14688 -9920
rect 15380 -10240 15700 -9920
rect 16392 -10240 16712 -9920
rect -17004 -10960 -16684 -10640
rect -15992 -10960 -15672 -10640
rect -14980 -10960 -14660 -10640
rect -13968 -10960 -13648 -10640
rect -12956 -10960 -12636 -10640
rect -11944 -10960 -11624 -10640
rect -10932 -10960 -10612 -10640
rect -9920 -10960 -9600 -10640
rect -8908 -10960 -8588 -10640
rect -7896 -10960 -7576 -10640
rect -6884 -10960 -6564 -10640
rect -5872 -10960 -5552 -10640
rect -4860 -10960 -4540 -10640
rect -3848 -10960 -3528 -10640
rect -2836 -10960 -2516 -10640
rect -1824 -10960 -1504 -10640
rect -812 -10960 -492 -10640
rect 200 -10960 520 -10640
rect 1212 -10960 1532 -10640
rect 2224 -10960 2544 -10640
rect 3236 -10960 3556 -10640
rect 4248 -10960 4568 -10640
rect 5260 -10960 5580 -10640
rect 6272 -10960 6592 -10640
rect 7284 -10960 7604 -10640
rect 8296 -10960 8616 -10640
rect 9308 -10960 9628 -10640
rect 10320 -10960 10640 -10640
rect 11332 -10960 11652 -10640
rect 12344 -10960 12664 -10640
rect 13356 -10960 13676 -10640
rect 14368 -10960 14688 -10640
rect 15380 -10960 15700 -10640
rect 16392 -10960 16712 -10640
rect -17004 -11680 -16684 -11360
rect -15992 -11680 -15672 -11360
rect -14980 -11680 -14660 -11360
rect -13968 -11680 -13648 -11360
rect -12956 -11680 -12636 -11360
rect -11944 -11680 -11624 -11360
rect -10932 -11680 -10612 -11360
rect -9920 -11680 -9600 -11360
rect -8908 -11680 -8588 -11360
rect -7896 -11680 -7576 -11360
rect -6884 -11680 -6564 -11360
rect -5872 -11680 -5552 -11360
rect -4860 -11680 -4540 -11360
rect -3848 -11680 -3528 -11360
rect -2836 -11680 -2516 -11360
rect -1824 -11680 -1504 -11360
rect -812 -11680 -492 -11360
rect 200 -11680 520 -11360
rect 1212 -11680 1532 -11360
rect 2224 -11680 2544 -11360
rect 3236 -11680 3556 -11360
rect 4248 -11680 4568 -11360
rect 5260 -11680 5580 -11360
rect 6272 -11680 6592 -11360
rect 7284 -11680 7604 -11360
rect 8296 -11680 8616 -11360
rect 9308 -11680 9628 -11360
rect 10320 -11680 10640 -11360
rect 11332 -11680 11652 -11360
rect 12344 -11680 12664 -11360
rect 13356 -11680 13676 -11360
rect 14368 -11680 14688 -11360
rect 15380 -11680 15700 -11360
rect 16392 -11680 16712 -11360
<< metal4 >>
rect -16412 11732 -16316 11748
rect -17005 11680 -16683 11681
rect -17005 11360 -17004 11680
rect -16684 11360 -16683 11680
rect -17005 11359 -16683 11360
rect -16412 11308 -16396 11732
rect -16332 11308 -16316 11732
rect -15400 11732 -15304 11748
rect -15993 11680 -15671 11681
rect -15993 11360 -15992 11680
rect -15672 11360 -15671 11680
rect -15993 11359 -15671 11360
rect -16412 11292 -16316 11308
rect -15400 11308 -15384 11732
rect -15320 11308 -15304 11732
rect -14388 11732 -14292 11748
rect -14981 11680 -14659 11681
rect -14981 11360 -14980 11680
rect -14660 11360 -14659 11680
rect -14981 11359 -14659 11360
rect -15400 11292 -15304 11308
rect -14388 11308 -14372 11732
rect -14308 11308 -14292 11732
rect -13376 11732 -13280 11748
rect -13969 11680 -13647 11681
rect -13969 11360 -13968 11680
rect -13648 11360 -13647 11680
rect -13969 11359 -13647 11360
rect -14388 11292 -14292 11308
rect -13376 11308 -13360 11732
rect -13296 11308 -13280 11732
rect -12364 11732 -12268 11748
rect -12957 11680 -12635 11681
rect -12957 11360 -12956 11680
rect -12636 11360 -12635 11680
rect -12957 11359 -12635 11360
rect -13376 11292 -13280 11308
rect -12364 11308 -12348 11732
rect -12284 11308 -12268 11732
rect -11352 11732 -11256 11748
rect -11945 11680 -11623 11681
rect -11945 11360 -11944 11680
rect -11624 11360 -11623 11680
rect -11945 11359 -11623 11360
rect -12364 11292 -12268 11308
rect -11352 11308 -11336 11732
rect -11272 11308 -11256 11732
rect -10340 11732 -10244 11748
rect -10933 11680 -10611 11681
rect -10933 11360 -10932 11680
rect -10612 11360 -10611 11680
rect -10933 11359 -10611 11360
rect -11352 11292 -11256 11308
rect -10340 11308 -10324 11732
rect -10260 11308 -10244 11732
rect -9328 11732 -9232 11748
rect -9921 11680 -9599 11681
rect -9921 11360 -9920 11680
rect -9600 11360 -9599 11680
rect -9921 11359 -9599 11360
rect -10340 11292 -10244 11308
rect -9328 11308 -9312 11732
rect -9248 11308 -9232 11732
rect -8316 11732 -8220 11748
rect -8909 11680 -8587 11681
rect -8909 11360 -8908 11680
rect -8588 11360 -8587 11680
rect -8909 11359 -8587 11360
rect -9328 11292 -9232 11308
rect -8316 11308 -8300 11732
rect -8236 11308 -8220 11732
rect -7304 11732 -7208 11748
rect -7897 11680 -7575 11681
rect -7897 11360 -7896 11680
rect -7576 11360 -7575 11680
rect -7897 11359 -7575 11360
rect -8316 11292 -8220 11308
rect -7304 11308 -7288 11732
rect -7224 11308 -7208 11732
rect -6292 11732 -6196 11748
rect -6885 11680 -6563 11681
rect -6885 11360 -6884 11680
rect -6564 11360 -6563 11680
rect -6885 11359 -6563 11360
rect -7304 11292 -7208 11308
rect -6292 11308 -6276 11732
rect -6212 11308 -6196 11732
rect -5280 11732 -5184 11748
rect -5873 11680 -5551 11681
rect -5873 11360 -5872 11680
rect -5552 11360 -5551 11680
rect -5873 11359 -5551 11360
rect -6292 11292 -6196 11308
rect -5280 11308 -5264 11732
rect -5200 11308 -5184 11732
rect -4268 11732 -4172 11748
rect -4861 11680 -4539 11681
rect -4861 11360 -4860 11680
rect -4540 11360 -4539 11680
rect -4861 11359 -4539 11360
rect -5280 11292 -5184 11308
rect -4268 11308 -4252 11732
rect -4188 11308 -4172 11732
rect -3256 11732 -3160 11748
rect -3849 11680 -3527 11681
rect -3849 11360 -3848 11680
rect -3528 11360 -3527 11680
rect -3849 11359 -3527 11360
rect -4268 11292 -4172 11308
rect -3256 11308 -3240 11732
rect -3176 11308 -3160 11732
rect -2244 11732 -2148 11748
rect -2837 11680 -2515 11681
rect -2837 11360 -2836 11680
rect -2516 11360 -2515 11680
rect -2837 11359 -2515 11360
rect -3256 11292 -3160 11308
rect -2244 11308 -2228 11732
rect -2164 11308 -2148 11732
rect -1232 11732 -1136 11748
rect -1825 11680 -1503 11681
rect -1825 11360 -1824 11680
rect -1504 11360 -1503 11680
rect -1825 11359 -1503 11360
rect -2244 11292 -2148 11308
rect -1232 11308 -1216 11732
rect -1152 11308 -1136 11732
rect -220 11732 -124 11748
rect -813 11680 -491 11681
rect -813 11360 -812 11680
rect -492 11360 -491 11680
rect -813 11359 -491 11360
rect -1232 11292 -1136 11308
rect -220 11308 -204 11732
rect -140 11308 -124 11732
rect 792 11732 888 11748
rect 199 11680 521 11681
rect 199 11360 200 11680
rect 520 11360 521 11680
rect 199 11359 521 11360
rect -220 11292 -124 11308
rect 792 11308 808 11732
rect 872 11308 888 11732
rect 1804 11732 1900 11748
rect 1211 11680 1533 11681
rect 1211 11360 1212 11680
rect 1532 11360 1533 11680
rect 1211 11359 1533 11360
rect 792 11292 888 11308
rect 1804 11308 1820 11732
rect 1884 11308 1900 11732
rect 2816 11732 2912 11748
rect 2223 11680 2545 11681
rect 2223 11360 2224 11680
rect 2544 11360 2545 11680
rect 2223 11359 2545 11360
rect 1804 11292 1900 11308
rect 2816 11308 2832 11732
rect 2896 11308 2912 11732
rect 3828 11732 3924 11748
rect 3235 11680 3557 11681
rect 3235 11360 3236 11680
rect 3556 11360 3557 11680
rect 3235 11359 3557 11360
rect 2816 11292 2912 11308
rect 3828 11308 3844 11732
rect 3908 11308 3924 11732
rect 4840 11732 4936 11748
rect 4247 11680 4569 11681
rect 4247 11360 4248 11680
rect 4568 11360 4569 11680
rect 4247 11359 4569 11360
rect 3828 11292 3924 11308
rect 4840 11308 4856 11732
rect 4920 11308 4936 11732
rect 5852 11732 5948 11748
rect 5259 11680 5581 11681
rect 5259 11360 5260 11680
rect 5580 11360 5581 11680
rect 5259 11359 5581 11360
rect 4840 11292 4936 11308
rect 5852 11308 5868 11732
rect 5932 11308 5948 11732
rect 6864 11732 6960 11748
rect 6271 11680 6593 11681
rect 6271 11360 6272 11680
rect 6592 11360 6593 11680
rect 6271 11359 6593 11360
rect 5852 11292 5948 11308
rect 6864 11308 6880 11732
rect 6944 11308 6960 11732
rect 7876 11732 7972 11748
rect 7283 11680 7605 11681
rect 7283 11360 7284 11680
rect 7604 11360 7605 11680
rect 7283 11359 7605 11360
rect 6864 11292 6960 11308
rect 7876 11308 7892 11732
rect 7956 11308 7972 11732
rect 8888 11732 8984 11748
rect 8295 11680 8617 11681
rect 8295 11360 8296 11680
rect 8616 11360 8617 11680
rect 8295 11359 8617 11360
rect 7876 11292 7972 11308
rect 8888 11308 8904 11732
rect 8968 11308 8984 11732
rect 9900 11732 9996 11748
rect 9307 11680 9629 11681
rect 9307 11360 9308 11680
rect 9628 11360 9629 11680
rect 9307 11359 9629 11360
rect 8888 11292 8984 11308
rect 9900 11308 9916 11732
rect 9980 11308 9996 11732
rect 10912 11732 11008 11748
rect 10319 11680 10641 11681
rect 10319 11360 10320 11680
rect 10640 11360 10641 11680
rect 10319 11359 10641 11360
rect 9900 11292 9996 11308
rect 10912 11308 10928 11732
rect 10992 11308 11008 11732
rect 11924 11732 12020 11748
rect 11331 11680 11653 11681
rect 11331 11360 11332 11680
rect 11652 11360 11653 11680
rect 11331 11359 11653 11360
rect 10912 11292 11008 11308
rect 11924 11308 11940 11732
rect 12004 11308 12020 11732
rect 12936 11732 13032 11748
rect 12343 11680 12665 11681
rect 12343 11360 12344 11680
rect 12664 11360 12665 11680
rect 12343 11359 12665 11360
rect 11924 11292 12020 11308
rect 12936 11308 12952 11732
rect 13016 11308 13032 11732
rect 13948 11732 14044 11748
rect 13355 11680 13677 11681
rect 13355 11360 13356 11680
rect 13676 11360 13677 11680
rect 13355 11359 13677 11360
rect 12936 11292 13032 11308
rect 13948 11308 13964 11732
rect 14028 11308 14044 11732
rect 14960 11732 15056 11748
rect 14367 11680 14689 11681
rect 14367 11360 14368 11680
rect 14688 11360 14689 11680
rect 14367 11359 14689 11360
rect 13948 11292 14044 11308
rect 14960 11308 14976 11732
rect 15040 11308 15056 11732
rect 15972 11732 16068 11748
rect 15379 11680 15701 11681
rect 15379 11360 15380 11680
rect 15700 11360 15701 11680
rect 15379 11359 15701 11360
rect 14960 11292 15056 11308
rect 15972 11308 15988 11732
rect 16052 11308 16068 11732
rect 16984 11732 17080 11748
rect 16391 11680 16713 11681
rect 16391 11360 16392 11680
rect 16712 11360 16713 11680
rect 16391 11359 16713 11360
rect 15972 11292 16068 11308
rect 16984 11308 17000 11732
rect 17064 11308 17080 11732
rect 16984 11292 17080 11308
rect -16412 11012 -16316 11028
rect -17005 10960 -16683 10961
rect -17005 10640 -17004 10960
rect -16684 10640 -16683 10960
rect -17005 10639 -16683 10640
rect -16412 10588 -16396 11012
rect -16332 10588 -16316 11012
rect -15400 11012 -15304 11028
rect -15993 10960 -15671 10961
rect -15993 10640 -15992 10960
rect -15672 10640 -15671 10960
rect -15993 10639 -15671 10640
rect -16412 10572 -16316 10588
rect -15400 10588 -15384 11012
rect -15320 10588 -15304 11012
rect -14388 11012 -14292 11028
rect -14981 10960 -14659 10961
rect -14981 10640 -14980 10960
rect -14660 10640 -14659 10960
rect -14981 10639 -14659 10640
rect -15400 10572 -15304 10588
rect -14388 10588 -14372 11012
rect -14308 10588 -14292 11012
rect -13376 11012 -13280 11028
rect -13969 10960 -13647 10961
rect -13969 10640 -13968 10960
rect -13648 10640 -13647 10960
rect -13969 10639 -13647 10640
rect -14388 10572 -14292 10588
rect -13376 10588 -13360 11012
rect -13296 10588 -13280 11012
rect -12364 11012 -12268 11028
rect -12957 10960 -12635 10961
rect -12957 10640 -12956 10960
rect -12636 10640 -12635 10960
rect -12957 10639 -12635 10640
rect -13376 10572 -13280 10588
rect -12364 10588 -12348 11012
rect -12284 10588 -12268 11012
rect -11352 11012 -11256 11028
rect -11945 10960 -11623 10961
rect -11945 10640 -11944 10960
rect -11624 10640 -11623 10960
rect -11945 10639 -11623 10640
rect -12364 10572 -12268 10588
rect -11352 10588 -11336 11012
rect -11272 10588 -11256 11012
rect -10340 11012 -10244 11028
rect -10933 10960 -10611 10961
rect -10933 10640 -10932 10960
rect -10612 10640 -10611 10960
rect -10933 10639 -10611 10640
rect -11352 10572 -11256 10588
rect -10340 10588 -10324 11012
rect -10260 10588 -10244 11012
rect -9328 11012 -9232 11028
rect -9921 10960 -9599 10961
rect -9921 10640 -9920 10960
rect -9600 10640 -9599 10960
rect -9921 10639 -9599 10640
rect -10340 10572 -10244 10588
rect -9328 10588 -9312 11012
rect -9248 10588 -9232 11012
rect -8316 11012 -8220 11028
rect -8909 10960 -8587 10961
rect -8909 10640 -8908 10960
rect -8588 10640 -8587 10960
rect -8909 10639 -8587 10640
rect -9328 10572 -9232 10588
rect -8316 10588 -8300 11012
rect -8236 10588 -8220 11012
rect -7304 11012 -7208 11028
rect -7897 10960 -7575 10961
rect -7897 10640 -7896 10960
rect -7576 10640 -7575 10960
rect -7897 10639 -7575 10640
rect -8316 10572 -8220 10588
rect -7304 10588 -7288 11012
rect -7224 10588 -7208 11012
rect -6292 11012 -6196 11028
rect -6885 10960 -6563 10961
rect -6885 10640 -6884 10960
rect -6564 10640 -6563 10960
rect -6885 10639 -6563 10640
rect -7304 10572 -7208 10588
rect -6292 10588 -6276 11012
rect -6212 10588 -6196 11012
rect -5280 11012 -5184 11028
rect -5873 10960 -5551 10961
rect -5873 10640 -5872 10960
rect -5552 10640 -5551 10960
rect -5873 10639 -5551 10640
rect -6292 10572 -6196 10588
rect -5280 10588 -5264 11012
rect -5200 10588 -5184 11012
rect -4268 11012 -4172 11028
rect -4861 10960 -4539 10961
rect -4861 10640 -4860 10960
rect -4540 10640 -4539 10960
rect -4861 10639 -4539 10640
rect -5280 10572 -5184 10588
rect -4268 10588 -4252 11012
rect -4188 10588 -4172 11012
rect -3256 11012 -3160 11028
rect -3849 10960 -3527 10961
rect -3849 10640 -3848 10960
rect -3528 10640 -3527 10960
rect -3849 10639 -3527 10640
rect -4268 10572 -4172 10588
rect -3256 10588 -3240 11012
rect -3176 10588 -3160 11012
rect -2244 11012 -2148 11028
rect -2837 10960 -2515 10961
rect -2837 10640 -2836 10960
rect -2516 10640 -2515 10960
rect -2837 10639 -2515 10640
rect -3256 10572 -3160 10588
rect -2244 10588 -2228 11012
rect -2164 10588 -2148 11012
rect -1232 11012 -1136 11028
rect -1825 10960 -1503 10961
rect -1825 10640 -1824 10960
rect -1504 10640 -1503 10960
rect -1825 10639 -1503 10640
rect -2244 10572 -2148 10588
rect -1232 10588 -1216 11012
rect -1152 10588 -1136 11012
rect -220 11012 -124 11028
rect -813 10960 -491 10961
rect -813 10640 -812 10960
rect -492 10640 -491 10960
rect -813 10639 -491 10640
rect -1232 10572 -1136 10588
rect -220 10588 -204 11012
rect -140 10588 -124 11012
rect 792 11012 888 11028
rect 199 10960 521 10961
rect 199 10640 200 10960
rect 520 10640 521 10960
rect 199 10639 521 10640
rect -220 10572 -124 10588
rect 792 10588 808 11012
rect 872 10588 888 11012
rect 1804 11012 1900 11028
rect 1211 10960 1533 10961
rect 1211 10640 1212 10960
rect 1532 10640 1533 10960
rect 1211 10639 1533 10640
rect 792 10572 888 10588
rect 1804 10588 1820 11012
rect 1884 10588 1900 11012
rect 2816 11012 2912 11028
rect 2223 10960 2545 10961
rect 2223 10640 2224 10960
rect 2544 10640 2545 10960
rect 2223 10639 2545 10640
rect 1804 10572 1900 10588
rect 2816 10588 2832 11012
rect 2896 10588 2912 11012
rect 3828 11012 3924 11028
rect 3235 10960 3557 10961
rect 3235 10640 3236 10960
rect 3556 10640 3557 10960
rect 3235 10639 3557 10640
rect 2816 10572 2912 10588
rect 3828 10588 3844 11012
rect 3908 10588 3924 11012
rect 4840 11012 4936 11028
rect 4247 10960 4569 10961
rect 4247 10640 4248 10960
rect 4568 10640 4569 10960
rect 4247 10639 4569 10640
rect 3828 10572 3924 10588
rect 4840 10588 4856 11012
rect 4920 10588 4936 11012
rect 5852 11012 5948 11028
rect 5259 10960 5581 10961
rect 5259 10640 5260 10960
rect 5580 10640 5581 10960
rect 5259 10639 5581 10640
rect 4840 10572 4936 10588
rect 5852 10588 5868 11012
rect 5932 10588 5948 11012
rect 6864 11012 6960 11028
rect 6271 10960 6593 10961
rect 6271 10640 6272 10960
rect 6592 10640 6593 10960
rect 6271 10639 6593 10640
rect 5852 10572 5948 10588
rect 6864 10588 6880 11012
rect 6944 10588 6960 11012
rect 7876 11012 7972 11028
rect 7283 10960 7605 10961
rect 7283 10640 7284 10960
rect 7604 10640 7605 10960
rect 7283 10639 7605 10640
rect 6864 10572 6960 10588
rect 7876 10588 7892 11012
rect 7956 10588 7972 11012
rect 8888 11012 8984 11028
rect 8295 10960 8617 10961
rect 8295 10640 8296 10960
rect 8616 10640 8617 10960
rect 8295 10639 8617 10640
rect 7876 10572 7972 10588
rect 8888 10588 8904 11012
rect 8968 10588 8984 11012
rect 9900 11012 9996 11028
rect 9307 10960 9629 10961
rect 9307 10640 9308 10960
rect 9628 10640 9629 10960
rect 9307 10639 9629 10640
rect 8888 10572 8984 10588
rect 9900 10588 9916 11012
rect 9980 10588 9996 11012
rect 10912 11012 11008 11028
rect 10319 10960 10641 10961
rect 10319 10640 10320 10960
rect 10640 10640 10641 10960
rect 10319 10639 10641 10640
rect 9900 10572 9996 10588
rect 10912 10588 10928 11012
rect 10992 10588 11008 11012
rect 11924 11012 12020 11028
rect 11331 10960 11653 10961
rect 11331 10640 11332 10960
rect 11652 10640 11653 10960
rect 11331 10639 11653 10640
rect 10912 10572 11008 10588
rect 11924 10588 11940 11012
rect 12004 10588 12020 11012
rect 12936 11012 13032 11028
rect 12343 10960 12665 10961
rect 12343 10640 12344 10960
rect 12664 10640 12665 10960
rect 12343 10639 12665 10640
rect 11924 10572 12020 10588
rect 12936 10588 12952 11012
rect 13016 10588 13032 11012
rect 13948 11012 14044 11028
rect 13355 10960 13677 10961
rect 13355 10640 13356 10960
rect 13676 10640 13677 10960
rect 13355 10639 13677 10640
rect 12936 10572 13032 10588
rect 13948 10588 13964 11012
rect 14028 10588 14044 11012
rect 14960 11012 15056 11028
rect 14367 10960 14689 10961
rect 14367 10640 14368 10960
rect 14688 10640 14689 10960
rect 14367 10639 14689 10640
rect 13948 10572 14044 10588
rect 14960 10588 14976 11012
rect 15040 10588 15056 11012
rect 15972 11012 16068 11028
rect 15379 10960 15701 10961
rect 15379 10640 15380 10960
rect 15700 10640 15701 10960
rect 15379 10639 15701 10640
rect 14960 10572 15056 10588
rect 15972 10588 15988 11012
rect 16052 10588 16068 11012
rect 16984 11012 17080 11028
rect 16391 10960 16713 10961
rect 16391 10640 16392 10960
rect 16712 10640 16713 10960
rect 16391 10639 16713 10640
rect 15972 10572 16068 10588
rect 16984 10588 17000 11012
rect 17064 10588 17080 11012
rect 16984 10572 17080 10588
rect -16412 10292 -16316 10308
rect -17005 10240 -16683 10241
rect -17005 9920 -17004 10240
rect -16684 9920 -16683 10240
rect -17005 9919 -16683 9920
rect -16412 9868 -16396 10292
rect -16332 9868 -16316 10292
rect -15400 10292 -15304 10308
rect -15993 10240 -15671 10241
rect -15993 9920 -15992 10240
rect -15672 9920 -15671 10240
rect -15993 9919 -15671 9920
rect -16412 9852 -16316 9868
rect -15400 9868 -15384 10292
rect -15320 9868 -15304 10292
rect -14388 10292 -14292 10308
rect -14981 10240 -14659 10241
rect -14981 9920 -14980 10240
rect -14660 9920 -14659 10240
rect -14981 9919 -14659 9920
rect -15400 9852 -15304 9868
rect -14388 9868 -14372 10292
rect -14308 9868 -14292 10292
rect -13376 10292 -13280 10308
rect -13969 10240 -13647 10241
rect -13969 9920 -13968 10240
rect -13648 9920 -13647 10240
rect -13969 9919 -13647 9920
rect -14388 9852 -14292 9868
rect -13376 9868 -13360 10292
rect -13296 9868 -13280 10292
rect -12364 10292 -12268 10308
rect -12957 10240 -12635 10241
rect -12957 9920 -12956 10240
rect -12636 9920 -12635 10240
rect -12957 9919 -12635 9920
rect -13376 9852 -13280 9868
rect -12364 9868 -12348 10292
rect -12284 9868 -12268 10292
rect -11352 10292 -11256 10308
rect -11945 10240 -11623 10241
rect -11945 9920 -11944 10240
rect -11624 9920 -11623 10240
rect -11945 9919 -11623 9920
rect -12364 9852 -12268 9868
rect -11352 9868 -11336 10292
rect -11272 9868 -11256 10292
rect -10340 10292 -10244 10308
rect -10933 10240 -10611 10241
rect -10933 9920 -10932 10240
rect -10612 9920 -10611 10240
rect -10933 9919 -10611 9920
rect -11352 9852 -11256 9868
rect -10340 9868 -10324 10292
rect -10260 9868 -10244 10292
rect -9328 10292 -9232 10308
rect -9921 10240 -9599 10241
rect -9921 9920 -9920 10240
rect -9600 9920 -9599 10240
rect -9921 9919 -9599 9920
rect -10340 9852 -10244 9868
rect -9328 9868 -9312 10292
rect -9248 9868 -9232 10292
rect -8316 10292 -8220 10308
rect -8909 10240 -8587 10241
rect -8909 9920 -8908 10240
rect -8588 9920 -8587 10240
rect -8909 9919 -8587 9920
rect -9328 9852 -9232 9868
rect -8316 9868 -8300 10292
rect -8236 9868 -8220 10292
rect -7304 10292 -7208 10308
rect -7897 10240 -7575 10241
rect -7897 9920 -7896 10240
rect -7576 9920 -7575 10240
rect -7897 9919 -7575 9920
rect -8316 9852 -8220 9868
rect -7304 9868 -7288 10292
rect -7224 9868 -7208 10292
rect -6292 10292 -6196 10308
rect -6885 10240 -6563 10241
rect -6885 9920 -6884 10240
rect -6564 9920 -6563 10240
rect -6885 9919 -6563 9920
rect -7304 9852 -7208 9868
rect -6292 9868 -6276 10292
rect -6212 9868 -6196 10292
rect -5280 10292 -5184 10308
rect -5873 10240 -5551 10241
rect -5873 9920 -5872 10240
rect -5552 9920 -5551 10240
rect -5873 9919 -5551 9920
rect -6292 9852 -6196 9868
rect -5280 9868 -5264 10292
rect -5200 9868 -5184 10292
rect -4268 10292 -4172 10308
rect -4861 10240 -4539 10241
rect -4861 9920 -4860 10240
rect -4540 9920 -4539 10240
rect -4861 9919 -4539 9920
rect -5280 9852 -5184 9868
rect -4268 9868 -4252 10292
rect -4188 9868 -4172 10292
rect -3256 10292 -3160 10308
rect -3849 10240 -3527 10241
rect -3849 9920 -3848 10240
rect -3528 9920 -3527 10240
rect -3849 9919 -3527 9920
rect -4268 9852 -4172 9868
rect -3256 9868 -3240 10292
rect -3176 9868 -3160 10292
rect -2244 10292 -2148 10308
rect -2837 10240 -2515 10241
rect -2837 9920 -2836 10240
rect -2516 9920 -2515 10240
rect -2837 9919 -2515 9920
rect -3256 9852 -3160 9868
rect -2244 9868 -2228 10292
rect -2164 9868 -2148 10292
rect -1232 10292 -1136 10308
rect -1825 10240 -1503 10241
rect -1825 9920 -1824 10240
rect -1504 9920 -1503 10240
rect -1825 9919 -1503 9920
rect -2244 9852 -2148 9868
rect -1232 9868 -1216 10292
rect -1152 9868 -1136 10292
rect -220 10292 -124 10308
rect -813 10240 -491 10241
rect -813 9920 -812 10240
rect -492 9920 -491 10240
rect -813 9919 -491 9920
rect -1232 9852 -1136 9868
rect -220 9868 -204 10292
rect -140 9868 -124 10292
rect 792 10292 888 10308
rect 199 10240 521 10241
rect 199 9920 200 10240
rect 520 9920 521 10240
rect 199 9919 521 9920
rect -220 9852 -124 9868
rect 792 9868 808 10292
rect 872 9868 888 10292
rect 1804 10292 1900 10308
rect 1211 10240 1533 10241
rect 1211 9920 1212 10240
rect 1532 9920 1533 10240
rect 1211 9919 1533 9920
rect 792 9852 888 9868
rect 1804 9868 1820 10292
rect 1884 9868 1900 10292
rect 2816 10292 2912 10308
rect 2223 10240 2545 10241
rect 2223 9920 2224 10240
rect 2544 9920 2545 10240
rect 2223 9919 2545 9920
rect 1804 9852 1900 9868
rect 2816 9868 2832 10292
rect 2896 9868 2912 10292
rect 3828 10292 3924 10308
rect 3235 10240 3557 10241
rect 3235 9920 3236 10240
rect 3556 9920 3557 10240
rect 3235 9919 3557 9920
rect 2816 9852 2912 9868
rect 3828 9868 3844 10292
rect 3908 9868 3924 10292
rect 4840 10292 4936 10308
rect 4247 10240 4569 10241
rect 4247 9920 4248 10240
rect 4568 9920 4569 10240
rect 4247 9919 4569 9920
rect 3828 9852 3924 9868
rect 4840 9868 4856 10292
rect 4920 9868 4936 10292
rect 5852 10292 5948 10308
rect 5259 10240 5581 10241
rect 5259 9920 5260 10240
rect 5580 9920 5581 10240
rect 5259 9919 5581 9920
rect 4840 9852 4936 9868
rect 5852 9868 5868 10292
rect 5932 9868 5948 10292
rect 6864 10292 6960 10308
rect 6271 10240 6593 10241
rect 6271 9920 6272 10240
rect 6592 9920 6593 10240
rect 6271 9919 6593 9920
rect 5852 9852 5948 9868
rect 6864 9868 6880 10292
rect 6944 9868 6960 10292
rect 7876 10292 7972 10308
rect 7283 10240 7605 10241
rect 7283 9920 7284 10240
rect 7604 9920 7605 10240
rect 7283 9919 7605 9920
rect 6864 9852 6960 9868
rect 7876 9868 7892 10292
rect 7956 9868 7972 10292
rect 8888 10292 8984 10308
rect 8295 10240 8617 10241
rect 8295 9920 8296 10240
rect 8616 9920 8617 10240
rect 8295 9919 8617 9920
rect 7876 9852 7972 9868
rect 8888 9868 8904 10292
rect 8968 9868 8984 10292
rect 9900 10292 9996 10308
rect 9307 10240 9629 10241
rect 9307 9920 9308 10240
rect 9628 9920 9629 10240
rect 9307 9919 9629 9920
rect 8888 9852 8984 9868
rect 9900 9868 9916 10292
rect 9980 9868 9996 10292
rect 10912 10292 11008 10308
rect 10319 10240 10641 10241
rect 10319 9920 10320 10240
rect 10640 9920 10641 10240
rect 10319 9919 10641 9920
rect 9900 9852 9996 9868
rect 10912 9868 10928 10292
rect 10992 9868 11008 10292
rect 11924 10292 12020 10308
rect 11331 10240 11653 10241
rect 11331 9920 11332 10240
rect 11652 9920 11653 10240
rect 11331 9919 11653 9920
rect 10912 9852 11008 9868
rect 11924 9868 11940 10292
rect 12004 9868 12020 10292
rect 12936 10292 13032 10308
rect 12343 10240 12665 10241
rect 12343 9920 12344 10240
rect 12664 9920 12665 10240
rect 12343 9919 12665 9920
rect 11924 9852 12020 9868
rect 12936 9868 12952 10292
rect 13016 9868 13032 10292
rect 13948 10292 14044 10308
rect 13355 10240 13677 10241
rect 13355 9920 13356 10240
rect 13676 9920 13677 10240
rect 13355 9919 13677 9920
rect 12936 9852 13032 9868
rect 13948 9868 13964 10292
rect 14028 9868 14044 10292
rect 14960 10292 15056 10308
rect 14367 10240 14689 10241
rect 14367 9920 14368 10240
rect 14688 9920 14689 10240
rect 14367 9919 14689 9920
rect 13948 9852 14044 9868
rect 14960 9868 14976 10292
rect 15040 9868 15056 10292
rect 15972 10292 16068 10308
rect 15379 10240 15701 10241
rect 15379 9920 15380 10240
rect 15700 9920 15701 10240
rect 15379 9919 15701 9920
rect 14960 9852 15056 9868
rect 15972 9868 15988 10292
rect 16052 9868 16068 10292
rect 16984 10292 17080 10308
rect 16391 10240 16713 10241
rect 16391 9920 16392 10240
rect 16712 9920 16713 10240
rect 16391 9919 16713 9920
rect 15972 9852 16068 9868
rect 16984 9868 17000 10292
rect 17064 9868 17080 10292
rect 16984 9852 17080 9868
rect -16412 9572 -16316 9588
rect -17005 9520 -16683 9521
rect -17005 9200 -17004 9520
rect -16684 9200 -16683 9520
rect -17005 9199 -16683 9200
rect -16412 9148 -16396 9572
rect -16332 9148 -16316 9572
rect -15400 9572 -15304 9588
rect -15993 9520 -15671 9521
rect -15993 9200 -15992 9520
rect -15672 9200 -15671 9520
rect -15993 9199 -15671 9200
rect -16412 9132 -16316 9148
rect -15400 9148 -15384 9572
rect -15320 9148 -15304 9572
rect -14388 9572 -14292 9588
rect -14981 9520 -14659 9521
rect -14981 9200 -14980 9520
rect -14660 9200 -14659 9520
rect -14981 9199 -14659 9200
rect -15400 9132 -15304 9148
rect -14388 9148 -14372 9572
rect -14308 9148 -14292 9572
rect -13376 9572 -13280 9588
rect -13969 9520 -13647 9521
rect -13969 9200 -13968 9520
rect -13648 9200 -13647 9520
rect -13969 9199 -13647 9200
rect -14388 9132 -14292 9148
rect -13376 9148 -13360 9572
rect -13296 9148 -13280 9572
rect -12364 9572 -12268 9588
rect -12957 9520 -12635 9521
rect -12957 9200 -12956 9520
rect -12636 9200 -12635 9520
rect -12957 9199 -12635 9200
rect -13376 9132 -13280 9148
rect -12364 9148 -12348 9572
rect -12284 9148 -12268 9572
rect -11352 9572 -11256 9588
rect -11945 9520 -11623 9521
rect -11945 9200 -11944 9520
rect -11624 9200 -11623 9520
rect -11945 9199 -11623 9200
rect -12364 9132 -12268 9148
rect -11352 9148 -11336 9572
rect -11272 9148 -11256 9572
rect -10340 9572 -10244 9588
rect -10933 9520 -10611 9521
rect -10933 9200 -10932 9520
rect -10612 9200 -10611 9520
rect -10933 9199 -10611 9200
rect -11352 9132 -11256 9148
rect -10340 9148 -10324 9572
rect -10260 9148 -10244 9572
rect -9328 9572 -9232 9588
rect -9921 9520 -9599 9521
rect -9921 9200 -9920 9520
rect -9600 9200 -9599 9520
rect -9921 9199 -9599 9200
rect -10340 9132 -10244 9148
rect -9328 9148 -9312 9572
rect -9248 9148 -9232 9572
rect -8316 9572 -8220 9588
rect -8909 9520 -8587 9521
rect -8909 9200 -8908 9520
rect -8588 9200 -8587 9520
rect -8909 9199 -8587 9200
rect -9328 9132 -9232 9148
rect -8316 9148 -8300 9572
rect -8236 9148 -8220 9572
rect -7304 9572 -7208 9588
rect -7897 9520 -7575 9521
rect -7897 9200 -7896 9520
rect -7576 9200 -7575 9520
rect -7897 9199 -7575 9200
rect -8316 9132 -8220 9148
rect -7304 9148 -7288 9572
rect -7224 9148 -7208 9572
rect -6292 9572 -6196 9588
rect -6885 9520 -6563 9521
rect -6885 9200 -6884 9520
rect -6564 9200 -6563 9520
rect -6885 9199 -6563 9200
rect -7304 9132 -7208 9148
rect -6292 9148 -6276 9572
rect -6212 9148 -6196 9572
rect -5280 9572 -5184 9588
rect -5873 9520 -5551 9521
rect -5873 9200 -5872 9520
rect -5552 9200 -5551 9520
rect -5873 9199 -5551 9200
rect -6292 9132 -6196 9148
rect -5280 9148 -5264 9572
rect -5200 9148 -5184 9572
rect -4268 9572 -4172 9588
rect -4861 9520 -4539 9521
rect -4861 9200 -4860 9520
rect -4540 9200 -4539 9520
rect -4861 9199 -4539 9200
rect -5280 9132 -5184 9148
rect -4268 9148 -4252 9572
rect -4188 9148 -4172 9572
rect -3256 9572 -3160 9588
rect -3849 9520 -3527 9521
rect -3849 9200 -3848 9520
rect -3528 9200 -3527 9520
rect -3849 9199 -3527 9200
rect -4268 9132 -4172 9148
rect -3256 9148 -3240 9572
rect -3176 9148 -3160 9572
rect -2244 9572 -2148 9588
rect -2837 9520 -2515 9521
rect -2837 9200 -2836 9520
rect -2516 9200 -2515 9520
rect -2837 9199 -2515 9200
rect -3256 9132 -3160 9148
rect -2244 9148 -2228 9572
rect -2164 9148 -2148 9572
rect -1232 9572 -1136 9588
rect -1825 9520 -1503 9521
rect -1825 9200 -1824 9520
rect -1504 9200 -1503 9520
rect -1825 9199 -1503 9200
rect -2244 9132 -2148 9148
rect -1232 9148 -1216 9572
rect -1152 9148 -1136 9572
rect -220 9572 -124 9588
rect -813 9520 -491 9521
rect -813 9200 -812 9520
rect -492 9200 -491 9520
rect -813 9199 -491 9200
rect -1232 9132 -1136 9148
rect -220 9148 -204 9572
rect -140 9148 -124 9572
rect 792 9572 888 9588
rect 199 9520 521 9521
rect 199 9200 200 9520
rect 520 9200 521 9520
rect 199 9199 521 9200
rect -220 9132 -124 9148
rect 792 9148 808 9572
rect 872 9148 888 9572
rect 1804 9572 1900 9588
rect 1211 9520 1533 9521
rect 1211 9200 1212 9520
rect 1532 9200 1533 9520
rect 1211 9199 1533 9200
rect 792 9132 888 9148
rect 1804 9148 1820 9572
rect 1884 9148 1900 9572
rect 2816 9572 2912 9588
rect 2223 9520 2545 9521
rect 2223 9200 2224 9520
rect 2544 9200 2545 9520
rect 2223 9199 2545 9200
rect 1804 9132 1900 9148
rect 2816 9148 2832 9572
rect 2896 9148 2912 9572
rect 3828 9572 3924 9588
rect 3235 9520 3557 9521
rect 3235 9200 3236 9520
rect 3556 9200 3557 9520
rect 3235 9199 3557 9200
rect 2816 9132 2912 9148
rect 3828 9148 3844 9572
rect 3908 9148 3924 9572
rect 4840 9572 4936 9588
rect 4247 9520 4569 9521
rect 4247 9200 4248 9520
rect 4568 9200 4569 9520
rect 4247 9199 4569 9200
rect 3828 9132 3924 9148
rect 4840 9148 4856 9572
rect 4920 9148 4936 9572
rect 5852 9572 5948 9588
rect 5259 9520 5581 9521
rect 5259 9200 5260 9520
rect 5580 9200 5581 9520
rect 5259 9199 5581 9200
rect 4840 9132 4936 9148
rect 5852 9148 5868 9572
rect 5932 9148 5948 9572
rect 6864 9572 6960 9588
rect 6271 9520 6593 9521
rect 6271 9200 6272 9520
rect 6592 9200 6593 9520
rect 6271 9199 6593 9200
rect 5852 9132 5948 9148
rect 6864 9148 6880 9572
rect 6944 9148 6960 9572
rect 7876 9572 7972 9588
rect 7283 9520 7605 9521
rect 7283 9200 7284 9520
rect 7604 9200 7605 9520
rect 7283 9199 7605 9200
rect 6864 9132 6960 9148
rect 7876 9148 7892 9572
rect 7956 9148 7972 9572
rect 8888 9572 8984 9588
rect 8295 9520 8617 9521
rect 8295 9200 8296 9520
rect 8616 9200 8617 9520
rect 8295 9199 8617 9200
rect 7876 9132 7972 9148
rect 8888 9148 8904 9572
rect 8968 9148 8984 9572
rect 9900 9572 9996 9588
rect 9307 9520 9629 9521
rect 9307 9200 9308 9520
rect 9628 9200 9629 9520
rect 9307 9199 9629 9200
rect 8888 9132 8984 9148
rect 9900 9148 9916 9572
rect 9980 9148 9996 9572
rect 10912 9572 11008 9588
rect 10319 9520 10641 9521
rect 10319 9200 10320 9520
rect 10640 9200 10641 9520
rect 10319 9199 10641 9200
rect 9900 9132 9996 9148
rect 10912 9148 10928 9572
rect 10992 9148 11008 9572
rect 11924 9572 12020 9588
rect 11331 9520 11653 9521
rect 11331 9200 11332 9520
rect 11652 9200 11653 9520
rect 11331 9199 11653 9200
rect 10912 9132 11008 9148
rect 11924 9148 11940 9572
rect 12004 9148 12020 9572
rect 12936 9572 13032 9588
rect 12343 9520 12665 9521
rect 12343 9200 12344 9520
rect 12664 9200 12665 9520
rect 12343 9199 12665 9200
rect 11924 9132 12020 9148
rect 12936 9148 12952 9572
rect 13016 9148 13032 9572
rect 13948 9572 14044 9588
rect 13355 9520 13677 9521
rect 13355 9200 13356 9520
rect 13676 9200 13677 9520
rect 13355 9199 13677 9200
rect 12936 9132 13032 9148
rect 13948 9148 13964 9572
rect 14028 9148 14044 9572
rect 14960 9572 15056 9588
rect 14367 9520 14689 9521
rect 14367 9200 14368 9520
rect 14688 9200 14689 9520
rect 14367 9199 14689 9200
rect 13948 9132 14044 9148
rect 14960 9148 14976 9572
rect 15040 9148 15056 9572
rect 15972 9572 16068 9588
rect 15379 9520 15701 9521
rect 15379 9200 15380 9520
rect 15700 9200 15701 9520
rect 15379 9199 15701 9200
rect 14960 9132 15056 9148
rect 15972 9148 15988 9572
rect 16052 9148 16068 9572
rect 16984 9572 17080 9588
rect 16391 9520 16713 9521
rect 16391 9200 16392 9520
rect 16712 9200 16713 9520
rect 16391 9199 16713 9200
rect 15972 9132 16068 9148
rect 16984 9148 17000 9572
rect 17064 9148 17080 9572
rect 16984 9132 17080 9148
rect -16412 8852 -16316 8868
rect -17005 8800 -16683 8801
rect -17005 8480 -17004 8800
rect -16684 8480 -16683 8800
rect -17005 8479 -16683 8480
rect -16412 8428 -16396 8852
rect -16332 8428 -16316 8852
rect -15400 8852 -15304 8868
rect -15993 8800 -15671 8801
rect -15993 8480 -15992 8800
rect -15672 8480 -15671 8800
rect -15993 8479 -15671 8480
rect -16412 8412 -16316 8428
rect -15400 8428 -15384 8852
rect -15320 8428 -15304 8852
rect -14388 8852 -14292 8868
rect -14981 8800 -14659 8801
rect -14981 8480 -14980 8800
rect -14660 8480 -14659 8800
rect -14981 8479 -14659 8480
rect -15400 8412 -15304 8428
rect -14388 8428 -14372 8852
rect -14308 8428 -14292 8852
rect -13376 8852 -13280 8868
rect -13969 8800 -13647 8801
rect -13969 8480 -13968 8800
rect -13648 8480 -13647 8800
rect -13969 8479 -13647 8480
rect -14388 8412 -14292 8428
rect -13376 8428 -13360 8852
rect -13296 8428 -13280 8852
rect -12364 8852 -12268 8868
rect -12957 8800 -12635 8801
rect -12957 8480 -12956 8800
rect -12636 8480 -12635 8800
rect -12957 8479 -12635 8480
rect -13376 8412 -13280 8428
rect -12364 8428 -12348 8852
rect -12284 8428 -12268 8852
rect -11352 8852 -11256 8868
rect -11945 8800 -11623 8801
rect -11945 8480 -11944 8800
rect -11624 8480 -11623 8800
rect -11945 8479 -11623 8480
rect -12364 8412 -12268 8428
rect -11352 8428 -11336 8852
rect -11272 8428 -11256 8852
rect -10340 8852 -10244 8868
rect -10933 8800 -10611 8801
rect -10933 8480 -10932 8800
rect -10612 8480 -10611 8800
rect -10933 8479 -10611 8480
rect -11352 8412 -11256 8428
rect -10340 8428 -10324 8852
rect -10260 8428 -10244 8852
rect -9328 8852 -9232 8868
rect -9921 8800 -9599 8801
rect -9921 8480 -9920 8800
rect -9600 8480 -9599 8800
rect -9921 8479 -9599 8480
rect -10340 8412 -10244 8428
rect -9328 8428 -9312 8852
rect -9248 8428 -9232 8852
rect -8316 8852 -8220 8868
rect -8909 8800 -8587 8801
rect -8909 8480 -8908 8800
rect -8588 8480 -8587 8800
rect -8909 8479 -8587 8480
rect -9328 8412 -9232 8428
rect -8316 8428 -8300 8852
rect -8236 8428 -8220 8852
rect -7304 8852 -7208 8868
rect -7897 8800 -7575 8801
rect -7897 8480 -7896 8800
rect -7576 8480 -7575 8800
rect -7897 8479 -7575 8480
rect -8316 8412 -8220 8428
rect -7304 8428 -7288 8852
rect -7224 8428 -7208 8852
rect -6292 8852 -6196 8868
rect -6885 8800 -6563 8801
rect -6885 8480 -6884 8800
rect -6564 8480 -6563 8800
rect -6885 8479 -6563 8480
rect -7304 8412 -7208 8428
rect -6292 8428 -6276 8852
rect -6212 8428 -6196 8852
rect -5280 8852 -5184 8868
rect -5873 8800 -5551 8801
rect -5873 8480 -5872 8800
rect -5552 8480 -5551 8800
rect -5873 8479 -5551 8480
rect -6292 8412 -6196 8428
rect -5280 8428 -5264 8852
rect -5200 8428 -5184 8852
rect -4268 8852 -4172 8868
rect -4861 8800 -4539 8801
rect -4861 8480 -4860 8800
rect -4540 8480 -4539 8800
rect -4861 8479 -4539 8480
rect -5280 8412 -5184 8428
rect -4268 8428 -4252 8852
rect -4188 8428 -4172 8852
rect -3256 8852 -3160 8868
rect -3849 8800 -3527 8801
rect -3849 8480 -3848 8800
rect -3528 8480 -3527 8800
rect -3849 8479 -3527 8480
rect -4268 8412 -4172 8428
rect -3256 8428 -3240 8852
rect -3176 8428 -3160 8852
rect -2244 8852 -2148 8868
rect -2837 8800 -2515 8801
rect -2837 8480 -2836 8800
rect -2516 8480 -2515 8800
rect -2837 8479 -2515 8480
rect -3256 8412 -3160 8428
rect -2244 8428 -2228 8852
rect -2164 8428 -2148 8852
rect -1232 8852 -1136 8868
rect -1825 8800 -1503 8801
rect -1825 8480 -1824 8800
rect -1504 8480 -1503 8800
rect -1825 8479 -1503 8480
rect -2244 8412 -2148 8428
rect -1232 8428 -1216 8852
rect -1152 8428 -1136 8852
rect -220 8852 -124 8868
rect -813 8800 -491 8801
rect -813 8480 -812 8800
rect -492 8480 -491 8800
rect -813 8479 -491 8480
rect -1232 8412 -1136 8428
rect -220 8428 -204 8852
rect -140 8428 -124 8852
rect 792 8852 888 8868
rect 199 8800 521 8801
rect 199 8480 200 8800
rect 520 8480 521 8800
rect 199 8479 521 8480
rect -220 8412 -124 8428
rect 792 8428 808 8852
rect 872 8428 888 8852
rect 1804 8852 1900 8868
rect 1211 8800 1533 8801
rect 1211 8480 1212 8800
rect 1532 8480 1533 8800
rect 1211 8479 1533 8480
rect 792 8412 888 8428
rect 1804 8428 1820 8852
rect 1884 8428 1900 8852
rect 2816 8852 2912 8868
rect 2223 8800 2545 8801
rect 2223 8480 2224 8800
rect 2544 8480 2545 8800
rect 2223 8479 2545 8480
rect 1804 8412 1900 8428
rect 2816 8428 2832 8852
rect 2896 8428 2912 8852
rect 3828 8852 3924 8868
rect 3235 8800 3557 8801
rect 3235 8480 3236 8800
rect 3556 8480 3557 8800
rect 3235 8479 3557 8480
rect 2816 8412 2912 8428
rect 3828 8428 3844 8852
rect 3908 8428 3924 8852
rect 4840 8852 4936 8868
rect 4247 8800 4569 8801
rect 4247 8480 4248 8800
rect 4568 8480 4569 8800
rect 4247 8479 4569 8480
rect 3828 8412 3924 8428
rect 4840 8428 4856 8852
rect 4920 8428 4936 8852
rect 5852 8852 5948 8868
rect 5259 8800 5581 8801
rect 5259 8480 5260 8800
rect 5580 8480 5581 8800
rect 5259 8479 5581 8480
rect 4840 8412 4936 8428
rect 5852 8428 5868 8852
rect 5932 8428 5948 8852
rect 6864 8852 6960 8868
rect 6271 8800 6593 8801
rect 6271 8480 6272 8800
rect 6592 8480 6593 8800
rect 6271 8479 6593 8480
rect 5852 8412 5948 8428
rect 6864 8428 6880 8852
rect 6944 8428 6960 8852
rect 7876 8852 7972 8868
rect 7283 8800 7605 8801
rect 7283 8480 7284 8800
rect 7604 8480 7605 8800
rect 7283 8479 7605 8480
rect 6864 8412 6960 8428
rect 7876 8428 7892 8852
rect 7956 8428 7972 8852
rect 8888 8852 8984 8868
rect 8295 8800 8617 8801
rect 8295 8480 8296 8800
rect 8616 8480 8617 8800
rect 8295 8479 8617 8480
rect 7876 8412 7972 8428
rect 8888 8428 8904 8852
rect 8968 8428 8984 8852
rect 9900 8852 9996 8868
rect 9307 8800 9629 8801
rect 9307 8480 9308 8800
rect 9628 8480 9629 8800
rect 9307 8479 9629 8480
rect 8888 8412 8984 8428
rect 9900 8428 9916 8852
rect 9980 8428 9996 8852
rect 10912 8852 11008 8868
rect 10319 8800 10641 8801
rect 10319 8480 10320 8800
rect 10640 8480 10641 8800
rect 10319 8479 10641 8480
rect 9900 8412 9996 8428
rect 10912 8428 10928 8852
rect 10992 8428 11008 8852
rect 11924 8852 12020 8868
rect 11331 8800 11653 8801
rect 11331 8480 11332 8800
rect 11652 8480 11653 8800
rect 11331 8479 11653 8480
rect 10912 8412 11008 8428
rect 11924 8428 11940 8852
rect 12004 8428 12020 8852
rect 12936 8852 13032 8868
rect 12343 8800 12665 8801
rect 12343 8480 12344 8800
rect 12664 8480 12665 8800
rect 12343 8479 12665 8480
rect 11924 8412 12020 8428
rect 12936 8428 12952 8852
rect 13016 8428 13032 8852
rect 13948 8852 14044 8868
rect 13355 8800 13677 8801
rect 13355 8480 13356 8800
rect 13676 8480 13677 8800
rect 13355 8479 13677 8480
rect 12936 8412 13032 8428
rect 13948 8428 13964 8852
rect 14028 8428 14044 8852
rect 14960 8852 15056 8868
rect 14367 8800 14689 8801
rect 14367 8480 14368 8800
rect 14688 8480 14689 8800
rect 14367 8479 14689 8480
rect 13948 8412 14044 8428
rect 14960 8428 14976 8852
rect 15040 8428 15056 8852
rect 15972 8852 16068 8868
rect 15379 8800 15701 8801
rect 15379 8480 15380 8800
rect 15700 8480 15701 8800
rect 15379 8479 15701 8480
rect 14960 8412 15056 8428
rect 15972 8428 15988 8852
rect 16052 8428 16068 8852
rect 16984 8852 17080 8868
rect 16391 8800 16713 8801
rect 16391 8480 16392 8800
rect 16712 8480 16713 8800
rect 16391 8479 16713 8480
rect 15972 8412 16068 8428
rect 16984 8428 17000 8852
rect 17064 8428 17080 8852
rect 16984 8412 17080 8428
rect -16412 8132 -16316 8148
rect -17005 8080 -16683 8081
rect -17005 7760 -17004 8080
rect -16684 7760 -16683 8080
rect -17005 7759 -16683 7760
rect -16412 7708 -16396 8132
rect -16332 7708 -16316 8132
rect -15400 8132 -15304 8148
rect -15993 8080 -15671 8081
rect -15993 7760 -15992 8080
rect -15672 7760 -15671 8080
rect -15993 7759 -15671 7760
rect -16412 7692 -16316 7708
rect -15400 7708 -15384 8132
rect -15320 7708 -15304 8132
rect -14388 8132 -14292 8148
rect -14981 8080 -14659 8081
rect -14981 7760 -14980 8080
rect -14660 7760 -14659 8080
rect -14981 7759 -14659 7760
rect -15400 7692 -15304 7708
rect -14388 7708 -14372 8132
rect -14308 7708 -14292 8132
rect -13376 8132 -13280 8148
rect -13969 8080 -13647 8081
rect -13969 7760 -13968 8080
rect -13648 7760 -13647 8080
rect -13969 7759 -13647 7760
rect -14388 7692 -14292 7708
rect -13376 7708 -13360 8132
rect -13296 7708 -13280 8132
rect -12364 8132 -12268 8148
rect -12957 8080 -12635 8081
rect -12957 7760 -12956 8080
rect -12636 7760 -12635 8080
rect -12957 7759 -12635 7760
rect -13376 7692 -13280 7708
rect -12364 7708 -12348 8132
rect -12284 7708 -12268 8132
rect -11352 8132 -11256 8148
rect -11945 8080 -11623 8081
rect -11945 7760 -11944 8080
rect -11624 7760 -11623 8080
rect -11945 7759 -11623 7760
rect -12364 7692 -12268 7708
rect -11352 7708 -11336 8132
rect -11272 7708 -11256 8132
rect -10340 8132 -10244 8148
rect -10933 8080 -10611 8081
rect -10933 7760 -10932 8080
rect -10612 7760 -10611 8080
rect -10933 7759 -10611 7760
rect -11352 7692 -11256 7708
rect -10340 7708 -10324 8132
rect -10260 7708 -10244 8132
rect -9328 8132 -9232 8148
rect -9921 8080 -9599 8081
rect -9921 7760 -9920 8080
rect -9600 7760 -9599 8080
rect -9921 7759 -9599 7760
rect -10340 7692 -10244 7708
rect -9328 7708 -9312 8132
rect -9248 7708 -9232 8132
rect -8316 8132 -8220 8148
rect -8909 8080 -8587 8081
rect -8909 7760 -8908 8080
rect -8588 7760 -8587 8080
rect -8909 7759 -8587 7760
rect -9328 7692 -9232 7708
rect -8316 7708 -8300 8132
rect -8236 7708 -8220 8132
rect -7304 8132 -7208 8148
rect -7897 8080 -7575 8081
rect -7897 7760 -7896 8080
rect -7576 7760 -7575 8080
rect -7897 7759 -7575 7760
rect -8316 7692 -8220 7708
rect -7304 7708 -7288 8132
rect -7224 7708 -7208 8132
rect -6292 8132 -6196 8148
rect -6885 8080 -6563 8081
rect -6885 7760 -6884 8080
rect -6564 7760 -6563 8080
rect -6885 7759 -6563 7760
rect -7304 7692 -7208 7708
rect -6292 7708 -6276 8132
rect -6212 7708 -6196 8132
rect -5280 8132 -5184 8148
rect -5873 8080 -5551 8081
rect -5873 7760 -5872 8080
rect -5552 7760 -5551 8080
rect -5873 7759 -5551 7760
rect -6292 7692 -6196 7708
rect -5280 7708 -5264 8132
rect -5200 7708 -5184 8132
rect -4268 8132 -4172 8148
rect -4861 8080 -4539 8081
rect -4861 7760 -4860 8080
rect -4540 7760 -4539 8080
rect -4861 7759 -4539 7760
rect -5280 7692 -5184 7708
rect -4268 7708 -4252 8132
rect -4188 7708 -4172 8132
rect -3256 8132 -3160 8148
rect -3849 8080 -3527 8081
rect -3849 7760 -3848 8080
rect -3528 7760 -3527 8080
rect -3849 7759 -3527 7760
rect -4268 7692 -4172 7708
rect -3256 7708 -3240 8132
rect -3176 7708 -3160 8132
rect -2244 8132 -2148 8148
rect -2837 8080 -2515 8081
rect -2837 7760 -2836 8080
rect -2516 7760 -2515 8080
rect -2837 7759 -2515 7760
rect -3256 7692 -3160 7708
rect -2244 7708 -2228 8132
rect -2164 7708 -2148 8132
rect -1232 8132 -1136 8148
rect -1825 8080 -1503 8081
rect -1825 7760 -1824 8080
rect -1504 7760 -1503 8080
rect -1825 7759 -1503 7760
rect -2244 7692 -2148 7708
rect -1232 7708 -1216 8132
rect -1152 7708 -1136 8132
rect -220 8132 -124 8148
rect -813 8080 -491 8081
rect -813 7760 -812 8080
rect -492 7760 -491 8080
rect -813 7759 -491 7760
rect -1232 7692 -1136 7708
rect -220 7708 -204 8132
rect -140 7708 -124 8132
rect 792 8132 888 8148
rect 199 8080 521 8081
rect 199 7760 200 8080
rect 520 7760 521 8080
rect 199 7759 521 7760
rect -220 7692 -124 7708
rect 792 7708 808 8132
rect 872 7708 888 8132
rect 1804 8132 1900 8148
rect 1211 8080 1533 8081
rect 1211 7760 1212 8080
rect 1532 7760 1533 8080
rect 1211 7759 1533 7760
rect 792 7692 888 7708
rect 1804 7708 1820 8132
rect 1884 7708 1900 8132
rect 2816 8132 2912 8148
rect 2223 8080 2545 8081
rect 2223 7760 2224 8080
rect 2544 7760 2545 8080
rect 2223 7759 2545 7760
rect 1804 7692 1900 7708
rect 2816 7708 2832 8132
rect 2896 7708 2912 8132
rect 3828 8132 3924 8148
rect 3235 8080 3557 8081
rect 3235 7760 3236 8080
rect 3556 7760 3557 8080
rect 3235 7759 3557 7760
rect 2816 7692 2912 7708
rect 3828 7708 3844 8132
rect 3908 7708 3924 8132
rect 4840 8132 4936 8148
rect 4247 8080 4569 8081
rect 4247 7760 4248 8080
rect 4568 7760 4569 8080
rect 4247 7759 4569 7760
rect 3828 7692 3924 7708
rect 4840 7708 4856 8132
rect 4920 7708 4936 8132
rect 5852 8132 5948 8148
rect 5259 8080 5581 8081
rect 5259 7760 5260 8080
rect 5580 7760 5581 8080
rect 5259 7759 5581 7760
rect 4840 7692 4936 7708
rect 5852 7708 5868 8132
rect 5932 7708 5948 8132
rect 6864 8132 6960 8148
rect 6271 8080 6593 8081
rect 6271 7760 6272 8080
rect 6592 7760 6593 8080
rect 6271 7759 6593 7760
rect 5852 7692 5948 7708
rect 6864 7708 6880 8132
rect 6944 7708 6960 8132
rect 7876 8132 7972 8148
rect 7283 8080 7605 8081
rect 7283 7760 7284 8080
rect 7604 7760 7605 8080
rect 7283 7759 7605 7760
rect 6864 7692 6960 7708
rect 7876 7708 7892 8132
rect 7956 7708 7972 8132
rect 8888 8132 8984 8148
rect 8295 8080 8617 8081
rect 8295 7760 8296 8080
rect 8616 7760 8617 8080
rect 8295 7759 8617 7760
rect 7876 7692 7972 7708
rect 8888 7708 8904 8132
rect 8968 7708 8984 8132
rect 9900 8132 9996 8148
rect 9307 8080 9629 8081
rect 9307 7760 9308 8080
rect 9628 7760 9629 8080
rect 9307 7759 9629 7760
rect 8888 7692 8984 7708
rect 9900 7708 9916 8132
rect 9980 7708 9996 8132
rect 10912 8132 11008 8148
rect 10319 8080 10641 8081
rect 10319 7760 10320 8080
rect 10640 7760 10641 8080
rect 10319 7759 10641 7760
rect 9900 7692 9996 7708
rect 10912 7708 10928 8132
rect 10992 7708 11008 8132
rect 11924 8132 12020 8148
rect 11331 8080 11653 8081
rect 11331 7760 11332 8080
rect 11652 7760 11653 8080
rect 11331 7759 11653 7760
rect 10912 7692 11008 7708
rect 11924 7708 11940 8132
rect 12004 7708 12020 8132
rect 12936 8132 13032 8148
rect 12343 8080 12665 8081
rect 12343 7760 12344 8080
rect 12664 7760 12665 8080
rect 12343 7759 12665 7760
rect 11924 7692 12020 7708
rect 12936 7708 12952 8132
rect 13016 7708 13032 8132
rect 13948 8132 14044 8148
rect 13355 8080 13677 8081
rect 13355 7760 13356 8080
rect 13676 7760 13677 8080
rect 13355 7759 13677 7760
rect 12936 7692 13032 7708
rect 13948 7708 13964 8132
rect 14028 7708 14044 8132
rect 14960 8132 15056 8148
rect 14367 8080 14689 8081
rect 14367 7760 14368 8080
rect 14688 7760 14689 8080
rect 14367 7759 14689 7760
rect 13948 7692 14044 7708
rect 14960 7708 14976 8132
rect 15040 7708 15056 8132
rect 15972 8132 16068 8148
rect 15379 8080 15701 8081
rect 15379 7760 15380 8080
rect 15700 7760 15701 8080
rect 15379 7759 15701 7760
rect 14960 7692 15056 7708
rect 15972 7708 15988 8132
rect 16052 7708 16068 8132
rect 16984 8132 17080 8148
rect 16391 8080 16713 8081
rect 16391 7760 16392 8080
rect 16712 7760 16713 8080
rect 16391 7759 16713 7760
rect 15972 7692 16068 7708
rect 16984 7708 17000 8132
rect 17064 7708 17080 8132
rect 16984 7692 17080 7708
rect -16412 7412 -16316 7428
rect -17005 7360 -16683 7361
rect -17005 7040 -17004 7360
rect -16684 7040 -16683 7360
rect -17005 7039 -16683 7040
rect -16412 6988 -16396 7412
rect -16332 6988 -16316 7412
rect -15400 7412 -15304 7428
rect -15993 7360 -15671 7361
rect -15993 7040 -15992 7360
rect -15672 7040 -15671 7360
rect -15993 7039 -15671 7040
rect -16412 6972 -16316 6988
rect -15400 6988 -15384 7412
rect -15320 6988 -15304 7412
rect -14388 7412 -14292 7428
rect -14981 7360 -14659 7361
rect -14981 7040 -14980 7360
rect -14660 7040 -14659 7360
rect -14981 7039 -14659 7040
rect -15400 6972 -15304 6988
rect -14388 6988 -14372 7412
rect -14308 6988 -14292 7412
rect -13376 7412 -13280 7428
rect -13969 7360 -13647 7361
rect -13969 7040 -13968 7360
rect -13648 7040 -13647 7360
rect -13969 7039 -13647 7040
rect -14388 6972 -14292 6988
rect -13376 6988 -13360 7412
rect -13296 6988 -13280 7412
rect -12364 7412 -12268 7428
rect -12957 7360 -12635 7361
rect -12957 7040 -12956 7360
rect -12636 7040 -12635 7360
rect -12957 7039 -12635 7040
rect -13376 6972 -13280 6988
rect -12364 6988 -12348 7412
rect -12284 6988 -12268 7412
rect -11352 7412 -11256 7428
rect -11945 7360 -11623 7361
rect -11945 7040 -11944 7360
rect -11624 7040 -11623 7360
rect -11945 7039 -11623 7040
rect -12364 6972 -12268 6988
rect -11352 6988 -11336 7412
rect -11272 6988 -11256 7412
rect -10340 7412 -10244 7428
rect -10933 7360 -10611 7361
rect -10933 7040 -10932 7360
rect -10612 7040 -10611 7360
rect -10933 7039 -10611 7040
rect -11352 6972 -11256 6988
rect -10340 6988 -10324 7412
rect -10260 6988 -10244 7412
rect -9328 7412 -9232 7428
rect -9921 7360 -9599 7361
rect -9921 7040 -9920 7360
rect -9600 7040 -9599 7360
rect -9921 7039 -9599 7040
rect -10340 6972 -10244 6988
rect -9328 6988 -9312 7412
rect -9248 6988 -9232 7412
rect -8316 7412 -8220 7428
rect -8909 7360 -8587 7361
rect -8909 7040 -8908 7360
rect -8588 7040 -8587 7360
rect -8909 7039 -8587 7040
rect -9328 6972 -9232 6988
rect -8316 6988 -8300 7412
rect -8236 6988 -8220 7412
rect -7304 7412 -7208 7428
rect -7897 7360 -7575 7361
rect -7897 7040 -7896 7360
rect -7576 7040 -7575 7360
rect -7897 7039 -7575 7040
rect -8316 6972 -8220 6988
rect -7304 6988 -7288 7412
rect -7224 6988 -7208 7412
rect -6292 7412 -6196 7428
rect -6885 7360 -6563 7361
rect -6885 7040 -6884 7360
rect -6564 7040 -6563 7360
rect -6885 7039 -6563 7040
rect -7304 6972 -7208 6988
rect -6292 6988 -6276 7412
rect -6212 6988 -6196 7412
rect -5280 7412 -5184 7428
rect -5873 7360 -5551 7361
rect -5873 7040 -5872 7360
rect -5552 7040 -5551 7360
rect -5873 7039 -5551 7040
rect -6292 6972 -6196 6988
rect -5280 6988 -5264 7412
rect -5200 6988 -5184 7412
rect -4268 7412 -4172 7428
rect -4861 7360 -4539 7361
rect -4861 7040 -4860 7360
rect -4540 7040 -4539 7360
rect -4861 7039 -4539 7040
rect -5280 6972 -5184 6988
rect -4268 6988 -4252 7412
rect -4188 6988 -4172 7412
rect -3256 7412 -3160 7428
rect -3849 7360 -3527 7361
rect -3849 7040 -3848 7360
rect -3528 7040 -3527 7360
rect -3849 7039 -3527 7040
rect -4268 6972 -4172 6988
rect -3256 6988 -3240 7412
rect -3176 6988 -3160 7412
rect -2244 7412 -2148 7428
rect -2837 7360 -2515 7361
rect -2837 7040 -2836 7360
rect -2516 7040 -2515 7360
rect -2837 7039 -2515 7040
rect -3256 6972 -3160 6988
rect -2244 6988 -2228 7412
rect -2164 6988 -2148 7412
rect -1232 7412 -1136 7428
rect -1825 7360 -1503 7361
rect -1825 7040 -1824 7360
rect -1504 7040 -1503 7360
rect -1825 7039 -1503 7040
rect -2244 6972 -2148 6988
rect -1232 6988 -1216 7412
rect -1152 6988 -1136 7412
rect -220 7412 -124 7428
rect -813 7360 -491 7361
rect -813 7040 -812 7360
rect -492 7040 -491 7360
rect -813 7039 -491 7040
rect -1232 6972 -1136 6988
rect -220 6988 -204 7412
rect -140 6988 -124 7412
rect 792 7412 888 7428
rect 199 7360 521 7361
rect 199 7040 200 7360
rect 520 7040 521 7360
rect 199 7039 521 7040
rect -220 6972 -124 6988
rect 792 6988 808 7412
rect 872 6988 888 7412
rect 1804 7412 1900 7428
rect 1211 7360 1533 7361
rect 1211 7040 1212 7360
rect 1532 7040 1533 7360
rect 1211 7039 1533 7040
rect 792 6972 888 6988
rect 1804 6988 1820 7412
rect 1884 6988 1900 7412
rect 2816 7412 2912 7428
rect 2223 7360 2545 7361
rect 2223 7040 2224 7360
rect 2544 7040 2545 7360
rect 2223 7039 2545 7040
rect 1804 6972 1900 6988
rect 2816 6988 2832 7412
rect 2896 6988 2912 7412
rect 3828 7412 3924 7428
rect 3235 7360 3557 7361
rect 3235 7040 3236 7360
rect 3556 7040 3557 7360
rect 3235 7039 3557 7040
rect 2816 6972 2912 6988
rect 3828 6988 3844 7412
rect 3908 6988 3924 7412
rect 4840 7412 4936 7428
rect 4247 7360 4569 7361
rect 4247 7040 4248 7360
rect 4568 7040 4569 7360
rect 4247 7039 4569 7040
rect 3828 6972 3924 6988
rect 4840 6988 4856 7412
rect 4920 6988 4936 7412
rect 5852 7412 5948 7428
rect 5259 7360 5581 7361
rect 5259 7040 5260 7360
rect 5580 7040 5581 7360
rect 5259 7039 5581 7040
rect 4840 6972 4936 6988
rect 5852 6988 5868 7412
rect 5932 6988 5948 7412
rect 6864 7412 6960 7428
rect 6271 7360 6593 7361
rect 6271 7040 6272 7360
rect 6592 7040 6593 7360
rect 6271 7039 6593 7040
rect 5852 6972 5948 6988
rect 6864 6988 6880 7412
rect 6944 6988 6960 7412
rect 7876 7412 7972 7428
rect 7283 7360 7605 7361
rect 7283 7040 7284 7360
rect 7604 7040 7605 7360
rect 7283 7039 7605 7040
rect 6864 6972 6960 6988
rect 7876 6988 7892 7412
rect 7956 6988 7972 7412
rect 8888 7412 8984 7428
rect 8295 7360 8617 7361
rect 8295 7040 8296 7360
rect 8616 7040 8617 7360
rect 8295 7039 8617 7040
rect 7876 6972 7972 6988
rect 8888 6988 8904 7412
rect 8968 6988 8984 7412
rect 9900 7412 9996 7428
rect 9307 7360 9629 7361
rect 9307 7040 9308 7360
rect 9628 7040 9629 7360
rect 9307 7039 9629 7040
rect 8888 6972 8984 6988
rect 9900 6988 9916 7412
rect 9980 6988 9996 7412
rect 10912 7412 11008 7428
rect 10319 7360 10641 7361
rect 10319 7040 10320 7360
rect 10640 7040 10641 7360
rect 10319 7039 10641 7040
rect 9900 6972 9996 6988
rect 10912 6988 10928 7412
rect 10992 6988 11008 7412
rect 11924 7412 12020 7428
rect 11331 7360 11653 7361
rect 11331 7040 11332 7360
rect 11652 7040 11653 7360
rect 11331 7039 11653 7040
rect 10912 6972 11008 6988
rect 11924 6988 11940 7412
rect 12004 6988 12020 7412
rect 12936 7412 13032 7428
rect 12343 7360 12665 7361
rect 12343 7040 12344 7360
rect 12664 7040 12665 7360
rect 12343 7039 12665 7040
rect 11924 6972 12020 6988
rect 12936 6988 12952 7412
rect 13016 6988 13032 7412
rect 13948 7412 14044 7428
rect 13355 7360 13677 7361
rect 13355 7040 13356 7360
rect 13676 7040 13677 7360
rect 13355 7039 13677 7040
rect 12936 6972 13032 6988
rect 13948 6988 13964 7412
rect 14028 6988 14044 7412
rect 14960 7412 15056 7428
rect 14367 7360 14689 7361
rect 14367 7040 14368 7360
rect 14688 7040 14689 7360
rect 14367 7039 14689 7040
rect 13948 6972 14044 6988
rect 14960 6988 14976 7412
rect 15040 6988 15056 7412
rect 15972 7412 16068 7428
rect 15379 7360 15701 7361
rect 15379 7040 15380 7360
rect 15700 7040 15701 7360
rect 15379 7039 15701 7040
rect 14960 6972 15056 6988
rect 15972 6988 15988 7412
rect 16052 6988 16068 7412
rect 16984 7412 17080 7428
rect 16391 7360 16713 7361
rect 16391 7040 16392 7360
rect 16712 7040 16713 7360
rect 16391 7039 16713 7040
rect 15972 6972 16068 6988
rect 16984 6988 17000 7412
rect 17064 6988 17080 7412
rect 16984 6972 17080 6988
rect -16412 6692 -16316 6708
rect -17005 6640 -16683 6641
rect -17005 6320 -17004 6640
rect -16684 6320 -16683 6640
rect -17005 6319 -16683 6320
rect -16412 6268 -16396 6692
rect -16332 6268 -16316 6692
rect -15400 6692 -15304 6708
rect -15993 6640 -15671 6641
rect -15993 6320 -15992 6640
rect -15672 6320 -15671 6640
rect -15993 6319 -15671 6320
rect -16412 6252 -16316 6268
rect -15400 6268 -15384 6692
rect -15320 6268 -15304 6692
rect -14388 6692 -14292 6708
rect -14981 6640 -14659 6641
rect -14981 6320 -14980 6640
rect -14660 6320 -14659 6640
rect -14981 6319 -14659 6320
rect -15400 6252 -15304 6268
rect -14388 6268 -14372 6692
rect -14308 6268 -14292 6692
rect -13376 6692 -13280 6708
rect -13969 6640 -13647 6641
rect -13969 6320 -13968 6640
rect -13648 6320 -13647 6640
rect -13969 6319 -13647 6320
rect -14388 6252 -14292 6268
rect -13376 6268 -13360 6692
rect -13296 6268 -13280 6692
rect -12364 6692 -12268 6708
rect -12957 6640 -12635 6641
rect -12957 6320 -12956 6640
rect -12636 6320 -12635 6640
rect -12957 6319 -12635 6320
rect -13376 6252 -13280 6268
rect -12364 6268 -12348 6692
rect -12284 6268 -12268 6692
rect -11352 6692 -11256 6708
rect -11945 6640 -11623 6641
rect -11945 6320 -11944 6640
rect -11624 6320 -11623 6640
rect -11945 6319 -11623 6320
rect -12364 6252 -12268 6268
rect -11352 6268 -11336 6692
rect -11272 6268 -11256 6692
rect -10340 6692 -10244 6708
rect -10933 6640 -10611 6641
rect -10933 6320 -10932 6640
rect -10612 6320 -10611 6640
rect -10933 6319 -10611 6320
rect -11352 6252 -11256 6268
rect -10340 6268 -10324 6692
rect -10260 6268 -10244 6692
rect -9328 6692 -9232 6708
rect -9921 6640 -9599 6641
rect -9921 6320 -9920 6640
rect -9600 6320 -9599 6640
rect -9921 6319 -9599 6320
rect -10340 6252 -10244 6268
rect -9328 6268 -9312 6692
rect -9248 6268 -9232 6692
rect -8316 6692 -8220 6708
rect -8909 6640 -8587 6641
rect -8909 6320 -8908 6640
rect -8588 6320 -8587 6640
rect -8909 6319 -8587 6320
rect -9328 6252 -9232 6268
rect -8316 6268 -8300 6692
rect -8236 6268 -8220 6692
rect -7304 6692 -7208 6708
rect -7897 6640 -7575 6641
rect -7897 6320 -7896 6640
rect -7576 6320 -7575 6640
rect -7897 6319 -7575 6320
rect -8316 6252 -8220 6268
rect -7304 6268 -7288 6692
rect -7224 6268 -7208 6692
rect -6292 6692 -6196 6708
rect -6885 6640 -6563 6641
rect -6885 6320 -6884 6640
rect -6564 6320 -6563 6640
rect -6885 6319 -6563 6320
rect -7304 6252 -7208 6268
rect -6292 6268 -6276 6692
rect -6212 6268 -6196 6692
rect -5280 6692 -5184 6708
rect -5873 6640 -5551 6641
rect -5873 6320 -5872 6640
rect -5552 6320 -5551 6640
rect -5873 6319 -5551 6320
rect -6292 6252 -6196 6268
rect -5280 6268 -5264 6692
rect -5200 6268 -5184 6692
rect -4268 6692 -4172 6708
rect -4861 6640 -4539 6641
rect -4861 6320 -4860 6640
rect -4540 6320 -4539 6640
rect -4861 6319 -4539 6320
rect -5280 6252 -5184 6268
rect -4268 6268 -4252 6692
rect -4188 6268 -4172 6692
rect -3256 6692 -3160 6708
rect -3849 6640 -3527 6641
rect -3849 6320 -3848 6640
rect -3528 6320 -3527 6640
rect -3849 6319 -3527 6320
rect -4268 6252 -4172 6268
rect -3256 6268 -3240 6692
rect -3176 6268 -3160 6692
rect -2244 6692 -2148 6708
rect -2837 6640 -2515 6641
rect -2837 6320 -2836 6640
rect -2516 6320 -2515 6640
rect -2837 6319 -2515 6320
rect -3256 6252 -3160 6268
rect -2244 6268 -2228 6692
rect -2164 6268 -2148 6692
rect -1232 6692 -1136 6708
rect -1825 6640 -1503 6641
rect -1825 6320 -1824 6640
rect -1504 6320 -1503 6640
rect -1825 6319 -1503 6320
rect -2244 6252 -2148 6268
rect -1232 6268 -1216 6692
rect -1152 6268 -1136 6692
rect -220 6692 -124 6708
rect -813 6640 -491 6641
rect -813 6320 -812 6640
rect -492 6320 -491 6640
rect -813 6319 -491 6320
rect -1232 6252 -1136 6268
rect -220 6268 -204 6692
rect -140 6268 -124 6692
rect 792 6692 888 6708
rect 199 6640 521 6641
rect 199 6320 200 6640
rect 520 6320 521 6640
rect 199 6319 521 6320
rect -220 6252 -124 6268
rect 792 6268 808 6692
rect 872 6268 888 6692
rect 1804 6692 1900 6708
rect 1211 6640 1533 6641
rect 1211 6320 1212 6640
rect 1532 6320 1533 6640
rect 1211 6319 1533 6320
rect 792 6252 888 6268
rect 1804 6268 1820 6692
rect 1884 6268 1900 6692
rect 2816 6692 2912 6708
rect 2223 6640 2545 6641
rect 2223 6320 2224 6640
rect 2544 6320 2545 6640
rect 2223 6319 2545 6320
rect 1804 6252 1900 6268
rect 2816 6268 2832 6692
rect 2896 6268 2912 6692
rect 3828 6692 3924 6708
rect 3235 6640 3557 6641
rect 3235 6320 3236 6640
rect 3556 6320 3557 6640
rect 3235 6319 3557 6320
rect 2816 6252 2912 6268
rect 3828 6268 3844 6692
rect 3908 6268 3924 6692
rect 4840 6692 4936 6708
rect 4247 6640 4569 6641
rect 4247 6320 4248 6640
rect 4568 6320 4569 6640
rect 4247 6319 4569 6320
rect 3828 6252 3924 6268
rect 4840 6268 4856 6692
rect 4920 6268 4936 6692
rect 5852 6692 5948 6708
rect 5259 6640 5581 6641
rect 5259 6320 5260 6640
rect 5580 6320 5581 6640
rect 5259 6319 5581 6320
rect 4840 6252 4936 6268
rect 5852 6268 5868 6692
rect 5932 6268 5948 6692
rect 6864 6692 6960 6708
rect 6271 6640 6593 6641
rect 6271 6320 6272 6640
rect 6592 6320 6593 6640
rect 6271 6319 6593 6320
rect 5852 6252 5948 6268
rect 6864 6268 6880 6692
rect 6944 6268 6960 6692
rect 7876 6692 7972 6708
rect 7283 6640 7605 6641
rect 7283 6320 7284 6640
rect 7604 6320 7605 6640
rect 7283 6319 7605 6320
rect 6864 6252 6960 6268
rect 7876 6268 7892 6692
rect 7956 6268 7972 6692
rect 8888 6692 8984 6708
rect 8295 6640 8617 6641
rect 8295 6320 8296 6640
rect 8616 6320 8617 6640
rect 8295 6319 8617 6320
rect 7876 6252 7972 6268
rect 8888 6268 8904 6692
rect 8968 6268 8984 6692
rect 9900 6692 9996 6708
rect 9307 6640 9629 6641
rect 9307 6320 9308 6640
rect 9628 6320 9629 6640
rect 9307 6319 9629 6320
rect 8888 6252 8984 6268
rect 9900 6268 9916 6692
rect 9980 6268 9996 6692
rect 10912 6692 11008 6708
rect 10319 6640 10641 6641
rect 10319 6320 10320 6640
rect 10640 6320 10641 6640
rect 10319 6319 10641 6320
rect 9900 6252 9996 6268
rect 10912 6268 10928 6692
rect 10992 6268 11008 6692
rect 11924 6692 12020 6708
rect 11331 6640 11653 6641
rect 11331 6320 11332 6640
rect 11652 6320 11653 6640
rect 11331 6319 11653 6320
rect 10912 6252 11008 6268
rect 11924 6268 11940 6692
rect 12004 6268 12020 6692
rect 12936 6692 13032 6708
rect 12343 6640 12665 6641
rect 12343 6320 12344 6640
rect 12664 6320 12665 6640
rect 12343 6319 12665 6320
rect 11924 6252 12020 6268
rect 12936 6268 12952 6692
rect 13016 6268 13032 6692
rect 13948 6692 14044 6708
rect 13355 6640 13677 6641
rect 13355 6320 13356 6640
rect 13676 6320 13677 6640
rect 13355 6319 13677 6320
rect 12936 6252 13032 6268
rect 13948 6268 13964 6692
rect 14028 6268 14044 6692
rect 14960 6692 15056 6708
rect 14367 6640 14689 6641
rect 14367 6320 14368 6640
rect 14688 6320 14689 6640
rect 14367 6319 14689 6320
rect 13948 6252 14044 6268
rect 14960 6268 14976 6692
rect 15040 6268 15056 6692
rect 15972 6692 16068 6708
rect 15379 6640 15701 6641
rect 15379 6320 15380 6640
rect 15700 6320 15701 6640
rect 15379 6319 15701 6320
rect 14960 6252 15056 6268
rect 15972 6268 15988 6692
rect 16052 6268 16068 6692
rect 16984 6692 17080 6708
rect 16391 6640 16713 6641
rect 16391 6320 16392 6640
rect 16712 6320 16713 6640
rect 16391 6319 16713 6320
rect 15972 6252 16068 6268
rect 16984 6268 17000 6692
rect 17064 6268 17080 6692
rect 16984 6252 17080 6268
rect -16412 5972 -16316 5988
rect -17005 5920 -16683 5921
rect -17005 5600 -17004 5920
rect -16684 5600 -16683 5920
rect -17005 5599 -16683 5600
rect -16412 5548 -16396 5972
rect -16332 5548 -16316 5972
rect -15400 5972 -15304 5988
rect -15993 5920 -15671 5921
rect -15993 5600 -15992 5920
rect -15672 5600 -15671 5920
rect -15993 5599 -15671 5600
rect -16412 5532 -16316 5548
rect -15400 5548 -15384 5972
rect -15320 5548 -15304 5972
rect -14388 5972 -14292 5988
rect -14981 5920 -14659 5921
rect -14981 5600 -14980 5920
rect -14660 5600 -14659 5920
rect -14981 5599 -14659 5600
rect -15400 5532 -15304 5548
rect -14388 5548 -14372 5972
rect -14308 5548 -14292 5972
rect -13376 5972 -13280 5988
rect -13969 5920 -13647 5921
rect -13969 5600 -13968 5920
rect -13648 5600 -13647 5920
rect -13969 5599 -13647 5600
rect -14388 5532 -14292 5548
rect -13376 5548 -13360 5972
rect -13296 5548 -13280 5972
rect -12364 5972 -12268 5988
rect -12957 5920 -12635 5921
rect -12957 5600 -12956 5920
rect -12636 5600 -12635 5920
rect -12957 5599 -12635 5600
rect -13376 5532 -13280 5548
rect -12364 5548 -12348 5972
rect -12284 5548 -12268 5972
rect -11352 5972 -11256 5988
rect -11945 5920 -11623 5921
rect -11945 5600 -11944 5920
rect -11624 5600 -11623 5920
rect -11945 5599 -11623 5600
rect -12364 5532 -12268 5548
rect -11352 5548 -11336 5972
rect -11272 5548 -11256 5972
rect -10340 5972 -10244 5988
rect -10933 5920 -10611 5921
rect -10933 5600 -10932 5920
rect -10612 5600 -10611 5920
rect -10933 5599 -10611 5600
rect -11352 5532 -11256 5548
rect -10340 5548 -10324 5972
rect -10260 5548 -10244 5972
rect -9328 5972 -9232 5988
rect -9921 5920 -9599 5921
rect -9921 5600 -9920 5920
rect -9600 5600 -9599 5920
rect -9921 5599 -9599 5600
rect -10340 5532 -10244 5548
rect -9328 5548 -9312 5972
rect -9248 5548 -9232 5972
rect -8316 5972 -8220 5988
rect -8909 5920 -8587 5921
rect -8909 5600 -8908 5920
rect -8588 5600 -8587 5920
rect -8909 5599 -8587 5600
rect -9328 5532 -9232 5548
rect -8316 5548 -8300 5972
rect -8236 5548 -8220 5972
rect -7304 5972 -7208 5988
rect -7897 5920 -7575 5921
rect -7897 5600 -7896 5920
rect -7576 5600 -7575 5920
rect -7897 5599 -7575 5600
rect -8316 5532 -8220 5548
rect -7304 5548 -7288 5972
rect -7224 5548 -7208 5972
rect -6292 5972 -6196 5988
rect -6885 5920 -6563 5921
rect -6885 5600 -6884 5920
rect -6564 5600 -6563 5920
rect -6885 5599 -6563 5600
rect -7304 5532 -7208 5548
rect -6292 5548 -6276 5972
rect -6212 5548 -6196 5972
rect -5280 5972 -5184 5988
rect -5873 5920 -5551 5921
rect -5873 5600 -5872 5920
rect -5552 5600 -5551 5920
rect -5873 5599 -5551 5600
rect -6292 5532 -6196 5548
rect -5280 5548 -5264 5972
rect -5200 5548 -5184 5972
rect -4268 5972 -4172 5988
rect -4861 5920 -4539 5921
rect -4861 5600 -4860 5920
rect -4540 5600 -4539 5920
rect -4861 5599 -4539 5600
rect -5280 5532 -5184 5548
rect -4268 5548 -4252 5972
rect -4188 5548 -4172 5972
rect -3256 5972 -3160 5988
rect -3849 5920 -3527 5921
rect -3849 5600 -3848 5920
rect -3528 5600 -3527 5920
rect -3849 5599 -3527 5600
rect -4268 5532 -4172 5548
rect -3256 5548 -3240 5972
rect -3176 5548 -3160 5972
rect -2244 5972 -2148 5988
rect -2837 5920 -2515 5921
rect -2837 5600 -2836 5920
rect -2516 5600 -2515 5920
rect -2837 5599 -2515 5600
rect -3256 5532 -3160 5548
rect -2244 5548 -2228 5972
rect -2164 5548 -2148 5972
rect -1232 5972 -1136 5988
rect -1825 5920 -1503 5921
rect -1825 5600 -1824 5920
rect -1504 5600 -1503 5920
rect -1825 5599 -1503 5600
rect -2244 5532 -2148 5548
rect -1232 5548 -1216 5972
rect -1152 5548 -1136 5972
rect -220 5972 -124 5988
rect -813 5920 -491 5921
rect -813 5600 -812 5920
rect -492 5600 -491 5920
rect -813 5599 -491 5600
rect -1232 5532 -1136 5548
rect -220 5548 -204 5972
rect -140 5548 -124 5972
rect 792 5972 888 5988
rect 199 5920 521 5921
rect 199 5600 200 5920
rect 520 5600 521 5920
rect 199 5599 521 5600
rect -220 5532 -124 5548
rect 792 5548 808 5972
rect 872 5548 888 5972
rect 1804 5972 1900 5988
rect 1211 5920 1533 5921
rect 1211 5600 1212 5920
rect 1532 5600 1533 5920
rect 1211 5599 1533 5600
rect 792 5532 888 5548
rect 1804 5548 1820 5972
rect 1884 5548 1900 5972
rect 2816 5972 2912 5988
rect 2223 5920 2545 5921
rect 2223 5600 2224 5920
rect 2544 5600 2545 5920
rect 2223 5599 2545 5600
rect 1804 5532 1900 5548
rect 2816 5548 2832 5972
rect 2896 5548 2912 5972
rect 3828 5972 3924 5988
rect 3235 5920 3557 5921
rect 3235 5600 3236 5920
rect 3556 5600 3557 5920
rect 3235 5599 3557 5600
rect 2816 5532 2912 5548
rect 3828 5548 3844 5972
rect 3908 5548 3924 5972
rect 4840 5972 4936 5988
rect 4247 5920 4569 5921
rect 4247 5600 4248 5920
rect 4568 5600 4569 5920
rect 4247 5599 4569 5600
rect 3828 5532 3924 5548
rect 4840 5548 4856 5972
rect 4920 5548 4936 5972
rect 5852 5972 5948 5988
rect 5259 5920 5581 5921
rect 5259 5600 5260 5920
rect 5580 5600 5581 5920
rect 5259 5599 5581 5600
rect 4840 5532 4936 5548
rect 5852 5548 5868 5972
rect 5932 5548 5948 5972
rect 6864 5972 6960 5988
rect 6271 5920 6593 5921
rect 6271 5600 6272 5920
rect 6592 5600 6593 5920
rect 6271 5599 6593 5600
rect 5852 5532 5948 5548
rect 6864 5548 6880 5972
rect 6944 5548 6960 5972
rect 7876 5972 7972 5988
rect 7283 5920 7605 5921
rect 7283 5600 7284 5920
rect 7604 5600 7605 5920
rect 7283 5599 7605 5600
rect 6864 5532 6960 5548
rect 7876 5548 7892 5972
rect 7956 5548 7972 5972
rect 8888 5972 8984 5988
rect 8295 5920 8617 5921
rect 8295 5600 8296 5920
rect 8616 5600 8617 5920
rect 8295 5599 8617 5600
rect 7876 5532 7972 5548
rect 8888 5548 8904 5972
rect 8968 5548 8984 5972
rect 9900 5972 9996 5988
rect 9307 5920 9629 5921
rect 9307 5600 9308 5920
rect 9628 5600 9629 5920
rect 9307 5599 9629 5600
rect 8888 5532 8984 5548
rect 9900 5548 9916 5972
rect 9980 5548 9996 5972
rect 10912 5972 11008 5988
rect 10319 5920 10641 5921
rect 10319 5600 10320 5920
rect 10640 5600 10641 5920
rect 10319 5599 10641 5600
rect 9900 5532 9996 5548
rect 10912 5548 10928 5972
rect 10992 5548 11008 5972
rect 11924 5972 12020 5988
rect 11331 5920 11653 5921
rect 11331 5600 11332 5920
rect 11652 5600 11653 5920
rect 11331 5599 11653 5600
rect 10912 5532 11008 5548
rect 11924 5548 11940 5972
rect 12004 5548 12020 5972
rect 12936 5972 13032 5988
rect 12343 5920 12665 5921
rect 12343 5600 12344 5920
rect 12664 5600 12665 5920
rect 12343 5599 12665 5600
rect 11924 5532 12020 5548
rect 12936 5548 12952 5972
rect 13016 5548 13032 5972
rect 13948 5972 14044 5988
rect 13355 5920 13677 5921
rect 13355 5600 13356 5920
rect 13676 5600 13677 5920
rect 13355 5599 13677 5600
rect 12936 5532 13032 5548
rect 13948 5548 13964 5972
rect 14028 5548 14044 5972
rect 14960 5972 15056 5988
rect 14367 5920 14689 5921
rect 14367 5600 14368 5920
rect 14688 5600 14689 5920
rect 14367 5599 14689 5600
rect 13948 5532 14044 5548
rect 14960 5548 14976 5972
rect 15040 5548 15056 5972
rect 15972 5972 16068 5988
rect 15379 5920 15701 5921
rect 15379 5600 15380 5920
rect 15700 5600 15701 5920
rect 15379 5599 15701 5600
rect 14960 5532 15056 5548
rect 15972 5548 15988 5972
rect 16052 5548 16068 5972
rect 16984 5972 17080 5988
rect 16391 5920 16713 5921
rect 16391 5600 16392 5920
rect 16712 5600 16713 5920
rect 16391 5599 16713 5600
rect 15972 5532 16068 5548
rect 16984 5548 17000 5972
rect 17064 5548 17080 5972
rect 16984 5532 17080 5548
rect -16412 5252 -16316 5268
rect -17005 5200 -16683 5201
rect -17005 4880 -17004 5200
rect -16684 4880 -16683 5200
rect -17005 4879 -16683 4880
rect -16412 4828 -16396 5252
rect -16332 4828 -16316 5252
rect -15400 5252 -15304 5268
rect -15993 5200 -15671 5201
rect -15993 4880 -15992 5200
rect -15672 4880 -15671 5200
rect -15993 4879 -15671 4880
rect -16412 4812 -16316 4828
rect -15400 4828 -15384 5252
rect -15320 4828 -15304 5252
rect -14388 5252 -14292 5268
rect -14981 5200 -14659 5201
rect -14981 4880 -14980 5200
rect -14660 4880 -14659 5200
rect -14981 4879 -14659 4880
rect -15400 4812 -15304 4828
rect -14388 4828 -14372 5252
rect -14308 4828 -14292 5252
rect -13376 5252 -13280 5268
rect -13969 5200 -13647 5201
rect -13969 4880 -13968 5200
rect -13648 4880 -13647 5200
rect -13969 4879 -13647 4880
rect -14388 4812 -14292 4828
rect -13376 4828 -13360 5252
rect -13296 4828 -13280 5252
rect -12364 5252 -12268 5268
rect -12957 5200 -12635 5201
rect -12957 4880 -12956 5200
rect -12636 4880 -12635 5200
rect -12957 4879 -12635 4880
rect -13376 4812 -13280 4828
rect -12364 4828 -12348 5252
rect -12284 4828 -12268 5252
rect -11352 5252 -11256 5268
rect -11945 5200 -11623 5201
rect -11945 4880 -11944 5200
rect -11624 4880 -11623 5200
rect -11945 4879 -11623 4880
rect -12364 4812 -12268 4828
rect -11352 4828 -11336 5252
rect -11272 4828 -11256 5252
rect -10340 5252 -10244 5268
rect -10933 5200 -10611 5201
rect -10933 4880 -10932 5200
rect -10612 4880 -10611 5200
rect -10933 4879 -10611 4880
rect -11352 4812 -11256 4828
rect -10340 4828 -10324 5252
rect -10260 4828 -10244 5252
rect -9328 5252 -9232 5268
rect -9921 5200 -9599 5201
rect -9921 4880 -9920 5200
rect -9600 4880 -9599 5200
rect -9921 4879 -9599 4880
rect -10340 4812 -10244 4828
rect -9328 4828 -9312 5252
rect -9248 4828 -9232 5252
rect -8316 5252 -8220 5268
rect -8909 5200 -8587 5201
rect -8909 4880 -8908 5200
rect -8588 4880 -8587 5200
rect -8909 4879 -8587 4880
rect -9328 4812 -9232 4828
rect -8316 4828 -8300 5252
rect -8236 4828 -8220 5252
rect -7304 5252 -7208 5268
rect -7897 5200 -7575 5201
rect -7897 4880 -7896 5200
rect -7576 4880 -7575 5200
rect -7897 4879 -7575 4880
rect -8316 4812 -8220 4828
rect -7304 4828 -7288 5252
rect -7224 4828 -7208 5252
rect -6292 5252 -6196 5268
rect -6885 5200 -6563 5201
rect -6885 4880 -6884 5200
rect -6564 4880 -6563 5200
rect -6885 4879 -6563 4880
rect -7304 4812 -7208 4828
rect -6292 4828 -6276 5252
rect -6212 4828 -6196 5252
rect -5280 5252 -5184 5268
rect -5873 5200 -5551 5201
rect -5873 4880 -5872 5200
rect -5552 4880 -5551 5200
rect -5873 4879 -5551 4880
rect -6292 4812 -6196 4828
rect -5280 4828 -5264 5252
rect -5200 4828 -5184 5252
rect -4268 5252 -4172 5268
rect -4861 5200 -4539 5201
rect -4861 4880 -4860 5200
rect -4540 4880 -4539 5200
rect -4861 4879 -4539 4880
rect -5280 4812 -5184 4828
rect -4268 4828 -4252 5252
rect -4188 4828 -4172 5252
rect -3256 5252 -3160 5268
rect -3849 5200 -3527 5201
rect -3849 4880 -3848 5200
rect -3528 4880 -3527 5200
rect -3849 4879 -3527 4880
rect -4268 4812 -4172 4828
rect -3256 4828 -3240 5252
rect -3176 4828 -3160 5252
rect -2244 5252 -2148 5268
rect -2837 5200 -2515 5201
rect -2837 4880 -2836 5200
rect -2516 4880 -2515 5200
rect -2837 4879 -2515 4880
rect -3256 4812 -3160 4828
rect -2244 4828 -2228 5252
rect -2164 4828 -2148 5252
rect -1232 5252 -1136 5268
rect -1825 5200 -1503 5201
rect -1825 4880 -1824 5200
rect -1504 4880 -1503 5200
rect -1825 4879 -1503 4880
rect -2244 4812 -2148 4828
rect -1232 4828 -1216 5252
rect -1152 4828 -1136 5252
rect -220 5252 -124 5268
rect -813 5200 -491 5201
rect -813 4880 -812 5200
rect -492 4880 -491 5200
rect -813 4879 -491 4880
rect -1232 4812 -1136 4828
rect -220 4828 -204 5252
rect -140 4828 -124 5252
rect 792 5252 888 5268
rect 199 5200 521 5201
rect 199 4880 200 5200
rect 520 4880 521 5200
rect 199 4879 521 4880
rect -220 4812 -124 4828
rect 792 4828 808 5252
rect 872 4828 888 5252
rect 1804 5252 1900 5268
rect 1211 5200 1533 5201
rect 1211 4880 1212 5200
rect 1532 4880 1533 5200
rect 1211 4879 1533 4880
rect 792 4812 888 4828
rect 1804 4828 1820 5252
rect 1884 4828 1900 5252
rect 2816 5252 2912 5268
rect 2223 5200 2545 5201
rect 2223 4880 2224 5200
rect 2544 4880 2545 5200
rect 2223 4879 2545 4880
rect 1804 4812 1900 4828
rect 2816 4828 2832 5252
rect 2896 4828 2912 5252
rect 3828 5252 3924 5268
rect 3235 5200 3557 5201
rect 3235 4880 3236 5200
rect 3556 4880 3557 5200
rect 3235 4879 3557 4880
rect 2816 4812 2912 4828
rect 3828 4828 3844 5252
rect 3908 4828 3924 5252
rect 4840 5252 4936 5268
rect 4247 5200 4569 5201
rect 4247 4880 4248 5200
rect 4568 4880 4569 5200
rect 4247 4879 4569 4880
rect 3828 4812 3924 4828
rect 4840 4828 4856 5252
rect 4920 4828 4936 5252
rect 5852 5252 5948 5268
rect 5259 5200 5581 5201
rect 5259 4880 5260 5200
rect 5580 4880 5581 5200
rect 5259 4879 5581 4880
rect 4840 4812 4936 4828
rect 5852 4828 5868 5252
rect 5932 4828 5948 5252
rect 6864 5252 6960 5268
rect 6271 5200 6593 5201
rect 6271 4880 6272 5200
rect 6592 4880 6593 5200
rect 6271 4879 6593 4880
rect 5852 4812 5948 4828
rect 6864 4828 6880 5252
rect 6944 4828 6960 5252
rect 7876 5252 7972 5268
rect 7283 5200 7605 5201
rect 7283 4880 7284 5200
rect 7604 4880 7605 5200
rect 7283 4879 7605 4880
rect 6864 4812 6960 4828
rect 7876 4828 7892 5252
rect 7956 4828 7972 5252
rect 8888 5252 8984 5268
rect 8295 5200 8617 5201
rect 8295 4880 8296 5200
rect 8616 4880 8617 5200
rect 8295 4879 8617 4880
rect 7876 4812 7972 4828
rect 8888 4828 8904 5252
rect 8968 4828 8984 5252
rect 9900 5252 9996 5268
rect 9307 5200 9629 5201
rect 9307 4880 9308 5200
rect 9628 4880 9629 5200
rect 9307 4879 9629 4880
rect 8888 4812 8984 4828
rect 9900 4828 9916 5252
rect 9980 4828 9996 5252
rect 10912 5252 11008 5268
rect 10319 5200 10641 5201
rect 10319 4880 10320 5200
rect 10640 4880 10641 5200
rect 10319 4879 10641 4880
rect 9900 4812 9996 4828
rect 10912 4828 10928 5252
rect 10992 4828 11008 5252
rect 11924 5252 12020 5268
rect 11331 5200 11653 5201
rect 11331 4880 11332 5200
rect 11652 4880 11653 5200
rect 11331 4879 11653 4880
rect 10912 4812 11008 4828
rect 11924 4828 11940 5252
rect 12004 4828 12020 5252
rect 12936 5252 13032 5268
rect 12343 5200 12665 5201
rect 12343 4880 12344 5200
rect 12664 4880 12665 5200
rect 12343 4879 12665 4880
rect 11924 4812 12020 4828
rect 12936 4828 12952 5252
rect 13016 4828 13032 5252
rect 13948 5252 14044 5268
rect 13355 5200 13677 5201
rect 13355 4880 13356 5200
rect 13676 4880 13677 5200
rect 13355 4879 13677 4880
rect 12936 4812 13032 4828
rect 13948 4828 13964 5252
rect 14028 4828 14044 5252
rect 14960 5252 15056 5268
rect 14367 5200 14689 5201
rect 14367 4880 14368 5200
rect 14688 4880 14689 5200
rect 14367 4879 14689 4880
rect 13948 4812 14044 4828
rect 14960 4828 14976 5252
rect 15040 4828 15056 5252
rect 15972 5252 16068 5268
rect 15379 5200 15701 5201
rect 15379 4880 15380 5200
rect 15700 4880 15701 5200
rect 15379 4879 15701 4880
rect 14960 4812 15056 4828
rect 15972 4828 15988 5252
rect 16052 4828 16068 5252
rect 16984 5252 17080 5268
rect 16391 5200 16713 5201
rect 16391 4880 16392 5200
rect 16712 4880 16713 5200
rect 16391 4879 16713 4880
rect 15972 4812 16068 4828
rect 16984 4828 17000 5252
rect 17064 4828 17080 5252
rect 16984 4812 17080 4828
rect -16412 4532 -16316 4548
rect -17005 4480 -16683 4481
rect -17005 4160 -17004 4480
rect -16684 4160 -16683 4480
rect -17005 4159 -16683 4160
rect -16412 4108 -16396 4532
rect -16332 4108 -16316 4532
rect -15400 4532 -15304 4548
rect -15993 4480 -15671 4481
rect -15993 4160 -15992 4480
rect -15672 4160 -15671 4480
rect -15993 4159 -15671 4160
rect -16412 4092 -16316 4108
rect -15400 4108 -15384 4532
rect -15320 4108 -15304 4532
rect -14388 4532 -14292 4548
rect -14981 4480 -14659 4481
rect -14981 4160 -14980 4480
rect -14660 4160 -14659 4480
rect -14981 4159 -14659 4160
rect -15400 4092 -15304 4108
rect -14388 4108 -14372 4532
rect -14308 4108 -14292 4532
rect -13376 4532 -13280 4548
rect -13969 4480 -13647 4481
rect -13969 4160 -13968 4480
rect -13648 4160 -13647 4480
rect -13969 4159 -13647 4160
rect -14388 4092 -14292 4108
rect -13376 4108 -13360 4532
rect -13296 4108 -13280 4532
rect -12364 4532 -12268 4548
rect -12957 4480 -12635 4481
rect -12957 4160 -12956 4480
rect -12636 4160 -12635 4480
rect -12957 4159 -12635 4160
rect -13376 4092 -13280 4108
rect -12364 4108 -12348 4532
rect -12284 4108 -12268 4532
rect -11352 4532 -11256 4548
rect -11945 4480 -11623 4481
rect -11945 4160 -11944 4480
rect -11624 4160 -11623 4480
rect -11945 4159 -11623 4160
rect -12364 4092 -12268 4108
rect -11352 4108 -11336 4532
rect -11272 4108 -11256 4532
rect -10340 4532 -10244 4548
rect -10933 4480 -10611 4481
rect -10933 4160 -10932 4480
rect -10612 4160 -10611 4480
rect -10933 4159 -10611 4160
rect -11352 4092 -11256 4108
rect -10340 4108 -10324 4532
rect -10260 4108 -10244 4532
rect -9328 4532 -9232 4548
rect -9921 4480 -9599 4481
rect -9921 4160 -9920 4480
rect -9600 4160 -9599 4480
rect -9921 4159 -9599 4160
rect -10340 4092 -10244 4108
rect -9328 4108 -9312 4532
rect -9248 4108 -9232 4532
rect -8316 4532 -8220 4548
rect -8909 4480 -8587 4481
rect -8909 4160 -8908 4480
rect -8588 4160 -8587 4480
rect -8909 4159 -8587 4160
rect -9328 4092 -9232 4108
rect -8316 4108 -8300 4532
rect -8236 4108 -8220 4532
rect -7304 4532 -7208 4548
rect -7897 4480 -7575 4481
rect -7897 4160 -7896 4480
rect -7576 4160 -7575 4480
rect -7897 4159 -7575 4160
rect -8316 4092 -8220 4108
rect -7304 4108 -7288 4532
rect -7224 4108 -7208 4532
rect -6292 4532 -6196 4548
rect -6885 4480 -6563 4481
rect -6885 4160 -6884 4480
rect -6564 4160 -6563 4480
rect -6885 4159 -6563 4160
rect -7304 4092 -7208 4108
rect -6292 4108 -6276 4532
rect -6212 4108 -6196 4532
rect -5280 4532 -5184 4548
rect -5873 4480 -5551 4481
rect -5873 4160 -5872 4480
rect -5552 4160 -5551 4480
rect -5873 4159 -5551 4160
rect -6292 4092 -6196 4108
rect -5280 4108 -5264 4532
rect -5200 4108 -5184 4532
rect -4268 4532 -4172 4548
rect -4861 4480 -4539 4481
rect -4861 4160 -4860 4480
rect -4540 4160 -4539 4480
rect -4861 4159 -4539 4160
rect -5280 4092 -5184 4108
rect -4268 4108 -4252 4532
rect -4188 4108 -4172 4532
rect -3256 4532 -3160 4548
rect -3849 4480 -3527 4481
rect -3849 4160 -3848 4480
rect -3528 4160 -3527 4480
rect -3849 4159 -3527 4160
rect -4268 4092 -4172 4108
rect -3256 4108 -3240 4532
rect -3176 4108 -3160 4532
rect -2244 4532 -2148 4548
rect -2837 4480 -2515 4481
rect -2837 4160 -2836 4480
rect -2516 4160 -2515 4480
rect -2837 4159 -2515 4160
rect -3256 4092 -3160 4108
rect -2244 4108 -2228 4532
rect -2164 4108 -2148 4532
rect -1232 4532 -1136 4548
rect -1825 4480 -1503 4481
rect -1825 4160 -1824 4480
rect -1504 4160 -1503 4480
rect -1825 4159 -1503 4160
rect -2244 4092 -2148 4108
rect -1232 4108 -1216 4532
rect -1152 4108 -1136 4532
rect -220 4532 -124 4548
rect -813 4480 -491 4481
rect -813 4160 -812 4480
rect -492 4160 -491 4480
rect -813 4159 -491 4160
rect -1232 4092 -1136 4108
rect -220 4108 -204 4532
rect -140 4108 -124 4532
rect 792 4532 888 4548
rect 199 4480 521 4481
rect 199 4160 200 4480
rect 520 4160 521 4480
rect 199 4159 521 4160
rect -220 4092 -124 4108
rect 792 4108 808 4532
rect 872 4108 888 4532
rect 1804 4532 1900 4548
rect 1211 4480 1533 4481
rect 1211 4160 1212 4480
rect 1532 4160 1533 4480
rect 1211 4159 1533 4160
rect 792 4092 888 4108
rect 1804 4108 1820 4532
rect 1884 4108 1900 4532
rect 2816 4532 2912 4548
rect 2223 4480 2545 4481
rect 2223 4160 2224 4480
rect 2544 4160 2545 4480
rect 2223 4159 2545 4160
rect 1804 4092 1900 4108
rect 2816 4108 2832 4532
rect 2896 4108 2912 4532
rect 3828 4532 3924 4548
rect 3235 4480 3557 4481
rect 3235 4160 3236 4480
rect 3556 4160 3557 4480
rect 3235 4159 3557 4160
rect 2816 4092 2912 4108
rect 3828 4108 3844 4532
rect 3908 4108 3924 4532
rect 4840 4532 4936 4548
rect 4247 4480 4569 4481
rect 4247 4160 4248 4480
rect 4568 4160 4569 4480
rect 4247 4159 4569 4160
rect 3828 4092 3924 4108
rect 4840 4108 4856 4532
rect 4920 4108 4936 4532
rect 5852 4532 5948 4548
rect 5259 4480 5581 4481
rect 5259 4160 5260 4480
rect 5580 4160 5581 4480
rect 5259 4159 5581 4160
rect 4840 4092 4936 4108
rect 5852 4108 5868 4532
rect 5932 4108 5948 4532
rect 6864 4532 6960 4548
rect 6271 4480 6593 4481
rect 6271 4160 6272 4480
rect 6592 4160 6593 4480
rect 6271 4159 6593 4160
rect 5852 4092 5948 4108
rect 6864 4108 6880 4532
rect 6944 4108 6960 4532
rect 7876 4532 7972 4548
rect 7283 4480 7605 4481
rect 7283 4160 7284 4480
rect 7604 4160 7605 4480
rect 7283 4159 7605 4160
rect 6864 4092 6960 4108
rect 7876 4108 7892 4532
rect 7956 4108 7972 4532
rect 8888 4532 8984 4548
rect 8295 4480 8617 4481
rect 8295 4160 8296 4480
rect 8616 4160 8617 4480
rect 8295 4159 8617 4160
rect 7876 4092 7972 4108
rect 8888 4108 8904 4532
rect 8968 4108 8984 4532
rect 9900 4532 9996 4548
rect 9307 4480 9629 4481
rect 9307 4160 9308 4480
rect 9628 4160 9629 4480
rect 9307 4159 9629 4160
rect 8888 4092 8984 4108
rect 9900 4108 9916 4532
rect 9980 4108 9996 4532
rect 10912 4532 11008 4548
rect 10319 4480 10641 4481
rect 10319 4160 10320 4480
rect 10640 4160 10641 4480
rect 10319 4159 10641 4160
rect 9900 4092 9996 4108
rect 10912 4108 10928 4532
rect 10992 4108 11008 4532
rect 11924 4532 12020 4548
rect 11331 4480 11653 4481
rect 11331 4160 11332 4480
rect 11652 4160 11653 4480
rect 11331 4159 11653 4160
rect 10912 4092 11008 4108
rect 11924 4108 11940 4532
rect 12004 4108 12020 4532
rect 12936 4532 13032 4548
rect 12343 4480 12665 4481
rect 12343 4160 12344 4480
rect 12664 4160 12665 4480
rect 12343 4159 12665 4160
rect 11924 4092 12020 4108
rect 12936 4108 12952 4532
rect 13016 4108 13032 4532
rect 13948 4532 14044 4548
rect 13355 4480 13677 4481
rect 13355 4160 13356 4480
rect 13676 4160 13677 4480
rect 13355 4159 13677 4160
rect 12936 4092 13032 4108
rect 13948 4108 13964 4532
rect 14028 4108 14044 4532
rect 14960 4532 15056 4548
rect 14367 4480 14689 4481
rect 14367 4160 14368 4480
rect 14688 4160 14689 4480
rect 14367 4159 14689 4160
rect 13948 4092 14044 4108
rect 14960 4108 14976 4532
rect 15040 4108 15056 4532
rect 15972 4532 16068 4548
rect 15379 4480 15701 4481
rect 15379 4160 15380 4480
rect 15700 4160 15701 4480
rect 15379 4159 15701 4160
rect 14960 4092 15056 4108
rect 15972 4108 15988 4532
rect 16052 4108 16068 4532
rect 16984 4532 17080 4548
rect 16391 4480 16713 4481
rect 16391 4160 16392 4480
rect 16712 4160 16713 4480
rect 16391 4159 16713 4160
rect 15972 4092 16068 4108
rect 16984 4108 17000 4532
rect 17064 4108 17080 4532
rect 16984 4092 17080 4108
rect -16412 3812 -16316 3828
rect -17005 3760 -16683 3761
rect -17005 3440 -17004 3760
rect -16684 3440 -16683 3760
rect -17005 3439 -16683 3440
rect -16412 3388 -16396 3812
rect -16332 3388 -16316 3812
rect -15400 3812 -15304 3828
rect -15993 3760 -15671 3761
rect -15993 3440 -15992 3760
rect -15672 3440 -15671 3760
rect -15993 3439 -15671 3440
rect -16412 3372 -16316 3388
rect -15400 3388 -15384 3812
rect -15320 3388 -15304 3812
rect -14388 3812 -14292 3828
rect -14981 3760 -14659 3761
rect -14981 3440 -14980 3760
rect -14660 3440 -14659 3760
rect -14981 3439 -14659 3440
rect -15400 3372 -15304 3388
rect -14388 3388 -14372 3812
rect -14308 3388 -14292 3812
rect -13376 3812 -13280 3828
rect -13969 3760 -13647 3761
rect -13969 3440 -13968 3760
rect -13648 3440 -13647 3760
rect -13969 3439 -13647 3440
rect -14388 3372 -14292 3388
rect -13376 3388 -13360 3812
rect -13296 3388 -13280 3812
rect -12364 3812 -12268 3828
rect -12957 3760 -12635 3761
rect -12957 3440 -12956 3760
rect -12636 3440 -12635 3760
rect -12957 3439 -12635 3440
rect -13376 3372 -13280 3388
rect -12364 3388 -12348 3812
rect -12284 3388 -12268 3812
rect -11352 3812 -11256 3828
rect -11945 3760 -11623 3761
rect -11945 3440 -11944 3760
rect -11624 3440 -11623 3760
rect -11945 3439 -11623 3440
rect -12364 3372 -12268 3388
rect -11352 3388 -11336 3812
rect -11272 3388 -11256 3812
rect -10340 3812 -10244 3828
rect -10933 3760 -10611 3761
rect -10933 3440 -10932 3760
rect -10612 3440 -10611 3760
rect -10933 3439 -10611 3440
rect -11352 3372 -11256 3388
rect -10340 3388 -10324 3812
rect -10260 3388 -10244 3812
rect -9328 3812 -9232 3828
rect -9921 3760 -9599 3761
rect -9921 3440 -9920 3760
rect -9600 3440 -9599 3760
rect -9921 3439 -9599 3440
rect -10340 3372 -10244 3388
rect -9328 3388 -9312 3812
rect -9248 3388 -9232 3812
rect -8316 3812 -8220 3828
rect -8909 3760 -8587 3761
rect -8909 3440 -8908 3760
rect -8588 3440 -8587 3760
rect -8909 3439 -8587 3440
rect -9328 3372 -9232 3388
rect -8316 3388 -8300 3812
rect -8236 3388 -8220 3812
rect -7304 3812 -7208 3828
rect -7897 3760 -7575 3761
rect -7897 3440 -7896 3760
rect -7576 3440 -7575 3760
rect -7897 3439 -7575 3440
rect -8316 3372 -8220 3388
rect -7304 3388 -7288 3812
rect -7224 3388 -7208 3812
rect -6292 3812 -6196 3828
rect -6885 3760 -6563 3761
rect -6885 3440 -6884 3760
rect -6564 3440 -6563 3760
rect -6885 3439 -6563 3440
rect -7304 3372 -7208 3388
rect -6292 3388 -6276 3812
rect -6212 3388 -6196 3812
rect -5280 3812 -5184 3828
rect -5873 3760 -5551 3761
rect -5873 3440 -5872 3760
rect -5552 3440 -5551 3760
rect -5873 3439 -5551 3440
rect -6292 3372 -6196 3388
rect -5280 3388 -5264 3812
rect -5200 3388 -5184 3812
rect -4268 3812 -4172 3828
rect -4861 3760 -4539 3761
rect -4861 3440 -4860 3760
rect -4540 3440 -4539 3760
rect -4861 3439 -4539 3440
rect -5280 3372 -5184 3388
rect -4268 3388 -4252 3812
rect -4188 3388 -4172 3812
rect -3256 3812 -3160 3828
rect -3849 3760 -3527 3761
rect -3849 3440 -3848 3760
rect -3528 3440 -3527 3760
rect -3849 3439 -3527 3440
rect -4268 3372 -4172 3388
rect -3256 3388 -3240 3812
rect -3176 3388 -3160 3812
rect -2244 3812 -2148 3828
rect -2837 3760 -2515 3761
rect -2837 3440 -2836 3760
rect -2516 3440 -2515 3760
rect -2837 3439 -2515 3440
rect -3256 3372 -3160 3388
rect -2244 3388 -2228 3812
rect -2164 3388 -2148 3812
rect -1232 3812 -1136 3828
rect -1825 3760 -1503 3761
rect -1825 3440 -1824 3760
rect -1504 3440 -1503 3760
rect -1825 3439 -1503 3440
rect -2244 3372 -2148 3388
rect -1232 3388 -1216 3812
rect -1152 3388 -1136 3812
rect -220 3812 -124 3828
rect -813 3760 -491 3761
rect -813 3440 -812 3760
rect -492 3440 -491 3760
rect -813 3439 -491 3440
rect -1232 3372 -1136 3388
rect -220 3388 -204 3812
rect -140 3388 -124 3812
rect 792 3812 888 3828
rect 199 3760 521 3761
rect 199 3440 200 3760
rect 520 3440 521 3760
rect 199 3439 521 3440
rect -220 3372 -124 3388
rect 792 3388 808 3812
rect 872 3388 888 3812
rect 1804 3812 1900 3828
rect 1211 3760 1533 3761
rect 1211 3440 1212 3760
rect 1532 3440 1533 3760
rect 1211 3439 1533 3440
rect 792 3372 888 3388
rect 1804 3388 1820 3812
rect 1884 3388 1900 3812
rect 2816 3812 2912 3828
rect 2223 3760 2545 3761
rect 2223 3440 2224 3760
rect 2544 3440 2545 3760
rect 2223 3439 2545 3440
rect 1804 3372 1900 3388
rect 2816 3388 2832 3812
rect 2896 3388 2912 3812
rect 3828 3812 3924 3828
rect 3235 3760 3557 3761
rect 3235 3440 3236 3760
rect 3556 3440 3557 3760
rect 3235 3439 3557 3440
rect 2816 3372 2912 3388
rect 3828 3388 3844 3812
rect 3908 3388 3924 3812
rect 4840 3812 4936 3828
rect 4247 3760 4569 3761
rect 4247 3440 4248 3760
rect 4568 3440 4569 3760
rect 4247 3439 4569 3440
rect 3828 3372 3924 3388
rect 4840 3388 4856 3812
rect 4920 3388 4936 3812
rect 5852 3812 5948 3828
rect 5259 3760 5581 3761
rect 5259 3440 5260 3760
rect 5580 3440 5581 3760
rect 5259 3439 5581 3440
rect 4840 3372 4936 3388
rect 5852 3388 5868 3812
rect 5932 3388 5948 3812
rect 6864 3812 6960 3828
rect 6271 3760 6593 3761
rect 6271 3440 6272 3760
rect 6592 3440 6593 3760
rect 6271 3439 6593 3440
rect 5852 3372 5948 3388
rect 6864 3388 6880 3812
rect 6944 3388 6960 3812
rect 7876 3812 7972 3828
rect 7283 3760 7605 3761
rect 7283 3440 7284 3760
rect 7604 3440 7605 3760
rect 7283 3439 7605 3440
rect 6864 3372 6960 3388
rect 7876 3388 7892 3812
rect 7956 3388 7972 3812
rect 8888 3812 8984 3828
rect 8295 3760 8617 3761
rect 8295 3440 8296 3760
rect 8616 3440 8617 3760
rect 8295 3439 8617 3440
rect 7876 3372 7972 3388
rect 8888 3388 8904 3812
rect 8968 3388 8984 3812
rect 9900 3812 9996 3828
rect 9307 3760 9629 3761
rect 9307 3440 9308 3760
rect 9628 3440 9629 3760
rect 9307 3439 9629 3440
rect 8888 3372 8984 3388
rect 9900 3388 9916 3812
rect 9980 3388 9996 3812
rect 10912 3812 11008 3828
rect 10319 3760 10641 3761
rect 10319 3440 10320 3760
rect 10640 3440 10641 3760
rect 10319 3439 10641 3440
rect 9900 3372 9996 3388
rect 10912 3388 10928 3812
rect 10992 3388 11008 3812
rect 11924 3812 12020 3828
rect 11331 3760 11653 3761
rect 11331 3440 11332 3760
rect 11652 3440 11653 3760
rect 11331 3439 11653 3440
rect 10912 3372 11008 3388
rect 11924 3388 11940 3812
rect 12004 3388 12020 3812
rect 12936 3812 13032 3828
rect 12343 3760 12665 3761
rect 12343 3440 12344 3760
rect 12664 3440 12665 3760
rect 12343 3439 12665 3440
rect 11924 3372 12020 3388
rect 12936 3388 12952 3812
rect 13016 3388 13032 3812
rect 13948 3812 14044 3828
rect 13355 3760 13677 3761
rect 13355 3440 13356 3760
rect 13676 3440 13677 3760
rect 13355 3439 13677 3440
rect 12936 3372 13032 3388
rect 13948 3388 13964 3812
rect 14028 3388 14044 3812
rect 14960 3812 15056 3828
rect 14367 3760 14689 3761
rect 14367 3440 14368 3760
rect 14688 3440 14689 3760
rect 14367 3439 14689 3440
rect 13948 3372 14044 3388
rect 14960 3388 14976 3812
rect 15040 3388 15056 3812
rect 15972 3812 16068 3828
rect 15379 3760 15701 3761
rect 15379 3440 15380 3760
rect 15700 3440 15701 3760
rect 15379 3439 15701 3440
rect 14960 3372 15056 3388
rect 15972 3388 15988 3812
rect 16052 3388 16068 3812
rect 16984 3812 17080 3828
rect 16391 3760 16713 3761
rect 16391 3440 16392 3760
rect 16712 3440 16713 3760
rect 16391 3439 16713 3440
rect 15972 3372 16068 3388
rect 16984 3388 17000 3812
rect 17064 3388 17080 3812
rect 16984 3372 17080 3388
rect -16412 3092 -16316 3108
rect -17005 3040 -16683 3041
rect -17005 2720 -17004 3040
rect -16684 2720 -16683 3040
rect -17005 2719 -16683 2720
rect -16412 2668 -16396 3092
rect -16332 2668 -16316 3092
rect -15400 3092 -15304 3108
rect -15993 3040 -15671 3041
rect -15993 2720 -15992 3040
rect -15672 2720 -15671 3040
rect -15993 2719 -15671 2720
rect -16412 2652 -16316 2668
rect -15400 2668 -15384 3092
rect -15320 2668 -15304 3092
rect -14388 3092 -14292 3108
rect -14981 3040 -14659 3041
rect -14981 2720 -14980 3040
rect -14660 2720 -14659 3040
rect -14981 2719 -14659 2720
rect -15400 2652 -15304 2668
rect -14388 2668 -14372 3092
rect -14308 2668 -14292 3092
rect -13376 3092 -13280 3108
rect -13969 3040 -13647 3041
rect -13969 2720 -13968 3040
rect -13648 2720 -13647 3040
rect -13969 2719 -13647 2720
rect -14388 2652 -14292 2668
rect -13376 2668 -13360 3092
rect -13296 2668 -13280 3092
rect -12364 3092 -12268 3108
rect -12957 3040 -12635 3041
rect -12957 2720 -12956 3040
rect -12636 2720 -12635 3040
rect -12957 2719 -12635 2720
rect -13376 2652 -13280 2668
rect -12364 2668 -12348 3092
rect -12284 2668 -12268 3092
rect -11352 3092 -11256 3108
rect -11945 3040 -11623 3041
rect -11945 2720 -11944 3040
rect -11624 2720 -11623 3040
rect -11945 2719 -11623 2720
rect -12364 2652 -12268 2668
rect -11352 2668 -11336 3092
rect -11272 2668 -11256 3092
rect -10340 3092 -10244 3108
rect -10933 3040 -10611 3041
rect -10933 2720 -10932 3040
rect -10612 2720 -10611 3040
rect -10933 2719 -10611 2720
rect -11352 2652 -11256 2668
rect -10340 2668 -10324 3092
rect -10260 2668 -10244 3092
rect -9328 3092 -9232 3108
rect -9921 3040 -9599 3041
rect -9921 2720 -9920 3040
rect -9600 2720 -9599 3040
rect -9921 2719 -9599 2720
rect -10340 2652 -10244 2668
rect -9328 2668 -9312 3092
rect -9248 2668 -9232 3092
rect -8316 3092 -8220 3108
rect -8909 3040 -8587 3041
rect -8909 2720 -8908 3040
rect -8588 2720 -8587 3040
rect -8909 2719 -8587 2720
rect -9328 2652 -9232 2668
rect -8316 2668 -8300 3092
rect -8236 2668 -8220 3092
rect -7304 3092 -7208 3108
rect -7897 3040 -7575 3041
rect -7897 2720 -7896 3040
rect -7576 2720 -7575 3040
rect -7897 2719 -7575 2720
rect -8316 2652 -8220 2668
rect -7304 2668 -7288 3092
rect -7224 2668 -7208 3092
rect -6292 3092 -6196 3108
rect -6885 3040 -6563 3041
rect -6885 2720 -6884 3040
rect -6564 2720 -6563 3040
rect -6885 2719 -6563 2720
rect -7304 2652 -7208 2668
rect -6292 2668 -6276 3092
rect -6212 2668 -6196 3092
rect -5280 3092 -5184 3108
rect -5873 3040 -5551 3041
rect -5873 2720 -5872 3040
rect -5552 2720 -5551 3040
rect -5873 2719 -5551 2720
rect -6292 2652 -6196 2668
rect -5280 2668 -5264 3092
rect -5200 2668 -5184 3092
rect -4268 3092 -4172 3108
rect -4861 3040 -4539 3041
rect -4861 2720 -4860 3040
rect -4540 2720 -4539 3040
rect -4861 2719 -4539 2720
rect -5280 2652 -5184 2668
rect -4268 2668 -4252 3092
rect -4188 2668 -4172 3092
rect -3256 3092 -3160 3108
rect -3849 3040 -3527 3041
rect -3849 2720 -3848 3040
rect -3528 2720 -3527 3040
rect -3849 2719 -3527 2720
rect -4268 2652 -4172 2668
rect -3256 2668 -3240 3092
rect -3176 2668 -3160 3092
rect -2244 3092 -2148 3108
rect -2837 3040 -2515 3041
rect -2837 2720 -2836 3040
rect -2516 2720 -2515 3040
rect -2837 2719 -2515 2720
rect -3256 2652 -3160 2668
rect -2244 2668 -2228 3092
rect -2164 2668 -2148 3092
rect -1232 3092 -1136 3108
rect -1825 3040 -1503 3041
rect -1825 2720 -1824 3040
rect -1504 2720 -1503 3040
rect -1825 2719 -1503 2720
rect -2244 2652 -2148 2668
rect -1232 2668 -1216 3092
rect -1152 2668 -1136 3092
rect -220 3092 -124 3108
rect -813 3040 -491 3041
rect -813 2720 -812 3040
rect -492 2720 -491 3040
rect -813 2719 -491 2720
rect -1232 2652 -1136 2668
rect -220 2668 -204 3092
rect -140 2668 -124 3092
rect 792 3092 888 3108
rect 199 3040 521 3041
rect 199 2720 200 3040
rect 520 2720 521 3040
rect 199 2719 521 2720
rect -220 2652 -124 2668
rect 792 2668 808 3092
rect 872 2668 888 3092
rect 1804 3092 1900 3108
rect 1211 3040 1533 3041
rect 1211 2720 1212 3040
rect 1532 2720 1533 3040
rect 1211 2719 1533 2720
rect 792 2652 888 2668
rect 1804 2668 1820 3092
rect 1884 2668 1900 3092
rect 2816 3092 2912 3108
rect 2223 3040 2545 3041
rect 2223 2720 2224 3040
rect 2544 2720 2545 3040
rect 2223 2719 2545 2720
rect 1804 2652 1900 2668
rect 2816 2668 2832 3092
rect 2896 2668 2912 3092
rect 3828 3092 3924 3108
rect 3235 3040 3557 3041
rect 3235 2720 3236 3040
rect 3556 2720 3557 3040
rect 3235 2719 3557 2720
rect 2816 2652 2912 2668
rect 3828 2668 3844 3092
rect 3908 2668 3924 3092
rect 4840 3092 4936 3108
rect 4247 3040 4569 3041
rect 4247 2720 4248 3040
rect 4568 2720 4569 3040
rect 4247 2719 4569 2720
rect 3828 2652 3924 2668
rect 4840 2668 4856 3092
rect 4920 2668 4936 3092
rect 5852 3092 5948 3108
rect 5259 3040 5581 3041
rect 5259 2720 5260 3040
rect 5580 2720 5581 3040
rect 5259 2719 5581 2720
rect 4840 2652 4936 2668
rect 5852 2668 5868 3092
rect 5932 2668 5948 3092
rect 6864 3092 6960 3108
rect 6271 3040 6593 3041
rect 6271 2720 6272 3040
rect 6592 2720 6593 3040
rect 6271 2719 6593 2720
rect 5852 2652 5948 2668
rect 6864 2668 6880 3092
rect 6944 2668 6960 3092
rect 7876 3092 7972 3108
rect 7283 3040 7605 3041
rect 7283 2720 7284 3040
rect 7604 2720 7605 3040
rect 7283 2719 7605 2720
rect 6864 2652 6960 2668
rect 7876 2668 7892 3092
rect 7956 2668 7972 3092
rect 8888 3092 8984 3108
rect 8295 3040 8617 3041
rect 8295 2720 8296 3040
rect 8616 2720 8617 3040
rect 8295 2719 8617 2720
rect 7876 2652 7972 2668
rect 8888 2668 8904 3092
rect 8968 2668 8984 3092
rect 9900 3092 9996 3108
rect 9307 3040 9629 3041
rect 9307 2720 9308 3040
rect 9628 2720 9629 3040
rect 9307 2719 9629 2720
rect 8888 2652 8984 2668
rect 9900 2668 9916 3092
rect 9980 2668 9996 3092
rect 10912 3092 11008 3108
rect 10319 3040 10641 3041
rect 10319 2720 10320 3040
rect 10640 2720 10641 3040
rect 10319 2719 10641 2720
rect 9900 2652 9996 2668
rect 10912 2668 10928 3092
rect 10992 2668 11008 3092
rect 11924 3092 12020 3108
rect 11331 3040 11653 3041
rect 11331 2720 11332 3040
rect 11652 2720 11653 3040
rect 11331 2719 11653 2720
rect 10912 2652 11008 2668
rect 11924 2668 11940 3092
rect 12004 2668 12020 3092
rect 12936 3092 13032 3108
rect 12343 3040 12665 3041
rect 12343 2720 12344 3040
rect 12664 2720 12665 3040
rect 12343 2719 12665 2720
rect 11924 2652 12020 2668
rect 12936 2668 12952 3092
rect 13016 2668 13032 3092
rect 13948 3092 14044 3108
rect 13355 3040 13677 3041
rect 13355 2720 13356 3040
rect 13676 2720 13677 3040
rect 13355 2719 13677 2720
rect 12936 2652 13032 2668
rect 13948 2668 13964 3092
rect 14028 2668 14044 3092
rect 14960 3092 15056 3108
rect 14367 3040 14689 3041
rect 14367 2720 14368 3040
rect 14688 2720 14689 3040
rect 14367 2719 14689 2720
rect 13948 2652 14044 2668
rect 14960 2668 14976 3092
rect 15040 2668 15056 3092
rect 15972 3092 16068 3108
rect 15379 3040 15701 3041
rect 15379 2720 15380 3040
rect 15700 2720 15701 3040
rect 15379 2719 15701 2720
rect 14960 2652 15056 2668
rect 15972 2668 15988 3092
rect 16052 2668 16068 3092
rect 16984 3092 17080 3108
rect 16391 3040 16713 3041
rect 16391 2720 16392 3040
rect 16712 2720 16713 3040
rect 16391 2719 16713 2720
rect 15972 2652 16068 2668
rect 16984 2668 17000 3092
rect 17064 2668 17080 3092
rect 16984 2652 17080 2668
rect -16412 2372 -16316 2388
rect -17005 2320 -16683 2321
rect -17005 2000 -17004 2320
rect -16684 2000 -16683 2320
rect -17005 1999 -16683 2000
rect -16412 1948 -16396 2372
rect -16332 1948 -16316 2372
rect -15400 2372 -15304 2388
rect -15993 2320 -15671 2321
rect -15993 2000 -15992 2320
rect -15672 2000 -15671 2320
rect -15993 1999 -15671 2000
rect -16412 1932 -16316 1948
rect -15400 1948 -15384 2372
rect -15320 1948 -15304 2372
rect -14388 2372 -14292 2388
rect -14981 2320 -14659 2321
rect -14981 2000 -14980 2320
rect -14660 2000 -14659 2320
rect -14981 1999 -14659 2000
rect -15400 1932 -15304 1948
rect -14388 1948 -14372 2372
rect -14308 1948 -14292 2372
rect -13376 2372 -13280 2388
rect -13969 2320 -13647 2321
rect -13969 2000 -13968 2320
rect -13648 2000 -13647 2320
rect -13969 1999 -13647 2000
rect -14388 1932 -14292 1948
rect -13376 1948 -13360 2372
rect -13296 1948 -13280 2372
rect -12364 2372 -12268 2388
rect -12957 2320 -12635 2321
rect -12957 2000 -12956 2320
rect -12636 2000 -12635 2320
rect -12957 1999 -12635 2000
rect -13376 1932 -13280 1948
rect -12364 1948 -12348 2372
rect -12284 1948 -12268 2372
rect -11352 2372 -11256 2388
rect -11945 2320 -11623 2321
rect -11945 2000 -11944 2320
rect -11624 2000 -11623 2320
rect -11945 1999 -11623 2000
rect -12364 1932 -12268 1948
rect -11352 1948 -11336 2372
rect -11272 1948 -11256 2372
rect -10340 2372 -10244 2388
rect -10933 2320 -10611 2321
rect -10933 2000 -10932 2320
rect -10612 2000 -10611 2320
rect -10933 1999 -10611 2000
rect -11352 1932 -11256 1948
rect -10340 1948 -10324 2372
rect -10260 1948 -10244 2372
rect -9328 2372 -9232 2388
rect -9921 2320 -9599 2321
rect -9921 2000 -9920 2320
rect -9600 2000 -9599 2320
rect -9921 1999 -9599 2000
rect -10340 1932 -10244 1948
rect -9328 1948 -9312 2372
rect -9248 1948 -9232 2372
rect -8316 2372 -8220 2388
rect -8909 2320 -8587 2321
rect -8909 2000 -8908 2320
rect -8588 2000 -8587 2320
rect -8909 1999 -8587 2000
rect -9328 1932 -9232 1948
rect -8316 1948 -8300 2372
rect -8236 1948 -8220 2372
rect -7304 2372 -7208 2388
rect -7897 2320 -7575 2321
rect -7897 2000 -7896 2320
rect -7576 2000 -7575 2320
rect -7897 1999 -7575 2000
rect -8316 1932 -8220 1948
rect -7304 1948 -7288 2372
rect -7224 1948 -7208 2372
rect -6292 2372 -6196 2388
rect -6885 2320 -6563 2321
rect -6885 2000 -6884 2320
rect -6564 2000 -6563 2320
rect -6885 1999 -6563 2000
rect -7304 1932 -7208 1948
rect -6292 1948 -6276 2372
rect -6212 1948 -6196 2372
rect -5280 2372 -5184 2388
rect -5873 2320 -5551 2321
rect -5873 2000 -5872 2320
rect -5552 2000 -5551 2320
rect -5873 1999 -5551 2000
rect -6292 1932 -6196 1948
rect -5280 1948 -5264 2372
rect -5200 1948 -5184 2372
rect -4268 2372 -4172 2388
rect -4861 2320 -4539 2321
rect -4861 2000 -4860 2320
rect -4540 2000 -4539 2320
rect -4861 1999 -4539 2000
rect -5280 1932 -5184 1948
rect -4268 1948 -4252 2372
rect -4188 1948 -4172 2372
rect -3256 2372 -3160 2388
rect -3849 2320 -3527 2321
rect -3849 2000 -3848 2320
rect -3528 2000 -3527 2320
rect -3849 1999 -3527 2000
rect -4268 1932 -4172 1948
rect -3256 1948 -3240 2372
rect -3176 1948 -3160 2372
rect -2244 2372 -2148 2388
rect -2837 2320 -2515 2321
rect -2837 2000 -2836 2320
rect -2516 2000 -2515 2320
rect -2837 1999 -2515 2000
rect -3256 1932 -3160 1948
rect -2244 1948 -2228 2372
rect -2164 1948 -2148 2372
rect -1232 2372 -1136 2388
rect -1825 2320 -1503 2321
rect -1825 2000 -1824 2320
rect -1504 2000 -1503 2320
rect -1825 1999 -1503 2000
rect -2244 1932 -2148 1948
rect -1232 1948 -1216 2372
rect -1152 1948 -1136 2372
rect -220 2372 -124 2388
rect -813 2320 -491 2321
rect -813 2000 -812 2320
rect -492 2000 -491 2320
rect -813 1999 -491 2000
rect -1232 1932 -1136 1948
rect -220 1948 -204 2372
rect -140 1948 -124 2372
rect 792 2372 888 2388
rect 199 2320 521 2321
rect 199 2000 200 2320
rect 520 2000 521 2320
rect 199 1999 521 2000
rect -220 1932 -124 1948
rect 792 1948 808 2372
rect 872 1948 888 2372
rect 1804 2372 1900 2388
rect 1211 2320 1533 2321
rect 1211 2000 1212 2320
rect 1532 2000 1533 2320
rect 1211 1999 1533 2000
rect 792 1932 888 1948
rect 1804 1948 1820 2372
rect 1884 1948 1900 2372
rect 2816 2372 2912 2388
rect 2223 2320 2545 2321
rect 2223 2000 2224 2320
rect 2544 2000 2545 2320
rect 2223 1999 2545 2000
rect 1804 1932 1900 1948
rect 2816 1948 2832 2372
rect 2896 1948 2912 2372
rect 3828 2372 3924 2388
rect 3235 2320 3557 2321
rect 3235 2000 3236 2320
rect 3556 2000 3557 2320
rect 3235 1999 3557 2000
rect 2816 1932 2912 1948
rect 3828 1948 3844 2372
rect 3908 1948 3924 2372
rect 4840 2372 4936 2388
rect 4247 2320 4569 2321
rect 4247 2000 4248 2320
rect 4568 2000 4569 2320
rect 4247 1999 4569 2000
rect 3828 1932 3924 1948
rect 4840 1948 4856 2372
rect 4920 1948 4936 2372
rect 5852 2372 5948 2388
rect 5259 2320 5581 2321
rect 5259 2000 5260 2320
rect 5580 2000 5581 2320
rect 5259 1999 5581 2000
rect 4840 1932 4936 1948
rect 5852 1948 5868 2372
rect 5932 1948 5948 2372
rect 6864 2372 6960 2388
rect 6271 2320 6593 2321
rect 6271 2000 6272 2320
rect 6592 2000 6593 2320
rect 6271 1999 6593 2000
rect 5852 1932 5948 1948
rect 6864 1948 6880 2372
rect 6944 1948 6960 2372
rect 7876 2372 7972 2388
rect 7283 2320 7605 2321
rect 7283 2000 7284 2320
rect 7604 2000 7605 2320
rect 7283 1999 7605 2000
rect 6864 1932 6960 1948
rect 7876 1948 7892 2372
rect 7956 1948 7972 2372
rect 8888 2372 8984 2388
rect 8295 2320 8617 2321
rect 8295 2000 8296 2320
rect 8616 2000 8617 2320
rect 8295 1999 8617 2000
rect 7876 1932 7972 1948
rect 8888 1948 8904 2372
rect 8968 1948 8984 2372
rect 9900 2372 9996 2388
rect 9307 2320 9629 2321
rect 9307 2000 9308 2320
rect 9628 2000 9629 2320
rect 9307 1999 9629 2000
rect 8888 1932 8984 1948
rect 9900 1948 9916 2372
rect 9980 1948 9996 2372
rect 10912 2372 11008 2388
rect 10319 2320 10641 2321
rect 10319 2000 10320 2320
rect 10640 2000 10641 2320
rect 10319 1999 10641 2000
rect 9900 1932 9996 1948
rect 10912 1948 10928 2372
rect 10992 1948 11008 2372
rect 11924 2372 12020 2388
rect 11331 2320 11653 2321
rect 11331 2000 11332 2320
rect 11652 2000 11653 2320
rect 11331 1999 11653 2000
rect 10912 1932 11008 1948
rect 11924 1948 11940 2372
rect 12004 1948 12020 2372
rect 12936 2372 13032 2388
rect 12343 2320 12665 2321
rect 12343 2000 12344 2320
rect 12664 2000 12665 2320
rect 12343 1999 12665 2000
rect 11924 1932 12020 1948
rect 12936 1948 12952 2372
rect 13016 1948 13032 2372
rect 13948 2372 14044 2388
rect 13355 2320 13677 2321
rect 13355 2000 13356 2320
rect 13676 2000 13677 2320
rect 13355 1999 13677 2000
rect 12936 1932 13032 1948
rect 13948 1948 13964 2372
rect 14028 1948 14044 2372
rect 14960 2372 15056 2388
rect 14367 2320 14689 2321
rect 14367 2000 14368 2320
rect 14688 2000 14689 2320
rect 14367 1999 14689 2000
rect 13948 1932 14044 1948
rect 14960 1948 14976 2372
rect 15040 1948 15056 2372
rect 15972 2372 16068 2388
rect 15379 2320 15701 2321
rect 15379 2000 15380 2320
rect 15700 2000 15701 2320
rect 15379 1999 15701 2000
rect 14960 1932 15056 1948
rect 15972 1948 15988 2372
rect 16052 1948 16068 2372
rect 16984 2372 17080 2388
rect 16391 2320 16713 2321
rect 16391 2000 16392 2320
rect 16712 2000 16713 2320
rect 16391 1999 16713 2000
rect 15972 1932 16068 1948
rect 16984 1948 17000 2372
rect 17064 1948 17080 2372
rect 16984 1932 17080 1948
rect -16412 1652 -16316 1668
rect -17005 1600 -16683 1601
rect -17005 1280 -17004 1600
rect -16684 1280 -16683 1600
rect -17005 1279 -16683 1280
rect -16412 1228 -16396 1652
rect -16332 1228 -16316 1652
rect -15400 1652 -15304 1668
rect -15993 1600 -15671 1601
rect -15993 1280 -15992 1600
rect -15672 1280 -15671 1600
rect -15993 1279 -15671 1280
rect -16412 1212 -16316 1228
rect -15400 1228 -15384 1652
rect -15320 1228 -15304 1652
rect -14388 1652 -14292 1668
rect -14981 1600 -14659 1601
rect -14981 1280 -14980 1600
rect -14660 1280 -14659 1600
rect -14981 1279 -14659 1280
rect -15400 1212 -15304 1228
rect -14388 1228 -14372 1652
rect -14308 1228 -14292 1652
rect -13376 1652 -13280 1668
rect -13969 1600 -13647 1601
rect -13969 1280 -13968 1600
rect -13648 1280 -13647 1600
rect -13969 1279 -13647 1280
rect -14388 1212 -14292 1228
rect -13376 1228 -13360 1652
rect -13296 1228 -13280 1652
rect -12364 1652 -12268 1668
rect -12957 1600 -12635 1601
rect -12957 1280 -12956 1600
rect -12636 1280 -12635 1600
rect -12957 1279 -12635 1280
rect -13376 1212 -13280 1228
rect -12364 1228 -12348 1652
rect -12284 1228 -12268 1652
rect -11352 1652 -11256 1668
rect -11945 1600 -11623 1601
rect -11945 1280 -11944 1600
rect -11624 1280 -11623 1600
rect -11945 1279 -11623 1280
rect -12364 1212 -12268 1228
rect -11352 1228 -11336 1652
rect -11272 1228 -11256 1652
rect -10340 1652 -10244 1668
rect -10933 1600 -10611 1601
rect -10933 1280 -10932 1600
rect -10612 1280 -10611 1600
rect -10933 1279 -10611 1280
rect -11352 1212 -11256 1228
rect -10340 1228 -10324 1652
rect -10260 1228 -10244 1652
rect -9328 1652 -9232 1668
rect -9921 1600 -9599 1601
rect -9921 1280 -9920 1600
rect -9600 1280 -9599 1600
rect -9921 1279 -9599 1280
rect -10340 1212 -10244 1228
rect -9328 1228 -9312 1652
rect -9248 1228 -9232 1652
rect -8316 1652 -8220 1668
rect -8909 1600 -8587 1601
rect -8909 1280 -8908 1600
rect -8588 1280 -8587 1600
rect -8909 1279 -8587 1280
rect -9328 1212 -9232 1228
rect -8316 1228 -8300 1652
rect -8236 1228 -8220 1652
rect -7304 1652 -7208 1668
rect -7897 1600 -7575 1601
rect -7897 1280 -7896 1600
rect -7576 1280 -7575 1600
rect -7897 1279 -7575 1280
rect -8316 1212 -8220 1228
rect -7304 1228 -7288 1652
rect -7224 1228 -7208 1652
rect -6292 1652 -6196 1668
rect -6885 1600 -6563 1601
rect -6885 1280 -6884 1600
rect -6564 1280 -6563 1600
rect -6885 1279 -6563 1280
rect -7304 1212 -7208 1228
rect -6292 1228 -6276 1652
rect -6212 1228 -6196 1652
rect -5280 1652 -5184 1668
rect -5873 1600 -5551 1601
rect -5873 1280 -5872 1600
rect -5552 1280 -5551 1600
rect -5873 1279 -5551 1280
rect -6292 1212 -6196 1228
rect -5280 1228 -5264 1652
rect -5200 1228 -5184 1652
rect -4268 1652 -4172 1668
rect -4861 1600 -4539 1601
rect -4861 1280 -4860 1600
rect -4540 1280 -4539 1600
rect -4861 1279 -4539 1280
rect -5280 1212 -5184 1228
rect -4268 1228 -4252 1652
rect -4188 1228 -4172 1652
rect -3256 1652 -3160 1668
rect -3849 1600 -3527 1601
rect -3849 1280 -3848 1600
rect -3528 1280 -3527 1600
rect -3849 1279 -3527 1280
rect -4268 1212 -4172 1228
rect -3256 1228 -3240 1652
rect -3176 1228 -3160 1652
rect -2244 1652 -2148 1668
rect -2837 1600 -2515 1601
rect -2837 1280 -2836 1600
rect -2516 1280 -2515 1600
rect -2837 1279 -2515 1280
rect -3256 1212 -3160 1228
rect -2244 1228 -2228 1652
rect -2164 1228 -2148 1652
rect -1232 1652 -1136 1668
rect -1825 1600 -1503 1601
rect -1825 1280 -1824 1600
rect -1504 1280 -1503 1600
rect -1825 1279 -1503 1280
rect -2244 1212 -2148 1228
rect -1232 1228 -1216 1652
rect -1152 1228 -1136 1652
rect -220 1652 -124 1668
rect -813 1600 -491 1601
rect -813 1280 -812 1600
rect -492 1280 -491 1600
rect -813 1279 -491 1280
rect -1232 1212 -1136 1228
rect -220 1228 -204 1652
rect -140 1228 -124 1652
rect 792 1652 888 1668
rect 199 1600 521 1601
rect 199 1280 200 1600
rect 520 1280 521 1600
rect 199 1279 521 1280
rect -220 1212 -124 1228
rect 792 1228 808 1652
rect 872 1228 888 1652
rect 1804 1652 1900 1668
rect 1211 1600 1533 1601
rect 1211 1280 1212 1600
rect 1532 1280 1533 1600
rect 1211 1279 1533 1280
rect 792 1212 888 1228
rect 1804 1228 1820 1652
rect 1884 1228 1900 1652
rect 2816 1652 2912 1668
rect 2223 1600 2545 1601
rect 2223 1280 2224 1600
rect 2544 1280 2545 1600
rect 2223 1279 2545 1280
rect 1804 1212 1900 1228
rect 2816 1228 2832 1652
rect 2896 1228 2912 1652
rect 3828 1652 3924 1668
rect 3235 1600 3557 1601
rect 3235 1280 3236 1600
rect 3556 1280 3557 1600
rect 3235 1279 3557 1280
rect 2816 1212 2912 1228
rect 3828 1228 3844 1652
rect 3908 1228 3924 1652
rect 4840 1652 4936 1668
rect 4247 1600 4569 1601
rect 4247 1280 4248 1600
rect 4568 1280 4569 1600
rect 4247 1279 4569 1280
rect 3828 1212 3924 1228
rect 4840 1228 4856 1652
rect 4920 1228 4936 1652
rect 5852 1652 5948 1668
rect 5259 1600 5581 1601
rect 5259 1280 5260 1600
rect 5580 1280 5581 1600
rect 5259 1279 5581 1280
rect 4840 1212 4936 1228
rect 5852 1228 5868 1652
rect 5932 1228 5948 1652
rect 6864 1652 6960 1668
rect 6271 1600 6593 1601
rect 6271 1280 6272 1600
rect 6592 1280 6593 1600
rect 6271 1279 6593 1280
rect 5852 1212 5948 1228
rect 6864 1228 6880 1652
rect 6944 1228 6960 1652
rect 7876 1652 7972 1668
rect 7283 1600 7605 1601
rect 7283 1280 7284 1600
rect 7604 1280 7605 1600
rect 7283 1279 7605 1280
rect 6864 1212 6960 1228
rect 7876 1228 7892 1652
rect 7956 1228 7972 1652
rect 8888 1652 8984 1668
rect 8295 1600 8617 1601
rect 8295 1280 8296 1600
rect 8616 1280 8617 1600
rect 8295 1279 8617 1280
rect 7876 1212 7972 1228
rect 8888 1228 8904 1652
rect 8968 1228 8984 1652
rect 9900 1652 9996 1668
rect 9307 1600 9629 1601
rect 9307 1280 9308 1600
rect 9628 1280 9629 1600
rect 9307 1279 9629 1280
rect 8888 1212 8984 1228
rect 9900 1228 9916 1652
rect 9980 1228 9996 1652
rect 10912 1652 11008 1668
rect 10319 1600 10641 1601
rect 10319 1280 10320 1600
rect 10640 1280 10641 1600
rect 10319 1279 10641 1280
rect 9900 1212 9996 1228
rect 10912 1228 10928 1652
rect 10992 1228 11008 1652
rect 11924 1652 12020 1668
rect 11331 1600 11653 1601
rect 11331 1280 11332 1600
rect 11652 1280 11653 1600
rect 11331 1279 11653 1280
rect 10912 1212 11008 1228
rect 11924 1228 11940 1652
rect 12004 1228 12020 1652
rect 12936 1652 13032 1668
rect 12343 1600 12665 1601
rect 12343 1280 12344 1600
rect 12664 1280 12665 1600
rect 12343 1279 12665 1280
rect 11924 1212 12020 1228
rect 12936 1228 12952 1652
rect 13016 1228 13032 1652
rect 13948 1652 14044 1668
rect 13355 1600 13677 1601
rect 13355 1280 13356 1600
rect 13676 1280 13677 1600
rect 13355 1279 13677 1280
rect 12936 1212 13032 1228
rect 13948 1228 13964 1652
rect 14028 1228 14044 1652
rect 14960 1652 15056 1668
rect 14367 1600 14689 1601
rect 14367 1280 14368 1600
rect 14688 1280 14689 1600
rect 14367 1279 14689 1280
rect 13948 1212 14044 1228
rect 14960 1228 14976 1652
rect 15040 1228 15056 1652
rect 15972 1652 16068 1668
rect 15379 1600 15701 1601
rect 15379 1280 15380 1600
rect 15700 1280 15701 1600
rect 15379 1279 15701 1280
rect 14960 1212 15056 1228
rect 15972 1228 15988 1652
rect 16052 1228 16068 1652
rect 16984 1652 17080 1668
rect 16391 1600 16713 1601
rect 16391 1280 16392 1600
rect 16712 1280 16713 1600
rect 16391 1279 16713 1280
rect 15972 1212 16068 1228
rect 16984 1228 17000 1652
rect 17064 1228 17080 1652
rect 16984 1212 17080 1228
rect -16412 932 -16316 948
rect -17005 880 -16683 881
rect -17005 560 -17004 880
rect -16684 560 -16683 880
rect -17005 559 -16683 560
rect -16412 508 -16396 932
rect -16332 508 -16316 932
rect -15400 932 -15304 948
rect -15993 880 -15671 881
rect -15993 560 -15992 880
rect -15672 560 -15671 880
rect -15993 559 -15671 560
rect -16412 492 -16316 508
rect -15400 508 -15384 932
rect -15320 508 -15304 932
rect -14388 932 -14292 948
rect -14981 880 -14659 881
rect -14981 560 -14980 880
rect -14660 560 -14659 880
rect -14981 559 -14659 560
rect -15400 492 -15304 508
rect -14388 508 -14372 932
rect -14308 508 -14292 932
rect -13376 932 -13280 948
rect -13969 880 -13647 881
rect -13969 560 -13968 880
rect -13648 560 -13647 880
rect -13969 559 -13647 560
rect -14388 492 -14292 508
rect -13376 508 -13360 932
rect -13296 508 -13280 932
rect -12364 932 -12268 948
rect -12957 880 -12635 881
rect -12957 560 -12956 880
rect -12636 560 -12635 880
rect -12957 559 -12635 560
rect -13376 492 -13280 508
rect -12364 508 -12348 932
rect -12284 508 -12268 932
rect -11352 932 -11256 948
rect -11945 880 -11623 881
rect -11945 560 -11944 880
rect -11624 560 -11623 880
rect -11945 559 -11623 560
rect -12364 492 -12268 508
rect -11352 508 -11336 932
rect -11272 508 -11256 932
rect -10340 932 -10244 948
rect -10933 880 -10611 881
rect -10933 560 -10932 880
rect -10612 560 -10611 880
rect -10933 559 -10611 560
rect -11352 492 -11256 508
rect -10340 508 -10324 932
rect -10260 508 -10244 932
rect -9328 932 -9232 948
rect -9921 880 -9599 881
rect -9921 560 -9920 880
rect -9600 560 -9599 880
rect -9921 559 -9599 560
rect -10340 492 -10244 508
rect -9328 508 -9312 932
rect -9248 508 -9232 932
rect -8316 932 -8220 948
rect -8909 880 -8587 881
rect -8909 560 -8908 880
rect -8588 560 -8587 880
rect -8909 559 -8587 560
rect -9328 492 -9232 508
rect -8316 508 -8300 932
rect -8236 508 -8220 932
rect -7304 932 -7208 948
rect -7897 880 -7575 881
rect -7897 560 -7896 880
rect -7576 560 -7575 880
rect -7897 559 -7575 560
rect -8316 492 -8220 508
rect -7304 508 -7288 932
rect -7224 508 -7208 932
rect -6292 932 -6196 948
rect -6885 880 -6563 881
rect -6885 560 -6884 880
rect -6564 560 -6563 880
rect -6885 559 -6563 560
rect -7304 492 -7208 508
rect -6292 508 -6276 932
rect -6212 508 -6196 932
rect -5280 932 -5184 948
rect -5873 880 -5551 881
rect -5873 560 -5872 880
rect -5552 560 -5551 880
rect -5873 559 -5551 560
rect -6292 492 -6196 508
rect -5280 508 -5264 932
rect -5200 508 -5184 932
rect -4268 932 -4172 948
rect -4861 880 -4539 881
rect -4861 560 -4860 880
rect -4540 560 -4539 880
rect -4861 559 -4539 560
rect -5280 492 -5184 508
rect -4268 508 -4252 932
rect -4188 508 -4172 932
rect -3256 932 -3160 948
rect -3849 880 -3527 881
rect -3849 560 -3848 880
rect -3528 560 -3527 880
rect -3849 559 -3527 560
rect -4268 492 -4172 508
rect -3256 508 -3240 932
rect -3176 508 -3160 932
rect -2244 932 -2148 948
rect -2837 880 -2515 881
rect -2837 560 -2836 880
rect -2516 560 -2515 880
rect -2837 559 -2515 560
rect -3256 492 -3160 508
rect -2244 508 -2228 932
rect -2164 508 -2148 932
rect -1232 932 -1136 948
rect -1825 880 -1503 881
rect -1825 560 -1824 880
rect -1504 560 -1503 880
rect -1825 559 -1503 560
rect -2244 492 -2148 508
rect -1232 508 -1216 932
rect -1152 508 -1136 932
rect -220 932 -124 948
rect -813 880 -491 881
rect -813 560 -812 880
rect -492 560 -491 880
rect -813 559 -491 560
rect -1232 492 -1136 508
rect -220 508 -204 932
rect -140 508 -124 932
rect 792 932 888 948
rect 199 880 521 881
rect 199 560 200 880
rect 520 560 521 880
rect 199 559 521 560
rect -220 492 -124 508
rect 792 508 808 932
rect 872 508 888 932
rect 1804 932 1900 948
rect 1211 880 1533 881
rect 1211 560 1212 880
rect 1532 560 1533 880
rect 1211 559 1533 560
rect 792 492 888 508
rect 1804 508 1820 932
rect 1884 508 1900 932
rect 2816 932 2912 948
rect 2223 880 2545 881
rect 2223 560 2224 880
rect 2544 560 2545 880
rect 2223 559 2545 560
rect 1804 492 1900 508
rect 2816 508 2832 932
rect 2896 508 2912 932
rect 3828 932 3924 948
rect 3235 880 3557 881
rect 3235 560 3236 880
rect 3556 560 3557 880
rect 3235 559 3557 560
rect 2816 492 2912 508
rect 3828 508 3844 932
rect 3908 508 3924 932
rect 4840 932 4936 948
rect 4247 880 4569 881
rect 4247 560 4248 880
rect 4568 560 4569 880
rect 4247 559 4569 560
rect 3828 492 3924 508
rect 4840 508 4856 932
rect 4920 508 4936 932
rect 5852 932 5948 948
rect 5259 880 5581 881
rect 5259 560 5260 880
rect 5580 560 5581 880
rect 5259 559 5581 560
rect 4840 492 4936 508
rect 5852 508 5868 932
rect 5932 508 5948 932
rect 6864 932 6960 948
rect 6271 880 6593 881
rect 6271 560 6272 880
rect 6592 560 6593 880
rect 6271 559 6593 560
rect 5852 492 5948 508
rect 6864 508 6880 932
rect 6944 508 6960 932
rect 7876 932 7972 948
rect 7283 880 7605 881
rect 7283 560 7284 880
rect 7604 560 7605 880
rect 7283 559 7605 560
rect 6864 492 6960 508
rect 7876 508 7892 932
rect 7956 508 7972 932
rect 8888 932 8984 948
rect 8295 880 8617 881
rect 8295 560 8296 880
rect 8616 560 8617 880
rect 8295 559 8617 560
rect 7876 492 7972 508
rect 8888 508 8904 932
rect 8968 508 8984 932
rect 9900 932 9996 948
rect 9307 880 9629 881
rect 9307 560 9308 880
rect 9628 560 9629 880
rect 9307 559 9629 560
rect 8888 492 8984 508
rect 9900 508 9916 932
rect 9980 508 9996 932
rect 10912 932 11008 948
rect 10319 880 10641 881
rect 10319 560 10320 880
rect 10640 560 10641 880
rect 10319 559 10641 560
rect 9900 492 9996 508
rect 10912 508 10928 932
rect 10992 508 11008 932
rect 11924 932 12020 948
rect 11331 880 11653 881
rect 11331 560 11332 880
rect 11652 560 11653 880
rect 11331 559 11653 560
rect 10912 492 11008 508
rect 11924 508 11940 932
rect 12004 508 12020 932
rect 12936 932 13032 948
rect 12343 880 12665 881
rect 12343 560 12344 880
rect 12664 560 12665 880
rect 12343 559 12665 560
rect 11924 492 12020 508
rect 12936 508 12952 932
rect 13016 508 13032 932
rect 13948 932 14044 948
rect 13355 880 13677 881
rect 13355 560 13356 880
rect 13676 560 13677 880
rect 13355 559 13677 560
rect 12936 492 13032 508
rect 13948 508 13964 932
rect 14028 508 14044 932
rect 14960 932 15056 948
rect 14367 880 14689 881
rect 14367 560 14368 880
rect 14688 560 14689 880
rect 14367 559 14689 560
rect 13948 492 14044 508
rect 14960 508 14976 932
rect 15040 508 15056 932
rect 15972 932 16068 948
rect 15379 880 15701 881
rect 15379 560 15380 880
rect 15700 560 15701 880
rect 15379 559 15701 560
rect 14960 492 15056 508
rect 15972 508 15988 932
rect 16052 508 16068 932
rect 16984 932 17080 948
rect 16391 880 16713 881
rect 16391 560 16392 880
rect 16712 560 16713 880
rect 16391 559 16713 560
rect 15972 492 16068 508
rect 16984 508 17000 932
rect 17064 508 17080 932
rect 16984 492 17080 508
rect -16412 212 -16316 228
rect -17005 160 -16683 161
rect -17005 -160 -17004 160
rect -16684 -160 -16683 160
rect -17005 -161 -16683 -160
rect -16412 -212 -16396 212
rect -16332 -212 -16316 212
rect -15400 212 -15304 228
rect -15993 160 -15671 161
rect -15993 -160 -15992 160
rect -15672 -160 -15671 160
rect -15993 -161 -15671 -160
rect -16412 -228 -16316 -212
rect -15400 -212 -15384 212
rect -15320 -212 -15304 212
rect -14388 212 -14292 228
rect -14981 160 -14659 161
rect -14981 -160 -14980 160
rect -14660 -160 -14659 160
rect -14981 -161 -14659 -160
rect -15400 -228 -15304 -212
rect -14388 -212 -14372 212
rect -14308 -212 -14292 212
rect -13376 212 -13280 228
rect -13969 160 -13647 161
rect -13969 -160 -13968 160
rect -13648 -160 -13647 160
rect -13969 -161 -13647 -160
rect -14388 -228 -14292 -212
rect -13376 -212 -13360 212
rect -13296 -212 -13280 212
rect -12364 212 -12268 228
rect -12957 160 -12635 161
rect -12957 -160 -12956 160
rect -12636 -160 -12635 160
rect -12957 -161 -12635 -160
rect -13376 -228 -13280 -212
rect -12364 -212 -12348 212
rect -12284 -212 -12268 212
rect -11352 212 -11256 228
rect -11945 160 -11623 161
rect -11945 -160 -11944 160
rect -11624 -160 -11623 160
rect -11945 -161 -11623 -160
rect -12364 -228 -12268 -212
rect -11352 -212 -11336 212
rect -11272 -212 -11256 212
rect -10340 212 -10244 228
rect -10933 160 -10611 161
rect -10933 -160 -10932 160
rect -10612 -160 -10611 160
rect -10933 -161 -10611 -160
rect -11352 -228 -11256 -212
rect -10340 -212 -10324 212
rect -10260 -212 -10244 212
rect -9328 212 -9232 228
rect -9921 160 -9599 161
rect -9921 -160 -9920 160
rect -9600 -160 -9599 160
rect -9921 -161 -9599 -160
rect -10340 -228 -10244 -212
rect -9328 -212 -9312 212
rect -9248 -212 -9232 212
rect -8316 212 -8220 228
rect -8909 160 -8587 161
rect -8909 -160 -8908 160
rect -8588 -160 -8587 160
rect -8909 -161 -8587 -160
rect -9328 -228 -9232 -212
rect -8316 -212 -8300 212
rect -8236 -212 -8220 212
rect -7304 212 -7208 228
rect -7897 160 -7575 161
rect -7897 -160 -7896 160
rect -7576 -160 -7575 160
rect -7897 -161 -7575 -160
rect -8316 -228 -8220 -212
rect -7304 -212 -7288 212
rect -7224 -212 -7208 212
rect -6292 212 -6196 228
rect -6885 160 -6563 161
rect -6885 -160 -6884 160
rect -6564 -160 -6563 160
rect -6885 -161 -6563 -160
rect -7304 -228 -7208 -212
rect -6292 -212 -6276 212
rect -6212 -212 -6196 212
rect -5280 212 -5184 228
rect -5873 160 -5551 161
rect -5873 -160 -5872 160
rect -5552 -160 -5551 160
rect -5873 -161 -5551 -160
rect -6292 -228 -6196 -212
rect -5280 -212 -5264 212
rect -5200 -212 -5184 212
rect -4268 212 -4172 228
rect -4861 160 -4539 161
rect -4861 -160 -4860 160
rect -4540 -160 -4539 160
rect -4861 -161 -4539 -160
rect -5280 -228 -5184 -212
rect -4268 -212 -4252 212
rect -4188 -212 -4172 212
rect -3256 212 -3160 228
rect -3849 160 -3527 161
rect -3849 -160 -3848 160
rect -3528 -160 -3527 160
rect -3849 -161 -3527 -160
rect -4268 -228 -4172 -212
rect -3256 -212 -3240 212
rect -3176 -212 -3160 212
rect -2244 212 -2148 228
rect -2837 160 -2515 161
rect -2837 -160 -2836 160
rect -2516 -160 -2515 160
rect -2837 -161 -2515 -160
rect -3256 -228 -3160 -212
rect -2244 -212 -2228 212
rect -2164 -212 -2148 212
rect -1232 212 -1136 228
rect -1825 160 -1503 161
rect -1825 -160 -1824 160
rect -1504 -160 -1503 160
rect -1825 -161 -1503 -160
rect -2244 -228 -2148 -212
rect -1232 -212 -1216 212
rect -1152 -212 -1136 212
rect -220 212 -124 228
rect -813 160 -491 161
rect -813 -160 -812 160
rect -492 -160 -491 160
rect -813 -161 -491 -160
rect -1232 -228 -1136 -212
rect -220 -212 -204 212
rect -140 -212 -124 212
rect 792 212 888 228
rect 199 160 521 161
rect 199 -160 200 160
rect 520 -160 521 160
rect 199 -161 521 -160
rect -220 -228 -124 -212
rect 792 -212 808 212
rect 872 -212 888 212
rect 1804 212 1900 228
rect 1211 160 1533 161
rect 1211 -160 1212 160
rect 1532 -160 1533 160
rect 1211 -161 1533 -160
rect 792 -228 888 -212
rect 1804 -212 1820 212
rect 1884 -212 1900 212
rect 2816 212 2912 228
rect 2223 160 2545 161
rect 2223 -160 2224 160
rect 2544 -160 2545 160
rect 2223 -161 2545 -160
rect 1804 -228 1900 -212
rect 2816 -212 2832 212
rect 2896 -212 2912 212
rect 3828 212 3924 228
rect 3235 160 3557 161
rect 3235 -160 3236 160
rect 3556 -160 3557 160
rect 3235 -161 3557 -160
rect 2816 -228 2912 -212
rect 3828 -212 3844 212
rect 3908 -212 3924 212
rect 4840 212 4936 228
rect 4247 160 4569 161
rect 4247 -160 4248 160
rect 4568 -160 4569 160
rect 4247 -161 4569 -160
rect 3828 -228 3924 -212
rect 4840 -212 4856 212
rect 4920 -212 4936 212
rect 5852 212 5948 228
rect 5259 160 5581 161
rect 5259 -160 5260 160
rect 5580 -160 5581 160
rect 5259 -161 5581 -160
rect 4840 -228 4936 -212
rect 5852 -212 5868 212
rect 5932 -212 5948 212
rect 6864 212 6960 228
rect 6271 160 6593 161
rect 6271 -160 6272 160
rect 6592 -160 6593 160
rect 6271 -161 6593 -160
rect 5852 -228 5948 -212
rect 6864 -212 6880 212
rect 6944 -212 6960 212
rect 7876 212 7972 228
rect 7283 160 7605 161
rect 7283 -160 7284 160
rect 7604 -160 7605 160
rect 7283 -161 7605 -160
rect 6864 -228 6960 -212
rect 7876 -212 7892 212
rect 7956 -212 7972 212
rect 8888 212 8984 228
rect 8295 160 8617 161
rect 8295 -160 8296 160
rect 8616 -160 8617 160
rect 8295 -161 8617 -160
rect 7876 -228 7972 -212
rect 8888 -212 8904 212
rect 8968 -212 8984 212
rect 9900 212 9996 228
rect 9307 160 9629 161
rect 9307 -160 9308 160
rect 9628 -160 9629 160
rect 9307 -161 9629 -160
rect 8888 -228 8984 -212
rect 9900 -212 9916 212
rect 9980 -212 9996 212
rect 10912 212 11008 228
rect 10319 160 10641 161
rect 10319 -160 10320 160
rect 10640 -160 10641 160
rect 10319 -161 10641 -160
rect 9900 -228 9996 -212
rect 10912 -212 10928 212
rect 10992 -212 11008 212
rect 11924 212 12020 228
rect 11331 160 11653 161
rect 11331 -160 11332 160
rect 11652 -160 11653 160
rect 11331 -161 11653 -160
rect 10912 -228 11008 -212
rect 11924 -212 11940 212
rect 12004 -212 12020 212
rect 12936 212 13032 228
rect 12343 160 12665 161
rect 12343 -160 12344 160
rect 12664 -160 12665 160
rect 12343 -161 12665 -160
rect 11924 -228 12020 -212
rect 12936 -212 12952 212
rect 13016 -212 13032 212
rect 13948 212 14044 228
rect 13355 160 13677 161
rect 13355 -160 13356 160
rect 13676 -160 13677 160
rect 13355 -161 13677 -160
rect 12936 -228 13032 -212
rect 13948 -212 13964 212
rect 14028 -212 14044 212
rect 14960 212 15056 228
rect 14367 160 14689 161
rect 14367 -160 14368 160
rect 14688 -160 14689 160
rect 14367 -161 14689 -160
rect 13948 -228 14044 -212
rect 14960 -212 14976 212
rect 15040 -212 15056 212
rect 15972 212 16068 228
rect 15379 160 15701 161
rect 15379 -160 15380 160
rect 15700 -160 15701 160
rect 15379 -161 15701 -160
rect 14960 -228 15056 -212
rect 15972 -212 15988 212
rect 16052 -212 16068 212
rect 16984 212 17080 228
rect 16391 160 16713 161
rect 16391 -160 16392 160
rect 16712 -160 16713 160
rect 16391 -161 16713 -160
rect 15972 -228 16068 -212
rect 16984 -212 17000 212
rect 17064 -212 17080 212
rect 16984 -228 17080 -212
rect -16412 -508 -16316 -492
rect -17005 -560 -16683 -559
rect -17005 -880 -17004 -560
rect -16684 -880 -16683 -560
rect -17005 -881 -16683 -880
rect -16412 -932 -16396 -508
rect -16332 -932 -16316 -508
rect -15400 -508 -15304 -492
rect -15993 -560 -15671 -559
rect -15993 -880 -15992 -560
rect -15672 -880 -15671 -560
rect -15993 -881 -15671 -880
rect -16412 -948 -16316 -932
rect -15400 -932 -15384 -508
rect -15320 -932 -15304 -508
rect -14388 -508 -14292 -492
rect -14981 -560 -14659 -559
rect -14981 -880 -14980 -560
rect -14660 -880 -14659 -560
rect -14981 -881 -14659 -880
rect -15400 -948 -15304 -932
rect -14388 -932 -14372 -508
rect -14308 -932 -14292 -508
rect -13376 -508 -13280 -492
rect -13969 -560 -13647 -559
rect -13969 -880 -13968 -560
rect -13648 -880 -13647 -560
rect -13969 -881 -13647 -880
rect -14388 -948 -14292 -932
rect -13376 -932 -13360 -508
rect -13296 -932 -13280 -508
rect -12364 -508 -12268 -492
rect -12957 -560 -12635 -559
rect -12957 -880 -12956 -560
rect -12636 -880 -12635 -560
rect -12957 -881 -12635 -880
rect -13376 -948 -13280 -932
rect -12364 -932 -12348 -508
rect -12284 -932 -12268 -508
rect -11352 -508 -11256 -492
rect -11945 -560 -11623 -559
rect -11945 -880 -11944 -560
rect -11624 -880 -11623 -560
rect -11945 -881 -11623 -880
rect -12364 -948 -12268 -932
rect -11352 -932 -11336 -508
rect -11272 -932 -11256 -508
rect -10340 -508 -10244 -492
rect -10933 -560 -10611 -559
rect -10933 -880 -10932 -560
rect -10612 -880 -10611 -560
rect -10933 -881 -10611 -880
rect -11352 -948 -11256 -932
rect -10340 -932 -10324 -508
rect -10260 -932 -10244 -508
rect -9328 -508 -9232 -492
rect -9921 -560 -9599 -559
rect -9921 -880 -9920 -560
rect -9600 -880 -9599 -560
rect -9921 -881 -9599 -880
rect -10340 -948 -10244 -932
rect -9328 -932 -9312 -508
rect -9248 -932 -9232 -508
rect -8316 -508 -8220 -492
rect -8909 -560 -8587 -559
rect -8909 -880 -8908 -560
rect -8588 -880 -8587 -560
rect -8909 -881 -8587 -880
rect -9328 -948 -9232 -932
rect -8316 -932 -8300 -508
rect -8236 -932 -8220 -508
rect -7304 -508 -7208 -492
rect -7897 -560 -7575 -559
rect -7897 -880 -7896 -560
rect -7576 -880 -7575 -560
rect -7897 -881 -7575 -880
rect -8316 -948 -8220 -932
rect -7304 -932 -7288 -508
rect -7224 -932 -7208 -508
rect -6292 -508 -6196 -492
rect -6885 -560 -6563 -559
rect -6885 -880 -6884 -560
rect -6564 -880 -6563 -560
rect -6885 -881 -6563 -880
rect -7304 -948 -7208 -932
rect -6292 -932 -6276 -508
rect -6212 -932 -6196 -508
rect -5280 -508 -5184 -492
rect -5873 -560 -5551 -559
rect -5873 -880 -5872 -560
rect -5552 -880 -5551 -560
rect -5873 -881 -5551 -880
rect -6292 -948 -6196 -932
rect -5280 -932 -5264 -508
rect -5200 -932 -5184 -508
rect -4268 -508 -4172 -492
rect -4861 -560 -4539 -559
rect -4861 -880 -4860 -560
rect -4540 -880 -4539 -560
rect -4861 -881 -4539 -880
rect -5280 -948 -5184 -932
rect -4268 -932 -4252 -508
rect -4188 -932 -4172 -508
rect -3256 -508 -3160 -492
rect -3849 -560 -3527 -559
rect -3849 -880 -3848 -560
rect -3528 -880 -3527 -560
rect -3849 -881 -3527 -880
rect -4268 -948 -4172 -932
rect -3256 -932 -3240 -508
rect -3176 -932 -3160 -508
rect -2244 -508 -2148 -492
rect -2837 -560 -2515 -559
rect -2837 -880 -2836 -560
rect -2516 -880 -2515 -560
rect -2837 -881 -2515 -880
rect -3256 -948 -3160 -932
rect -2244 -932 -2228 -508
rect -2164 -932 -2148 -508
rect -1232 -508 -1136 -492
rect -1825 -560 -1503 -559
rect -1825 -880 -1824 -560
rect -1504 -880 -1503 -560
rect -1825 -881 -1503 -880
rect -2244 -948 -2148 -932
rect -1232 -932 -1216 -508
rect -1152 -932 -1136 -508
rect -220 -508 -124 -492
rect -813 -560 -491 -559
rect -813 -880 -812 -560
rect -492 -880 -491 -560
rect -813 -881 -491 -880
rect -1232 -948 -1136 -932
rect -220 -932 -204 -508
rect -140 -932 -124 -508
rect 792 -508 888 -492
rect 199 -560 521 -559
rect 199 -880 200 -560
rect 520 -880 521 -560
rect 199 -881 521 -880
rect -220 -948 -124 -932
rect 792 -932 808 -508
rect 872 -932 888 -508
rect 1804 -508 1900 -492
rect 1211 -560 1533 -559
rect 1211 -880 1212 -560
rect 1532 -880 1533 -560
rect 1211 -881 1533 -880
rect 792 -948 888 -932
rect 1804 -932 1820 -508
rect 1884 -932 1900 -508
rect 2816 -508 2912 -492
rect 2223 -560 2545 -559
rect 2223 -880 2224 -560
rect 2544 -880 2545 -560
rect 2223 -881 2545 -880
rect 1804 -948 1900 -932
rect 2816 -932 2832 -508
rect 2896 -932 2912 -508
rect 3828 -508 3924 -492
rect 3235 -560 3557 -559
rect 3235 -880 3236 -560
rect 3556 -880 3557 -560
rect 3235 -881 3557 -880
rect 2816 -948 2912 -932
rect 3828 -932 3844 -508
rect 3908 -932 3924 -508
rect 4840 -508 4936 -492
rect 4247 -560 4569 -559
rect 4247 -880 4248 -560
rect 4568 -880 4569 -560
rect 4247 -881 4569 -880
rect 3828 -948 3924 -932
rect 4840 -932 4856 -508
rect 4920 -932 4936 -508
rect 5852 -508 5948 -492
rect 5259 -560 5581 -559
rect 5259 -880 5260 -560
rect 5580 -880 5581 -560
rect 5259 -881 5581 -880
rect 4840 -948 4936 -932
rect 5852 -932 5868 -508
rect 5932 -932 5948 -508
rect 6864 -508 6960 -492
rect 6271 -560 6593 -559
rect 6271 -880 6272 -560
rect 6592 -880 6593 -560
rect 6271 -881 6593 -880
rect 5852 -948 5948 -932
rect 6864 -932 6880 -508
rect 6944 -932 6960 -508
rect 7876 -508 7972 -492
rect 7283 -560 7605 -559
rect 7283 -880 7284 -560
rect 7604 -880 7605 -560
rect 7283 -881 7605 -880
rect 6864 -948 6960 -932
rect 7876 -932 7892 -508
rect 7956 -932 7972 -508
rect 8888 -508 8984 -492
rect 8295 -560 8617 -559
rect 8295 -880 8296 -560
rect 8616 -880 8617 -560
rect 8295 -881 8617 -880
rect 7876 -948 7972 -932
rect 8888 -932 8904 -508
rect 8968 -932 8984 -508
rect 9900 -508 9996 -492
rect 9307 -560 9629 -559
rect 9307 -880 9308 -560
rect 9628 -880 9629 -560
rect 9307 -881 9629 -880
rect 8888 -948 8984 -932
rect 9900 -932 9916 -508
rect 9980 -932 9996 -508
rect 10912 -508 11008 -492
rect 10319 -560 10641 -559
rect 10319 -880 10320 -560
rect 10640 -880 10641 -560
rect 10319 -881 10641 -880
rect 9900 -948 9996 -932
rect 10912 -932 10928 -508
rect 10992 -932 11008 -508
rect 11924 -508 12020 -492
rect 11331 -560 11653 -559
rect 11331 -880 11332 -560
rect 11652 -880 11653 -560
rect 11331 -881 11653 -880
rect 10912 -948 11008 -932
rect 11924 -932 11940 -508
rect 12004 -932 12020 -508
rect 12936 -508 13032 -492
rect 12343 -560 12665 -559
rect 12343 -880 12344 -560
rect 12664 -880 12665 -560
rect 12343 -881 12665 -880
rect 11924 -948 12020 -932
rect 12936 -932 12952 -508
rect 13016 -932 13032 -508
rect 13948 -508 14044 -492
rect 13355 -560 13677 -559
rect 13355 -880 13356 -560
rect 13676 -880 13677 -560
rect 13355 -881 13677 -880
rect 12936 -948 13032 -932
rect 13948 -932 13964 -508
rect 14028 -932 14044 -508
rect 14960 -508 15056 -492
rect 14367 -560 14689 -559
rect 14367 -880 14368 -560
rect 14688 -880 14689 -560
rect 14367 -881 14689 -880
rect 13948 -948 14044 -932
rect 14960 -932 14976 -508
rect 15040 -932 15056 -508
rect 15972 -508 16068 -492
rect 15379 -560 15701 -559
rect 15379 -880 15380 -560
rect 15700 -880 15701 -560
rect 15379 -881 15701 -880
rect 14960 -948 15056 -932
rect 15972 -932 15988 -508
rect 16052 -932 16068 -508
rect 16984 -508 17080 -492
rect 16391 -560 16713 -559
rect 16391 -880 16392 -560
rect 16712 -880 16713 -560
rect 16391 -881 16713 -880
rect 15972 -948 16068 -932
rect 16984 -932 17000 -508
rect 17064 -932 17080 -508
rect 16984 -948 17080 -932
rect -16412 -1228 -16316 -1212
rect -17005 -1280 -16683 -1279
rect -17005 -1600 -17004 -1280
rect -16684 -1600 -16683 -1280
rect -17005 -1601 -16683 -1600
rect -16412 -1652 -16396 -1228
rect -16332 -1652 -16316 -1228
rect -15400 -1228 -15304 -1212
rect -15993 -1280 -15671 -1279
rect -15993 -1600 -15992 -1280
rect -15672 -1600 -15671 -1280
rect -15993 -1601 -15671 -1600
rect -16412 -1668 -16316 -1652
rect -15400 -1652 -15384 -1228
rect -15320 -1652 -15304 -1228
rect -14388 -1228 -14292 -1212
rect -14981 -1280 -14659 -1279
rect -14981 -1600 -14980 -1280
rect -14660 -1600 -14659 -1280
rect -14981 -1601 -14659 -1600
rect -15400 -1668 -15304 -1652
rect -14388 -1652 -14372 -1228
rect -14308 -1652 -14292 -1228
rect -13376 -1228 -13280 -1212
rect -13969 -1280 -13647 -1279
rect -13969 -1600 -13968 -1280
rect -13648 -1600 -13647 -1280
rect -13969 -1601 -13647 -1600
rect -14388 -1668 -14292 -1652
rect -13376 -1652 -13360 -1228
rect -13296 -1652 -13280 -1228
rect -12364 -1228 -12268 -1212
rect -12957 -1280 -12635 -1279
rect -12957 -1600 -12956 -1280
rect -12636 -1600 -12635 -1280
rect -12957 -1601 -12635 -1600
rect -13376 -1668 -13280 -1652
rect -12364 -1652 -12348 -1228
rect -12284 -1652 -12268 -1228
rect -11352 -1228 -11256 -1212
rect -11945 -1280 -11623 -1279
rect -11945 -1600 -11944 -1280
rect -11624 -1600 -11623 -1280
rect -11945 -1601 -11623 -1600
rect -12364 -1668 -12268 -1652
rect -11352 -1652 -11336 -1228
rect -11272 -1652 -11256 -1228
rect -10340 -1228 -10244 -1212
rect -10933 -1280 -10611 -1279
rect -10933 -1600 -10932 -1280
rect -10612 -1600 -10611 -1280
rect -10933 -1601 -10611 -1600
rect -11352 -1668 -11256 -1652
rect -10340 -1652 -10324 -1228
rect -10260 -1652 -10244 -1228
rect -9328 -1228 -9232 -1212
rect -9921 -1280 -9599 -1279
rect -9921 -1600 -9920 -1280
rect -9600 -1600 -9599 -1280
rect -9921 -1601 -9599 -1600
rect -10340 -1668 -10244 -1652
rect -9328 -1652 -9312 -1228
rect -9248 -1652 -9232 -1228
rect -8316 -1228 -8220 -1212
rect -8909 -1280 -8587 -1279
rect -8909 -1600 -8908 -1280
rect -8588 -1600 -8587 -1280
rect -8909 -1601 -8587 -1600
rect -9328 -1668 -9232 -1652
rect -8316 -1652 -8300 -1228
rect -8236 -1652 -8220 -1228
rect -7304 -1228 -7208 -1212
rect -7897 -1280 -7575 -1279
rect -7897 -1600 -7896 -1280
rect -7576 -1600 -7575 -1280
rect -7897 -1601 -7575 -1600
rect -8316 -1668 -8220 -1652
rect -7304 -1652 -7288 -1228
rect -7224 -1652 -7208 -1228
rect -6292 -1228 -6196 -1212
rect -6885 -1280 -6563 -1279
rect -6885 -1600 -6884 -1280
rect -6564 -1600 -6563 -1280
rect -6885 -1601 -6563 -1600
rect -7304 -1668 -7208 -1652
rect -6292 -1652 -6276 -1228
rect -6212 -1652 -6196 -1228
rect -5280 -1228 -5184 -1212
rect -5873 -1280 -5551 -1279
rect -5873 -1600 -5872 -1280
rect -5552 -1600 -5551 -1280
rect -5873 -1601 -5551 -1600
rect -6292 -1668 -6196 -1652
rect -5280 -1652 -5264 -1228
rect -5200 -1652 -5184 -1228
rect -4268 -1228 -4172 -1212
rect -4861 -1280 -4539 -1279
rect -4861 -1600 -4860 -1280
rect -4540 -1600 -4539 -1280
rect -4861 -1601 -4539 -1600
rect -5280 -1668 -5184 -1652
rect -4268 -1652 -4252 -1228
rect -4188 -1652 -4172 -1228
rect -3256 -1228 -3160 -1212
rect -3849 -1280 -3527 -1279
rect -3849 -1600 -3848 -1280
rect -3528 -1600 -3527 -1280
rect -3849 -1601 -3527 -1600
rect -4268 -1668 -4172 -1652
rect -3256 -1652 -3240 -1228
rect -3176 -1652 -3160 -1228
rect -2244 -1228 -2148 -1212
rect -2837 -1280 -2515 -1279
rect -2837 -1600 -2836 -1280
rect -2516 -1600 -2515 -1280
rect -2837 -1601 -2515 -1600
rect -3256 -1668 -3160 -1652
rect -2244 -1652 -2228 -1228
rect -2164 -1652 -2148 -1228
rect -1232 -1228 -1136 -1212
rect -1825 -1280 -1503 -1279
rect -1825 -1600 -1824 -1280
rect -1504 -1600 -1503 -1280
rect -1825 -1601 -1503 -1600
rect -2244 -1668 -2148 -1652
rect -1232 -1652 -1216 -1228
rect -1152 -1652 -1136 -1228
rect -220 -1228 -124 -1212
rect -813 -1280 -491 -1279
rect -813 -1600 -812 -1280
rect -492 -1600 -491 -1280
rect -813 -1601 -491 -1600
rect -1232 -1668 -1136 -1652
rect -220 -1652 -204 -1228
rect -140 -1652 -124 -1228
rect 792 -1228 888 -1212
rect 199 -1280 521 -1279
rect 199 -1600 200 -1280
rect 520 -1600 521 -1280
rect 199 -1601 521 -1600
rect -220 -1668 -124 -1652
rect 792 -1652 808 -1228
rect 872 -1652 888 -1228
rect 1804 -1228 1900 -1212
rect 1211 -1280 1533 -1279
rect 1211 -1600 1212 -1280
rect 1532 -1600 1533 -1280
rect 1211 -1601 1533 -1600
rect 792 -1668 888 -1652
rect 1804 -1652 1820 -1228
rect 1884 -1652 1900 -1228
rect 2816 -1228 2912 -1212
rect 2223 -1280 2545 -1279
rect 2223 -1600 2224 -1280
rect 2544 -1600 2545 -1280
rect 2223 -1601 2545 -1600
rect 1804 -1668 1900 -1652
rect 2816 -1652 2832 -1228
rect 2896 -1652 2912 -1228
rect 3828 -1228 3924 -1212
rect 3235 -1280 3557 -1279
rect 3235 -1600 3236 -1280
rect 3556 -1600 3557 -1280
rect 3235 -1601 3557 -1600
rect 2816 -1668 2912 -1652
rect 3828 -1652 3844 -1228
rect 3908 -1652 3924 -1228
rect 4840 -1228 4936 -1212
rect 4247 -1280 4569 -1279
rect 4247 -1600 4248 -1280
rect 4568 -1600 4569 -1280
rect 4247 -1601 4569 -1600
rect 3828 -1668 3924 -1652
rect 4840 -1652 4856 -1228
rect 4920 -1652 4936 -1228
rect 5852 -1228 5948 -1212
rect 5259 -1280 5581 -1279
rect 5259 -1600 5260 -1280
rect 5580 -1600 5581 -1280
rect 5259 -1601 5581 -1600
rect 4840 -1668 4936 -1652
rect 5852 -1652 5868 -1228
rect 5932 -1652 5948 -1228
rect 6864 -1228 6960 -1212
rect 6271 -1280 6593 -1279
rect 6271 -1600 6272 -1280
rect 6592 -1600 6593 -1280
rect 6271 -1601 6593 -1600
rect 5852 -1668 5948 -1652
rect 6864 -1652 6880 -1228
rect 6944 -1652 6960 -1228
rect 7876 -1228 7972 -1212
rect 7283 -1280 7605 -1279
rect 7283 -1600 7284 -1280
rect 7604 -1600 7605 -1280
rect 7283 -1601 7605 -1600
rect 6864 -1668 6960 -1652
rect 7876 -1652 7892 -1228
rect 7956 -1652 7972 -1228
rect 8888 -1228 8984 -1212
rect 8295 -1280 8617 -1279
rect 8295 -1600 8296 -1280
rect 8616 -1600 8617 -1280
rect 8295 -1601 8617 -1600
rect 7876 -1668 7972 -1652
rect 8888 -1652 8904 -1228
rect 8968 -1652 8984 -1228
rect 9900 -1228 9996 -1212
rect 9307 -1280 9629 -1279
rect 9307 -1600 9308 -1280
rect 9628 -1600 9629 -1280
rect 9307 -1601 9629 -1600
rect 8888 -1668 8984 -1652
rect 9900 -1652 9916 -1228
rect 9980 -1652 9996 -1228
rect 10912 -1228 11008 -1212
rect 10319 -1280 10641 -1279
rect 10319 -1600 10320 -1280
rect 10640 -1600 10641 -1280
rect 10319 -1601 10641 -1600
rect 9900 -1668 9996 -1652
rect 10912 -1652 10928 -1228
rect 10992 -1652 11008 -1228
rect 11924 -1228 12020 -1212
rect 11331 -1280 11653 -1279
rect 11331 -1600 11332 -1280
rect 11652 -1600 11653 -1280
rect 11331 -1601 11653 -1600
rect 10912 -1668 11008 -1652
rect 11924 -1652 11940 -1228
rect 12004 -1652 12020 -1228
rect 12936 -1228 13032 -1212
rect 12343 -1280 12665 -1279
rect 12343 -1600 12344 -1280
rect 12664 -1600 12665 -1280
rect 12343 -1601 12665 -1600
rect 11924 -1668 12020 -1652
rect 12936 -1652 12952 -1228
rect 13016 -1652 13032 -1228
rect 13948 -1228 14044 -1212
rect 13355 -1280 13677 -1279
rect 13355 -1600 13356 -1280
rect 13676 -1600 13677 -1280
rect 13355 -1601 13677 -1600
rect 12936 -1668 13032 -1652
rect 13948 -1652 13964 -1228
rect 14028 -1652 14044 -1228
rect 14960 -1228 15056 -1212
rect 14367 -1280 14689 -1279
rect 14367 -1600 14368 -1280
rect 14688 -1600 14689 -1280
rect 14367 -1601 14689 -1600
rect 13948 -1668 14044 -1652
rect 14960 -1652 14976 -1228
rect 15040 -1652 15056 -1228
rect 15972 -1228 16068 -1212
rect 15379 -1280 15701 -1279
rect 15379 -1600 15380 -1280
rect 15700 -1600 15701 -1280
rect 15379 -1601 15701 -1600
rect 14960 -1668 15056 -1652
rect 15972 -1652 15988 -1228
rect 16052 -1652 16068 -1228
rect 16984 -1228 17080 -1212
rect 16391 -1280 16713 -1279
rect 16391 -1600 16392 -1280
rect 16712 -1600 16713 -1280
rect 16391 -1601 16713 -1600
rect 15972 -1668 16068 -1652
rect 16984 -1652 17000 -1228
rect 17064 -1652 17080 -1228
rect 16984 -1668 17080 -1652
rect -16412 -1948 -16316 -1932
rect -17005 -2000 -16683 -1999
rect -17005 -2320 -17004 -2000
rect -16684 -2320 -16683 -2000
rect -17005 -2321 -16683 -2320
rect -16412 -2372 -16396 -1948
rect -16332 -2372 -16316 -1948
rect -15400 -1948 -15304 -1932
rect -15993 -2000 -15671 -1999
rect -15993 -2320 -15992 -2000
rect -15672 -2320 -15671 -2000
rect -15993 -2321 -15671 -2320
rect -16412 -2388 -16316 -2372
rect -15400 -2372 -15384 -1948
rect -15320 -2372 -15304 -1948
rect -14388 -1948 -14292 -1932
rect -14981 -2000 -14659 -1999
rect -14981 -2320 -14980 -2000
rect -14660 -2320 -14659 -2000
rect -14981 -2321 -14659 -2320
rect -15400 -2388 -15304 -2372
rect -14388 -2372 -14372 -1948
rect -14308 -2372 -14292 -1948
rect -13376 -1948 -13280 -1932
rect -13969 -2000 -13647 -1999
rect -13969 -2320 -13968 -2000
rect -13648 -2320 -13647 -2000
rect -13969 -2321 -13647 -2320
rect -14388 -2388 -14292 -2372
rect -13376 -2372 -13360 -1948
rect -13296 -2372 -13280 -1948
rect -12364 -1948 -12268 -1932
rect -12957 -2000 -12635 -1999
rect -12957 -2320 -12956 -2000
rect -12636 -2320 -12635 -2000
rect -12957 -2321 -12635 -2320
rect -13376 -2388 -13280 -2372
rect -12364 -2372 -12348 -1948
rect -12284 -2372 -12268 -1948
rect -11352 -1948 -11256 -1932
rect -11945 -2000 -11623 -1999
rect -11945 -2320 -11944 -2000
rect -11624 -2320 -11623 -2000
rect -11945 -2321 -11623 -2320
rect -12364 -2388 -12268 -2372
rect -11352 -2372 -11336 -1948
rect -11272 -2372 -11256 -1948
rect -10340 -1948 -10244 -1932
rect -10933 -2000 -10611 -1999
rect -10933 -2320 -10932 -2000
rect -10612 -2320 -10611 -2000
rect -10933 -2321 -10611 -2320
rect -11352 -2388 -11256 -2372
rect -10340 -2372 -10324 -1948
rect -10260 -2372 -10244 -1948
rect -9328 -1948 -9232 -1932
rect -9921 -2000 -9599 -1999
rect -9921 -2320 -9920 -2000
rect -9600 -2320 -9599 -2000
rect -9921 -2321 -9599 -2320
rect -10340 -2388 -10244 -2372
rect -9328 -2372 -9312 -1948
rect -9248 -2372 -9232 -1948
rect -8316 -1948 -8220 -1932
rect -8909 -2000 -8587 -1999
rect -8909 -2320 -8908 -2000
rect -8588 -2320 -8587 -2000
rect -8909 -2321 -8587 -2320
rect -9328 -2388 -9232 -2372
rect -8316 -2372 -8300 -1948
rect -8236 -2372 -8220 -1948
rect -7304 -1948 -7208 -1932
rect -7897 -2000 -7575 -1999
rect -7897 -2320 -7896 -2000
rect -7576 -2320 -7575 -2000
rect -7897 -2321 -7575 -2320
rect -8316 -2388 -8220 -2372
rect -7304 -2372 -7288 -1948
rect -7224 -2372 -7208 -1948
rect -6292 -1948 -6196 -1932
rect -6885 -2000 -6563 -1999
rect -6885 -2320 -6884 -2000
rect -6564 -2320 -6563 -2000
rect -6885 -2321 -6563 -2320
rect -7304 -2388 -7208 -2372
rect -6292 -2372 -6276 -1948
rect -6212 -2372 -6196 -1948
rect -5280 -1948 -5184 -1932
rect -5873 -2000 -5551 -1999
rect -5873 -2320 -5872 -2000
rect -5552 -2320 -5551 -2000
rect -5873 -2321 -5551 -2320
rect -6292 -2388 -6196 -2372
rect -5280 -2372 -5264 -1948
rect -5200 -2372 -5184 -1948
rect -4268 -1948 -4172 -1932
rect -4861 -2000 -4539 -1999
rect -4861 -2320 -4860 -2000
rect -4540 -2320 -4539 -2000
rect -4861 -2321 -4539 -2320
rect -5280 -2388 -5184 -2372
rect -4268 -2372 -4252 -1948
rect -4188 -2372 -4172 -1948
rect -3256 -1948 -3160 -1932
rect -3849 -2000 -3527 -1999
rect -3849 -2320 -3848 -2000
rect -3528 -2320 -3527 -2000
rect -3849 -2321 -3527 -2320
rect -4268 -2388 -4172 -2372
rect -3256 -2372 -3240 -1948
rect -3176 -2372 -3160 -1948
rect -2244 -1948 -2148 -1932
rect -2837 -2000 -2515 -1999
rect -2837 -2320 -2836 -2000
rect -2516 -2320 -2515 -2000
rect -2837 -2321 -2515 -2320
rect -3256 -2388 -3160 -2372
rect -2244 -2372 -2228 -1948
rect -2164 -2372 -2148 -1948
rect -1232 -1948 -1136 -1932
rect -1825 -2000 -1503 -1999
rect -1825 -2320 -1824 -2000
rect -1504 -2320 -1503 -2000
rect -1825 -2321 -1503 -2320
rect -2244 -2388 -2148 -2372
rect -1232 -2372 -1216 -1948
rect -1152 -2372 -1136 -1948
rect -220 -1948 -124 -1932
rect -813 -2000 -491 -1999
rect -813 -2320 -812 -2000
rect -492 -2320 -491 -2000
rect -813 -2321 -491 -2320
rect -1232 -2388 -1136 -2372
rect -220 -2372 -204 -1948
rect -140 -2372 -124 -1948
rect 792 -1948 888 -1932
rect 199 -2000 521 -1999
rect 199 -2320 200 -2000
rect 520 -2320 521 -2000
rect 199 -2321 521 -2320
rect -220 -2388 -124 -2372
rect 792 -2372 808 -1948
rect 872 -2372 888 -1948
rect 1804 -1948 1900 -1932
rect 1211 -2000 1533 -1999
rect 1211 -2320 1212 -2000
rect 1532 -2320 1533 -2000
rect 1211 -2321 1533 -2320
rect 792 -2388 888 -2372
rect 1804 -2372 1820 -1948
rect 1884 -2372 1900 -1948
rect 2816 -1948 2912 -1932
rect 2223 -2000 2545 -1999
rect 2223 -2320 2224 -2000
rect 2544 -2320 2545 -2000
rect 2223 -2321 2545 -2320
rect 1804 -2388 1900 -2372
rect 2816 -2372 2832 -1948
rect 2896 -2372 2912 -1948
rect 3828 -1948 3924 -1932
rect 3235 -2000 3557 -1999
rect 3235 -2320 3236 -2000
rect 3556 -2320 3557 -2000
rect 3235 -2321 3557 -2320
rect 2816 -2388 2912 -2372
rect 3828 -2372 3844 -1948
rect 3908 -2372 3924 -1948
rect 4840 -1948 4936 -1932
rect 4247 -2000 4569 -1999
rect 4247 -2320 4248 -2000
rect 4568 -2320 4569 -2000
rect 4247 -2321 4569 -2320
rect 3828 -2388 3924 -2372
rect 4840 -2372 4856 -1948
rect 4920 -2372 4936 -1948
rect 5852 -1948 5948 -1932
rect 5259 -2000 5581 -1999
rect 5259 -2320 5260 -2000
rect 5580 -2320 5581 -2000
rect 5259 -2321 5581 -2320
rect 4840 -2388 4936 -2372
rect 5852 -2372 5868 -1948
rect 5932 -2372 5948 -1948
rect 6864 -1948 6960 -1932
rect 6271 -2000 6593 -1999
rect 6271 -2320 6272 -2000
rect 6592 -2320 6593 -2000
rect 6271 -2321 6593 -2320
rect 5852 -2388 5948 -2372
rect 6864 -2372 6880 -1948
rect 6944 -2372 6960 -1948
rect 7876 -1948 7972 -1932
rect 7283 -2000 7605 -1999
rect 7283 -2320 7284 -2000
rect 7604 -2320 7605 -2000
rect 7283 -2321 7605 -2320
rect 6864 -2388 6960 -2372
rect 7876 -2372 7892 -1948
rect 7956 -2372 7972 -1948
rect 8888 -1948 8984 -1932
rect 8295 -2000 8617 -1999
rect 8295 -2320 8296 -2000
rect 8616 -2320 8617 -2000
rect 8295 -2321 8617 -2320
rect 7876 -2388 7972 -2372
rect 8888 -2372 8904 -1948
rect 8968 -2372 8984 -1948
rect 9900 -1948 9996 -1932
rect 9307 -2000 9629 -1999
rect 9307 -2320 9308 -2000
rect 9628 -2320 9629 -2000
rect 9307 -2321 9629 -2320
rect 8888 -2388 8984 -2372
rect 9900 -2372 9916 -1948
rect 9980 -2372 9996 -1948
rect 10912 -1948 11008 -1932
rect 10319 -2000 10641 -1999
rect 10319 -2320 10320 -2000
rect 10640 -2320 10641 -2000
rect 10319 -2321 10641 -2320
rect 9900 -2388 9996 -2372
rect 10912 -2372 10928 -1948
rect 10992 -2372 11008 -1948
rect 11924 -1948 12020 -1932
rect 11331 -2000 11653 -1999
rect 11331 -2320 11332 -2000
rect 11652 -2320 11653 -2000
rect 11331 -2321 11653 -2320
rect 10912 -2388 11008 -2372
rect 11924 -2372 11940 -1948
rect 12004 -2372 12020 -1948
rect 12936 -1948 13032 -1932
rect 12343 -2000 12665 -1999
rect 12343 -2320 12344 -2000
rect 12664 -2320 12665 -2000
rect 12343 -2321 12665 -2320
rect 11924 -2388 12020 -2372
rect 12936 -2372 12952 -1948
rect 13016 -2372 13032 -1948
rect 13948 -1948 14044 -1932
rect 13355 -2000 13677 -1999
rect 13355 -2320 13356 -2000
rect 13676 -2320 13677 -2000
rect 13355 -2321 13677 -2320
rect 12936 -2388 13032 -2372
rect 13948 -2372 13964 -1948
rect 14028 -2372 14044 -1948
rect 14960 -1948 15056 -1932
rect 14367 -2000 14689 -1999
rect 14367 -2320 14368 -2000
rect 14688 -2320 14689 -2000
rect 14367 -2321 14689 -2320
rect 13948 -2388 14044 -2372
rect 14960 -2372 14976 -1948
rect 15040 -2372 15056 -1948
rect 15972 -1948 16068 -1932
rect 15379 -2000 15701 -1999
rect 15379 -2320 15380 -2000
rect 15700 -2320 15701 -2000
rect 15379 -2321 15701 -2320
rect 14960 -2388 15056 -2372
rect 15972 -2372 15988 -1948
rect 16052 -2372 16068 -1948
rect 16984 -1948 17080 -1932
rect 16391 -2000 16713 -1999
rect 16391 -2320 16392 -2000
rect 16712 -2320 16713 -2000
rect 16391 -2321 16713 -2320
rect 15972 -2388 16068 -2372
rect 16984 -2372 17000 -1948
rect 17064 -2372 17080 -1948
rect 16984 -2388 17080 -2372
rect -16412 -2668 -16316 -2652
rect -17005 -2720 -16683 -2719
rect -17005 -3040 -17004 -2720
rect -16684 -3040 -16683 -2720
rect -17005 -3041 -16683 -3040
rect -16412 -3092 -16396 -2668
rect -16332 -3092 -16316 -2668
rect -15400 -2668 -15304 -2652
rect -15993 -2720 -15671 -2719
rect -15993 -3040 -15992 -2720
rect -15672 -3040 -15671 -2720
rect -15993 -3041 -15671 -3040
rect -16412 -3108 -16316 -3092
rect -15400 -3092 -15384 -2668
rect -15320 -3092 -15304 -2668
rect -14388 -2668 -14292 -2652
rect -14981 -2720 -14659 -2719
rect -14981 -3040 -14980 -2720
rect -14660 -3040 -14659 -2720
rect -14981 -3041 -14659 -3040
rect -15400 -3108 -15304 -3092
rect -14388 -3092 -14372 -2668
rect -14308 -3092 -14292 -2668
rect -13376 -2668 -13280 -2652
rect -13969 -2720 -13647 -2719
rect -13969 -3040 -13968 -2720
rect -13648 -3040 -13647 -2720
rect -13969 -3041 -13647 -3040
rect -14388 -3108 -14292 -3092
rect -13376 -3092 -13360 -2668
rect -13296 -3092 -13280 -2668
rect -12364 -2668 -12268 -2652
rect -12957 -2720 -12635 -2719
rect -12957 -3040 -12956 -2720
rect -12636 -3040 -12635 -2720
rect -12957 -3041 -12635 -3040
rect -13376 -3108 -13280 -3092
rect -12364 -3092 -12348 -2668
rect -12284 -3092 -12268 -2668
rect -11352 -2668 -11256 -2652
rect -11945 -2720 -11623 -2719
rect -11945 -3040 -11944 -2720
rect -11624 -3040 -11623 -2720
rect -11945 -3041 -11623 -3040
rect -12364 -3108 -12268 -3092
rect -11352 -3092 -11336 -2668
rect -11272 -3092 -11256 -2668
rect -10340 -2668 -10244 -2652
rect -10933 -2720 -10611 -2719
rect -10933 -3040 -10932 -2720
rect -10612 -3040 -10611 -2720
rect -10933 -3041 -10611 -3040
rect -11352 -3108 -11256 -3092
rect -10340 -3092 -10324 -2668
rect -10260 -3092 -10244 -2668
rect -9328 -2668 -9232 -2652
rect -9921 -2720 -9599 -2719
rect -9921 -3040 -9920 -2720
rect -9600 -3040 -9599 -2720
rect -9921 -3041 -9599 -3040
rect -10340 -3108 -10244 -3092
rect -9328 -3092 -9312 -2668
rect -9248 -3092 -9232 -2668
rect -8316 -2668 -8220 -2652
rect -8909 -2720 -8587 -2719
rect -8909 -3040 -8908 -2720
rect -8588 -3040 -8587 -2720
rect -8909 -3041 -8587 -3040
rect -9328 -3108 -9232 -3092
rect -8316 -3092 -8300 -2668
rect -8236 -3092 -8220 -2668
rect -7304 -2668 -7208 -2652
rect -7897 -2720 -7575 -2719
rect -7897 -3040 -7896 -2720
rect -7576 -3040 -7575 -2720
rect -7897 -3041 -7575 -3040
rect -8316 -3108 -8220 -3092
rect -7304 -3092 -7288 -2668
rect -7224 -3092 -7208 -2668
rect -6292 -2668 -6196 -2652
rect -6885 -2720 -6563 -2719
rect -6885 -3040 -6884 -2720
rect -6564 -3040 -6563 -2720
rect -6885 -3041 -6563 -3040
rect -7304 -3108 -7208 -3092
rect -6292 -3092 -6276 -2668
rect -6212 -3092 -6196 -2668
rect -5280 -2668 -5184 -2652
rect -5873 -2720 -5551 -2719
rect -5873 -3040 -5872 -2720
rect -5552 -3040 -5551 -2720
rect -5873 -3041 -5551 -3040
rect -6292 -3108 -6196 -3092
rect -5280 -3092 -5264 -2668
rect -5200 -3092 -5184 -2668
rect -4268 -2668 -4172 -2652
rect -4861 -2720 -4539 -2719
rect -4861 -3040 -4860 -2720
rect -4540 -3040 -4539 -2720
rect -4861 -3041 -4539 -3040
rect -5280 -3108 -5184 -3092
rect -4268 -3092 -4252 -2668
rect -4188 -3092 -4172 -2668
rect -3256 -2668 -3160 -2652
rect -3849 -2720 -3527 -2719
rect -3849 -3040 -3848 -2720
rect -3528 -3040 -3527 -2720
rect -3849 -3041 -3527 -3040
rect -4268 -3108 -4172 -3092
rect -3256 -3092 -3240 -2668
rect -3176 -3092 -3160 -2668
rect -2244 -2668 -2148 -2652
rect -2837 -2720 -2515 -2719
rect -2837 -3040 -2836 -2720
rect -2516 -3040 -2515 -2720
rect -2837 -3041 -2515 -3040
rect -3256 -3108 -3160 -3092
rect -2244 -3092 -2228 -2668
rect -2164 -3092 -2148 -2668
rect -1232 -2668 -1136 -2652
rect -1825 -2720 -1503 -2719
rect -1825 -3040 -1824 -2720
rect -1504 -3040 -1503 -2720
rect -1825 -3041 -1503 -3040
rect -2244 -3108 -2148 -3092
rect -1232 -3092 -1216 -2668
rect -1152 -3092 -1136 -2668
rect -220 -2668 -124 -2652
rect -813 -2720 -491 -2719
rect -813 -3040 -812 -2720
rect -492 -3040 -491 -2720
rect -813 -3041 -491 -3040
rect -1232 -3108 -1136 -3092
rect -220 -3092 -204 -2668
rect -140 -3092 -124 -2668
rect 792 -2668 888 -2652
rect 199 -2720 521 -2719
rect 199 -3040 200 -2720
rect 520 -3040 521 -2720
rect 199 -3041 521 -3040
rect -220 -3108 -124 -3092
rect 792 -3092 808 -2668
rect 872 -3092 888 -2668
rect 1804 -2668 1900 -2652
rect 1211 -2720 1533 -2719
rect 1211 -3040 1212 -2720
rect 1532 -3040 1533 -2720
rect 1211 -3041 1533 -3040
rect 792 -3108 888 -3092
rect 1804 -3092 1820 -2668
rect 1884 -3092 1900 -2668
rect 2816 -2668 2912 -2652
rect 2223 -2720 2545 -2719
rect 2223 -3040 2224 -2720
rect 2544 -3040 2545 -2720
rect 2223 -3041 2545 -3040
rect 1804 -3108 1900 -3092
rect 2816 -3092 2832 -2668
rect 2896 -3092 2912 -2668
rect 3828 -2668 3924 -2652
rect 3235 -2720 3557 -2719
rect 3235 -3040 3236 -2720
rect 3556 -3040 3557 -2720
rect 3235 -3041 3557 -3040
rect 2816 -3108 2912 -3092
rect 3828 -3092 3844 -2668
rect 3908 -3092 3924 -2668
rect 4840 -2668 4936 -2652
rect 4247 -2720 4569 -2719
rect 4247 -3040 4248 -2720
rect 4568 -3040 4569 -2720
rect 4247 -3041 4569 -3040
rect 3828 -3108 3924 -3092
rect 4840 -3092 4856 -2668
rect 4920 -3092 4936 -2668
rect 5852 -2668 5948 -2652
rect 5259 -2720 5581 -2719
rect 5259 -3040 5260 -2720
rect 5580 -3040 5581 -2720
rect 5259 -3041 5581 -3040
rect 4840 -3108 4936 -3092
rect 5852 -3092 5868 -2668
rect 5932 -3092 5948 -2668
rect 6864 -2668 6960 -2652
rect 6271 -2720 6593 -2719
rect 6271 -3040 6272 -2720
rect 6592 -3040 6593 -2720
rect 6271 -3041 6593 -3040
rect 5852 -3108 5948 -3092
rect 6864 -3092 6880 -2668
rect 6944 -3092 6960 -2668
rect 7876 -2668 7972 -2652
rect 7283 -2720 7605 -2719
rect 7283 -3040 7284 -2720
rect 7604 -3040 7605 -2720
rect 7283 -3041 7605 -3040
rect 6864 -3108 6960 -3092
rect 7876 -3092 7892 -2668
rect 7956 -3092 7972 -2668
rect 8888 -2668 8984 -2652
rect 8295 -2720 8617 -2719
rect 8295 -3040 8296 -2720
rect 8616 -3040 8617 -2720
rect 8295 -3041 8617 -3040
rect 7876 -3108 7972 -3092
rect 8888 -3092 8904 -2668
rect 8968 -3092 8984 -2668
rect 9900 -2668 9996 -2652
rect 9307 -2720 9629 -2719
rect 9307 -3040 9308 -2720
rect 9628 -3040 9629 -2720
rect 9307 -3041 9629 -3040
rect 8888 -3108 8984 -3092
rect 9900 -3092 9916 -2668
rect 9980 -3092 9996 -2668
rect 10912 -2668 11008 -2652
rect 10319 -2720 10641 -2719
rect 10319 -3040 10320 -2720
rect 10640 -3040 10641 -2720
rect 10319 -3041 10641 -3040
rect 9900 -3108 9996 -3092
rect 10912 -3092 10928 -2668
rect 10992 -3092 11008 -2668
rect 11924 -2668 12020 -2652
rect 11331 -2720 11653 -2719
rect 11331 -3040 11332 -2720
rect 11652 -3040 11653 -2720
rect 11331 -3041 11653 -3040
rect 10912 -3108 11008 -3092
rect 11924 -3092 11940 -2668
rect 12004 -3092 12020 -2668
rect 12936 -2668 13032 -2652
rect 12343 -2720 12665 -2719
rect 12343 -3040 12344 -2720
rect 12664 -3040 12665 -2720
rect 12343 -3041 12665 -3040
rect 11924 -3108 12020 -3092
rect 12936 -3092 12952 -2668
rect 13016 -3092 13032 -2668
rect 13948 -2668 14044 -2652
rect 13355 -2720 13677 -2719
rect 13355 -3040 13356 -2720
rect 13676 -3040 13677 -2720
rect 13355 -3041 13677 -3040
rect 12936 -3108 13032 -3092
rect 13948 -3092 13964 -2668
rect 14028 -3092 14044 -2668
rect 14960 -2668 15056 -2652
rect 14367 -2720 14689 -2719
rect 14367 -3040 14368 -2720
rect 14688 -3040 14689 -2720
rect 14367 -3041 14689 -3040
rect 13948 -3108 14044 -3092
rect 14960 -3092 14976 -2668
rect 15040 -3092 15056 -2668
rect 15972 -2668 16068 -2652
rect 15379 -2720 15701 -2719
rect 15379 -3040 15380 -2720
rect 15700 -3040 15701 -2720
rect 15379 -3041 15701 -3040
rect 14960 -3108 15056 -3092
rect 15972 -3092 15988 -2668
rect 16052 -3092 16068 -2668
rect 16984 -2668 17080 -2652
rect 16391 -2720 16713 -2719
rect 16391 -3040 16392 -2720
rect 16712 -3040 16713 -2720
rect 16391 -3041 16713 -3040
rect 15972 -3108 16068 -3092
rect 16984 -3092 17000 -2668
rect 17064 -3092 17080 -2668
rect 16984 -3108 17080 -3092
rect -16412 -3388 -16316 -3372
rect -17005 -3440 -16683 -3439
rect -17005 -3760 -17004 -3440
rect -16684 -3760 -16683 -3440
rect -17005 -3761 -16683 -3760
rect -16412 -3812 -16396 -3388
rect -16332 -3812 -16316 -3388
rect -15400 -3388 -15304 -3372
rect -15993 -3440 -15671 -3439
rect -15993 -3760 -15992 -3440
rect -15672 -3760 -15671 -3440
rect -15993 -3761 -15671 -3760
rect -16412 -3828 -16316 -3812
rect -15400 -3812 -15384 -3388
rect -15320 -3812 -15304 -3388
rect -14388 -3388 -14292 -3372
rect -14981 -3440 -14659 -3439
rect -14981 -3760 -14980 -3440
rect -14660 -3760 -14659 -3440
rect -14981 -3761 -14659 -3760
rect -15400 -3828 -15304 -3812
rect -14388 -3812 -14372 -3388
rect -14308 -3812 -14292 -3388
rect -13376 -3388 -13280 -3372
rect -13969 -3440 -13647 -3439
rect -13969 -3760 -13968 -3440
rect -13648 -3760 -13647 -3440
rect -13969 -3761 -13647 -3760
rect -14388 -3828 -14292 -3812
rect -13376 -3812 -13360 -3388
rect -13296 -3812 -13280 -3388
rect -12364 -3388 -12268 -3372
rect -12957 -3440 -12635 -3439
rect -12957 -3760 -12956 -3440
rect -12636 -3760 -12635 -3440
rect -12957 -3761 -12635 -3760
rect -13376 -3828 -13280 -3812
rect -12364 -3812 -12348 -3388
rect -12284 -3812 -12268 -3388
rect -11352 -3388 -11256 -3372
rect -11945 -3440 -11623 -3439
rect -11945 -3760 -11944 -3440
rect -11624 -3760 -11623 -3440
rect -11945 -3761 -11623 -3760
rect -12364 -3828 -12268 -3812
rect -11352 -3812 -11336 -3388
rect -11272 -3812 -11256 -3388
rect -10340 -3388 -10244 -3372
rect -10933 -3440 -10611 -3439
rect -10933 -3760 -10932 -3440
rect -10612 -3760 -10611 -3440
rect -10933 -3761 -10611 -3760
rect -11352 -3828 -11256 -3812
rect -10340 -3812 -10324 -3388
rect -10260 -3812 -10244 -3388
rect -9328 -3388 -9232 -3372
rect -9921 -3440 -9599 -3439
rect -9921 -3760 -9920 -3440
rect -9600 -3760 -9599 -3440
rect -9921 -3761 -9599 -3760
rect -10340 -3828 -10244 -3812
rect -9328 -3812 -9312 -3388
rect -9248 -3812 -9232 -3388
rect -8316 -3388 -8220 -3372
rect -8909 -3440 -8587 -3439
rect -8909 -3760 -8908 -3440
rect -8588 -3760 -8587 -3440
rect -8909 -3761 -8587 -3760
rect -9328 -3828 -9232 -3812
rect -8316 -3812 -8300 -3388
rect -8236 -3812 -8220 -3388
rect -7304 -3388 -7208 -3372
rect -7897 -3440 -7575 -3439
rect -7897 -3760 -7896 -3440
rect -7576 -3760 -7575 -3440
rect -7897 -3761 -7575 -3760
rect -8316 -3828 -8220 -3812
rect -7304 -3812 -7288 -3388
rect -7224 -3812 -7208 -3388
rect -6292 -3388 -6196 -3372
rect -6885 -3440 -6563 -3439
rect -6885 -3760 -6884 -3440
rect -6564 -3760 -6563 -3440
rect -6885 -3761 -6563 -3760
rect -7304 -3828 -7208 -3812
rect -6292 -3812 -6276 -3388
rect -6212 -3812 -6196 -3388
rect -5280 -3388 -5184 -3372
rect -5873 -3440 -5551 -3439
rect -5873 -3760 -5872 -3440
rect -5552 -3760 -5551 -3440
rect -5873 -3761 -5551 -3760
rect -6292 -3828 -6196 -3812
rect -5280 -3812 -5264 -3388
rect -5200 -3812 -5184 -3388
rect -4268 -3388 -4172 -3372
rect -4861 -3440 -4539 -3439
rect -4861 -3760 -4860 -3440
rect -4540 -3760 -4539 -3440
rect -4861 -3761 -4539 -3760
rect -5280 -3828 -5184 -3812
rect -4268 -3812 -4252 -3388
rect -4188 -3812 -4172 -3388
rect -3256 -3388 -3160 -3372
rect -3849 -3440 -3527 -3439
rect -3849 -3760 -3848 -3440
rect -3528 -3760 -3527 -3440
rect -3849 -3761 -3527 -3760
rect -4268 -3828 -4172 -3812
rect -3256 -3812 -3240 -3388
rect -3176 -3812 -3160 -3388
rect -2244 -3388 -2148 -3372
rect -2837 -3440 -2515 -3439
rect -2837 -3760 -2836 -3440
rect -2516 -3760 -2515 -3440
rect -2837 -3761 -2515 -3760
rect -3256 -3828 -3160 -3812
rect -2244 -3812 -2228 -3388
rect -2164 -3812 -2148 -3388
rect -1232 -3388 -1136 -3372
rect -1825 -3440 -1503 -3439
rect -1825 -3760 -1824 -3440
rect -1504 -3760 -1503 -3440
rect -1825 -3761 -1503 -3760
rect -2244 -3828 -2148 -3812
rect -1232 -3812 -1216 -3388
rect -1152 -3812 -1136 -3388
rect -220 -3388 -124 -3372
rect -813 -3440 -491 -3439
rect -813 -3760 -812 -3440
rect -492 -3760 -491 -3440
rect -813 -3761 -491 -3760
rect -1232 -3828 -1136 -3812
rect -220 -3812 -204 -3388
rect -140 -3812 -124 -3388
rect 792 -3388 888 -3372
rect 199 -3440 521 -3439
rect 199 -3760 200 -3440
rect 520 -3760 521 -3440
rect 199 -3761 521 -3760
rect -220 -3828 -124 -3812
rect 792 -3812 808 -3388
rect 872 -3812 888 -3388
rect 1804 -3388 1900 -3372
rect 1211 -3440 1533 -3439
rect 1211 -3760 1212 -3440
rect 1532 -3760 1533 -3440
rect 1211 -3761 1533 -3760
rect 792 -3828 888 -3812
rect 1804 -3812 1820 -3388
rect 1884 -3812 1900 -3388
rect 2816 -3388 2912 -3372
rect 2223 -3440 2545 -3439
rect 2223 -3760 2224 -3440
rect 2544 -3760 2545 -3440
rect 2223 -3761 2545 -3760
rect 1804 -3828 1900 -3812
rect 2816 -3812 2832 -3388
rect 2896 -3812 2912 -3388
rect 3828 -3388 3924 -3372
rect 3235 -3440 3557 -3439
rect 3235 -3760 3236 -3440
rect 3556 -3760 3557 -3440
rect 3235 -3761 3557 -3760
rect 2816 -3828 2912 -3812
rect 3828 -3812 3844 -3388
rect 3908 -3812 3924 -3388
rect 4840 -3388 4936 -3372
rect 4247 -3440 4569 -3439
rect 4247 -3760 4248 -3440
rect 4568 -3760 4569 -3440
rect 4247 -3761 4569 -3760
rect 3828 -3828 3924 -3812
rect 4840 -3812 4856 -3388
rect 4920 -3812 4936 -3388
rect 5852 -3388 5948 -3372
rect 5259 -3440 5581 -3439
rect 5259 -3760 5260 -3440
rect 5580 -3760 5581 -3440
rect 5259 -3761 5581 -3760
rect 4840 -3828 4936 -3812
rect 5852 -3812 5868 -3388
rect 5932 -3812 5948 -3388
rect 6864 -3388 6960 -3372
rect 6271 -3440 6593 -3439
rect 6271 -3760 6272 -3440
rect 6592 -3760 6593 -3440
rect 6271 -3761 6593 -3760
rect 5852 -3828 5948 -3812
rect 6864 -3812 6880 -3388
rect 6944 -3812 6960 -3388
rect 7876 -3388 7972 -3372
rect 7283 -3440 7605 -3439
rect 7283 -3760 7284 -3440
rect 7604 -3760 7605 -3440
rect 7283 -3761 7605 -3760
rect 6864 -3828 6960 -3812
rect 7876 -3812 7892 -3388
rect 7956 -3812 7972 -3388
rect 8888 -3388 8984 -3372
rect 8295 -3440 8617 -3439
rect 8295 -3760 8296 -3440
rect 8616 -3760 8617 -3440
rect 8295 -3761 8617 -3760
rect 7876 -3828 7972 -3812
rect 8888 -3812 8904 -3388
rect 8968 -3812 8984 -3388
rect 9900 -3388 9996 -3372
rect 9307 -3440 9629 -3439
rect 9307 -3760 9308 -3440
rect 9628 -3760 9629 -3440
rect 9307 -3761 9629 -3760
rect 8888 -3828 8984 -3812
rect 9900 -3812 9916 -3388
rect 9980 -3812 9996 -3388
rect 10912 -3388 11008 -3372
rect 10319 -3440 10641 -3439
rect 10319 -3760 10320 -3440
rect 10640 -3760 10641 -3440
rect 10319 -3761 10641 -3760
rect 9900 -3828 9996 -3812
rect 10912 -3812 10928 -3388
rect 10992 -3812 11008 -3388
rect 11924 -3388 12020 -3372
rect 11331 -3440 11653 -3439
rect 11331 -3760 11332 -3440
rect 11652 -3760 11653 -3440
rect 11331 -3761 11653 -3760
rect 10912 -3828 11008 -3812
rect 11924 -3812 11940 -3388
rect 12004 -3812 12020 -3388
rect 12936 -3388 13032 -3372
rect 12343 -3440 12665 -3439
rect 12343 -3760 12344 -3440
rect 12664 -3760 12665 -3440
rect 12343 -3761 12665 -3760
rect 11924 -3828 12020 -3812
rect 12936 -3812 12952 -3388
rect 13016 -3812 13032 -3388
rect 13948 -3388 14044 -3372
rect 13355 -3440 13677 -3439
rect 13355 -3760 13356 -3440
rect 13676 -3760 13677 -3440
rect 13355 -3761 13677 -3760
rect 12936 -3828 13032 -3812
rect 13948 -3812 13964 -3388
rect 14028 -3812 14044 -3388
rect 14960 -3388 15056 -3372
rect 14367 -3440 14689 -3439
rect 14367 -3760 14368 -3440
rect 14688 -3760 14689 -3440
rect 14367 -3761 14689 -3760
rect 13948 -3828 14044 -3812
rect 14960 -3812 14976 -3388
rect 15040 -3812 15056 -3388
rect 15972 -3388 16068 -3372
rect 15379 -3440 15701 -3439
rect 15379 -3760 15380 -3440
rect 15700 -3760 15701 -3440
rect 15379 -3761 15701 -3760
rect 14960 -3828 15056 -3812
rect 15972 -3812 15988 -3388
rect 16052 -3812 16068 -3388
rect 16984 -3388 17080 -3372
rect 16391 -3440 16713 -3439
rect 16391 -3760 16392 -3440
rect 16712 -3760 16713 -3440
rect 16391 -3761 16713 -3760
rect 15972 -3828 16068 -3812
rect 16984 -3812 17000 -3388
rect 17064 -3812 17080 -3388
rect 16984 -3828 17080 -3812
rect -16412 -4108 -16316 -4092
rect -17005 -4160 -16683 -4159
rect -17005 -4480 -17004 -4160
rect -16684 -4480 -16683 -4160
rect -17005 -4481 -16683 -4480
rect -16412 -4532 -16396 -4108
rect -16332 -4532 -16316 -4108
rect -15400 -4108 -15304 -4092
rect -15993 -4160 -15671 -4159
rect -15993 -4480 -15992 -4160
rect -15672 -4480 -15671 -4160
rect -15993 -4481 -15671 -4480
rect -16412 -4548 -16316 -4532
rect -15400 -4532 -15384 -4108
rect -15320 -4532 -15304 -4108
rect -14388 -4108 -14292 -4092
rect -14981 -4160 -14659 -4159
rect -14981 -4480 -14980 -4160
rect -14660 -4480 -14659 -4160
rect -14981 -4481 -14659 -4480
rect -15400 -4548 -15304 -4532
rect -14388 -4532 -14372 -4108
rect -14308 -4532 -14292 -4108
rect -13376 -4108 -13280 -4092
rect -13969 -4160 -13647 -4159
rect -13969 -4480 -13968 -4160
rect -13648 -4480 -13647 -4160
rect -13969 -4481 -13647 -4480
rect -14388 -4548 -14292 -4532
rect -13376 -4532 -13360 -4108
rect -13296 -4532 -13280 -4108
rect -12364 -4108 -12268 -4092
rect -12957 -4160 -12635 -4159
rect -12957 -4480 -12956 -4160
rect -12636 -4480 -12635 -4160
rect -12957 -4481 -12635 -4480
rect -13376 -4548 -13280 -4532
rect -12364 -4532 -12348 -4108
rect -12284 -4532 -12268 -4108
rect -11352 -4108 -11256 -4092
rect -11945 -4160 -11623 -4159
rect -11945 -4480 -11944 -4160
rect -11624 -4480 -11623 -4160
rect -11945 -4481 -11623 -4480
rect -12364 -4548 -12268 -4532
rect -11352 -4532 -11336 -4108
rect -11272 -4532 -11256 -4108
rect -10340 -4108 -10244 -4092
rect -10933 -4160 -10611 -4159
rect -10933 -4480 -10932 -4160
rect -10612 -4480 -10611 -4160
rect -10933 -4481 -10611 -4480
rect -11352 -4548 -11256 -4532
rect -10340 -4532 -10324 -4108
rect -10260 -4532 -10244 -4108
rect -9328 -4108 -9232 -4092
rect -9921 -4160 -9599 -4159
rect -9921 -4480 -9920 -4160
rect -9600 -4480 -9599 -4160
rect -9921 -4481 -9599 -4480
rect -10340 -4548 -10244 -4532
rect -9328 -4532 -9312 -4108
rect -9248 -4532 -9232 -4108
rect -8316 -4108 -8220 -4092
rect -8909 -4160 -8587 -4159
rect -8909 -4480 -8908 -4160
rect -8588 -4480 -8587 -4160
rect -8909 -4481 -8587 -4480
rect -9328 -4548 -9232 -4532
rect -8316 -4532 -8300 -4108
rect -8236 -4532 -8220 -4108
rect -7304 -4108 -7208 -4092
rect -7897 -4160 -7575 -4159
rect -7897 -4480 -7896 -4160
rect -7576 -4480 -7575 -4160
rect -7897 -4481 -7575 -4480
rect -8316 -4548 -8220 -4532
rect -7304 -4532 -7288 -4108
rect -7224 -4532 -7208 -4108
rect -6292 -4108 -6196 -4092
rect -6885 -4160 -6563 -4159
rect -6885 -4480 -6884 -4160
rect -6564 -4480 -6563 -4160
rect -6885 -4481 -6563 -4480
rect -7304 -4548 -7208 -4532
rect -6292 -4532 -6276 -4108
rect -6212 -4532 -6196 -4108
rect -5280 -4108 -5184 -4092
rect -5873 -4160 -5551 -4159
rect -5873 -4480 -5872 -4160
rect -5552 -4480 -5551 -4160
rect -5873 -4481 -5551 -4480
rect -6292 -4548 -6196 -4532
rect -5280 -4532 -5264 -4108
rect -5200 -4532 -5184 -4108
rect -4268 -4108 -4172 -4092
rect -4861 -4160 -4539 -4159
rect -4861 -4480 -4860 -4160
rect -4540 -4480 -4539 -4160
rect -4861 -4481 -4539 -4480
rect -5280 -4548 -5184 -4532
rect -4268 -4532 -4252 -4108
rect -4188 -4532 -4172 -4108
rect -3256 -4108 -3160 -4092
rect -3849 -4160 -3527 -4159
rect -3849 -4480 -3848 -4160
rect -3528 -4480 -3527 -4160
rect -3849 -4481 -3527 -4480
rect -4268 -4548 -4172 -4532
rect -3256 -4532 -3240 -4108
rect -3176 -4532 -3160 -4108
rect -2244 -4108 -2148 -4092
rect -2837 -4160 -2515 -4159
rect -2837 -4480 -2836 -4160
rect -2516 -4480 -2515 -4160
rect -2837 -4481 -2515 -4480
rect -3256 -4548 -3160 -4532
rect -2244 -4532 -2228 -4108
rect -2164 -4532 -2148 -4108
rect -1232 -4108 -1136 -4092
rect -1825 -4160 -1503 -4159
rect -1825 -4480 -1824 -4160
rect -1504 -4480 -1503 -4160
rect -1825 -4481 -1503 -4480
rect -2244 -4548 -2148 -4532
rect -1232 -4532 -1216 -4108
rect -1152 -4532 -1136 -4108
rect -220 -4108 -124 -4092
rect -813 -4160 -491 -4159
rect -813 -4480 -812 -4160
rect -492 -4480 -491 -4160
rect -813 -4481 -491 -4480
rect -1232 -4548 -1136 -4532
rect -220 -4532 -204 -4108
rect -140 -4532 -124 -4108
rect 792 -4108 888 -4092
rect 199 -4160 521 -4159
rect 199 -4480 200 -4160
rect 520 -4480 521 -4160
rect 199 -4481 521 -4480
rect -220 -4548 -124 -4532
rect 792 -4532 808 -4108
rect 872 -4532 888 -4108
rect 1804 -4108 1900 -4092
rect 1211 -4160 1533 -4159
rect 1211 -4480 1212 -4160
rect 1532 -4480 1533 -4160
rect 1211 -4481 1533 -4480
rect 792 -4548 888 -4532
rect 1804 -4532 1820 -4108
rect 1884 -4532 1900 -4108
rect 2816 -4108 2912 -4092
rect 2223 -4160 2545 -4159
rect 2223 -4480 2224 -4160
rect 2544 -4480 2545 -4160
rect 2223 -4481 2545 -4480
rect 1804 -4548 1900 -4532
rect 2816 -4532 2832 -4108
rect 2896 -4532 2912 -4108
rect 3828 -4108 3924 -4092
rect 3235 -4160 3557 -4159
rect 3235 -4480 3236 -4160
rect 3556 -4480 3557 -4160
rect 3235 -4481 3557 -4480
rect 2816 -4548 2912 -4532
rect 3828 -4532 3844 -4108
rect 3908 -4532 3924 -4108
rect 4840 -4108 4936 -4092
rect 4247 -4160 4569 -4159
rect 4247 -4480 4248 -4160
rect 4568 -4480 4569 -4160
rect 4247 -4481 4569 -4480
rect 3828 -4548 3924 -4532
rect 4840 -4532 4856 -4108
rect 4920 -4532 4936 -4108
rect 5852 -4108 5948 -4092
rect 5259 -4160 5581 -4159
rect 5259 -4480 5260 -4160
rect 5580 -4480 5581 -4160
rect 5259 -4481 5581 -4480
rect 4840 -4548 4936 -4532
rect 5852 -4532 5868 -4108
rect 5932 -4532 5948 -4108
rect 6864 -4108 6960 -4092
rect 6271 -4160 6593 -4159
rect 6271 -4480 6272 -4160
rect 6592 -4480 6593 -4160
rect 6271 -4481 6593 -4480
rect 5852 -4548 5948 -4532
rect 6864 -4532 6880 -4108
rect 6944 -4532 6960 -4108
rect 7876 -4108 7972 -4092
rect 7283 -4160 7605 -4159
rect 7283 -4480 7284 -4160
rect 7604 -4480 7605 -4160
rect 7283 -4481 7605 -4480
rect 6864 -4548 6960 -4532
rect 7876 -4532 7892 -4108
rect 7956 -4532 7972 -4108
rect 8888 -4108 8984 -4092
rect 8295 -4160 8617 -4159
rect 8295 -4480 8296 -4160
rect 8616 -4480 8617 -4160
rect 8295 -4481 8617 -4480
rect 7876 -4548 7972 -4532
rect 8888 -4532 8904 -4108
rect 8968 -4532 8984 -4108
rect 9900 -4108 9996 -4092
rect 9307 -4160 9629 -4159
rect 9307 -4480 9308 -4160
rect 9628 -4480 9629 -4160
rect 9307 -4481 9629 -4480
rect 8888 -4548 8984 -4532
rect 9900 -4532 9916 -4108
rect 9980 -4532 9996 -4108
rect 10912 -4108 11008 -4092
rect 10319 -4160 10641 -4159
rect 10319 -4480 10320 -4160
rect 10640 -4480 10641 -4160
rect 10319 -4481 10641 -4480
rect 9900 -4548 9996 -4532
rect 10912 -4532 10928 -4108
rect 10992 -4532 11008 -4108
rect 11924 -4108 12020 -4092
rect 11331 -4160 11653 -4159
rect 11331 -4480 11332 -4160
rect 11652 -4480 11653 -4160
rect 11331 -4481 11653 -4480
rect 10912 -4548 11008 -4532
rect 11924 -4532 11940 -4108
rect 12004 -4532 12020 -4108
rect 12936 -4108 13032 -4092
rect 12343 -4160 12665 -4159
rect 12343 -4480 12344 -4160
rect 12664 -4480 12665 -4160
rect 12343 -4481 12665 -4480
rect 11924 -4548 12020 -4532
rect 12936 -4532 12952 -4108
rect 13016 -4532 13032 -4108
rect 13948 -4108 14044 -4092
rect 13355 -4160 13677 -4159
rect 13355 -4480 13356 -4160
rect 13676 -4480 13677 -4160
rect 13355 -4481 13677 -4480
rect 12936 -4548 13032 -4532
rect 13948 -4532 13964 -4108
rect 14028 -4532 14044 -4108
rect 14960 -4108 15056 -4092
rect 14367 -4160 14689 -4159
rect 14367 -4480 14368 -4160
rect 14688 -4480 14689 -4160
rect 14367 -4481 14689 -4480
rect 13948 -4548 14044 -4532
rect 14960 -4532 14976 -4108
rect 15040 -4532 15056 -4108
rect 15972 -4108 16068 -4092
rect 15379 -4160 15701 -4159
rect 15379 -4480 15380 -4160
rect 15700 -4480 15701 -4160
rect 15379 -4481 15701 -4480
rect 14960 -4548 15056 -4532
rect 15972 -4532 15988 -4108
rect 16052 -4532 16068 -4108
rect 16984 -4108 17080 -4092
rect 16391 -4160 16713 -4159
rect 16391 -4480 16392 -4160
rect 16712 -4480 16713 -4160
rect 16391 -4481 16713 -4480
rect 15972 -4548 16068 -4532
rect 16984 -4532 17000 -4108
rect 17064 -4532 17080 -4108
rect 16984 -4548 17080 -4532
rect -16412 -4828 -16316 -4812
rect -17005 -4880 -16683 -4879
rect -17005 -5200 -17004 -4880
rect -16684 -5200 -16683 -4880
rect -17005 -5201 -16683 -5200
rect -16412 -5252 -16396 -4828
rect -16332 -5252 -16316 -4828
rect -15400 -4828 -15304 -4812
rect -15993 -4880 -15671 -4879
rect -15993 -5200 -15992 -4880
rect -15672 -5200 -15671 -4880
rect -15993 -5201 -15671 -5200
rect -16412 -5268 -16316 -5252
rect -15400 -5252 -15384 -4828
rect -15320 -5252 -15304 -4828
rect -14388 -4828 -14292 -4812
rect -14981 -4880 -14659 -4879
rect -14981 -5200 -14980 -4880
rect -14660 -5200 -14659 -4880
rect -14981 -5201 -14659 -5200
rect -15400 -5268 -15304 -5252
rect -14388 -5252 -14372 -4828
rect -14308 -5252 -14292 -4828
rect -13376 -4828 -13280 -4812
rect -13969 -4880 -13647 -4879
rect -13969 -5200 -13968 -4880
rect -13648 -5200 -13647 -4880
rect -13969 -5201 -13647 -5200
rect -14388 -5268 -14292 -5252
rect -13376 -5252 -13360 -4828
rect -13296 -5252 -13280 -4828
rect -12364 -4828 -12268 -4812
rect -12957 -4880 -12635 -4879
rect -12957 -5200 -12956 -4880
rect -12636 -5200 -12635 -4880
rect -12957 -5201 -12635 -5200
rect -13376 -5268 -13280 -5252
rect -12364 -5252 -12348 -4828
rect -12284 -5252 -12268 -4828
rect -11352 -4828 -11256 -4812
rect -11945 -4880 -11623 -4879
rect -11945 -5200 -11944 -4880
rect -11624 -5200 -11623 -4880
rect -11945 -5201 -11623 -5200
rect -12364 -5268 -12268 -5252
rect -11352 -5252 -11336 -4828
rect -11272 -5252 -11256 -4828
rect -10340 -4828 -10244 -4812
rect -10933 -4880 -10611 -4879
rect -10933 -5200 -10932 -4880
rect -10612 -5200 -10611 -4880
rect -10933 -5201 -10611 -5200
rect -11352 -5268 -11256 -5252
rect -10340 -5252 -10324 -4828
rect -10260 -5252 -10244 -4828
rect -9328 -4828 -9232 -4812
rect -9921 -4880 -9599 -4879
rect -9921 -5200 -9920 -4880
rect -9600 -5200 -9599 -4880
rect -9921 -5201 -9599 -5200
rect -10340 -5268 -10244 -5252
rect -9328 -5252 -9312 -4828
rect -9248 -5252 -9232 -4828
rect -8316 -4828 -8220 -4812
rect -8909 -4880 -8587 -4879
rect -8909 -5200 -8908 -4880
rect -8588 -5200 -8587 -4880
rect -8909 -5201 -8587 -5200
rect -9328 -5268 -9232 -5252
rect -8316 -5252 -8300 -4828
rect -8236 -5252 -8220 -4828
rect -7304 -4828 -7208 -4812
rect -7897 -4880 -7575 -4879
rect -7897 -5200 -7896 -4880
rect -7576 -5200 -7575 -4880
rect -7897 -5201 -7575 -5200
rect -8316 -5268 -8220 -5252
rect -7304 -5252 -7288 -4828
rect -7224 -5252 -7208 -4828
rect -6292 -4828 -6196 -4812
rect -6885 -4880 -6563 -4879
rect -6885 -5200 -6884 -4880
rect -6564 -5200 -6563 -4880
rect -6885 -5201 -6563 -5200
rect -7304 -5268 -7208 -5252
rect -6292 -5252 -6276 -4828
rect -6212 -5252 -6196 -4828
rect -5280 -4828 -5184 -4812
rect -5873 -4880 -5551 -4879
rect -5873 -5200 -5872 -4880
rect -5552 -5200 -5551 -4880
rect -5873 -5201 -5551 -5200
rect -6292 -5268 -6196 -5252
rect -5280 -5252 -5264 -4828
rect -5200 -5252 -5184 -4828
rect -4268 -4828 -4172 -4812
rect -4861 -4880 -4539 -4879
rect -4861 -5200 -4860 -4880
rect -4540 -5200 -4539 -4880
rect -4861 -5201 -4539 -5200
rect -5280 -5268 -5184 -5252
rect -4268 -5252 -4252 -4828
rect -4188 -5252 -4172 -4828
rect -3256 -4828 -3160 -4812
rect -3849 -4880 -3527 -4879
rect -3849 -5200 -3848 -4880
rect -3528 -5200 -3527 -4880
rect -3849 -5201 -3527 -5200
rect -4268 -5268 -4172 -5252
rect -3256 -5252 -3240 -4828
rect -3176 -5252 -3160 -4828
rect -2244 -4828 -2148 -4812
rect -2837 -4880 -2515 -4879
rect -2837 -5200 -2836 -4880
rect -2516 -5200 -2515 -4880
rect -2837 -5201 -2515 -5200
rect -3256 -5268 -3160 -5252
rect -2244 -5252 -2228 -4828
rect -2164 -5252 -2148 -4828
rect -1232 -4828 -1136 -4812
rect -1825 -4880 -1503 -4879
rect -1825 -5200 -1824 -4880
rect -1504 -5200 -1503 -4880
rect -1825 -5201 -1503 -5200
rect -2244 -5268 -2148 -5252
rect -1232 -5252 -1216 -4828
rect -1152 -5252 -1136 -4828
rect -220 -4828 -124 -4812
rect -813 -4880 -491 -4879
rect -813 -5200 -812 -4880
rect -492 -5200 -491 -4880
rect -813 -5201 -491 -5200
rect -1232 -5268 -1136 -5252
rect -220 -5252 -204 -4828
rect -140 -5252 -124 -4828
rect 792 -4828 888 -4812
rect 199 -4880 521 -4879
rect 199 -5200 200 -4880
rect 520 -5200 521 -4880
rect 199 -5201 521 -5200
rect -220 -5268 -124 -5252
rect 792 -5252 808 -4828
rect 872 -5252 888 -4828
rect 1804 -4828 1900 -4812
rect 1211 -4880 1533 -4879
rect 1211 -5200 1212 -4880
rect 1532 -5200 1533 -4880
rect 1211 -5201 1533 -5200
rect 792 -5268 888 -5252
rect 1804 -5252 1820 -4828
rect 1884 -5252 1900 -4828
rect 2816 -4828 2912 -4812
rect 2223 -4880 2545 -4879
rect 2223 -5200 2224 -4880
rect 2544 -5200 2545 -4880
rect 2223 -5201 2545 -5200
rect 1804 -5268 1900 -5252
rect 2816 -5252 2832 -4828
rect 2896 -5252 2912 -4828
rect 3828 -4828 3924 -4812
rect 3235 -4880 3557 -4879
rect 3235 -5200 3236 -4880
rect 3556 -5200 3557 -4880
rect 3235 -5201 3557 -5200
rect 2816 -5268 2912 -5252
rect 3828 -5252 3844 -4828
rect 3908 -5252 3924 -4828
rect 4840 -4828 4936 -4812
rect 4247 -4880 4569 -4879
rect 4247 -5200 4248 -4880
rect 4568 -5200 4569 -4880
rect 4247 -5201 4569 -5200
rect 3828 -5268 3924 -5252
rect 4840 -5252 4856 -4828
rect 4920 -5252 4936 -4828
rect 5852 -4828 5948 -4812
rect 5259 -4880 5581 -4879
rect 5259 -5200 5260 -4880
rect 5580 -5200 5581 -4880
rect 5259 -5201 5581 -5200
rect 4840 -5268 4936 -5252
rect 5852 -5252 5868 -4828
rect 5932 -5252 5948 -4828
rect 6864 -4828 6960 -4812
rect 6271 -4880 6593 -4879
rect 6271 -5200 6272 -4880
rect 6592 -5200 6593 -4880
rect 6271 -5201 6593 -5200
rect 5852 -5268 5948 -5252
rect 6864 -5252 6880 -4828
rect 6944 -5252 6960 -4828
rect 7876 -4828 7972 -4812
rect 7283 -4880 7605 -4879
rect 7283 -5200 7284 -4880
rect 7604 -5200 7605 -4880
rect 7283 -5201 7605 -5200
rect 6864 -5268 6960 -5252
rect 7876 -5252 7892 -4828
rect 7956 -5252 7972 -4828
rect 8888 -4828 8984 -4812
rect 8295 -4880 8617 -4879
rect 8295 -5200 8296 -4880
rect 8616 -5200 8617 -4880
rect 8295 -5201 8617 -5200
rect 7876 -5268 7972 -5252
rect 8888 -5252 8904 -4828
rect 8968 -5252 8984 -4828
rect 9900 -4828 9996 -4812
rect 9307 -4880 9629 -4879
rect 9307 -5200 9308 -4880
rect 9628 -5200 9629 -4880
rect 9307 -5201 9629 -5200
rect 8888 -5268 8984 -5252
rect 9900 -5252 9916 -4828
rect 9980 -5252 9996 -4828
rect 10912 -4828 11008 -4812
rect 10319 -4880 10641 -4879
rect 10319 -5200 10320 -4880
rect 10640 -5200 10641 -4880
rect 10319 -5201 10641 -5200
rect 9900 -5268 9996 -5252
rect 10912 -5252 10928 -4828
rect 10992 -5252 11008 -4828
rect 11924 -4828 12020 -4812
rect 11331 -4880 11653 -4879
rect 11331 -5200 11332 -4880
rect 11652 -5200 11653 -4880
rect 11331 -5201 11653 -5200
rect 10912 -5268 11008 -5252
rect 11924 -5252 11940 -4828
rect 12004 -5252 12020 -4828
rect 12936 -4828 13032 -4812
rect 12343 -4880 12665 -4879
rect 12343 -5200 12344 -4880
rect 12664 -5200 12665 -4880
rect 12343 -5201 12665 -5200
rect 11924 -5268 12020 -5252
rect 12936 -5252 12952 -4828
rect 13016 -5252 13032 -4828
rect 13948 -4828 14044 -4812
rect 13355 -4880 13677 -4879
rect 13355 -5200 13356 -4880
rect 13676 -5200 13677 -4880
rect 13355 -5201 13677 -5200
rect 12936 -5268 13032 -5252
rect 13948 -5252 13964 -4828
rect 14028 -5252 14044 -4828
rect 14960 -4828 15056 -4812
rect 14367 -4880 14689 -4879
rect 14367 -5200 14368 -4880
rect 14688 -5200 14689 -4880
rect 14367 -5201 14689 -5200
rect 13948 -5268 14044 -5252
rect 14960 -5252 14976 -4828
rect 15040 -5252 15056 -4828
rect 15972 -4828 16068 -4812
rect 15379 -4880 15701 -4879
rect 15379 -5200 15380 -4880
rect 15700 -5200 15701 -4880
rect 15379 -5201 15701 -5200
rect 14960 -5268 15056 -5252
rect 15972 -5252 15988 -4828
rect 16052 -5252 16068 -4828
rect 16984 -4828 17080 -4812
rect 16391 -4880 16713 -4879
rect 16391 -5200 16392 -4880
rect 16712 -5200 16713 -4880
rect 16391 -5201 16713 -5200
rect 15972 -5268 16068 -5252
rect 16984 -5252 17000 -4828
rect 17064 -5252 17080 -4828
rect 16984 -5268 17080 -5252
rect -16412 -5548 -16316 -5532
rect -17005 -5600 -16683 -5599
rect -17005 -5920 -17004 -5600
rect -16684 -5920 -16683 -5600
rect -17005 -5921 -16683 -5920
rect -16412 -5972 -16396 -5548
rect -16332 -5972 -16316 -5548
rect -15400 -5548 -15304 -5532
rect -15993 -5600 -15671 -5599
rect -15993 -5920 -15992 -5600
rect -15672 -5920 -15671 -5600
rect -15993 -5921 -15671 -5920
rect -16412 -5988 -16316 -5972
rect -15400 -5972 -15384 -5548
rect -15320 -5972 -15304 -5548
rect -14388 -5548 -14292 -5532
rect -14981 -5600 -14659 -5599
rect -14981 -5920 -14980 -5600
rect -14660 -5920 -14659 -5600
rect -14981 -5921 -14659 -5920
rect -15400 -5988 -15304 -5972
rect -14388 -5972 -14372 -5548
rect -14308 -5972 -14292 -5548
rect -13376 -5548 -13280 -5532
rect -13969 -5600 -13647 -5599
rect -13969 -5920 -13968 -5600
rect -13648 -5920 -13647 -5600
rect -13969 -5921 -13647 -5920
rect -14388 -5988 -14292 -5972
rect -13376 -5972 -13360 -5548
rect -13296 -5972 -13280 -5548
rect -12364 -5548 -12268 -5532
rect -12957 -5600 -12635 -5599
rect -12957 -5920 -12956 -5600
rect -12636 -5920 -12635 -5600
rect -12957 -5921 -12635 -5920
rect -13376 -5988 -13280 -5972
rect -12364 -5972 -12348 -5548
rect -12284 -5972 -12268 -5548
rect -11352 -5548 -11256 -5532
rect -11945 -5600 -11623 -5599
rect -11945 -5920 -11944 -5600
rect -11624 -5920 -11623 -5600
rect -11945 -5921 -11623 -5920
rect -12364 -5988 -12268 -5972
rect -11352 -5972 -11336 -5548
rect -11272 -5972 -11256 -5548
rect -10340 -5548 -10244 -5532
rect -10933 -5600 -10611 -5599
rect -10933 -5920 -10932 -5600
rect -10612 -5920 -10611 -5600
rect -10933 -5921 -10611 -5920
rect -11352 -5988 -11256 -5972
rect -10340 -5972 -10324 -5548
rect -10260 -5972 -10244 -5548
rect -9328 -5548 -9232 -5532
rect -9921 -5600 -9599 -5599
rect -9921 -5920 -9920 -5600
rect -9600 -5920 -9599 -5600
rect -9921 -5921 -9599 -5920
rect -10340 -5988 -10244 -5972
rect -9328 -5972 -9312 -5548
rect -9248 -5972 -9232 -5548
rect -8316 -5548 -8220 -5532
rect -8909 -5600 -8587 -5599
rect -8909 -5920 -8908 -5600
rect -8588 -5920 -8587 -5600
rect -8909 -5921 -8587 -5920
rect -9328 -5988 -9232 -5972
rect -8316 -5972 -8300 -5548
rect -8236 -5972 -8220 -5548
rect -7304 -5548 -7208 -5532
rect -7897 -5600 -7575 -5599
rect -7897 -5920 -7896 -5600
rect -7576 -5920 -7575 -5600
rect -7897 -5921 -7575 -5920
rect -8316 -5988 -8220 -5972
rect -7304 -5972 -7288 -5548
rect -7224 -5972 -7208 -5548
rect -6292 -5548 -6196 -5532
rect -6885 -5600 -6563 -5599
rect -6885 -5920 -6884 -5600
rect -6564 -5920 -6563 -5600
rect -6885 -5921 -6563 -5920
rect -7304 -5988 -7208 -5972
rect -6292 -5972 -6276 -5548
rect -6212 -5972 -6196 -5548
rect -5280 -5548 -5184 -5532
rect -5873 -5600 -5551 -5599
rect -5873 -5920 -5872 -5600
rect -5552 -5920 -5551 -5600
rect -5873 -5921 -5551 -5920
rect -6292 -5988 -6196 -5972
rect -5280 -5972 -5264 -5548
rect -5200 -5972 -5184 -5548
rect -4268 -5548 -4172 -5532
rect -4861 -5600 -4539 -5599
rect -4861 -5920 -4860 -5600
rect -4540 -5920 -4539 -5600
rect -4861 -5921 -4539 -5920
rect -5280 -5988 -5184 -5972
rect -4268 -5972 -4252 -5548
rect -4188 -5972 -4172 -5548
rect -3256 -5548 -3160 -5532
rect -3849 -5600 -3527 -5599
rect -3849 -5920 -3848 -5600
rect -3528 -5920 -3527 -5600
rect -3849 -5921 -3527 -5920
rect -4268 -5988 -4172 -5972
rect -3256 -5972 -3240 -5548
rect -3176 -5972 -3160 -5548
rect -2244 -5548 -2148 -5532
rect -2837 -5600 -2515 -5599
rect -2837 -5920 -2836 -5600
rect -2516 -5920 -2515 -5600
rect -2837 -5921 -2515 -5920
rect -3256 -5988 -3160 -5972
rect -2244 -5972 -2228 -5548
rect -2164 -5972 -2148 -5548
rect -1232 -5548 -1136 -5532
rect -1825 -5600 -1503 -5599
rect -1825 -5920 -1824 -5600
rect -1504 -5920 -1503 -5600
rect -1825 -5921 -1503 -5920
rect -2244 -5988 -2148 -5972
rect -1232 -5972 -1216 -5548
rect -1152 -5972 -1136 -5548
rect -220 -5548 -124 -5532
rect -813 -5600 -491 -5599
rect -813 -5920 -812 -5600
rect -492 -5920 -491 -5600
rect -813 -5921 -491 -5920
rect -1232 -5988 -1136 -5972
rect -220 -5972 -204 -5548
rect -140 -5972 -124 -5548
rect 792 -5548 888 -5532
rect 199 -5600 521 -5599
rect 199 -5920 200 -5600
rect 520 -5920 521 -5600
rect 199 -5921 521 -5920
rect -220 -5988 -124 -5972
rect 792 -5972 808 -5548
rect 872 -5972 888 -5548
rect 1804 -5548 1900 -5532
rect 1211 -5600 1533 -5599
rect 1211 -5920 1212 -5600
rect 1532 -5920 1533 -5600
rect 1211 -5921 1533 -5920
rect 792 -5988 888 -5972
rect 1804 -5972 1820 -5548
rect 1884 -5972 1900 -5548
rect 2816 -5548 2912 -5532
rect 2223 -5600 2545 -5599
rect 2223 -5920 2224 -5600
rect 2544 -5920 2545 -5600
rect 2223 -5921 2545 -5920
rect 1804 -5988 1900 -5972
rect 2816 -5972 2832 -5548
rect 2896 -5972 2912 -5548
rect 3828 -5548 3924 -5532
rect 3235 -5600 3557 -5599
rect 3235 -5920 3236 -5600
rect 3556 -5920 3557 -5600
rect 3235 -5921 3557 -5920
rect 2816 -5988 2912 -5972
rect 3828 -5972 3844 -5548
rect 3908 -5972 3924 -5548
rect 4840 -5548 4936 -5532
rect 4247 -5600 4569 -5599
rect 4247 -5920 4248 -5600
rect 4568 -5920 4569 -5600
rect 4247 -5921 4569 -5920
rect 3828 -5988 3924 -5972
rect 4840 -5972 4856 -5548
rect 4920 -5972 4936 -5548
rect 5852 -5548 5948 -5532
rect 5259 -5600 5581 -5599
rect 5259 -5920 5260 -5600
rect 5580 -5920 5581 -5600
rect 5259 -5921 5581 -5920
rect 4840 -5988 4936 -5972
rect 5852 -5972 5868 -5548
rect 5932 -5972 5948 -5548
rect 6864 -5548 6960 -5532
rect 6271 -5600 6593 -5599
rect 6271 -5920 6272 -5600
rect 6592 -5920 6593 -5600
rect 6271 -5921 6593 -5920
rect 5852 -5988 5948 -5972
rect 6864 -5972 6880 -5548
rect 6944 -5972 6960 -5548
rect 7876 -5548 7972 -5532
rect 7283 -5600 7605 -5599
rect 7283 -5920 7284 -5600
rect 7604 -5920 7605 -5600
rect 7283 -5921 7605 -5920
rect 6864 -5988 6960 -5972
rect 7876 -5972 7892 -5548
rect 7956 -5972 7972 -5548
rect 8888 -5548 8984 -5532
rect 8295 -5600 8617 -5599
rect 8295 -5920 8296 -5600
rect 8616 -5920 8617 -5600
rect 8295 -5921 8617 -5920
rect 7876 -5988 7972 -5972
rect 8888 -5972 8904 -5548
rect 8968 -5972 8984 -5548
rect 9900 -5548 9996 -5532
rect 9307 -5600 9629 -5599
rect 9307 -5920 9308 -5600
rect 9628 -5920 9629 -5600
rect 9307 -5921 9629 -5920
rect 8888 -5988 8984 -5972
rect 9900 -5972 9916 -5548
rect 9980 -5972 9996 -5548
rect 10912 -5548 11008 -5532
rect 10319 -5600 10641 -5599
rect 10319 -5920 10320 -5600
rect 10640 -5920 10641 -5600
rect 10319 -5921 10641 -5920
rect 9900 -5988 9996 -5972
rect 10912 -5972 10928 -5548
rect 10992 -5972 11008 -5548
rect 11924 -5548 12020 -5532
rect 11331 -5600 11653 -5599
rect 11331 -5920 11332 -5600
rect 11652 -5920 11653 -5600
rect 11331 -5921 11653 -5920
rect 10912 -5988 11008 -5972
rect 11924 -5972 11940 -5548
rect 12004 -5972 12020 -5548
rect 12936 -5548 13032 -5532
rect 12343 -5600 12665 -5599
rect 12343 -5920 12344 -5600
rect 12664 -5920 12665 -5600
rect 12343 -5921 12665 -5920
rect 11924 -5988 12020 -5972
rect 12936 -5972 12952 -5548
rect 13016 -5972 13032 -5548
rect 13948 -5548 14044 -5532
rect 13355 -5600 13677 -5599
rect 13355 -5920 13356 -5600
rect 13676 -5920 13677 -5600
rect 13355 -5921 13677 -5920
rect 12936 -5988 13032 -5972
rect 13948 -5972 13964 -5548
rect 14028 -5972 14044 -5548
rect 14960 -5548 15056 -5532
rect 14367 -5600 14689 -5599
rect 14367 -5920 14368 -5600
rect 14688 -5920 14689 -5600
rect 14367 -5921 14689 -5920
rect 13948 -5988 14044 -5972
rect 14960 -5972 14976 -5548
rect 15040 -5972 15056 -5548
rect 15972 -5548 16068 -5532
rect 15379 -5600 15701 -5599
rect 15379 -5920 15380 -5600
rect 15700 -5920 15701 -5600
rect 15379 -5921 15701 -5920
rect 14960 -5988 15056 -5972
rect 15972 -5972 15988 -5548
rect 16052 -5972 16068 -5548
rect 16984 -5548 17080 -5532
rect 16391 -5600 16713 -5599
rect 16391 -5920 16392 -5600
rect 16712 -5920 16713 -5600
rect 16391 -5921 16713 -5920
rect 15972 -5988 16068 -5972
rect 16984 -5972 17000 -5548
rect 17064 -5972 17080 -5548
rect 16984 -5988 17080 -5972
rect -16412 -6268 -16316 -6252
rect -17005 -6320 -16683 -6319
rect -17005 -6640 -17004 -6320
rect -16684 -6640 -16683 -6320
rect -17005 -6641 -16683 -6640
rect -16412 -6692 -16396 -6268
rect -16332 -6692 -16316 -6268
rect -15400 -6268 -15304 -6252
rect -15993 -6320 -15671 -6319
rect -15993 -6640 -15992 -6320
rect -15672 -6640 -15671 -6320
rect -15993 -6641 -15671 -6640
rect -16412 -6708 -16316 -6692
rect -15400 -6692 -15384 -6268
rect -15320 -6692 -15304 -6268
rect -14388 -6268 -14292 -6252
rect -14981 -6320 -14659 -6319
rect -14981 -6640 -14980 -6320
rect -14660 -6640 -14659 -6320
rect -14981 -6641 -14659 -6640
rect -15400 -6708 -15304 -6692
rect -14388 -6692 -14372 -6268
rect -14308 -6692 -14292 -6268
rect -13376 -6268 -13280 -6252
rect -13969 -6320 -13647 -6319
rect -13969 -6640 -13968 -6320
rect -13648 -6640 -13647 -6320
rect -13969 -6641 -13647 -6640
rect -14388 -6708 -14292 -6692
rect -13376 -6692 -13360 -6268
rect -13296 -6692 -13280 -6268
rect -12364 -6268 -12268 -6252
rect -12957 -6320 -12635 -6319
rect -12957 -6640 -12956 -6320
rect -12636 -6640 -12635 -6320
rect -12957 -6641 -12635 -6640
rect -13376 -6708 -13280 -6692
rect -12364 -6692 -12348 -6268
rect -12284 -6692 -12268 -6268
rect -11352 -6268 -11256 -6252
rect -11945 -6320 -11623 -6319
rect -11945 -6640 -11944 -6320
rect -11624 -6640 -11623 -6320
rect -11945 -6641 -11623 -6640
rect -12364 -6708 -12268 -6692
rect -11352 -6692 -11336 -6268
rect -11272 -6692 -11256 -6268
rect -10340 -6268 -10244 -6252
rect -10933 -6320 -10611 -6319
rect -10933 -6640 -10932 -6320
rect -10612 -6640 -10611 -6320
rect -10933 -6641 -10611 -6640
rect -11352 -6708 -11256 -6692
rect -10340 -6692 -10324 -6268
rect -10260 -6692 -10244 -6268
rect -9328 -6268 -9232 -6252
rect -9921 -6320 -9599 -6319
rect -9921 -6640 -9920 -6320
rect -9600 -6640 -9599 -6320
rect -9921 -6641 -9599 -6640
rect -10340 -6708 -10244 -6692
rect -9328 -6692 -9312 -6268
rect -9248 -6692 -9232 -6268
rect -8316 -6268 -8220 -6252
rect -8909 -6320 -8587 -6319
rect -8909 -6640 -8908 -6320
rect -8588 -6640 -8587 -6320
rect -8909 -6641 -8587 -6640
rect -9328 -6708 -9232 -6692
rect -8316 -6692 -8300 -6268
rect -8236 -6692 -8220 -6268
rect -7304 -6268 -7208 -6252
rect -7897 -6320 -7575 -6319
rect -7897 -6640 -7896 -6320
rect -7576 -6640 -7575 -6320
rect -7897 -6641 -7575 -6640
rect -8316 -6708 -8220 -6692
rect -7304 -6692 -7288 -6268
rect -7224 -6692 -7208 -6268
rect -6292 -6268 -6196 -6252
rect -6885 -6320 -6563 -6319
rect -6885 -6640 -6884 -6320
rect -6564 -6640 -6563 -6320
rect -6885 -6641 -6563 -6640
rect -7304 -6708 -7208 -6692
rect -6292 -6692 -6276 -6268
rect -6212 -6692 -6196 -6268
rect -5280 -6268 -5184 -6252
rect -5873 -6320 -5551 -6319
rect -5873 -6640 -5872 -6320
rect -5552 -6640 -5551 -6320
rect -5873 -6641 -5551 -6640
rect -6292 -6708 -6196 -6692
rect -5280 -6692 -5264 -6268
rect -5200 -6692 -5184 -6268
rect -4268 -6268 -4172 -6252
rect -4861 -6320 -4539 -6319
rect -4861 -6640 -4860 -6320
rect -4540 -6640 -4539 -6320
rect -4861 -6641 -4539 -6640
rect -5280 -6708 -5184 -6692
rect -4268 -6692 -4252 -6268
rect -4188 -6692 -4172 -6268
rect -3256 -6268 -3160 -6252
rect -3849 -6320 -3527 -6319
rect -3849 -6640 -3848 -6320
rect -3528 -6640 -3527 -6320
rect -3849 -6641 -3527 -6640
rect -4268 -6708 -4172 -6692
rect -3256 -6692 -3240 -6268
rect -3176 -6692 -3160 -6268
rect -2244 -6268 -2148 -6252
rect -2837 -6320 -2515 -6319
rect -2837 -6640 -2836 -6320
rect -2516 -6640 -2515 -6320
rect -2837 -6641 -2515 -6640
rect -3256 -6708 -3160 -6692
rect -2244 -6692 -2228 -6268
rect -2164 -6692 -2148 -6268
rect -1232 -6268 -1136 -6252
rect -1825 -6320 -1503 -6319
rect -1825 -6640 -1824 -6320
rect -1504 -6640 -1503 -6320
rect -1825 -6641 -1503 -6640
rect -2244 -6708 -2148 -6692
rect -1232 -6692 -1216 -6268
rect -1152 -6692 -1136 -6268
rect -220 -6268 -124 -6252
rect -813 -6320 -491 -6319
rect -813 -6640 -812 -6320
rect -492 -6640 -491 -6320
rect -813 -6641 -491 -6640
rect -1232 -6708 -1136 -6692
rect -220 -6692 -204 -6268
rect -140 -6692 -124 -6268
rect 792 -6268 888 -6252
rect 199 -6320 521 -6319
rect 199 -6640 200 -6320
rect 520 -6640 521 -6320
rect 199 -6641 521 -6640
rect -220 -6708 -124 -6692
rect 792 -6692 808 -6268
rect 872 -6692 888 -6268
rect 1804 -6268 1900 -6252
rect 1211 -6320 1533 -6319
rect 1211 -6640 1212 -6320
rect 1532 -6640 1533 -6320
rect 1211 -6641 1533 -6640
rect 792 -6708 888 -6692
rect 1804 -6692 1820 -6268
rect 1884 -6692 1900 -6268
rect 2816 -6268 2912 -6252
rect 2223 -6320 2545 -6319
rect 2223 -6640 2224 -6320
rect 2544 -6640 2545 -6320
rect 2223 -6641 2545 -6640
rect 1804 -6708 1900 -6692
rect 2816 -6692 2832 -6268
rect 2896 -6692 2912 -6268
rect 3828 -6268 3924 -6252
rect 3235 -6320 3557 -6319
rect 3235 -6640 3236 -6320
rect 3556 -6640 3557 -6320
rect 3235 -6641 3557 -6640
rect 2816 -6708 2912 -6692
rect 3828 -6692 3844 -6268
rect 3908 -6692 3924 -6268
rect 4840 -6268 4936 -6252
rect 4247 -6320 4569 -6319
rect 4247 -6640 4248 -6320
rect 4568 -6640 4569 -6320
rect 4247 -6641 4569 -6640
rect 3828 -6708 3924 -6692
rect 4840 -6692 4856 -6268
rect 4920 -6692 4936 -6268
rect 5852 -6268 5948 -6252
rect 5259 -6320 5581 -6319
rect 5259 -6640 5260 -6320
rect 5580 -6640 5581 -6320
rect 5259 -6641 5581 -6640
rect 4840 -6708 4936 -6692
rect 5852 -6692 5868 -6268
rect 5932 -6692 5948 -6268
rect 6864 -6268 6960 -6252
rect 6271 -6320 6593 -6319
rect 6271 -6640 6272 -6320
rect 6592 -6640 6593 -6320
rect 6271 -6641 6593 -6640
rect 5852 -6708 5948 -6692
rect 6864 -6692 6880 -6268
rect 6944 -6692 6960 -6268
rect 7876 -6268 7972 -6252
rect 7283 -6320 7605 -6319
rect 7283 -6640 7284 -6320
rect 7604 -6640 7605 -6320
rect 7283 -6641 7605 -6640
rect 6864 -6708 6960 -6692
rect 7876 -6692 7892 -6268
rect 7956 -6692 7972 -6268
rect 8888 -6268 8984 -6252
rect 8295 -6320 8617 -6319
rect 8295 -6640 8296 -6320
rect 8616 -6640 8617 -6320
rect 8295 -6641 8617 -6640
rect 7876 -6708 7972 -6692
rect 8888 -6692 8904 -6268
rect 8968 -6692 8984 -6268
rect 9900 -6268 9996 -6252
rect 9307 -6320 9629 -6319
rect 9307 -6640 9308 -6320
rect 9628 -6640 9629 -6320
rect 9307 -6641 9629 -6640
rect 8888 -6708 8984 -6692
rect 9900 -6692 9916 -6268
rect 9980 -6692 9996 -6268
rect 10912 -6268 11008 -6252
rect 10319 -6320 10641 -6319
rect 10319 -6640 10320 -6320
rect 10640 -6640 10641 -6320
rect 10319 -6641 10641 -6640
rect 9900 -6708 9996 -6692
rect 10912 -6692 10928 -6268
rect 10992 -6692 11008 -6268
rect 11924 -6268 12020 -6252
rect 11331 -6320 11653 -6319
rect 11331 -6640 11332 -6320
rect 11652 -6640 11653 -6320
rect 11331 -6641 11653 -6640
rect 10912 -6708 11008 -6692
rect 11924 -6692 11940 -6268
rect 12004 -6692 12020 -6268
rect 12936 -6268 13032 -6252
rect 12343 -6320 12665 -6319
rect 12343 -6640 12344 -6320
rect 12664 -6640 12665 -6320
rect 12343 -6641 12665 -6640
rect 11924 -6708 12020 -6692
rect 12936 -6692 12952 -6268
rect 13016 -6692 13032 -6268
rect 13948 -6268 14044 -6252
rect 13355 -6320 13677 -6319
rect 13355 -6640 13356 -6320
rect 13676 -6640 13677 -6320
rect 13355 -6641 13677 -6640
rect 12936 -6708 13032 -6692
rect 13948 -6692 13964 -6268
rect 14028 -6692 14044 -6268
rect 14960 -6268 15056 -6252
rect 14367 -6320 14689 -6319
rect 14367 -6640 14368 -6320
rect 14688 -6640 14689 -6320
rect 14367 -6641 14689 -6640
rect 13948 -6708 14044 -6692
rect 14960 -6692 14976 -6268
rect 15040 -6692 15056 -6268
rect 15972 -6268 16068 -6252
rect 15379 -6320 15701 -6319
rect 15379 -6640 15380 -6320
rect 15700 -6640 15701 -6320
rect 15379 -6641 15701 -6640
rect 14960 -6708 15056 -6692
rect 15972 -6692 15988 -6268
rect 16052 -6692 16068 -6268
rect 16984 -6268 17080 -6252
rect 16391 -6320 16713 -6319
rect 16391 -6640 16392 -6320
rect 16712 -6640 16713 -6320
rect 16391 -6641 16713 -6640
rect 15972 -6708 16068 -6692
rect 16984 -6692 17000 -6268
rect 17064 -6692 17080 -6268
rect 16984 -6708 17080 -6692
rect -16412 -6988 -16316 -6972
rect -17005 -7040 -16683 -7039
rect -17005 -7360 -17004 -7040
rect -16684 -7360 -16683 -7040
rect -17005 -7361 -16683 -7360
rect -16412 -7412 -16396 -6988
rect -16332 -7412 -16316 -6988
rect -15400 -6988 -15304 -6972
rect -15993 -7040 -15671 -7039
rect -15993 -7360 -15992 -7040
rect -15672 -7360 -15671 -7040
rect -15993 -7361 -15671 -7360
rect -16412 -7428 -16316 -7412
rect -15400 -7412 -15384 -6988
rect -15320 -7412 -15304 -6988
rect -14388 -6988 -14292 -6972
rect -14981 -7040 -14659 -7039
rect -14981 -7360 -14980 -7040
rect -14660 -7360 -14659 -7040
rect -14981 -7361 -14659 -7360
rect -15400 -7428 -15304 -7412
rect -14388 -7412 -14372 -6988
rect -14308 -7412 -14292 -6988
rect -13376 -6988 -13280 -6972
rect -13969 -7040 -13647 -7039
rect -13969 -7360 -13968 -7040
rect -13648 -7360 -13647 -7040
rect -13969 -7361 -13647 -7360
rect -14388 -7428 -14292 -7412
rect -13376 -7412 -13360 -6988
rect -13296 -7412 -13280 -6988
rect -12364 -6988 -12268 -6972
rect -12957 -7040 -12635 -7039
rect -12957 -7360 -12956 -7040
rect -12636 -7360 -12635 -7040
rect -12957 -7361 -12635 -7360
rect -13376 -7428 -13280 -7412
rect -12364 -7412 -12348 -6988
rect -12284 -7412 -12268 -6988
rect -11352 -6988 -11256 -6972
rect -11945 -7040 -11623 -7039
rect -11945 -7360 -11944 -7040
rect -11624 -7360 -11623 -7040
rect -11945 -7361 -11623 -7360
rect -12364 -7428 -12268 -7412
rect -11352 -7412 -11336 -6988
rect -11272 -7412 -11256 -6988
rect -10340 -6988 -10244 -6972
rect -10933 -7040 -10611 -7039
rect -10933 -7360 -10932 -7040
rect -10612 -7360 -10611 -7040
rect -10933 -7361 -10611 -7360
rect -11352 -7428 -11256 -7412
rect -10340 -7412 -10324 -6988
rect -10260 -7412 -10244 -6988
rect -9328 -6988 -9232 -6972
rect -9921 -7040 -9599 -7039
rect -9921 -7360 -9920 -7040
rect -9600 -7360 -9599 -7040
rect -9921 -7361 -9599 -7360
rect -10340 -7428 -10244 -7412
rect -9328 -7412 -9312 -6988
rect -9248 -7412 -9232 -6988
rect -8316 -6988 -8220 -6972
rect -8909 -7040 -8587 -7039
rect -8909 -7360 -8908 -7040
rect -8588 -7360 -8587 -7040
rect -8909 -7361 -8587 -7360
rect -9328 -7428 -9232 -7412
rect -8316 -7412 -8300 -6988
rect -8236 -7412 -8220 -6988
rect -7304 -6988 -7208 -6972
rect -7897 -7040 -7575 -7039
rect -7897 -7360 -7896 -7040
rect -7576 -7360 -7575 -7040
rect -7897 -7361 -7575 -7360
rect -8316 -7428 -8220 -7412
rect -7304 -7412 -7288 -6988
rect -7224 -7412 -7208 -6988
rect -6292 -6988 -6196 -6972
rect -6885 -7040 -6563 -7039
rect -6885 -7360 -6884 -7040
rect -6564 -7360 -6563 -7040
rect -6885 -7361 -6563 -7360
rect -7304 -7428 -7208 -7412
rect -6292 -7412 -6276 -6988
rect -6212 -7412 -6196 -6988
rect -5280 -6988 -5184 -6972
rect -5873 -7040 -5551 -7039
rect -5873 -7360 -5872 -7040
rect -5552 -7360 -5551 -7040
rect -5873 -7361 -5551 -7360
rect -6292 -7428 -6196 -7412
rect -5280 -7412 -5264 -6988
rect -5200 -7412 -5184 -6988
rect -4268 -6988 -4172 -6972
rect -4861 -7040 -4539 -7039
rect -4861 -7360 -4860 -7040
rect -4540 -7360 -4539 -7040
rect -4861 -7361 -4539 -7360
rect -5280 -7428 -5184 -7412
rect -4268 -7412 -4252 -6988
rect -4188 -7412 -4172 -6988
rect -3256 -6988 -3160 -6972
rect -3849 -7040 -3527 -7039
rect -3849 -7360 -3848 -7040
rect -3528 -7360 -3527 -7040
rect -3849 -7361 -3527 -7360
rect -4268 -7428 -4172 -7412
rect -3256 -7412 -3240 -6988
rect -3176 -7412 -3160 -6988
rect -2244 -6988 -2148 -6972
rect -2837 -7040 -2515 -7039
rect -2837 -7360 -2836 -7040
rect -2516 -7360 -2515 -7040
rect -2837 -7361 -2515 -7360
rect -3256 -7428 -3160 -7412
rect -2244 -7412 -2228 -6988
rect -2164 -7412 -2148 -6988
rect -1232 -6988 -1136 -6972
rect -1825 -7040 -1503 -7039
rect -1825 -7360 -1824 -7040
rect -1504 -7360 -1503 -7040
rect -1825 -7361 -1503 -7360
rect -2244 -7428 -2148 -7412
rect -1232 -7412 -1216 -6988
rect -1152 -7412 -1136 -6988
rect -220 -6988 -124 -6972
rect -813 -7040 -491 -7039
rect -813 -7360 -812 -7040
rect -492 -7360 -491 -7040
rect -813 -7361 -491 -7360
rect -1232 -7428 -1136 -7412
rect -220 -7412 -204 -6988
rect -140 -7412 -124 -6988
rect 792 -6988 888 -6972
rect 199 -7040 521 -7039
rect 199 -7360 200 -7040
rect 520 -7360 521 -7040
rect 199 -7361 521 -7360
rect -220 -7428 -124 -7412
rect 792 -7412 808 -6988
rect 872 -7412 888 -6988
rect 1804 -6988 1900 -6972
rect 1211 -7040 1533 -7039
rect 1211 -7360 1212 -7040
rect 1532 -7360 1533 -7040
rect 1211 -7361 1533 -7360
rect 792 -7428 888 -7412
rect 1804 -7412 1820 -6988
rect 1884 -7412 1900 -6988
rect 2816 -6988 2912 -6972
rect 2223 -7040 2545 -7039
rect 2223 -7360 2224 -7040
rect 2544 -7360 2545 -7040
rect 2223 -7361 2545 -7360
rect 1804 -7428 1900 -7412
rect 2816 -7412 2832 -6988
rect 2896 -7412 2912 -6988
rect 3828 -6988 3924 -6972
rect 3235 -7040 3557 -7039
rect 3235 -7360 3236 -7040
rect 3556 -7360 3557 -7040
rect 3235 -7361 3557 -7360
rect 2816 -7428 2912 -7412
rect 3828 -7412 3844 -6988
rect 3908 -7412 3924 -6988
rect 4840 -6988 4936 -6972
rect 4247 -7040 4569 -7039
rect 4247 -7360 4248 -7040
rect 4568 -7360 4569 -7040
rect 4247 -7361 4569 -7360
rect 3828 -7428 3924 -7412
rect 4840 -7412 4856 -6988
rect 4920 -7412 4936 -6988
rect 5852 -6988 5948 -6972
rect 5259 -7040 5581 -7039
rect 5259 -7360 5260 -7040
rect 5580 -7360 5581 -7040
rect 5259 -7361 5581 -7360
rect 4840 -7428 4936 -7412
rect 5852 -7412 5868 -6988
rect 5932 -7412 5948 -6988
rect 6864 -6988 6960 -6972
rect 6271 -7040 6593 -7039
rect 6271 -7360 6272 -7040
rect 6592 -7360 6593 -7040
rect 6271 -7361 6593 -7360
rect 5852 -7428 5948 -7412
rect 6864 -7412 6880 -6988
rect 6944 -7412 6960 -6988
rect 7876 -6988 7972 -6972
rect 7283 -7040 7605 -7039
rect 7283 -7360 7284 -7040
rect 7604 -7360 7605 -7040
rect 7283 -7361 7605 -7360
rect 6864 -7428 6960 -7412
rect 7876 -7412 7892 -6988
rect 7956 -7412 7972 -6988
rect 8888 -6988 8984 -6972
rect 8295 -7040 8617 -7039
rect 8295 -7360 8296 -7040
rect 8616 -7360 8617 -7040
rect 8295 -7361 8617 -7360
rect 7876 -7428 7972 -7412
rect 8888 -7412 8904 -6988
rect 8968 -7412 8984 -6988
rect 9900 -6988 9996 -6972
rect 9307 -7040 9629 -7039
rect 9307 -7360 9308 -7040
rect 9628 -7360 9629 -7040
rect 9307 -7361 9629 -7360
rect 8888 -7428 8984 -7412
rect 9900 -7412 9916 -6988
rect 9980 -7412 9996 -6988
rect 10912 -6988 11008 -6972
rect 10319 -7040 10641 -7039
rect 10319 -7360 10320 -7040
rect 10640 -7360 10641 -7040
rect 10319 -7361 10641 -7360
rect 9900 -7428 9996 -7412
rect 10912 -7412 10928 -6988
rect 10992 -7412 11008 -6988
rect 11924 -6988 12020 -6972
rect 11331 -7040 11653 -7039
rect 11331 -7360 11332 -7040
rect 11652 -7360 11653 -7040
rect 11331 -7361 11653 -7360
rect 10912 -7428 11008 -7412
rect 11924 -7412 11940 -6988
rect 12004 -7412 12020 -6988
rect 12936 -6988 13032 -6972
rect 12343 -7040 12665 -7039
rect 12343 -7360 12344 -7040
rect 12664 -7360 12665 -7040
rect 12343 -7361 12665 -7360
rect 11924 -7428 12020 -7412
rect 12936 -7412 12952 -6988
rect 13016 -7412 13032 -6988
rect 13948 -6988 14044 -6972
rect 13355 -7040 13677 -7039
rect 13355 -7360 13356 -7040
rect 13676 -7360 13677 -7040
rect 13355 -7361 13677 -7360
rect 12936 -7428 13032 -7412
rect 13948 -7412 13964 -6988
rect 14028 -7412 14044 -6988
rect 14960 -6988 15056 -6972
rect 14367 -7040 14689 -7039
rect 14367 -7360 14368 -7040
rect 14688 -7360 14689 -7040
rect 14367 -7361 14689 -7360
rect 13948 -7428 14044 -7412
rect 14960 -7412 14976 -6988
rect 15040 -7412 15056 -6988
rect 15972 -6988 16068 -6972
rect 15379 -7040 15701 -7039
rect 15379 -7360 15380 -7040
rect 15700 -7360 15701 -7040
rect 15379 -7361 15701 -7360
rect 14960 -7428 15056 -7412
rect 15972 -7412 15988 -6988
rect 16052 -7412 16068 -6988
rect 16984 -6988 17080 -6972
rect 16391 -7040 16713 -7039
rect 16391 -7360 16392 -7040
rect 16712 -7360 16713 -7040
rect 16391 -7361 16713 -7360
rect 15972 -7428 16068 -7412
rect 16984 -7412 17000 -6988
rect 17064 -7412 17080 -6988
rect 16984 -7428 17080 -7412
rect -16412 -7708 -16316 -7692
rect -17005 -7760 -16683 -7759
rect -17005 -8080 -17004 -7760
rect -16684 -8080 -16683 -7760
rect -17005 -8081 -16683 -8080
rect -16412 -8132 -16396 -7708
rect -16332 -8132 -16316 -7708
rect -15400 -7708 -15304 -7692
rect -15993 -7760 -15671 -7759
rect -15993 -8080 -15992 -7760
rect -15672 -8080 -15671 -7760
rect -15993 -8081 -15671 -8080
rect -16412 -8148 -16316 -8132
rect -15400 -8132 -15384 -7708
rect -15320 -8132 -15304 -7708
rect -14388 -7708 -14292 -7692
rect -14981 -7760 -14659 -7759
rect -14981 -8080 -14980 -7760
rect -14660 -8080 -14659 -7760
rect -14981 -8081 -14659 -8080
rect -15400 -8148 -15304 -8132
rect -14388 -8132 -14372 -7708
rect -14308 -8132 -14292 -7708
rect -13376 -7708 -13280 -7692
rect -13969 -7760 -13647 -7759
rect -13969 -8080 -13968 -7760
rect -13648 -8080 -13647 -7760
rect -13969 -8081 -13647 -8080
rect -14388 -8148 -14292 -8132
rect -13376 -8132 -13360 -7708
rect -13296 -8132 -13280 -7708
rect -12364 -7708 -12268 -7692
rect -12957 -7760 -12635 -7759
rect -12957 -8080 -12956 -7760
rect -12636 -8080 -12635 -7760
rect -12957 -8081 -12635 -8080
rect -13376 -8148 -13280 -8132
rect -12364 -8132 -12348 -7708
rect -12284 -8132 -12268 -7708
rect -11352 -7708 -11256 -7692
rect -11945 -7760 -11623 -7759
rect -11945 -8080 -11944 -7760
rect -11624 -8080 -11623 -7760
rect -11945 -8081 -11623 -8080
rect -12364 -8148 -12268 -8132
rect -11352 -8132 -11336 -7708
rect -11272 -8132 -11256 -7708
rect -10340 -7708 -10244 -7692
rect -10933 -7760 -10611 -7759
rect -10933 -8080 -10932 -7760
rect -10612 -8080 -10611 -7760
rect -10933 -8081 -10611 -8080
rect -11352 -8148 -11256 -8132
rect -10340 -8132 -10324 -7708
rect -10260 -8132 -10244 -7708
rect -9328 -7708 -9232 -7692
rect -9921 -7760 -9599 -7759
rect -9921 -8080 -9920 -7760
rect -9600 -8080 -9599 -7760
rect -9921 -8081 -9599 -8080
rect -10340 -8148 -10244 -8132
rect -9328 -8132 -9312 -7708
rect -9248 -8132 -9232 -7708
rect -8316 -7708 -8220 -7692
rect -8909 -7760 -8587 -7759
rect -8909 -8080 -8908 -7760
rect -8588 -8080 -8587 -7760
rect -8909 -8081 -8587 -8080
rect -9328 -8148 -9232 -8132
rect -8316 -8132 -8300 -7708
rect -8236 -8132 -8220 -7708
rect -7304 -7708 -7208 -7692
rect -7897 -7760 -7575 -7759
rect -7897 -8080 -7896 -7760
rect -7576 -8080 -7575 -7760
rect -7897 -8081 -7575 -8080
rect -8316 -8148 -8220 -8132
rect -7304 -8132 -7288 -7708
rect -7224 -8132 -7208 -7708
rect -6292 -7708 -6196 -7692
rect -6885 -7760 -6563 -7759
rect -6885 -8080 -6884 -7760
rect -6564 -8080 -6563 -7760
rect -6885 -8081 -6563 -8080
rect -7304 -8148 -7208 -8132
rect -6292 -8132 -6276 -7708
rect -6212 -8132 -6196 -7708
rect -5280 -7708 -5184 -7692
rect -5873 -7760 -5551 -7759
rect -5873 -8080 -5872 -7760
rect -5552 -8080 -5551 -7760
rect -5873 -8081 -5551 -8080
rect -6292 -8148 -6196 -8132
rect -5280 -8132 -5264 -7708
rect -5200 -8132 -5184 -7708
rect -4268 -7708 -4172 -7692
rect -4861 -7760 -4539 -7759
rect -4861 -8080 -4860 -7760
rect -4540 -8080 -4539 -7760
rect -4861 -8081 -4539 -8080
rect -5280 -8148 -5184 -8132
rect -4268 -8132 -4252 -7708
rect -4188 -8132 -4172 -7708
rect -3256 -7708 -3160 -7692
rect -3849 -7760 -3527 -7759
rect -3849 -8080 -3848 -7760
rect -3528 -8080 -3527 -7760
rect -3849 -8081 -3527 -8080
rect -4268 -8148 -4172 -8132
rect -3256 -8132 -3240 -7708
rect -3176 -8132 -3160 -7708
rect -2244 -7708 -2148 -7692
rect -2837 -7760 -2515 -7759
rect -2837 -8080 -2836 -7760
rect -2516 -8080 -2515 -7760
rect -2837 -8081 -2515 -8080
rect -3256 -8148 -3160 -8132
rect -2244 -8132 -2228 -7708
rect -2164 -8132 -2148 -7708
rect -1232 -7708 -1136 -7692
rect -1825 -7760 -1503 -7759
rect -1825 -8080 -1824 -7760
rect -1504 -8080 -1503 -7760
rect -1825 -8081 -1503 -8080
rect -2244 -8148 -2148 -8132
rect -1232 -8132 -1216 -7708
rect -1152 -8132 -1136 -7708
rect -220 -7708 -124 -7692
rect -813 -7760 -491 -7759
rect -813 -8080 -812 -7760
rect -492 -8080 -491 -7760
rect -813 -8081 -491 -8080
rect -1232 -8148 -1136 -8132
rect -220 -8132 -204 -7708
rect -140 -8132 -124 -7708
rect 792 -7708 888 -7692
rect 199 -7760 521 -7759
rect 199 -8080 200 -7760
rect 520 -8080 521 -7760
rect 199 -8081 521 -8080
rect -220 -8148 -124 -8132
rect 792 -8132 808 -7708
rect 872 -8132 888 -7708
rect 1804 -7708 1900 -7692
rect 1211 -7760 1533 -7759
rect 1211 -8080 1212 -7760
rect 1532 -8080 1533 -7760
rect 1211 -8081 1533 -8080
rect 792 -8148 888 -8132
rect 1804 -8132 1820 -7708
rect 1884 -8132 1900 -7708
rect 2816 -7708 2912 -7692
rect 2223 -7760 2545 -7759
rect 2223 -8080 2224 -7760
rect 2544 -8080 2545 -7760
rect 2223 -8081 2545 -8080
rect 1804 -8148 1900 -8132
rect 2816 -8132 2832 -7708
rect 2896 -8132 2912 -7708
rect 3828 -7708 3924 -7692
rect 3235 -7760 3557 -7759
rect 3235 -8080 3236 -7760
rect 3556 -8080 3557 -7760
rect 3235 -8081 3557 -8080
rect 2816 -8148 2912 -8132
rect 3828 -8132 3844 -7708
rect 3908 -8132 3924 -7708
rect 4840 -7708 4936 -7692
rect 4247 -7760 4569 -7759
rect 4247 -8080 4248 -7760
rect 4568 -8080 4569 -7760
rect 4247 -8081 4569 -8080
rect 3828 -8148 3924 -8132
rect 4840 -8132 4856 -7708
rect 4920 -8132 4936 -7708
rect 5852 -7708 5948 -7692
rect 5259 -7760 5581 -7759
rect 5259 -8080 5260 -7760
rect 5580 -8080 5581 -7760
rect 5259 -8081 5581 -8080
rect 4840 -8148 4936 -8132
rect 5852 -8132 5868 -7708
rect 5932 -8132 5948 -7708
rect 6864 -7708 6960 -7692
rect 6271 -7760 6593 -7759
rect 6271 -8080 6272 -7760
rect 6592 -8080 6593 -7760
rect 6271 -8081 6593 -8080
rect 5852 -8148 5948 -8132
rect 6864 -8132 6880 -7708
rect 6944 -8132 6960 -7708
rect 7876 -7708 7972 -7692
rect 7283 -7760 7605 -7759
rect 7283 -8080 7284 -7760
rect 7604 -8080 7605 -7760
rect 7283 -8081 7605 -8080
rect 6864 -8148 6960 -8132
rect 7876 -8132 7892 -7708
rect 7956 -8132 7972 -7708
rect 8888 -7708 8984 -7692
rect 8295 -7760 8617 -7759
rect 8295 -8080 8296 -7760
rect 8616 -8080 8617 -7760
rect 8295 -8081 8617 -8080
rect 7876 -8148 7972 -8132
rect 8888 -8132 8904 -7708
rect 8968 -8132 8984 -7708
rect 9900 -7708 9996 -7692
rect 9307 -7760 9629 -7759
rect 9307 -8080 9308 -7760
rect 9628 -8080 9629 -7760
rect 9307 -8081 9629 -8080
rect 8888 -8148 8984 -8132
rect 9900 -8132 9916 -7708
rect 9980 -8132 9996 -7708
rect 10912 -7708 11008 -7692
rect 10319 -7760 10641 -7759
rect 10319 -8080 10320 -7760
rect 10640 -8080 10641 -7760
rect 10319 -8081 10641 -8080
rect 9900 -8148 9996 -8132
rect 10912 -8132 10928 -7708
rect 10992 -8132 11008 -7708
rect 11924 -7708 12020 -7692
rect 11331 -7760 11653 -7759
rect 11331 -8080 11332 -7760
rect 11652 -8080 11653 -7760
rect 11331 -8081 11653 -8080
rect 10912 -8148 11008 -8132
rect 11924 -8132 11940 -7708
rect 12004 -8132 12020 -7708
rect 12936 -7708 13032 -7692
rect 12343 -7760 12665 -7759
rect 12343 -8080 12344 -7760
rect 12664 -8080 12665 -7760
rect 12343 -8081 12665 -8080
rect 11924 -8148 12020 -8132
rect 12936 -8132 12952 -7708
rect 13016 -8132 13032 -7708
rect 13948 -7708 14044 -7692
rect 13355 -7760 13677 -7759
rect 13355 -8080 13356 -7760
rect 13676 -8080 13677 -7760
rect 13355 -8081 13677 -8080
rect 12936 -8148 13032 -8132
rect 13948 -8132 13964 -7708
rect 14028 -8132 14044 -7708
rect 14960 -7708 15056 -7692
rect 14367 -7760 14689 -7759
rect 14367 -8080 14368 -7760
rect 14688 -8080 14689 -7760
rect 14367 -8081 14689 -8080
rect 13948 -8148 14044 -8132
rect 14960 -8132 14976 -7708
rect 15040 -8132 15056 -7708
rect 15972 -7708 16068 -7692
rect 15379 -7760 15701 -7759
rect 15379 -8080 15380 -7760
rect 15700 -8080 15701 -7760
rect 15379 -8081 15701 -8080
rect 14960 -8148 15056 -8132
rect 15972 -8132 15988 -7708
rect 16052 -8132 16068 -7708
rect 16984 -7708 17080 -7692
rect 16391 -7760 16713 -7759
rect 16391 -8080 16392 -7760
rect 16712 -8080 16713 -7760
rect 16391 -8081 16713 -8080
rect 15972 -8148 16068 -8132
rect 16984 -8132 17000 -7708
rect 17064 -8132 17080 -7708
rect 16984 -8148 17080 -8132
rect -16412 -8428 -16316 -8412
rect -17005 -8480 -16683 -8479
rect -17005 -8800 -17004 -8480
rect -16684 -8800 -16683 -8480
rect -17005 -8801 -16683 -8800
rect -16412 -8852 -16396 -8428
rect -16332 -8852 -16316 -8428
rect -15400 -8428 -15304 -8412
rect -15993 -8480 -15671 -8479
rect -15993 -8800 -15992 -8480
rect -15672 -8800 -15671 -8480
rect -15993 -8801 -15671 -8800
rect -16412 -8868 -16316 -8852
rect -15400 -8852 -15384 -8428
rect -15320 -8852 -15304 -8428
rect -14388 -8428 -14292 -8412
rect -14981 -8480 -14659 -8479
rect -14981 -8800 -14980 -8480
rect -14660 -8800 -14659 -8480
rect -14981 -8801 -14659 -8800
rect -15400 -8868 -15304 -8852
rect -14388 -8852 -14372 -8428
rect -14308 -8852 -14292 -8428
rect -13376 -8428 -13280 -8412
rect -13969 -8480 -13647 -8479
rect -13969 -8800 -13968 -8480
rect -13648 -8800 -13647 -8480
rect -13969 -8801 -13647 -8800
rect -14388 -8868 -14292 -8852
rect -13376 -8852 -13360 -8428
rect -13296 -8852 -13280 -8428
rect -12364 -8428 -12268 -8412
rect -12957 -8480 -12635 -8479
rect -12957 -8800 -12956 -8480
rect -12636 -8800 -12635 -8480
rect -12957 -8801 -12635 -8800
rect -13376 -8868 -13280 -8852
rect -12364 -8852 -12348 -8428
rect -12284 -8852 -12268 -8428
rect -11352 -8428 -11256 -8412
rect -11945 -8480 -11623 -8479
rect -11945 -8800 -11944 -8480
rect -11624 -8800 -11623 -8480
rect -11945 -8801 -11623 -8800
rect -12364 -8868 -12268 -8852
rect -11352 -8852 -11336 -8428
rect -11272 -8852 -11256 -8428
rect -10340 -8428 -10244 -8412
rect -10933 -8480 -10611 -8479
rect -10933 -8800 -10932 -8480
rect -10612 -8800 -10611 -8480
rect -10933 -8801 -10611 -8800
rect -11352 -8868 -11256 -8852
rect -10340 -8852 -10324 -8428
rect -10260 -8852 -10244 -8428
rect -9328 -8428 -9232 -8412
rect -9921 -8480 -9599 -8479
rect -9921 -8800 -9920 -8480
rect -9600 -8800 -9599 -8480
rect -9921 -8801 -9599 -8800
rect -10340 -8868 -10244 -8852
rect -9328 -8852 -9312 -8428
rect -9248 -8852 -9232 -8428
rect -8316 -8428 -8220 -8412
rect -8909 -8480 -8587 -8479
rect -8909 -8800 -8908 -8480
rect -8588 -8800 -8587 -8480
rect -8909 -8801 -8587 -8800
rect -9328 -8868 -9232 -8852
rect -8316 -8852 -8300 -8428
rect -8236 -8852 -8220 -8428
rect -7304 -8428 -7208 -8412
rect -7897 -8480 -7575 -8479
rect -7897 -8800 -7896 -8480
rect -7576 -8800 -7575 -8480
rect -7897 -8801 -7575 -8800
rect -8316 -8868 -8220 -8852
rect -7304 -8852 -7288 -8428
rect -7224 -8852 -7208 -8428
rect -6292 -8428 -6196 -8412
rect -6885 -8480 -6563 -8479
rect -6885 -8800 -6884 -8480
rect -6564 -8800 -6563 -8480
rect -6885 -8801 -6563 -8800
rect -7304 -8868 -7208 -8852
rect -6292 -8852 -6276 -8428
rect -6212 -8852 -6196 -8428
rect -5280 -8428 -5184 -8412
rect -5873 -8480 -5551 -8479
rect -5873 -8800 -5872 -8480
rect -5552 -8800 -5551 -8480
rect -5873 -8801 -5551 -8800
rect -6292 -8868 -6196 -8852
rect -5280 -8852 -5264 -8428
rect -5200 -8852 -5184 -8428
rect -4268 -8428 -4172 -8412
rect -4861 -8480 -4539 -8479
rect -4861 -8800 -4860 -8480
rect -4540 -8800 -4539 -8480
rect -4861 -8801 -4539 -8800
rect -5280 -8868 -5184 -8852
rect -4268 -8852 -4252 -8428
rect -4188 -8852 -4172 -8428
rect -3256 -8428 -3160 -8412
rect -3849 -8480 -3527 -8479
rect -3849 -8800 -3848 -8480
rect -3528 -8800 -3527 -8480
rect -3849 -8801 -3527 -8800
rect -4268 -8868 -4172 -8852
rect -3256 -8852 -3240 -8428
rect -3176 -8852 -3160 -8428
rect -2244 -8428 -2148 -8412
rect -2837 -8480 -2515 -8479
rect -2837 -8800 -2836 -8480
rect -2516 -8800 -2515 -8480
rect -2837 -8801 -2515 -8800
rect -3256 -8868 -3160 -8852
rect -2244 -8852 -2228 -8428
rect -2164 -8852 -2148 -8428
rect -1232 -8428 -1136 -8412
rect -1825 -8480 -1503 -8479
rect -1825 -8800 -1824 -8480
rect -1504 -8800 -1503 -8480
rect -1825 -8801 -1503 -8800
rect -2244 -8868 -2148 -8852
rect -1232 -8852 -1216 -8428
rect -1152 -8852 -1136 -8428
rect -220 -8428 -124 -8412
rect -813 -8480 -491 -8479
rect -813 -8800 -812 -8480
rect -492 -8800 -491 -8480
rect -813 -8801 -491 -8800
rect -1232 -8868 -1136 -8852
rect -220 -8852 -204 -8428
rect -140 -8852 -124 -8428
rect 792 -8428 888 -8412
rect 199 -8480 521 -8479
rect 199 -8800 200 -8480
rect 520 -8800 521 -8480
rect 199 -8801 521 -8800
rect -220 -8868 -124 -8852
rect 792 -8852 808 -8428
rect 872 -8852 888 -8428
rect 1804 -8428 1900 -8412
rect 1211 -8480 1533 -8479
rect 1211 -8800 1212 -8480
rect 1532 -8800 1533 -8480
rect 1211 -8801 1533 -8800
rect 792 -8868 888 -8852
rect 1804 -8852 1820 -8428
rect 1884 -8852 1900 -8428
rect 2816 -8428 2912 -8412
rect 2223 -8480 2545 -8479
rect 2223 -8800 2224 -8480
rect 2544 -8800 2545 -8480
rect 2223 -8801 2545 -8800
rect 1804 -8868 1900 -8852
rect 2816 -8852 2832 -8428
rect 2896 -8852 2912 -8428
rect 3828 -8428 3924 -8412
rect 3235 -8480 3557 -8479
rect 3235 -8800 3236 -8480
rect 3556 -8800 3557 -8480
rect 3235 -8801 3557 -8800
rect 2816 -8868 2912 -8852
rect 3828 -8852 3844 -8428
rect 3908 -8852 3924 -8428
rect 4840 -8428 4936 -8412
rect 4247 -8480 4569 -8479
rect 4247 -8800 4248 -8480
rect 4568 -8800 4569 -8480
rect 4247 -8801 4569 -8800
rect 3828 -8868 3924 -8852
rect 4840 -8852 4856 -8428
rect 4920 -8852 4936 -8428
rect 5852 -8428 5948 -8412
rect 5259 -8480 5581 -8479
rect 5259 -8800 5260 -8480
rect 5580 -8800 5581 -8480
rect 5259 -8801 5581 -8800
rect 4840 -8868 4936 -8852
rect 5852 -8852 5868 -8428
rect 5932 -8852 5948 -8428
rect 6864 -8428 6960 -8412
rect 6271 -8480 6593 -8479
rect 6271 -8800 6272 -8480
rect 6592 -8800 6593 -8480
rect 6271 -8801 6593 -8800
rect 5852 -8868 5948 -8852
rect 6864 -8852 6880 -8428
rect 6944 -8852 6960 -8428
rect 7876 -8428 7972 -8412
rect 7283 -8480 7605 -8479
rect 7283 -8800 7284 -8480
rect 7604 -8800 7605 -8480
rect 7283 -8801 7605 -8800
rect 6864 -8868 6960 -8852
rect 7876 -8852 7892 -8428
rect 7956 -8852 7972 -8428
rect 8888 -8428 8984 -8412
rect 8295 -8480 8617 -8479
rect 8295 -8800 8296 -8480
rect 8616 -8800 8617 -8480
rect 8295 -8801 8617 -8800
rect 7876 -8868 7972 -8852
rect 8888 -8852 8904 -8428
rect 8968 -8852 8984 -8428
rect 9900 -8428 9996 -8412
rect 9307 -8480 9629 -8479
rect 9307 -8800 9308 -8480
rect 9628 -8800 9629 -8480
rect 9307 -8801 9629 -8800
rect 8888 -8868 8984 -8852
rect 9900 -8852 9916 -8428
rect 9980 -8852 9996 -8428
rect 10912 -8428 11008 -8412
rect 10319 -8480 10641 -8479
rect 10319 -8800 10320 -8480
rect 10640 -8800 10641 -8480
rect 10319 -8801 10641 -8800
rect 9900 -8868 9996 -8852
rect 10912 -8852 10928 -8428
rect 10992 -8852 11008 -8428
rect 11924 -8428 12020 -8412
rect 11331 -8480 11653 -8479
rect 11331 -8800 11332 -8480
rect 11652 -8800 11653 -8480
rect 11331 -8801 11653 -8800
rect 10912 -8868 11008 -8852
rect 11924 -8852 11940 -8428
rect 12004 -8852 12020 -8428
rect 12936 -8428 13032 -8412
rect 12343 -8480 12665 -8479
rect 12343 -8800 12344 -8480
rect 12664 -8800 12665 -8480
rect 12343 -8801 12665 -8800
rect 11924 -8868 12020 -8852
rect 12936 -8852 12952 -8428
rect 13016 -8852 13032 -8428
rect 13948 -8428 14044 -8412
rect 13355 -8480 13677 -8479
rect 13355 -8800 13356 -8480
rect 13676 -8800 13677 -8480
rect 13355 -8801 13677 -8800
rect 12936 -8868 13032 -8852
rect 13948 -8852 13964 -8428
rect 14028 -8852 14044 -8428
rect 14960 -8428 15056 -8412
rect 14367 -8480 14689 -8479
rect 14367 -8800 14368 -8480
rect 14688 -8800 14689 -8480
rect 14367 -8801 14689 -8800
rect 13948 -8868 14044 -8852
rect 14960 -8852 14976 -8428
rect 15040 -8852 15056 -8428
rect 15972 -8428 16068 -8412
rect 15379 -8480 15701 -8479
rect 15379 -8800 15380 -8480
rect 15700 -8800 15701 -8480
rect 15379 -8801 15701 -8800
rect 14960 -8868 15056 -8852
rect 15972 -8852 15988 -8428
rect 16052 -8852 16068 -8428
rect 16984 -8428 17080 -8412
rect 16391 -8480 16713 -8479
rect 16391 -8800 16392 -8480
rect 16712 -8800 16713 -8480
rect 16391 -8801 16713 -8800
rect 15972 -8868 16068 -8852
rect 16984 -8852 17000 -8428
rect 17064 -8852 17080 -8428
rect 16984 -8868 17080 -8852
rect -16412 -9148 -16316 -9132
rect -17005 -9200 -16683 -9199
rect -17005 -9520 -17004 -9200
rect -16684 -9520 -16683 -9200
rect -17005 -9521 -16683 -9520
rect -16412 -9572 -16396 -9148
rect -16332 -9572 -16316 -9148
rect -15400 -9148 -15304 -9132
rect -15993 -9200 -15671 -9199
rect -15993 -9520 -15992 -9200
rect -15672 -9520 -15671 -9200
rect -15993 -9521 -15671 -9520
rect -16412 -9588 -16316 -9572
rect -15400 -9572 -15384 -9148
rect -15320 -9572 -15304 -9148
rect -14388 -9148 -14292 -9132
rect -14981 -9200 -14659 -9199
rect -14981 -9520 -14980 -9200
rect -14660 -9520 -14659 -9200
rect -14981 -9521 -14659 -9520
rect -15400 -9588 -15304 -9572
rect -14388 -9572 -14372 -9148
rect -14308 -9572 -14292 -9148
rect -13376 -9148 -13280 -9132
rect -13969 -9200 -13647 -9199
rect -13969 -9520 -13968 -9200
rect -13648 -9520 -13647 -9200
rect -13969 -9521 -13647 -9520
rect -14388 -9588 -14292 -9572
rect -13376 -9572 -13360 -9148
rect -13296 -9572 -13280 -9148
rect -12364 -9148 -12268 -9132
rect -12957 -9200 -12635 -9199
rect -12957 -9520 -12956 -9200
rect -12636 -9520 -12635 -9200
rect -12957 -9521 -12635 -9520
rect -13376 -9588 -13280 -9572
rect -12364 -9572 -12348 -9148
rect -12284 -9572 -12268 -9148
rect -11352 -9148 -11256 -9132
rect -11945 -9200 -11623 -9199
rect -11945 -9520 -11944 -9200
rect -11624 -9520 -11623 -9200
rect -11945 -9521 -11623 -9520
rect -12364 -9588 -12268 -9572
rect -11352 -9572 -11336 -9148
rect -11272 -9572 -11256 -9148
rect -10340 -9148 -10244 -9132
rect -10933 -9200 -10611 -9199
rect -10933 -9520 -10932 -9200
rect -10612 -9520 -10611 -9200
rect -10933 -9521 -10611 -9520
rect -11352 -9588 -11256 -9572
rect -10340 -9572 -10324 -9148
rect -10260 -9572 -10244 -9148
rect -9328 -9148 -9232 -9132
rect -9921 -9200 -9599 -9199
rect -9921 -9520 -9920 -9200
rect -9600 -9520 -9599 -9200
rect -9921 -9521 -9599 -9520
rect -10340 -9588 -10244 -9572
rect -9328 -9572 -9312 -9148
rect -9248 -9572 -9232 -9148
rect -8316 -9148 -8220 -9132
rect -8909 -9200 -8587 -9199
rect -8909 -9520 -8908 -9200
rect -8588 -9520 -8587 -9200
rect -8909 -9521 -8587 -9520
rect -9328 -9588 -9232 -9572
rect -8316 -9572 -8300 -9148
rect -8236 -9572 -8220 -9148
rect -7304 -9148 -7208 -9132
rect -7897 -9200 -7575 -9199
rect -7897 -9520 -7896 -9200
rect -7576 -9520 -7575 -9200
rect -7897 -9521 -7575 -9520
rect -8316 -9588 -8220 -9572
rect -7304 -9572 -7288 -9148
rect -7224 -9572 -7208 -9148
rect -6292 -9148 -6196 -9132
rect -6885 -9200 -6563 -9199
rect -6885 -9520 -6884 -9200
rect -6564 -9520 -6563 -9200
rect -6885 -9521 -6563 -9520
rect -7304 -9588 -7208 -9572
rect -6292 -9572 -6276 -9148
rect -6212 -9572 -6196 -9148
rect -5280 -9148 -5184 -9132
rect -5873 -9200 -5551 -9199
rect -5873 -9520 -5872 -9200
rect -5552 -9520 -5551 -9200
rect -5873 -9521 -5551 -9520
rect -6292 -9588 -6196 -9572
rect -5280 -9572 -5264 -9148
rect -5200 -9572 -5184 -9148
rect -4268 -9148 -4172 -9132
rect -4861 -9200 -4539 -9199
rect -4861 -9520 -4860 -9200
rect -4540 -9520 -4539 -9200
rect -4861 -9521 -4539 -9520
rect -5280 -9588 -5184 -9572
rect -4268 -9572 -4252 -9148
rect -4188 -9572 -4172 -9148
rect -3256 -9148 -3160 -9132
rect -3849 -9200 -3527 -9199
rect -3849 -9520 -3848 -9200
rect -3528 -9520 -3527 -9200
rect -3849 -9521 -3527 -9520
rect -4268 -9588 -4172 -9572
rect -3256 -9572 -3240 -9148
rect -3176 -9572 -3160 -9148
rect -2244 -9148 -2148 -9132
rect -2837 -9200 -2515 -9199
rect -2837 -9520 -2836 -9200
rect -2516 -9520 -2515 -9200
rect -2837 -9521 -2515 -9520
rect -3256 -9588 -3160 -9572
rect -2244 -9572 -2228 -9148
rect -2164 -9572 -2148 -9148
rect -1232 -9148 -1136 -9132
rect -1825 -9200 -1503 -9199
rect -1825 -9520 -1824 -9200
rect -1504 -9520 -1503 -9200
rect -1825 -9521 -1503 -9520
rect -2244 -9588 -2148 -9572
rect -1232 -9572 -1216 -9148
rect -1152 -9572 -1136 -9148
rect -220 -9148 -124 -9132
rect -813 -9200 -491 -9199
rect -813 -9520 -812 -9200
rect -492 -9520 -491 -9200
rect -813 -9521 -491 -9520
rect -1232 -9588 -1136 -9572
rect -220 -9572 -204 -9148
rect -140 -9572 -124 -9148
rect 792 -9148 888 -9132
rect 199 -9200 521 -9199
rect 199 -9520 200 -9200
rect 520 -9520 521 -9200
rect 199 -9521 521 -9520
rect -220 -9588 -124 -9572
rect 792 -9572 808 -9148
rect 872 -9572 888 -9148
rect 1804 -9148 1900 -9132
rect 1211 -9200 1533 -9199
rect 1211 -9520 1212 -9200
rect 1532 -9520 1533 -9200
rect 1211 -9521 1533 -9520
rect 792 -9588 888 -9572
rect 1804 -9572 1820 -9148
rect 1884 -9572 1900 -9148
rect 2816 -9148 2912 -9132
rect 2223 -9200 2545 -9199
rect 2223 -9520 2224 -9200
rect 2544 -9520 2545 -9200
rect 2223 -9521 2545 -9520
rect 1804 -9588 1900 -9572
rect 2816 -9572 2832 -9148
rect 2896 -9572 2912 -9148
rect 3828 -9148 3924 -9132
rect 3235 -9200 3557 -9199
rect 3235 -9520 3236 -9200
rect 3556 -9520 3557 -9200
rect 3235 -9521 3557 -9520
rect 2816 -9588 2912 -9572
rect 3828 -9572 3844 -9148
rect 3908 -9572 3924 -9148
rect 4840 -9148 4936 -9132
rect 4247 -9200 4569 -9199
rect 4247 -9520 4248 -9200
rect 4568 -9520 4569 -9200
rect 4247 -9521 4569 -9520
rect 3828 -9588 3924 -9572
rect 4840 -9572 4856 -9148
rect 4920 -9572 4936 -9148
rect 5852 -9148 5948 -9132
rect 5259 -9200 5581 -9199
rect 5259 -9520 5260 -9200
rect 5580 -9520 5581 -9200
rect 5259 -9521 5581 -9520
rect 4840 -9588 4936 -9572
rect 5852 -9572 5868 -9148
rect 5932 -9572 5948 -9148
rect 6864 -9148 6960 -9132
rect 6271 -9200 6593 -9199
rect 6271 -9520 6272 -9200
rect 6592 -9520 6593 -9200
rect 6271 -9521 6593 -9520
rect 5852 -9588 5948 -9572
rect 6864 -9572 6880 -9148
rect 6944 -9572 6960 -9148
rect 7876 -9148 7972 -9132
rect 7283 -9200 7605 -9199
rect 7283 -9520 7284 -9200
rect 7604 -9520 7605 -9200
rect 7283 -9521 7605 -9520
rect 6864 -9588 6960 -9572
rect 7876 -9572 7892 -9148
rect 7956 -9572 7972 -9148
rect 8888 -9148 8984 -9132
rect 8295 -9200 8617 -9199
rect 8295 -9520 8296 -9200
rect 8616 -9520 8617 -9200
rect 8295 -9521 8617 -9520
rect 7876 -9588 7972 -9572
rect 8888 -9572 8904 -9148
rect 8968 -9572 8984 -9148
rect 9900 -9148 9996 -9132
rect 9307 -9200 9629 -9199
rect 9307 -9520 9308 -9200
rect 9628 -9520 9629 -9200
rect 9307 -9521 9629 -9520
rect 8888 -9588 8984 -9572
rect 9900 -9572 9916 -9148
rect 9980 -9572 9996 -9148
rect 10912 -9148 11008 -9132
rect 10319 -9200 10641 -9199
rect 10319 -9520 10320 -9200
rect 10640 -9520 10641 -9200
rect 10319 -9521 10641 -9520
rect 9900 -9588 9996 -9572
rect 10912 -9572 10928 -9148
rect 10992 -9572 11008 -9148
rect 11924 -9148 12020 -9132
rect 11331 -9200 11653 -9199
rect 11331 -9520 11332 -9200
rect 11652 -9520 11653 -9200
rect 11331 -9521 11653 -9520
rect 10912 -9588 11008 -9572
rect 11924 -9572 11940 -9148
rect 12004 -9572 12020 -9148
rect 12936 -9148 13032 -9132
rect 12343 -9200 12665 -9199
rect 12343 -9520 12344 -9200
rect 12664 -9520 12665 -9200
rect 12343 -9521 12665 -9520
rect 11924 -9588 12020 -9572
rect 12936 -9572 12952 -9148
rect 13016 -9572 13032 -9148
rect 13948 -9148 14044 -9132
rect 13355 -9200 13677 -9199
rect 13355 -9520 13356 -9200
rect 13676 -9520 13677 -9200
rect 13355 -9521 13677 -9520
rect 12936 -9588 13032 -9572
rect 13948 -9572 13964 -9148
rect 14028 -9572 14044 -9148
rect 14960 -9148 15056 -9132
rect 14367 -9200 14689 -9199
rect 14367 -9520 14368 -9200
rect 14688 -9520 14689 -9200
rect 14367 -9521 14689 -9520
rect 13948 -9588 14044 -9572
rect 14960 -9572 14976 -9148
rect 15040 -9572 15056 -9148
rect 15972 -9148 16068 -9132
rect 15379 -9200 15701 -9199
rect 15379 -9520 15380 -9200
rect 15700 -9520 15701 -9200
rect 15379 -9521 15701 -9520
rect 14960 -9588 15056 -9572
rect 15972 -9572 15988 -9148
rect 16052 -9572 16068 -9148
rect 16984 -9148 17080 -9132
rect 16391 -9200 16713 -9199
rect 16391 -9520 16392 -9200
rect 16712 -9520 16713 -9200
rect 16391 -9521 16713 -9520
rect 15972 -9588 16068 -9572
rect 16984 -9572 17000 -9148
rect 17064 -9572 17080 -9148
rect 16984 -9588 17080 -9572
rect -16412 -9868 -16316 -9852
rect -17005 -9920 -16683 -9919
rect -17005 -10240 -17004 -9920
rect -16684 -10240 -16683 -9920
rect -17005 -10241 -16683 -10240
rect -16412 -10292 -16396 -9868
rect -16332 -10292 -16316 -9868
rect -15400 -9868 -15304 -9852
rect -15993 -9920 -15671 -9919
rect -15993 -10240 -15992 -9920
rect -15672 -10240 -15671 -9920
rect -15993 -10241 -15671 -10240
rect -16412 -10308 -16316 -10292
rect -15400 -10292 -15384 -9868
rect -15320 -10292 -15304 -9868
rect -14388 -9868 -14292 -9852
rect -14981 -9920 -14659 -9919
rect -14981 -10240 -14980 -9920
rect -14660 -10240 -14659 -9920
rect -14981 -10241 -14659 -10240
rect -15400 -10308 -15304 -10292
rect -14388 -10292 -14372 -9868
rect -14308 -10292 -14292 -9868
rect -13376 -9868 -13280 -9852
rect -13969 -9920 -13647 -9919
rect -13969 -10240 -13968 -9920
rect -13648 -10240 -13647 -9920
rect -13969 -10241 -13647 -10240
rect -14388 -10308 -14292 -10292
rect -13376 -10292 -13360 -9868
rect -13296 -10292 -13280 -9868
rect -12364 -9868 -12268 -9852
rect -12957 -9920 -12635 -9919
rect -12957 -10240 -12956 -9920
rect -12636 -10240 -12635 -9920
rect -12957 -10241 -12635 -10240
rect -13376 -10308 -13280 -10292
rect -12364 -10292 -12348 -9868
rect -12284 -10292 -12268 -9868
rect -11352 -9868 -11256 -9852
rect -11945 -9920 -11623 -9919
rect -11945 -10240 -11944 -9920
rect -11624 -10240 -11623 -9920
rect -11945 -10241 -11623 -10240
rect -12364 -10308 -12268 -10292
rect -11352 -10292 -11336 -9868
rect -11272 -10292 -11256 -9868
rect -10340 -9868 -10244 -9852
rect -10933 -9920 -10611 -9919
rect -10933 -10240 -10932 -9920
rect -10612 -10240 -10611 -9920
rect -10933 -10241 -10611 -10240
rect -11352 -10308 -11256 -10292
rect -10340 -10292 -10324 -9868
rect -10260 -10292 -10244 -9868
rect -9328 -9868 -9232 -9852
rect -9921 -9920 -9599 -9919
rect -9921 -10240 -9920 -9920
rect -9600 -10240 -9599 -9920
rect -9921 -10241 -9599 -10240
rect -10340 -10308 -10244 -10292
rect -9328 -10292 -9312 -9868
rect -9248 -10292 -9232 -9868
rect -8316 -9868 -8220 -9852
rect -8909 -9920 -8587 -9919
rect -8909 -10240 -8908 -9920
rect -8588 -10240 -8587 -9920
rect -8909 -10241 -8587 -10240
rect -9328 -10308 -9232 -10292
rect -8316 -10292 -8300 -9868
rect -8236 -10292 -8220 -9868
rect -7304 -9868 -7208 -9852
rect -7897 -9920 -7575 -9919
rect -7897 -10240 -7896 -9920
rect -7576 -10240 -7575 -9920
rect -7897 -10241 -7575 -10240
rect -8316 -10308 -8220 -10292
rect -7304 -10292 -7288 -9868
rect -7224 -10292 -7208 -9868
rect -6292 -9868 -6196 -9852
rect -6885 -9920 -6563 -9919
rect -6885 -10240 -6884 -9920
rect -6564 -10240 -6563 -9920
rect -6885 -10241 -6563 -10240
rect -7304 -10308 -7208 -10292
rect -6292 -10292 -6276 -9868
rect -6212 -10292 -6196 -9868
rect -5280 -9868 -5184 -9852
rect -5873 -9920 -5551 -9919
rect -5873 -10240 -5872 -9920
rect -5552 -10240 -5551 -9920
rect -5873 -10241 -5551 -10240
rect -6292 -10308 -6196 -10292
rect -5280 -10292 -5264 -9868
rect -5200 -10292 -5184 -9868
rect -4268 -9868 -4172 -9852
rect -4861 -9920 -4539 -9919
rect -4861 -10240 -4860 -9920
rect -4540 -10240 -4539 -9920
rect -4861 -10241 -4539 -10240
rect -5280 -10308 -5184 -10292
rect -4268 -10292 -4252 -9868
rect -4188 -10292 -4172 -9868
rect -3256 -9868 -3160 -9852
rect -3849 -9920 -3527 -9919
rect -3849 -10240 -3848 -9920
rect -3528 -10240 -3527 -9920
rect -3849 -10241 -3527 -10240
rect -4268 -10308 -4172 -10292
rect -3256 -10292 -3240 -9868
rect -3176 -10292 -3160 -9868
rect -2244 -9868 -2148 -9852
rect -2837 -9920 -2515 -9919
rect -2837 -10240 -2836 -9920
rect -2516 -10240 -2515 -9920
rect -2837 -10241 -2515 -10240
rect -3256 -10308 -3160 -10292
rect -2244 -10292 -2228 -9868
rect -2164 -10292 -2148 -9868
rect -1232 -9868 -1136 -9852
rect -1825 -9920 -1503 -9919
rect -1825 -10240 -1824 -9920
rect -1504 -10240 -1503 -9920
rect -1825 -10241 -1503 -10240
rect -2244 -10308 -2148 -10292
rect -1232 -10292 -1216 -9868
rect -1152 -10292 -1136 -9868
rect -220 -9868 -124 -9852
rect -813 -9920 -491 -9919
rect -813 -10240 -812 -9920
rect -492 -10240 -491 -9920
rect -813 -10241 -491 -10240
rect -1232 -10308 -1136 -10292
rect -220 -10292 -204 -9868
rect -140 -10292 -124 -9868
rect 792 -9868 888 -9852
rect 199 -9920 521 -9919
rect 199 -10240 200 -9920
rect 520 -10240 521 -9920
rect 199 -10241 521 -10240
rect -220 -10308 -124 -10292
rect 792 -10292 808 -9868
rect 872 -10292 888 -9868
rect 1804 -9868 1900 -9852
rect 1211 -9920 1533 -9919
rect 1211 -10240 1212 -9920
rect 1532 -10240 1533 -9920
rect 1211 -10241 1533 -10240
rect 792 -10308 888 -10292
rect 1804 -10292 1820 -9868
rect 1884 -10292 1900 -9868
rect 2816 -9868 2912 -9852
rect 2223 -9920 2545 -9919
rect 2223 -10240 2224 -9920
rect 2544 -10240 2545 -9920
rect 2223 -10241 2545 -10240
rect 1804 -10308 1900 -10292
rect 2816 -10292 2832 -9868
rect 2896 -10292 2912 -9868
rect 3828 -9868 3924 -9852
rect 3235 -9920 3557 -9919
rect 3235 -10240 3236 -9920
rect 3556 -10240 3557 -9920
rect 3235 -10241 3557 -10240
rect 2816 -10308 2912 -10292
rect 3828 -10292 3844 -9868
rect 3908 -10292 3924 -9868
rect 4840 -9868 4936 -9852
rect 4247 -9920 4569 -9919
rect 4247 -10240 4248 -9920
rect 4568 -10240 4569 -9920
rect 4247 -10241 4569 -10240
rect 3828 -10308 3924 -10292
rect 4840 -10292 4856 -9868
rect 4920 -10292 4936 -9868
rect 5852 -9868 5948 -9852
rect 5259 -9920 5581 -9919
rect 5259 -10240 5260 -9920
rect 5580 -10240 5581 -9920
rect 5259 -10241 5581 -10240
rect 4840 -10308 4936 -10292
rect 5852 -10292 5868 -9868
rect 5932 -10292 5948 -9868
rect 6864 -9868 6960 -9852
rect 6271 -9920 6593 -9919
rect 6271 -10240 6272 -9920
rect 6592 -10240 6593 -9920
rect 6271 -10241 6593 -10240
rect 5852 -10308 5948 -10292
rect 6864 -10292 6880 -9868
rect 6944 -10292 6960 -9868
rect 7876 -9868 7972 -9852
rect 7283 -9920 7605 -9919
rect 7283 -10240 7284 -9920
rect 7604 -10240 7605 -9920
rect 7283 -10241 7605 -10240
rect 6864 -10308 6960 -10292
rect 7876 -10292 7892 -9868
rect 7956 -10292 7972 -9868
rect 8888 -9868 8984 -9852
rect 8295 -9920 8617 -9919
rect 8295 -10240 8296 -9920
rect 8616 -10240 8617 -9920
rect 8295 -10241 8617 -10240
rect 7876 -10308 7972 -10292
rect 8888 -10292 8904 -9868
rect 8968 -10292 8984 -9868
rect 9900 -9868 9996 -9852
rect 9307 -9920 9629 -9919
rect 9307 -10240 9308 -9920
rect 9628 -10240 9629 -9920
rect 9307 -10241 9629 -10240
rect 8888 -10308 8984 -10292
rect 9900 -10292 9916 -9868
rect 9980 -10292 9996 -9868
rect 10912 -9868 11008 -9852
rect 10319 -9920 10641 -9919
rect 10319 -10240 10320 -9920
rect 10640 -10240 10641 -9920
rect 10319 -10241 10641 -10240
rect 9900 -10308 9996 -10292
rect 10912 -10292 10928 -9868
rect 10992 -10292 11008 -9868
rect 11924 -9868 12020 -9852
rect 11331 -9920 11653 -9919
rect 11331 -10240 11332 -9920
rect 11652 -10240 11653 -9920
rect 11331 -10241 11653 -10240
rect 10912 -10308 11008 -10292
rect 11924 -10292 11940 -9868
rect 12004 -10292 12020 -9868
rect 12936 -9868 13032 -9852
rect 12343 -9920 12665 -9919
rect 12343 -10240 12344 -9920
rect 12664 -10240 12665 -9920
rect 12343 -10241 12665 -10240
rect 11924 -10308 12020 -10292
rect 12936 -10292 12952 -9868
rect 13016 -10292 13032 -9868
rect 13948 -9868 14044 -9852
rect 13355 -9920 13677 -9919
rect 13355 -10240 13356 -9920
rect 13676 -10240 13677 -9920
rect 13355 -10241 13677 -10240
rect 12936 -10308 13032 -10292
rect 13948 -10292 13964 -9868
rect 14028 -10292 14044 -9868
rect 14960 -9868 15056 -9852
rect 14367 -9920 14689 -9919
rect 14367 -10240 14368 -9920
rect 14688 -10240 14689 -9920
rect 14367 -10241 14689 -10240
rect 13948 -10308 14044 -10292
rect 14960 -10292 14976 -9868
rect 15040 -10292 15056 -9868
rect 15972 -9868 16068 -9852
rect 15379 -9920 15701 -9919
rect 15379 -10240 15380 -9920
rect 15700 -10240 15701 -9920
rect 15379 -10241 15701 -10240
rect 14960 -10308 15056 -10292
rect 15972 -10292 15988 -9868
rect 16052 -10292 16068 -9868
rect 16984 -9868 17080 -9852
rect 16391 -9920 16713 -9919
rect 16391 -10240 16392 -9920
rect 16712 -10240 16713 -9920
rect 16391 -10241 16713 -10240
rect 15972 -10308 16068 -10292
rect 16984 -10292 17000 -9868
rect 17064 -10292 17080 -9868
rect 16984 -10308 17080 -10292
rect -16412 -10588 -16316 -10572
rect -17005 -10640 -16683 -10639
rect -17005 -10960 -17004 -10640
rect -16684 -10960 -16683 -10640
rect -17005 -10961 -16683 -10960
rect -16412 -11012 -16396 -10588
rect -16332 -11012 -16316 -10588
rect -15400 -10588 -15304 -10572
rect -15993 -10640 -15671 -10639
rect -15993 -10960 -15992 -10640
rect -15672 -10960 -15671 -10640
rect -15993 -10961 -15671 -10960
rect -16412 -11028 -16316 -11012
rect -15400 -11012 -15384 -10588
rect -15320 -11012 -15304 -10588
rect -14388 -10588 -14292 -10572
rect -14981 -10640 -14659 -10639
rect -14981 -10960 -14980 -10640
rect -14660 -10960 -14659 -10640
rect -14981 -10961 -14659 -10960
rect -15400 -11028 -15304 -11012
rect -14388 -11012 -14372 -10588
rect -14308 -11012 -14292 -10588
rect -13376 -10588 -13280 -10572
rect -13969 -10640 -13647 -10639
rect -13969 -10960 -13968 -10640
rect -13648 -10960 -13647 -10640
rect -13969 -10961 -13647 -10960
rect -14388 -11028 -14292 -11012
rect -13376 -11012 -13360 -10588
rect -13296 -11012 -13280 -10588
rect -12364 -10588 -12268 -10572
rect -12957 -10640 -12635 -10639
rect -12957 -10960 -12956 -10640
rect -12636 -10960 -12635 -10640
rect -12957 -10961 -12635 -10960
rect -13376 -11028 -13280 -11012
rect -12364 -11012 -12348 -10588
rect -12284 -11012 -12268 -10588
rect -11352 -10588 -11256 -10572
rect -11945 -10640 -11623 -10639
rect -11945 -10960 -11944 -10640
rect -11624 -10960 -11623 -10640
rect -11945 -10961 -11623 -10960
rect -12364 -11028 -12268 -11012
rect -11352 -11012 -11336 -10588
rect -11272 -11012 -11256 -10588
rect -10340 -10588 -10244 -10572
rect -10933 -10640 -10611 -10639
rect -10933 -10960 -10932 -10640
rect -10612 -10960 -10611 -10640
rect -10933 -10961 -10611 -10960
rect -11352 -11028 -11256 -11012
rect -10340 -11012 -10324 -10588
rect -10260 -11012 -10244 -10588
rect -9328 -10588 -9232 -10572
rect -9921 -10640 -9599 -10639
rect -9921 -10960 -9920 -10640
rect -9600 -10960 -9599 -10640
rect -9921 -10961 -9599 -10960
rect -10340 -11028 -10244 -11012
rect -9328 -11012 -9312 -10588
rect -9248 -11012 -9232 -10588
rect -8316 -10588 -8220 -10572
rect -8909 -10640 -8587 -10639
rect -8909 -10960 -8908 -10640
rect -8588 -10960 -8587 -10640
rect -8909 -10961 -8587 -10960
rect -9328 -11028 -9232 -11012
rect -8316 -11012 -8300 -10588
rect -8236 -11012 -8220 -10588
rect -7304 -10588 -7208 -10572
rect -7897 -10640 -7575 -10639
rect -7897 -10960 -7896 -10640
rect -7576 -10960 -7575 -10640
rect -7897 -10961 -7575 -10960
rect -8316 -11028 -8220 -11012
rect -7304 -11012 -7288 -10588
rect -7224 -11012 -7208 -10588
rect -6292 -10588 -6196 -10572
rect -6885 -10640 -6563 -10639
rect -6885 -10960 -6884 -10640
rect -6564 -10960 -6563 -10640
rect -6885 -10961 -6563 -10960
rect -7304 -11028 -7208 -11012
rect -6292 -11012 -6276 -10588
rect -6212 -11012 -6196 -10588
rect -5280 -10588 -5184 -10572
rect -5873 -10640 -5551 -10639
rect -5873 -10960 -5872 -10640
rect -5552 -10960 -5551 -10640
rect -5873 -10961 -5551 -10960
rect -6292 -11028 -6196 -11012
rect -5280 -11012 -5264 -10588
rect -5200 -11012 -5184 -10588
rect -4268 -10588 -4172 -10572
rect -4861 -10640 -4539 -10639
rect -4861 -10960 -4860 -10640
rect -4540 -10960 -4539 -10640
rect -4861 -10961 -4539 -10960
rect -5280 -11028 -5184 -11012
rect -4268 -11012 -4252 -10588
rect -4188 -11012 -4172 -10588
rect -3256 -10588 -3160 -10572
rect -3849 -10640 -3527 -10639
rect -3849 -10960 -3848 -10640
rect -3528 -10960 -3527 -10640
rect -3849 -10961 -3527 -10960
rect -4268 -11028 -4172 -11012
rect -3256 -11012 -3240 -10588
rect -3176 -11012 -3160 -10588
rect -2244 -10588 -2148 -10572
rect -2837 -10640 -2515 -10639
rect -2837 -10960 -2836 -10640
rect -2516 -10960 -2515 -10640
rect -2837 -10961 -2515 -10960
rect -3256 -11028 -3160 -11012
rect -2244 -11012 -2228 -10588
rect -2164 -11012 -2148 -10588
rect -1232 -10588 -1136 -10572
rect -1825 -10640 -1503 -10639
rect -1825 -10960 -1824 -10640
rect -1504 -10960 -1503 -10640
rect -1825 -10961 -1503 -10960
rect -2244 -11028 -2148 -11012
rect -1232 -11012 -1216 -10588
rect -1152 -11012 -1136 -10588
rect -220 -10588 -124 -10572
rect -813 -10640 -491 -10639
rect -813 -10960 -812 -10640
rect -492 -10960 -491 -10640
rect -813 -10961 -491 -10960
rect -1232 -11028 -1136 -11012
rect -220 -11012 -204 -10588
rect -140 -11012 -124 -10588
rect 792 -10588 888 -10572
rect 199 -10640 521 -10639
rect 199 -10960 200 -10640
rect 520 -10960 521 -10640
rect 199 -10961 521 -10960
rect -220 -11028 -124 -11012
rect 792 -11012 808 -10588
rect 872 -11012 888 -10588
rect 1804 -10588 1900 -10572
rect 1211 -10640 1533 -10639
rect 1211 -10960 1212 -10640
rect 1532 -10960 1533 -10640
rect 1211 -10961 1533 -10960
rect 792 -11028 888 -11012
rect 1804 -11012 1820 -10588
rect 1884 -11012 1900 -10588
rect 2816 -10588 2912 -10572
rect 2223 -10640 2545 -10639
rect 2223 -10960 2224 -10640
rect 2544 -10960 2545 -10640
rect 2223 -10961 2545 -10960
rect 1804 -11028 1900 -11012
rect 2816 -11012 2832 -10588
rect 2896 -11012 2912 -10588
rect 3828 -10588 3924 -10572
rect 3235 -10640 3557 -10639
rect 3235 -10960 3236 -10640
rect 3556 -10960 3557 -10640
rect 3235 -10961 3557 -10960
rect 2816 -11028 2912 -11012
rect 3828 -11012 3844 -10588
rect 3908 -11012 3924 -10588
rect 4840 -10588 4936 -10572
rect 4247 -10640 4569 -10639
rect 4247 -10960 4248 -10640
rect 4568 -10960 4569 -10640
rect 4247 -10961 4569 -10960
rect 3828 -11028 3924 -11012
rect 4840 -11012 4856 -10588
rect 4920 -11012 4936 -10588
rect 5852 -10588 5948 -10572
rect 5259 -10640 5581 -10639
rect 5259 -10960 5260 -10640
rect 5580 -10960 5581 -10640
rect 5259 -10961 5581 -10960
rect 4840 -11028 4936 -11012
rect 5852 -11012 5868 -10588
rect 5932 -11012 5948 -10588
rect 6864 -10588 6960 -10572
rect 6271 -10640 6593 -10639
rect 6271 -10960 6272 -10640
rect 6592 -10960 6593 -10640
rect 6271 -10961 6593 -10960
rect 5852 -11028 5948 -11012
rect 6864 -11012 6880 -10588
rect 6944 -11012 6960 -10588
rect 7876 -10588 7972 -10572
rect 7283 -10640 7605 -10639
rect 7283 -10960 7284 -10640
rect 7604 -10960 7605 -10640
rect 7283 -10961 7605 -10960
rect 6864 -11028 6960 -11012
rect 7876 -11012 7892 -10588
rect 7956 -11012 7972 -10588
rect 8888 -10588 8984 -10572
rect 8295 -10640 8617 -10639
rect 8295 -10960 8296 -10640
rect 8616 -10960 8617 -10640
rect 8295 -10961 8617 -10960
rect 7876 -11028 7972 -11012
rect 8888 -11012 8904 -10588
rect 8968 -11012 8984 -10588
rect 9900 -10588 9996 -10572
rect 9307 -10640 9629 -10639
rect 9307 -10960 9308 -10640
rect 9628 -10960 9629 -10640
rect 9307 -10961 9629 -10960
rect 8888 -11028 8984 -11012
rect 9900 -11012 9916 -10588
rect 9980 -11012 9996 -10588
rect 10912 -10588 11008 -10572
rect 10319 -10640 10641 -10639
rect 10319 -10960 10320 -10640
rect 10640 -10960 10641 -10640
rect 10319 -10961 10641 -10960
rect 9900 -11028 9996 -11012
rect 10912 -11012 10928 -10588
rect 10992 -11012 11008 -10588
rect 11924 -10588 12020 -10572
rect 11331 -10640 11653 -10639
rect 11331 -10960 11332 -10640
rect 11652 -10960 11653 -10640
rect 11331 -10961 11653 -10960
rect 10912 -11028 11008 -11012
rect 11924 -11012 11940 -10588
rect 12004 -11012 12020 -10588
rect 12936 -10588 13032 -10572
rect 12343 -10640 12665 -10639
rect 12343 -10960 12344 -10640
rect 12664 -10960 12665 -10640
rect 12343 -10961 12665 -10960
rect 11924 -11028 12020 -11012
rect 12936 -11012 12952 -10588
rect 13016 -11012 13032 -10588
rect 13948 -10588 14044 -10572
rect 13355 -10640 13677 -10639
rect 13355 -10960 13356 -10640
rect 13676 -10960 13677 -10640
rect 13355 -10961 13677 -10960
rect 12936 -11028 13032 -11012
rect 13948 -11012 13964 -10588
rect 14028 -11012 14044 -10588
rect 14960 -10588 15056 -10572
rect 14367 -10640 14689 -10639
rect 14367 -10960 14368 -10640
rect 14688 -10960 14689 -10640
rect 14367 -10961 14689 -10960
rect 13948 -11028 14044 -11012
rect 14960 -11012 14976 -10588
rect 15040 -11012 15056 -10588
rect 15972 -10588 16068 -10572
rect 15379 -10640 15701 -10639
rect 15379 -10960 15380 -10640
rect 15700 -10960 15701 -10640
rect 15379 -10961 15701 -10960
rect 14960 -11028 15056 -11012
rect 15972 -11012 15988 -10588
rect 16052 -11012 16068 -10588
rect 16984 -10588 17080 -10572
rect 16391 -10640 16713 -10639
rect 16391 -10960 16392 -10640
rect 16712 -10960 16713 -10640
rect 16391 -10961 16713 -10960
rect 15972 -11028 16068 -11012
rect 16984 -11012 17000 -10588
rect 17064 -11012 17080 -10588
rect 16984 -11028 17080 -11012
rect -16412 -11308 -16316 -11292
rect -17005 -11360 -16683 -11359
rect -17005 -11680 -17004 -11360
rect -16684 -11680 -16683 -11360
rect -17005 -11681 -16683 -11680
rect -16412 -11732 -16396 -11308
rect -16332 -11732 -16316 -11308
rect -15400 -11308 -15304 -11292
rect -15993 -11360 -15671 -11359
rect -15993 -11680 -15992 -11360
rect -15672 -11680 -15671 -11360
rect -15993 -11681 -15671 -11680
rect -16412 -11748 -16316 -11732
rect -15400 -11732 -15384 -11308
rect -15320 -11732 -15304 -11308
rect -14388 -11308 -14292 -11292
rect -14981 -11360 -14659 -11359
rect -14981 -11680 -14980 -11360
rect -14660 -11680 -14659 -11360
rect -14981 -11681 -14659 -11680
rect -15400 -11748 -15304 -11732
rect -14388 -11732 -14372 -11308
rect -14308 -11732 -14292 -11308
rect -13376 -11308 -13280 -11292
rect -13969 -11360 -13647 -11359
rect -13969 -11680 -13968 -11360
rect -13648 -11680 -13647 -11360
rect -13969 -11681 -13647 -11680
rect -14388 -11748 -14292 -11732
rect -13376 -11732 -13360 -11308
rect -13296 -11732 -13280 -11308
rect -12364 -11308 -12268 -11292
rect -12957 -11360 -12635 -11359
rect -12957 -11680 -12956 -11360
rect -12636 -11680 -12635 -11360
rect -12957 -11681 -12635 -11680
rect -13376 -11748 -13280 -11732
rect -12364 -11732 -12348 -11308
rect -12284 -11732 -12268 -11308
rect -11352 -11308 -11256 -11292
rect -11945 -11360 -11623 -11359
rect -11945 -11680 -11944 -11360
rect -11624 -11680 -11623 -11360
rect -11945 -11681 -11623 -11680
rect -12364 -11748 -12268 -11732
rect -11352 -11732 -11336 -11308
rect -11272 -11732 -11256 -11308
rect -10340 -11308 -10244 -11292
rect -10933 -11360 -10611 -11359
rect -10933 -11680 -10932 -11360
rect -10612 -11680 -10611 -11360
rect -10933 -11681 -10611 -11680
rect -11352 -11748 -11256 -11732
rect -10340 -11732 -10324 -11308
rect -10260 -11732 -10244 -11308
rect -9328 -11308 -9232 -11292
rect -9921 -11360 -9599 -11359
rect -9921 -11680 -9920 -11360
rect -9600 -11680 -9599 -11360
rect -9921 -11681 -9599 -11680
rect -10340 -11748 -10244 -11732
rect -9328 -11732 -9312 -11308
rect -9248 -11732 -9232 -11308
rect -8316 -11308 -8220 -11292
rect -8909 -11360 -8587 -11359
rect -8909 -11680 -8908 -11360
rect -8588 -11680 -8587 -11360
rect -8909 -11681 -8587 -11680
rect -9328 -11748 -9232 -11732
rect -8316 -11732 -8300 -11308
rect -8236 -11732 -8220 -11308
rect -7304 -11308 -7208 -11292
rect -7897 -11360 -7575 -11359
rect -7897 -11680 -7896 -11360
rect -7576 -11680 -7575 -11360
rect -7897 -11681 -7575 -11680
rect -8316 -11748 -8220 -11732
rect -7304 -11732 -7288 -11308
rect -7224 -11732 -7208 -11308
rect -6292 -11308 -6196 -11292
rect -6885 -11360 -6563 -11359
rect -6885 -11680 -6884 -11360
rect -6564 -11680 -6563 -11360
rect -6885 -11681 -6563 -11680
rect -7304 -11748 -7208 -11732
rect -6292 -11732 -6276 -11308
rect -6212 -11732 -6196 -11308
rect -5280 -11308 -5184 -11292
rect -5873 -11360 -5551 -11359
rect -5873 -11680 -5872 -11360
rect -5552 -11680 -5551 -11360
rect -5873 -11681 -5551 -11680
rect -6292 -11748 -6196 -11732
rect -5280 -11732 -5264 -11308
rect -5200 -11732 -5184 -11308
rect -4268 -11308 -4172 -11292
rect -4861 -11360 -4539 -11359
rect -4861 -11680 -4860 -11360
rect -4540 -11680 -4539 -11360
rect -4861 -11681 -4539 -11680
rect -5280 -11748 -5184 -11732
rect -4268 -11732 -4252 -11308
rect -4188 -11732 -4172 -11308
rect -3256 -11308 -3160 -11292
rect -3849 -11360 -3527 -11359
rect -3849 -11680 -3848 -11360
rect -3528 -11680 -3527 -11360
rect -3849 -11681 -3527 -11680
rect -4268 -11748 -4172 -11732
rect -3256 -11732 -3240 -11308
rect -3176 -11732 -3160 -11308
rect -2244 -11308 -2148 -11292
rect -2837 -11360 -2515 -11359
rect -2837 -11680 -2836 -11360
rect -2516 -11680 -2515 -11360
rect -2837 -11681 -2515 -11680
rect -3256 -11748 -3160 -11732
rect -2244 -11732 -2228 -11308
rect -2164 -11732 -2148 -11308
rect -1232 -11308 -1136 -11292
rect -1825 -11360 -1503 -11359
rect -1825 -11680 -1824 -11360
rect -1504 -11680 -1503 -11360
rect -1825 -11681 -1503 -11680
rect -2244 -11748 -2148 -11732
rect -1232 -11732 -1216 -11308
rect -1152 -11732 -1136 -11308
rect -220 -11308 -124 -11292
rect -813 -11360 -491 -11359
rect -813 -11680 -812 -11360
rect -492 -11680 -491 -11360
rect -813 -11681 -491 -11680
rect -1232 -11748 -1136 -11732
rect -220 -11732 -204 -11308
rect -140 -11732 -124 -11308
rect 792 -11308 888 -11292
rect 199 -11360 521 -11359
rect 199 -11680 200 -11360
rect 520 -11680 521 -11360
rect 199 -11681 521 -11680
rect -220 -11748 -124 -11732
rect 792 -11732 808 -11308
rect 872 -11732 888 -11308
rect 1804 -11308 1900 -11292
rect 1211 -11360 1533 -11359
rect 1211 -11680 1212 -11360
rect 1532 -11680 1533 -11360
rect 1211 -11681 1533 -11680
rect 792 -11748 888 -11732
rect 1804 -11732 1820 -11308
rect 1884 -11732 1900 -11308
rect 2816 -11308 2912 -11292
rect 2223 -11360 2545 -11359
rect 2223 -11680 2224 -11360
rect 2544 -11680 2545 -11360
rect 2223 -11681 2545 -11680
rect 1804 -11748 1900 -11732
rect 2816 -11732 2832 -11308
rect 2896 -11732 2912 -11308
rect 3828 -11308 3924 -11292
rect 3235 -11360 3557 -11359
rect 3235 -11680 3236 -11360
rect 3556 -11680 3557 -11360
rect 3235 -11681 3557 -11680
rect 2816 -11748 2912 -11732
rect 3828 -11732 3844 -11308
rect 3908 -11732 3924 -11308
rect 4840 -11308 4936 -11292
rect 4247 -11360 4569 -11359
rect 4247 -11680 4248 -11360
rect 4568 -11680 4569 -11360
rect 4247 -11681 4569 -11680
rect 3828 -11748 3924 -11732
rect 4840 -11732 4856 -11308
rect 4920 -11732 4936 -11308
rect 5852 -11308 5948 -11292
rect 5259 -11360 5581 -11359
rect 5259 -11680 5260 -11360
rect 5580 -11680 5581 -11360
rect 5259 -11681 5581 -11680
rect 4840 -11748 4936 -11732
rect 5852 -11732 5868 -11308
rect 5932 -11732 5948 -11308
rect 6864 -11308 6960 -11292
rect 6271 -11360 6593 -11359
rect 6271 -11680 6272 -11360
rect 6592 -11680 6593 -11360
rect 6271 -11681 6593 -11680
rect 5852 -11748 5948 -11732
rect 6864 -11732 6880 -11308
rect 6944 -11732 6960 -11308
rect 7876 -11308 7972 -11292
rect 7283 -11360 7605 -11359
rect 7283 -11680 7284 -11360
rect 7604 -11680 7605 -11360
rect 7283 -11681 7605 -11680
rect 6864 -11748 6960 -11732
rect 7876 -11732 7892 -11308
rect 7956 -11732 7972 -11308
rect 8888 -11308 8984 -11292
rect 8295 -11360 8617 -11359
rect 8295 -11680 8296 -11360
rect 8616 -11680 8617 -11360
rect 8295 -11681 8617 -11680
rect 7876 -11748 7972 -11732
rect 8888 -11732 8904 -11308
rect 8968 -11732 8984 -11308
rect 9900 -11308 9996 -11292
rect 9307 -11360 9629 -11359
rect 9307 -11680 9308 -11360
rect 9628 -11680 9629 -11360
rect 9307 -11681 9629 -11680
rect 8888 -11748 8984 -11732
rect 9900 -11732 9916 -11308
rect 9980 -11732 9996 -11308
rect 10912 -11308 11008 -11292
rect 10319 -11360 10641 -11359
rect 10319 -11680 10320 -11360
rect 10640 -11680 10641 -11360
rect 10319 -11681 10641 -11680
rect 9900 -11748 9996 -11732
rect 10912 -11732 10928 -11308
rect 10992 -11732 11008 -11308
rect 11924 -11308 12020 -11292
rect 11331 -11360 11653 -11359
rect 11331 -11680 11332 -11360
rect 11652 -11680 11653 -11360
rect 11331 -11681 11653 -11680
rect 10912 -11748 11008 -11732
rect 11924 -11732 11940 -11308
rect 12004 -11732 12020 -11308
rect 12936 -11308 13032 -11292
rect 12343 -11360 12665 -11359
rect 12343 -11680 12344 -11360
rect 12664 -11680 12665 -11360
rect 12343 -11681 12665 -11680
rect 11924 -11748 12020 -11732
rect 12936 -11732 12952 -11308
rect 13016 -11732 13032 -11308
rect 13948 -11308 14044 -11292
rect 13355 -11360 13677 -11359
rect 13355 -11680 13356 -11360
rect 13676 -11680 13677 -11360
rect 13355 -11681 13677 -11680
rect 12936 -11748 13032 -11732
rect 13948 -11732 13964 -11308
rect 14028 -11732 14044 -11308
rect 14960 -11308 15056 -11292
rect 14367 -11360 14689 -11359
rect 14367 -11680 14368 -11360
rect 14688 -11680 14689 -11360
rect 14367 -11681 14689 -11680
rect 13948 -11748 14044 -11732
rect 14960 -11732 14976 -11308
rect 15040 -11732 15056 -11308
rect 15972 -11308 16068 -11292
rect 15379 -11360 15701 -11359
rect 15379 -11680 15380 -11360
rect 15700 -11680 15701 -11360
rect 15379 -11681 15701 -11680
rect 14960 -11748 15056 -11732
rect 15972 -11732 15988 -11308
rect 16052 -11732 16068 -11308
rect 16984 -11308 17080 -11292
rect 16391 -11360 16713 -11359
rect 16391 -11680 16392 -11360
rect 16712 -11680 16713 -11360
rect 16391 -11681 16713 -11680
rect 15972 -11748 16068 -11732
rect 16984 -11732 17000 -11308
rect 17064 -11732 17080 -11308
rect 16984 -11748 17080 -11732
<< properties >>
string FIXED_BBOX 16312 11280 16792 11760
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 34 ny 33 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
