magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -38 332 134 704
<< pwell >>
rect 5 38 91 255
<< psubdiff >>
rect 31 205 65 229
rect 31 122 65 171
rect 31 64 65 88
<< nsubdiff >>
rect 31 578 65 602
rect 31 492 65 544
rect 31 434 65 458
<< psubdiffcont >>
rect 31 171 65 205
rect 31 88 65 122
<< nsubdiffcont >>
rect 31 544 65 578
rect 31 458 65 492
<< locali >>
rect 0 649 31 683
rect 65 649 96 683
rect 18 578 78 649
rect 18 544 31 578
rect 65 544 78 578
rect 18 492 78 544
rect 18 458 31 492
rect 65 458 78 492
rect 18 441 78 458
rect 18 205 78 221
rect 18 171 31 205
rect 65 171 78 205
rect 18 122 78 171
rect 18 88 31 122
rect 65 88 78 122
rect 18 17 78 88
rect 0 -17 31 17
rect 65 -17 96 17
<< viali >>
rect 31 649 65 683
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
flabel metal1 s 0 617 96 666 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 0 0 96 49 0 FreeSans 200 0 0 0 VGND
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 96 666
<< end >>
