VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tsar_adc
  CLASS BLOCK ;
  FOREIGN tt_um_tsar_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.368000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 125.279999 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 18.559999 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 18.559999 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 31.230000 ;
    ANTENNADIFFAREA 830.561707 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 31.230000 ;
    ANTENNADIFFAREA 830.561707 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 69.000000 ;
    ANTENNADIFFAREA 555.876160 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 129.205 151.475 129.450 151.850 ;
        RECT 129.205 150.425 130.445 151.475 ;
      LAYER nwell ;
        RECT 130.865 150.600 132.725 152.040 ;
      LAYER pwell ;
        RECT 153.215 151.475 153.460 151.850 ;
        RECT 129.205 150.390 129.450 150.425 ;
      LAYER nwell ;
        RECT 112.800 144.015 115.260 149.765 ;
      LAYER pwell ;
        RECT 115.310 144.065 117.670 149.715 ;
      LAYER nwell ;
        RECT 117.720 144.015 120.180 149.760 ;
      LAYER pwell ;
        RECT 129.205 149.020 130.445 150.390 ;
        RECT 129.205 148.595 129.450 149.020 ;
        RECT 129.205 147.545 130.445 148.595 ;
        RECT 129.205 147.530 129.450 147.545 ;
        RECT 129.395 147.075 130.480 147.505 ;
      LAYER nwell ;
        RECT 112.800 144.010 120.180 144.015 ;
      LAYER pwell ;
        RECT 129.205 146.675 129.450 147.050 ;
        RECT 129.205 145.625 130.445 146.675 ;
        RECT 129.205 145.605 129.450 145.625 ;
        RECT 10.200 143.375 23.160 143.620 ;
        RECT 10.280 142.645 12.090 143.375 ;
        RECT 12.605 142.700 14.515 143.375 ;
        RECT 14.525 142.700 17.380 143.375 ;
        RECT 17.885 142.380 19.875 143.375 ;
        RECT 20.285 142.700 23.140 143.375 ;
        RECT 23.185 142.345 23.615 143.430 ;
        RECT 23.640 143.375 36.120 143.620 ;
        RECT 23.645 142.680 34.660 143.375 ;
        RECT 23.645 142.665 33.280 142.680 ;
        RECT 23.645 142.570 25.615 142.665 ;
        RECT 23.645 142.380 24.625 142.570 ;
        RECT 27.970 142.380 33.280 142.665 ;
        RECT 36.145 142.345 36.575 143.430 ;
        RECT 36.600 143.375 49.080 143.620 ;
        RECT 37.565 142.700 40.420 143.375 ;
        RECT 40.445 142.700 43.300 143.375 ;
        RECT 43.325 142.700 46.180 143.375 ;
        RECT 46.220 142.700 49.075 143.375 ;
        RECT 49.105 142.345 49.535 143.430 ;
        RECT 49.560 143.375 62.040 143.620 ;
        RECT 49.565 142.700 52.420 143.375 ;
        RECT 52.520 142.645 54.330 143.375 ;
        RECT 54.845 142.700 57.700 143.375 ;
        RECT 59.180 142.700 62.035 143.375 ;
        RECT 62.065 142.345 62.495 143.430 ;
        RECT 62.520 143.375 69.720 143.620 ;
        RECT 62.525 142.700 65.380 143.375 ;
        RECT 65.405 142.720 67.315 143.375 ;
        RECT 65.440 142.700 67.315 142.720 ;
        RECT 67.830 142.645 69.640 143.375 ;
      LAYER nwell ;
        RECT 28.280 141.970 29.360 142.065 ;
        RECT 28.280 141.960 33.290 141.970 ;
        RECT 10.010 138.620 69.910 141.960 ;
        RECT 112.800 139.655 124.570 144.010 ;
      LAYER pwell ;
        RECT 129.205 143.215 130.445 145.605 ;
        RECT 129.205 143.210 129.450 143.215 ;
        RECT 129.395 142.755 130.480 143.185 ;
      LAYER nwell ;
        RECT 115.260 139.650 124.570 139.655 ;
        RECT 16.760 138.610 21.770 138.620 ;
        RECT 34.630 138.610 39.640 138.620 ;
        RECT 50.950 138.610 55.960 138.620 ;
        RECT 16.760 138.515 17.840 138.610 ;
        RECT 38.560 138.515 39.640 138.610 ;
        RECT 54.880 138.515 55.960 138.610 ;
      LAYER pwell ;
        RECT 12.125 138.010 13.105 138.200 ;
        RECT 10.280 137.205 12.090 137.935 ;
        RECT 12.125 137.915 14.095 138.010 ;
        RECT 16.450 137.915 21.760 138.200 ;
        RECT 12.125 137.900 21.760 137.915 ;
        RECT 12.125 137.205 23.140 137.900 ;
        RECT 10.200 136.960 23.160 137.205 ;
        RECT 23.185 137.150 23.615 138.235 ;
        RECT 24.045 137.205 26.035 138.200 ;
        RECT 26.045 137.205 28.900 137.880 ;
        RECT 29.000 137.205 30.810 137.935 ;
        RECT 34.640 137.915 39.950 138.200 ;
        RECT 43.295 138.010 44.275 138.200 ;
        RECT 42.305 137.915 44.275 138.010 ;
        RECT 34.640 137.900 44.275 137.915 ;
        RECT 31.325 137.205 33.235 137.880 ;
        RECT 33.260 137.205 44.275 137.900 ;
        RECT 44.285 137.205 46.195 137.880 ;
        RECT 46.220 137.205 49.075 137.880 ;
        RECT 23.640 136.960 49.080 137.205 ;
        RECT 49.105 137.150 49.535 138.235 ;
        RECT 50.960 137.915 56.270 138.200 ;
        RECT 59.615 138.010 60.595 138.200 ;
        RECT 58.625 137.915 60.595 138.010 ;
        RECT 50.960 137.900 60.595 137.915 ;
        RECT 49.580 137.205 60.595 137.900 ;
        RECT 62.060 137.205 64.915 137.880 ;
        RECT 64.940 137.205 67.795 137.880 ;
        RECT 67.830 137.205 69.640 137.935 ;
        RECT 49.560 136.960 69.720 137.205 ;
        RECT 10.200 136.715 36.120 136.960 ;
        RECT 10.280 135.985 12.090 136.715 ;
        RECT 12.125 136.060 14.035 136.715 ;
        RECT 12.125 136.040 14.000 136.060 ;
        RECT 14.045 136.020 25.060 136.715 ;
        RECT 25.100 136.020 36.115 136.715 ;
        RECT 14.045 136.005 23.680 136.020 ;
        RECT 14.045 135.910 16.015 136.005 ;
        RECT 14.045 135.720 15.025 135.910 ;
        RECT 18.370 135.720 23.680 136.005 ;
        RECT 26.480 136.005 36.115 136.020 ;
        RECT 26.480 135.720 31.790 136.005 ;
        RECT 34.145 135.910 36.115 136.005 ;
        RECT 35.135 135.720 36.115 135.910 ;
        RECT 36.145 135.685 36.575 136.770 ;
        RECT 36.600 136.715 62.040 136.960 ;
        RECT 44.285 136.020 55.300 136.715 ;
        RECT 56.300 136.040 59.155 136.715 ;
        RECT 59.180 136.040 62.035 136.715 ;
        RECT 44.285 136.005 53.920 136.020 ;
        RECT 44.285 135.910 46.255 136.005 ;
        RECT 44.285 135.720 45.265 135.910 ;
        RECT 48.610 135.720 53.920 136.005 ;
        RECT 62.065 135.685 62.495 136.770 ;
        RECT 62.520 136.715 69.720 136.960 ;
        RECT 62.670 135.590 64.800 136.715 ;
        RECT 64.925 136.040 67.780 136.715 ;
        RECT 67.830 135.985 69.640 136.715 ;
        RECT 62.670 135.510 63.615 135.590 ;
      LAYER nwell ;
        RECT 18.680 135.310 19.760 135.405 ;
        RECT 30.400 135.310 31.480 135.405 ;
        RECT 18.680 135.300 23.690 135.310 ;
        RECT 26.470 135.300 31.480 135.310 ;
        RECT 48.920 135.310 50.000 135.405 ;
        RECT 48.920 135.300 53.930 135.310 ;
        RECT 10.010 131.960 69.910 135.300 ;
      LAYER pwell ;
        RECT 112.850 133.955 115.210 139.605 ;
      LAYER nwell ;
        RECT 115.260 133.905 117.720 139.650 ;
      LAYER pwell ;
        RECT 117.770 133.950 120.130 139.600 ;
      LAYER nwell ;
        RECT 120.180 133.900 124.570 139.650 ;
      LAYER pwell ;
        RECT 129.205 142.710 129.450 142.730 ;
        RECT 124.620 133.950 128.910 139.600 ;
        RECT 129.205 138.505 130.445 142.710 ;
        RECT 129.205 138.390 129.450 138.505 ;
        RECT 129.205 134.185 130.445 138.390 ;
        RECT 129.205 134.090 129.450 134.185 ;
      LAYER nwell ;
        RECT 130.865 133.900 134.205 150.600 ;
      LAYER pwell ;
        RECT 153.215 150.425 154.455 151.475 ;
      LAYER nwell ;
        RECT 154.875 150.600 156.735 152.040 ;
      LAYER pwell ;
        RECT 177.225 151.475 177.470 151.850 ;
        RECT 135.620 150.360 135.865 150.410 ;
        RECT 134.625 148.990 135.865 150.360 ;
        RECT 153.215 150.390 153.460 150.425 ;
        RECT 135.620 148.595 135.865 148.990 ;
        RECT 134.625 147.545 135.865 148.595 ;
        RECT 135.620 147.530 135.865 147.545 ;
        RECT 134.590 147.075 135.675 147.505 ;
        RECT 135.620 146.675 135.865 147.050 ;
        RECT 134.625 145.625 135.865 146.675 ;
        RECT 135.620 145.605 135.865 145.625 ;
        RECT 134.625 143.215 135.865 145.605 ;
        RECT 135.620 143.210 135.865 143.215 ;
      LAYER nwell ;
        RECT 136.810 144.015 139.270 149.765 ;
      LAYER pwell ;
        RECT 139.320 144.065 141.680 149.715 ;
      LAYER nwell ;
        RECT 141.730 144.015 144.190 149.760 ;
      LAYER pwell ;
        RECT 153.215 149.020 154.455 150.390 ;
        RECT 153.215 148.595 153.460 149.020 ;
        RECT 153.215 147.545 154.455 148.595 ;
        RECT 153.215 147.530 153.460 147.545 ;
        RECT 153.405 147.075 154.490 147.505 ;
      LAYER nwell ;
        RECT 136.810 144.010 144.190 144.015 ;
      LAYER pwell ;
        RECT 153.215 146.675 153.460 147.050 ;
        RECT 153.215 145.625 154.455 146.675 ;
        RECT 153.215 145.605 153.460 145.625 ;
        RECT 134.590 142.755 135.675 143.185 ;
        RECT 135.620 142.710 135.865 142.730 ;
        RECT 134.625 138.505 135.865 142.710 ;
      LAYER nwell ;
        RECT 136.810 139.655 148.580 144.010 ;
      LAYER pwell ;
        RECT 153.215 143.215 154.455 145.605 ;
        RECT 153.215 143.210 153.460 143.215 ;
        RECT 153.405 142.755 154.490 143.185 ;
      LAYER nwell ;
        RECT 139.270 139.650 148.580 139.655 ;
      LAYER pwell ;
        RECT 135.620 138.390 135.865 138.505 ;
        RECT 134.625 134.185 135.865 138.390 ;
        RECT 135.620 134.090 135.865 134.185 ;
        RECT 136.860 133.955 139.220 139.605 ;
      LAYER nwell ;
        RECT 139.270 133.905 141.730 139.650 ;
      LAYER pwell ;
        RECT 141.780 133.950 144.140 139.600 ;
      LAYER nwell ;
        RECT 144.190 133.900 148.580 139.650 ;
      LAYER pwell ;
        RECT 153.215 142.710 153.460 142.730 ;
        RECT 148.630 133.950 152.920 139.600 ;
        RECT 153.215 138.505 154.455 142.710 ;
        RECT 153.215 138.390 153.460 138.505 ;
        RECT 153.215 134.185 154.455 138.390 ;
        RECT 153.215 134.090 153.460 134.185 ;
      LAYER nwell ;
        RECT 154.875 133.900 158.215 150.600 ;
      LAYER pwell ;
        RECT 177.225 150.425 178.465 151.475 ;
      LAYER nwell ;
        RECT 178.885 150.600 180.745 152.040 ;
      LAYER pwell ;
        RECT 201.235 151.475 201.480 151.850 ;
        RECT 159.630 150.360 159.875 150.410 ;
        RECT 158.635 148.990 159.875 150.360 ;
        RECT 177.225 150.390 177.470 150.425 ;
        RECT 159.630 148.595 159.875 148.990 ;
        RECT 158.635 147.545 159.875 148.595 ;
        RECT 159.630 147.530 159.875 147.545 ;
        RECT 158.600 147.075 159.685 147.505 ;
        RECT 159.630 146.675 159.875 147.050 ;
        RECT 158.635 145.625 159.875 146.675 ;
        RECT 159.630 145.605 159.875 145.625 ;
        RECT 158.635 143.215 159.875 145.605 ;
        RECT 159.630 143.210 159.875 143.215 ;
      LAYER nwell ;
        RECT 160.820 144.015 163.280 149.765 ;
      LAYER pwell ;
        RECT 163.330 144.065 165.690 149.715 ;
      LAYER nwell ;
        RECT 165.740 144.015 168.200 149.760 ;
      LAYER pwell ;
        RECT 177.225 149.020 178.465 150.390 ;
        RECT 177.225 148.595 177.470 149.020 ;
        RECT 177.225 147.545 178.465 148.595 ;
        RECT 177.225 147.530 177.470 147.545 ;
        RECT 177.415 147.075 178.500 147.505 ;
      LAYER nwell ;
        RECT 160.820 144.010 168.200 144.015 ;
      LAYER pwell ;
        RECT 177.225 146.675 177.470 147.050 ;
        RECT 177.225 145.625 178.465 146.675 ;
        RECT 177.225 145.605 177.470 145.625 ;
        RECT 158.600 142.755 159.685 143.185 ;
        RECT 159.630 142.710 159.875 142.730 ;
        RECT 158.635 138.505 159.875 142.710 ;
      LAYER nwell ;
        RECT 160.820 139.655 172.590 144.010 ;
      LAYER pwell ;
        RECT 177.225 143.215 178.465 145.605 ;
        RECT 177.225 143.210 177.470 143.215 ;
        RECT 177.415 142.755 178.500 143.185 ;
      LAYER nwell ;
        RECT 163.280 139.650 172.590 139.655 ;
      LAYER pwell ;
        RECT 159.630 138.390 159.875 138.505 ;
        RECT 158.635 134.185 159.875 138.390 ;
        RECT 159.630 134.090 159.875 134.185 ;
        RECT 160.870 133.955 163.230 139.605 ;
      LAYER nwell ;
        RECT 163.280 133.905 165.740 139.650 ;
      LAYER pwell ;
        RECT 165.790 133.950 168.150 139.600 ;
      LAYER nwell ;
        RECT 168.200 133.900 172.590 139.650 ;
      LAYER pwell ;
        RECT 177.225 142.710 177.470 142.730 ;
        RECT 172.640 133.950 176.930 139.600 ;
        RECT 177.225 138.505 178.465 142.710 ;
        RECT 177.225 138.390 177.470 138.505 ;
        RECT 177.225 134.185 178.465 138.390 ;
        RECT 177.225 134.090 177.470 134.185 ;
      LAYER nwell ;
        RECT 178.885 133.900 182.225 150.600 ;
      LAYER pwell ;
        RECT 201.235 150.425 202.475 151.475 ;
      LAYER nwell ;
        RECT 202.895 150.600 204.755 152.040 ;
      LAYER pwell ;
        RECT 225.245 151.475 225.490 151.850 ;
        RECT 183.640 150.360 183.885 150.410 ;
        RECT 182.645 148.990 183.885 150.360 ;
        RECT 201.235 150.390 201.480 150.425 ;
        RECT 183.640 148.595 183.885 148.990 ;
        RECT 182.645 147.545 183.885 148.595 ;
        RECT 183.640 147.530 183.885 147.545 ;
        RECT 182.610 147.075 183.695 147.505 ;
        RECT 183.640 146.675 183.885 147.050 ;
        RECT 182.645 145.625 183.885 146.675 ;
        RECT 183.640 145.605 183.885 145.625 ;
        RECT 182.645 143.215 183.885 145.605 ;
        RECT 183.640 143.210 183.885 143.215 ;
      LAYER nwell ;
        RECT 184.830 144.015 187.290 149.765 ;
      LAYER pwell ;
        RECT 187.340 144.065 189.700 149.715 ;
      LAYER nwell ;
        RECT 189.750 144.015 192.210 149.760 ;
      LAYER pwell ;
        RECT 201.235 149.020 202.475 150.390 ;
        RECT 201.235 148.595 201.480 149.020 ;
        RECT 201.235 147.545 202.475 148.595 ;
        RECT 201.235 147.530 201.480 147.545 ;
        RECT 201.425 147.075 202.510 147.505 ;
      LAYER nwell ;
        RECT 184.830 144.010 192.210 144.015 ;
      LAYER pwell ;
        RECT 201.235 146.675 201.480 147.050 ;
        RECT 201.235 145.625 202.475 146.675 ;
        RECT 201.235 145.605 201.480 145.625 ;
        RECT 182.610 142.755 183.695 143.185 ;
        RECT 183.640 142.710 183.885 142.730 ;
        RECT 182.645 138.505 183.885 142.710 ;
      LAYER nwell ;
        RECT 184.830 139.655 196.600 144.010 ;
      LAYER pwell ;
        RECT 201.235 143.215 202.475 145.605 ;
        RECT 201.235 143.210 201.480 143.215 ;
        RECT 201.425 142.755 202.510 143.185 ;
      LAYER nwell ;
        RECT 187.290 139.650 196.600 139.655 ;
      LAYER pwell ;
        RECT 183.640 138.390 183.885 138.505 ;
        RECT 182.645 134.185 183.885 138.390 ;
        RECT 183.640 134.090 183.885 134.185 ;
        RECT 184.880 133.955 187.240 139.605 ;
      LAYER nwell ;
        RECT 187.290 133.905 189.750 139.650 ;
      LAYER pwell ;
        RECT 189.800 133.950 192.160 139.600 ;
      LAYER nwell ;
        RECT 192.210 133.900 196.600 139.650 ;
      LAYER pwell ;
        RECT 201.235 142.710 201.480 142.730 ;
        RECT 196.650 133.950 200.940 139.600 ;
        RECT 201.235 138.505 202.475 142.710 ;
        RECT 201.235 138.390 201.480 138.505 ;
        RECT 201.235 134.185 202.475 138.390 ;
        RECT 201.235 134.090 201.480 134.185 ;
      LAYER nwell ;
        RECT 202.895 133.900 206.235 150.600 ;
      LAYER pwell ;
        RECT 225.245 150.425 226.485 151.475 ;
      LAYER nwell ;
        RECT 226.905 150.600 228.765 152.040 ;
      LAYER pwell ;
        RECT 249.260 151.475 249.505 151.850 ;
        RECT 207.650 150.360 207.895 150.410 ;
        RECT 206.655 148.990 207.895 150.360 ;
        RECT 225.245 150.390 225.490 150.425 ;
        RECT 207.650 148.595 207.895 148.990 ;
        RECT 206.655 147.545 207.895 148.595 ;
        RECT 207.650 147.530 207.895 147.545 ;
        RECT 206.620 147.075 207.705 147.505 ;
        RECT 207.650 146.675 207.895 147.050 ;
        RECT 206.655 145.625 207.895 146.675 ;
        RECT 207.650 145.605 207.895 145.625 ;
        RECT 206.655 143.215 207.895 145.605 ;
        RECT 207.650 143.210 207.895 143.215 ;
      LAYER nwell ;
        RECT 208.840 144.015 211.300 149.765 ;
      LAYER pwell ;
        RECT 211.350 144.065 213.710 149.715 ;
      LAYER nwell ;
        RECT 213.760 144.015 216.220 149.760 ;
      LAYER pwell ;
        RECT 225.245 149.020 226.485 150.390 ;
        RECT 225.245 148.595 225.490 149.020 ;
        RECT 225.245 147.545 226.485 148.595 ;
        RECT 225.245 147.530 225.490 147.545 ;
        RECT 225.435 147.075 226.520 147.505 ;
      LAYER nwell ;
        RECT 208.840 144.010 216.220 144.015 ;
      LAYER pwell ;
        RECT 225.245 146.675 225.490 147.050 ;
        RECT 225.245 145.625 226.485 146.675 ;
        RECT 225.245 145.605 225.490 145.625 ;
        RECT 206.620 142.755 207.705 143.185 ;
        RECT 207.650 142.710 207.895 142.730 ;
        RECT 206.655 138.505 207.895 142.710 ;
      LAYER nwell ;
        RECT 208.840 139.655 220.610 144.010 ;
      LAYER pwell ;
        RECT 225.245 143.215 226.485 145.605 ;
        RECT 225.245 143.210 225.490 143.215 ;
        RECT 225.435 142.755 226.520 143.185 ;
      LAYER nwell ;
        RECT 211.300 139.650 220.610 139.655 ;
      LAYER pwell ;
        RECT 207.650 138.390 207.895 138.505 ;
        RECT 206.655 134.185 207.895 138.390 ;
        RECT 207.650 134.090 207.895 134.185 ;
        RECT 208.890 133.955 211.250 139.605 ;
      LAYER nwell ;
        RECT 211.300 133.905 213.760 139.650 ;
      LAYER pwell ;
        RECT 213.810 133.950 216.170 139.600 ;
      LAYER nwell ;
        RECT 216.220 133.900 220.610 139.650 ;
      LAYER pwell ;
        RECT 225.245 142.710 225.490 142.730 ;
        RECT 220.660 133.950 224.950 139.600 ;
        RECT 225.245 138.505 226.485 142.710 ;
        RECT 225.245 138.390 225.490 138.505 ;
        RECT 225.245 134.185 226.485 138.390 ;
        RECT 225.245 134.090 225.490 134.185 ;
      LAYER nwell ;
        RECT 226.905 133.900 230.245 150.600 ;
      LAYER pwell ;
        RECT 249.260 150.425 250.500 151.475 ;
      LAYER nwell ;
        RECT 250.920 150.600 252.780 152.040 ;
      LAYER pwell ;
        RECT 273.315 151.475 273.560 151.850 ;
        RECT 231.660 150.360 231.905 150.410 ;
        RECT 230.665 148.990 231.905 150.360 ;
        RECT 249.260 150.390 249.505 150.425 ;
        RECT 231.660 148.595 231.905 148.990 ;
        RECT 230.665 147.545 231.905 148.595 ;
        RECT 231.660 147.530 231.905 147.545 ;
        RECT 230.630 147.075 231.715 147.505 ;
        RECT 231.660 146.675 231.905 147.050 ;
        RECT 230.665 145.625 231.905 146.675 ;
        RECT 231.660 145.605 231.905 145.625 ;
        RECT 230.665 143.215 231.905 145.605 ;
        RECT 231.660 143.210 231.905 143.215 ;
      LAYER nwell ;
        RECT 232.855 144.015 235.315 149.765 ;
      LAYER pwell ;
        RECT 235.365 144.065 237.725 149.715 ;
      LAYER nwell ;
        RECT 237.775 144.015 240.235 149.760 ;
      LAYER pwell ;
        RECT 249.260 149.020 250.500 150.390 ;
        RECT 249.260 148.595 249.505 149.020 ;
        RECT 249.260 147.545 250.500 148.595 ;
        RECT 249.260 147.530 249.505 147.545 ;
        RECT 249.450 147.075 250.535 147.505 ;
      LAYER nwell ;
        RECT 232.855 144.010 240.235 144.015 ;
      LAYER pwell ;
        RECT 249.260 146.675 249.505 147.050 ;
        RECT 249.260 145.625 250.500 146.675 ;
        RECT 249.260 145.605 249.505 145.625 ;
        RECT 230.630 142.755 231.715 143.185 ;
        RECT 231.660 142.710 231.905 142.730 ;
        RECT 230.665 138.505 231.905 142.710 ;
      LAYER nwell ;
        RECT 232.855 139.655 244.625 144.010 ;
      LAYER pwell ;
        RECT 249.260 143.215 250.500 145.605 ;
        RECT 249.260 143.210 249.505 143.215 ;
        RECT 249.450 142.755 250.535 143.185 ;
      LAYER nwell ;
        RECT 235.315 139.650 244.625 139.655 ;
      LAYER pwell ;
        RECT 231.660 138.390 231.905 138.505 ;
        RECT 230.665 134.185 231.905 138.390 ;
        RECT 231.660 134.090 231.905 134.185 ;
        RECT 232.905 133.955 235.265 139.605 ;
      LAYER nwell ;
        RECT 235.315 133.905 237.775 139.650 ;
      LAYER pwell ;
        RECT 237.825 133.950 240.185 139.600 ;
      LAYER nwell ;
        RECT 240.235 133.900 244.625 139.650 ;
      LAYER pwell ;
        RECT 249.260 142.710 249.505 142.730 ;
        RECT 244.675 133.950 248.965 139.600 ;
        RECT 249.260 138.505 250.500 142.710 ;
        RECT 249.260 138.390 249.505 138.505 ;
        RECT 249.260 134.185 250.500 138.390 ;
        RECT 249.260 134.090 249.505 134.185 ;
      LAYER nwell ;
        RECT 250.920 133.900 254.260 150.600 ;
      LAYER pwell ;
        RECT 273.315 150.425 274.555 151.475 ;
      LAYER nwell ;
        RECT 274.975 150.600 276.835 152.040 ;
      LAYER pwell ;
        RECT 297.275 151.475 297.520 151.850 ;
        RECT 255.675 150.360 255.920 150.410 ;
        RECT 254.680 148.990 255.920 150.360 ;
        RECT 273.315 150.390 273.560 150.425 ;
        RECT 255.675 148.595 255.920 148.990 ;
        RECT 254.680 147.545 255.920 148.595 ;
        RECT 255.675 147.530 255.920 147.545 ;
        RECT 254.645 147.075 255.730 147.505 ;
        RECT 255.675 146.675 255.920 147.050 ;
        RECT 254.680 145.625 255.920 146.675 ;
        RECT 255.675 145.605 255.920 145.625 ;
        RECT 254.680 143.215 255.920 145.605 ;
        RECT 255.675 143.210 255.920 143.215 ;
      LAYER nwell ;
        RECT 256.910 144.015 259.370 149.765 ;
      LAYER pwell ;
        RECT 259.420 144.065 261.780 149.715 ;
      LAYER nwell ;
        RECT 261.830 144.015 264.290 149.760 ;
      LAYER pwell ;
        RECT 273.315 149.020 274.555 150.390 ;
        RECT 273.315 148.595 273.560 149.020 ;
        RECT 273.315 147.545 274.555 148.595 ;
        RECT 273.315 147.530 273.560 147.545 ;
        RECT 273.505 147.075 274.590 147.505 ;
      LAYER nwell ;
        RECT 256.910 144.010 264.290 144.015 ;
      LAYER pwell ;
        RECT 273.315 146.675 273.560 147.050 ;
        RECT 273.315 145.625 274.555 146.675 ;
        RECT 273.315 145.605 273.560 145.625 ;
        RECT 254.645 142.755 255.730 143.185 ;
        RECT 255.675 142.710 255.920 142.730 ;
        RECT 254.680 138.505 255.920 142.710 ;
      LAYER nwell ;
        RECT 256.910 139.655 268.680 144.010 ;
      LAYER pwell ;
        RECT 273.315 143.215 274.555 145.605 ;
        RECT 273.315 143.210 273.560 143.215 ;
        RECT 273.505 142.755 274.590 143.185 ;
      LAYER nwell ;
        RECT 259.370 139.650 268.680 139.655 ;
      LAYER pwell ;
        RECT 255.675 138.390 255.920 138.505 ;
        RECT 254.680 134.185 255.920 138.390 ;
        RECT 255.675 134.090 255.920 134.185 ;
        RECT 256.960 133.955 259.320 139.605 ;
      LAYER nwell ;
        RECT 259.370 133.905 261.830 139.650 ;
      LAYER pwell ;
        RECT 261.880 133.950 264.240 139.600 ;
      LAYER nwell ;
        RECT 264.290 133.900 268.680 139.650 ;
      LAYER pwell ;
        RECT 273.315 142.710 273.560 142.730 ;
        RECT 268.730 133.950 273.020 139.600 ;
        RECT 273.315 138.505 274.555 142.710 ;
        RECT 273.315 138.390 273.560 138.505 ;
        RECT 273.315 134.185 274.555 138.390 ;
        RECT 273.315 134.090 273.560 134.185 ;
      LAYER nwell ;
        RECT 274.975 133.900 278.315 150.600 ;
      LAYER pwell ;
        RECT 297.275 150.425 298.515 151.475 ;
      LAYER nwell ;
        RECT 298.935 150.600 300.795 152.040 ;
      LAYER pwell ;
        RECT 321.285 151.475 321.530 151.850 ;
        RECT 279.730 150.360 279.975 150.410 ;
        RECT 278.735 148.990 279.975 150.360 ;
        RECT 297.275 150.390 297.520 150.425 ;
        RECT 279.730 148.595 279.975 148.990 ;
        RECT 278.735 147.545 279.975 148.595 ;
        RECT 279.730 147.530 279.975 147.545 ;
        RECT 278.700 147.075 279.785 147.505 ;
        RECT 279.730 146.675 279.975 147.050 ;
        RECT 278.735 145.625 279.975 146.675 ;
        RECT 279.730 145.605 279.975 145.625 ;
        RECT 278.735 143.215 279.975 145.605 ;
        RECT 279.730 143.210 279.975 143.215 ;
      LAYER nwell ;
        RECT 280.870 144.015 283.330 149.765 ;
      LAYER pwell ;
        RECT 283.380 144.065 285.740 149.715 ;
      LAYER nwell ;
        RECT 285.790 144.015 288.250 149.760 ;
      LAYER pwell ;
        RECT 297.275 149.020 298.515 150.390 ;
        RECT 297.275 148.595 297.520 149.020 ;
        RECT 297.275 147.545 298.515 148.595 ;
        RECT 297.275 147.530 297.520 147.545 ;
        RECT 297.465 147.075 298.550 147.505 ;
      LAYER nwell ;
        RECT 280.870 144.010 288.250 144.015 ;
      LAYER pwell ;
        RECT 297.275 146.675 297.520 147.050 ;
        RECT 297.275 145.625 298.515 146.675 ;
        RECT 297.275 145.605 297.520 145.625 ;
        RECT 278.700 142.755 279.785 143.185 ;
        RECT 279.730 142.710 279.975 142.730 ;
        RECT 278.735 138.505 279.975 142.710 ;
      LAYER nwell ;
        RECT 280.870 139.655 292.640 144.010 ;
      LAYER pwell ;
        RECT 297.275 143.215 298.515 145.605 ;
        RECT 297.275 143.210 297.520 143.215 ;
        RECT 297.465 142.755 298.550 143.185 ;
      LAYER nwell ;
        RECT 283.330 139.650 292.640 139.655 ;
      LAYER pwell ;
        RECT 279.730 138.390 279.975 138.505 ;
        RECT 278.735 134.185 279.975 138.390 ;
        RECT 279.730 134.090 279.975 134.185 ;
        RECT 280.920 133.955 283.280 139.605 ;
      LAYER nwell ;
        RECT 283.330 133.905 285.790 139.650 ;
      LAYER pwell ;
        RECT 285.840 133.950 288.200 139.600 ;
      LAYER nwell ;
        RECT 288.250 133.900 292.640 139.650 ;
      LAYER pwell ;
        RECT 297.275 142.710 297.520 142.730 ;
        RECT 292.690 133.950 296.980 139.600 ;
        RECT 297.275 138.505 298.515 142.710 ;
        RECT 297.275 138.390 297.520 138.505 ;
        RECT 297.275 134.185 298.515 138.390 ;
        RECT 297.275 134.090 297.520 134.185 ;
      LAYER nwell ;
        RECT 298.935 133.900 302.275 150.600 ;
      LAYER pwell ;
        RECT 321.285 150.425 322.525 151.475 ;
      LAYER nwell ;
        RECT 322.945 150.600 324.805 152.040 ;
      LAYER pwell ;
        RECT 303.690 150.360 303.935 150.410 ;
        RECT 302.695 148.990 303.935 150.360 ;
        RECT 321.285 150.390 321.530 150.425 ;
        RECT 303.690 148.595 303.935 148.990 ;
        RECT 302.695 147.545 303.935 148.595 ;
        RECT 303.690 147.530 303.935 147.545 ;
        RECT 302.660 147.075 303.745 147.505 ;
        RECT 303.690 146.675 303.935 147.050 ;
        RECT 302.695 145.625 303.935 146.675 ;
        RECT 303.690 145.605 303.935 145.625 ;
        RECT 302.695 143.215 303.935 145.605 ;
        RECT 303.690 143.210 303.935 143.215 ;
      LAYER nwell ;
        RECT 304.880 144.015 307.340 149.765 ;
      LAYER pwell ;
        RECT 307.390 144.065 309.750 149.715 ;
      LAYER nwell ;
        RECT 309.800 144.015 312.260 149.760 ;
      LAYER pwell ;
        RECT 321.285 149.020 322.525 150.390 ;
        RECT 321.285 148.595 321.530 149.020 ;
        RECT 321.285 147.545 322.525 148.595 ;
        RECT 321.285 147.530 321.530 147.545 ;
        RECT 321.475 147.075 322.560 147.505 ;
      LAYER nwell ;
        RECT 304.880 144.010 312.260 144.015 ;
      LAYER pwell ;
        RECT 321.285 146.675 321.530 147.050 ;
        RECT 321.285 145.625 322.525 146.675 ;
        RECT 321.285 145.605 321.530 145.625 ;
        RECT 302.660 142.755 303.745 143.185 ;
        RECT 303.690 142.710 303.935 142.730 ;
        RECT 302.695 138.505 303.935 142.710 ;
      LAYER nwell ;
        RECT 304.880 139.655 316.650 144.010 ;
      LAYER pwell ;
        RECT 321.285 143.215 322.525 145.605 ;
        RECT 321.285 143.210 321.530 143.215 ;
        RECT 321.475 142.755 322.560 143.185 ;
      LAYER nwell ;
        RECT 307.340 139.650 316.650 139.655 ;
      LAYER pwell ;
        RECT 303.690 138.390 303.935 138.505 ;
        RECT 302.695 134.185 303.935 138.390 ;
        RECT 303.690 134.090 303.935 134.185 ;
        RECT 304.930 133.955 307.290 139.605 ;
      LAYER nwell ;
        RECT 307.340 133.905 309.800 139.650 ;
      LAYER pwell ;
        RECT 309.850 133.950 312.210 139.600 ;
      LAYER nwell ;
        RECT 312.260 133.900 316.650 139.650 ;
      LAYER pwell ;
        RECT 321.285 142.710 321.530 142.730 ;
        RECT 316.700 133.950 320.990 139.600 ;
        RECT 321.285 138.505 322.525 142.710 ;
        RECT 321.285 138.390 321.530 138.505 ;
        RECT 321.285 134.185 322.525 138.390 ;
        RECT 321.285 134.090 321.530 134.185 ;
      LAYER nwell ;
        RECT 322.945 133.900 326.285 150.600 ;
      LAYER pwell ;
        RECT 327.700 150.360 327.945 150.410 ;
        RECT 326.705 148.990 327.945 150.360 ;
        RECT 327.700 148.595 327.945 148.990 ;
        RECT 326.705 147.545 327.945 148.595 ;
        RECT 327.700 147.530 327.945 147.545 ;
        RECT 326.670 147.075 327.755 147.505 ;
        RECT 327.700 146.675 327.945 147.050 ;
        RECT 326.705 145.625 327.945 146.675 ;
        RECT 327.700 145.605 327.945 145.625 ;
        RECT 326.705 143.215 327.945 145.605 ;
        RECT 327.700 143.210 327.945 143.215 ;
        RECT 326.670 142.755 327.755 143.185 ;
        RECT 327.700 142.710 327.945 142.730 ;
        RECT 326.705 138.505 327.945 142.710 ;
        RECT 327.700 138.390 327.945 138.505 ;
        RECT 326.705 134.185 327.945 138.390 ;
        RECT 327.700 134.090 327.945 134.185 ;
      LAYER nwell ;
        RECT 16.760 131.950 21.770 131.960 ;
        RECT 42.680 131.950 47.690 131.960 ;
        RECT 58.150 131.950 63.160 131.960 ;
        RECT 16.760 131.855 17.840 131.950 ;
        RECT 42.680 131.855 43.760 131.950 ;
        RECT 62.080 131.855 63.160 131.950 ;
      LAYER pwell ;
        RECT 12.125 131.350 13.105 131.540 ;
        RECT 10.280 130.545 12.090 131.275 ;
        RECT 12.125 131.255 14.095 131.350 ;
        RECT 16.450 131.255 21.760 131.540 ;
        RECT 12.125 131.240 21.760 131.255 ;
        RECT 12.125 130.545 23.140 131.240 ;
        RECT 10.200 130.300 23.160 130.545 ;
        RECT 23.185 130.490 23.615 131.575 ;
        RECT 38.045 131.350 39.025 131.540 ;
        RECT 35.240 130.545 37.050 131.275 ;
        RECT 38.045 131.255 40.015 131.350 ;
        RECT 42.370 131.255 47.680 131.540 ;
        RECT 38.045 131.240 47.680 131.255 ;
        RECT 38.045 130.545 49.060 131.240 ;
        RECT 23.640 130.300 49.080 130.545 ;
        RECT 49.105 130.490 49.535 131.575 ;
        RECT 58.160 131.255 63.470 131.540 ;
        RECT 66.815 131.350 67.795 131.540 ;
        RECT 65.825 131.255 67.795 131.350 ;
        RECT 58.160 131.240 67.795 131.255 ;
        RECT 53.900 130.545 56.755 131.220 ;
        RECT 56.780 130.545 67.795 131.240 ;
        RECT 67.830 130.545 69.640 131.275 ;
        RECT 49.560 130.300 69.720 130.545 ;
        RECT 10.200 130.055 36.120 130.300 ;
        RECT 10.280 129.325 12.090 130.055 ;
        RECT 16.445 129.400 18.355 130.055 ;
        RECT 16.480 129.380 18.355 129.400 ;
        RECT 18.365 129.245 26.515 130.055 ;
        RECT 34.280 129.325 36.090 130.055 ;
        RECT 18.365 129.130 21.880 129.245 ;
        RECT 18.365 129.060 19.310 129.130 ;
        RECT 22.960 129.125 26.515 129.245 ;
        RECT 23.435 129.060 26.515 129.125 ;
        RECT 23.435 128.870 24.055 129.060 ;
        RECT 36.145 129.025 36.575 130.110 ;
        RECT 36.600 130.055 62.040 130.300 ;
        RECT 48.200 129.325 50.010 130.055 ;
        RECT 51.005 129.360 62.020 130.055 ;
        RECT 51.005 129.345 60.640 129.360 ;
        RECT 51.005 129.250 52.975 129.345 ;
        RECT 51.005 129.060 51.985 129.250 ;
        RECT 55.330 129.060 60.640 129.345 ;
        RECT 62.065 129.025 62.495 130.110 ;
        RECT 62.520 130.055 69.720 130.300 ;
        RECT 62.600 129.325 64.410 130.055 ;
        RECT 64.925 129.380 67.780 130.055 ;
        RECT 67.830 129.325 69.640 130.055 ;
      LAYER nwell ;
        RECT 55.640 128.650 56.720 128.745 ;
        RECT 55.640 128.640 60.650 128.650 ;
        RECT 10.010 125.300 69.910 128.640 ;
        RECT 31.750 125.290 36.760 125.300 ;
        RECT 50.950 125.290 55.960 125.300 ;
        RECT 35.680 125.195 36.760 125.290 ;
        RECT 54.880 125.195 55.960 125.290 ;
      LAYER pwell ;
        RECT 10.280 123.885 12.090 124.615 ;
        RECT 12.620 123.885 13.990 124.880 ;
        RECT 14.110 123.885 17.795 124.945 ;
        RECT 17.960 123.885 19.770 124.615 ;
        RECT 19.840 124.540 21.715 124.560 ;
        RECT 19.805 123.885 21.715 124.540 ;
        RECT 10.200 123.640 23.160 123.885 ;
        RECT 23.185 123.830 23.615 124.915 ;
        RECT 23.720 123.885 25.530 124.615 ;
        RECT 31.760 124.595 37.070 124.880 ;
        RECT 40.415 124.690 41.395 124.880 ;
        RECT 39.425 124.595 41.395 124.690 ;
        RECT 31.760 124.580 41.395 124.595 ;
        RECT 25.600 124.540 27.475 124.560 ;
        RECT 27.520 124.540 29.395 124.560 ;
        RECT 25.565 123.885 27.475 124.540 ;
        RECT 27.485 123.885 29.395 124.540 ;
        RECT 30.380 123.885 41.395 124.580 ;
        RECT 46.125 123.885 48.115 124.880 ;
        RECT 23.640 123.640 49.080 123.885 ;
        RECT 49.105 123.830 49.535 124.915 ;
        RECT 50.960 124.595 56.270 124.880 ;
        RECT 59.615 124.690 60.595 124.880 ;
        RECT 58.625 124.595 60.595 124.690 ;
        RECT 50.960 124.580 60.595 124.595 ;
        RECT 49.580 123.885 60.595 124.580 ;
        RECT 62.045 123.885 64.900 124.560 ;
        RECT 64.925 123.885 67.780 124.560 ;
        RECT 67.830 123.885 69.640 124.615 ;
        RECT 49.560 123.640 69.720 123.885 ;
        RECT 10.200 123.395 36.120 123.640 ;
        RECT 10.280 122.665 12.090 123.395 ;
        RECT 12.200 122.665 14.010 123.395 ;
        RECT 14.045 122.585 22.195 123.395 ;
        RECT 14.045 122.465 17.600 122.585 ;
        RECT 18.680 122.470 22.195 122.585 ;
        RECT 14.045 122.400 17.125 122.465 ;
        RECT 21.250 122.400 22.195 122.470 ;
        RECT 16.505 122.210 17.125 122.400 ;
        RECT 22.240 122.270 24.835 123.395 ;
        RECT 25.085 122.700 36.100 123.395 ;
        RECT 25.085 122.685 34.720 122.700 ;
        RECT 25.085 122.590 27.055 122.685 ;
        RECT 25.085 122.400 26.065 122.590 ;
        RECT 29.410 122.400 34.720 122.685 ;
        RECT 36.145 122.365 36.575 123.450 ;
        RECT 36.600 123.395 62.040 123.640 ;
        RECT 36.605 122.400 38.595 123.395 ;
        RECT 44.285 122.740 46.195 123.395 ;
        RECT 44.320 122.720 46.195 122.740 ;
        RECT 46.220 122.700 57.235 123.395 ;
        RECT 47.600 122.685 57.235 122.700 ;
        RECT 47.600 122.400 52.910 122.685 ;
        RECT 55.265 122.590 57.235 122.685 ;
        RECT 56.255 122.400 57.235 122.590 ;
        RECT 62.065 122.365 62.495 123.450 ;
        RECT 62.520 123.395 69.720 123.640 ;
        RECT 62.600 122.665 64.410 123.395 ;
        RECT 64.925 122.720 67.780 123.395 ;
        RECT 67.830 122.665 69.640 123.395 ;
        RECT 22.240 122.190 23.745 122.270 ;
      LAYER nwell ;
        RECT 29.720 121.990 30.800 122.085 ;
        RECT 51.520 121.990 52.600 122.085 ;
        RECT 29.720 121.980 34.730 121.990 ;
        RECT 47.590 121.980 52.600 121.990 ;
        RECT 10.010 118.640 69.910 121.980 ;
        RECT 31.640 118.630 36.650 118.640 ;
        RECT 39.430 118.630 44.440 118.640 ;
        RECT 58.150 118.630 63.160 118.640 ;
        RECT 31.640 118.535 32.720 118.630 ;
        RECT 43.360 118.535 44.440 118.630 ;
        RECT 62.080 118.535 63.160 118.630 ;
      LAYER pwell ;
        RECT 10.280 117.225 12.090 117.955 ;
        RECT 12.125 117.225 21.715 117.900 ;
        RECT 10.200 116.980 23.160 117.225 ;
        RECT 23.185 117.170 23.615 118.255 ;
        RECT 23.645 117.225 26.035 118.220 ;
        RECT 27.005 118.030 27.985 118.220 ;
        RECT 27.005 117.935 28.975 118.030 ;
        RECT 31.330 117.935 36.640 118.220 ;
        RECT 27.005 117.920 36.640 117.935 ;
        RECT 39.440 117.935 44.750 118.220 ;
        RECT 48.095 118.030 49.075 118.220 ;
        RECT 47.105 117.935 49.075 118.030 ;
        RECT 39.440 117.920 49.075 117.935 ;
        RECT 27.005 117.225 38.020 117.920 ;
        RECT 38.060 117.225 49.075 117.920 ;
        RECT 23.640 116.980 49.080 117.225 ;
        RECT 49.105 117.170 49.535 118.255 ;
        RECT 51.005 117.225 52.995 118.220 ;
        RECT 58.160 117.935 63.470 118.220 ;
        RECT 66.815 118.030 67.795 118.220 ;
        RECT 65.825 117.935 67.795 118.030 ;
        RECT 58.160 117.920 67.795 117.935 ;
        RECT 53.405 117.880 55.280 117.900 ;
        RECT 53.405 117.225 55.315 117.880 ;
        RECT 56.780 117.225 67.795 117.920 ;
        RECT 67.830 117.225 69.640 117.955 ;
        RECT 49.560 116.980 69.720 117.225 ;
        RECT 10.200 116.735 36.120 116.980 ;
        RECT 10.280 116.005 12.090 116.735 ;
        RECT 12.200 116.005 14.010 116.735 ;
        RECT 14.045 116.080 15.955 116.735 ;
        RECT 14.080 116.060 15.955 116.080 ;
        RECT 15.965 115.930 20.755 116.735 ;
        RECT 21.245 116.060 30.835 116.735 ;
        RECT 16.475 115.840 20.755 115.930 ;
        RECT 16.475 115.740 17.420 115.840 ;
        RECT 30.845 115.740 32.255 116.735 ;
        RECT 32.290 116.060 35.955 116.735 ;
        RECT 34.175 115.740 35.955 116.060 ;
        RECT 36.145 115.705 36.575 116.790 ;
        RECT 36.600 116.735 62.040 116.980 ;
        RECT 36.850 115.740 38.790 116.735 ;
        RECT 39.500 116.040 50.515 116.735 ;
        RECT 51.020 116.040 62.035 116.735 ;
        RECT 40.880 116.025 50.515 116.040 ;
        RECT 40.880 115.740 46.190 116.025 ;
        RECT 48.545 115.930 50.515 116.025 ;
        RECT 49.535 115.740 50.515 115.930 ;
        RECT 52.400 116.025 62.035 116.040 ;
        RECT 52.400 115.740 57.710 116.025 ;
        RECT 60.065 115.930 62.035 116.025 ;
        RECT 61.055 115.740 62.035 115.930 ;
        RECT 62.065 115.705 62.495 116.790 ;
        RECT 62.520 116.735 69.720 116.980 ;
        RECT 62.600 116.005 64.410 116.735 ;
        RECT 64.925 116.060 67.780 116.735 ;
        RECT 67.830 116.005 69.640 116.735 ;
      LAYER nwell ;
        RECT 44.800 115.330 45.880 115.425 ;
        RECT 56.320 115.330 57.400 115.425 ;
        RECT 40.870 115.320 45.880 115.330 ;
        RECT 52.390 115.320 57.400 115.330 ;
        RECT 10.010 111.980 69.910 115.320 ;
        RECT 36.920 111.970 41.930 111.980 ;
        RECT 58.150 111.970 63.160 111.980 ;
        RECT 36.920 111.875 38.000 111.970 ;
        RECT 62.080 111.875 63.160 111.970 ;
      LAYER pwell ;
        RECT 17.465 111.560 18.085 111.750 ;
        RECT 10.280 110.565 12.090 111.295 ;
        RECT 12.145 110.565 13.555 111.560 ;
        RECT 13.585 110.565 14.995 111.560 ;
        RECT 15.005 111.495 18.085 111.560 ;
        RECT 15.005 111.375 18.560 111.495 ;
        RECT 22.210 111.490 23.155 111.560 ;
        RECT 19.640 111.375 23.155 111.490 ;
        RECT 15.005 110.565 23.155 111.375 ;
        RECT 10.200 110.320 23.160 110.565 ;
        RECT 23.185 110.510 23.615 111.595 ;
        RECT 26.105 111.560 26.725 111.750 ;
        RECT 23.645 111.495 26.725 111.560 ;
        RECT 23.645 111.375 27.200 111.495 ;
        RECT 30.850 111.490 31.795 111.560 ;
        RECT 28.280 111.375 31.795 111.490 ;
        RECT 23.645 110.565 31.795 111.375 ;
        RECT 32.285 111.370 33.265 111.560 ;
        RECT 32.285 111.275 34.255 111.370 ;
        RECT 36.610 111.275 41.920 111.560 ;
        RECT 32.285 111.260 41.920 111.275 ;
        RECT 32.285 110.565 43.300 111.260 ;
        RECT 47.240 110.565 49.050 111.295 ;
        RECT 23.640 110.320 49.080 110.565 ;
        RECT 49.105 110.510 49.535 111.595 ;
        RECT 53.480 110.565 55.290 111.295 ;
        RECT 58.160 111.275 63.470 111.560 ;
        RECT 66.815 111.370 67.795 111.560 ;
        RECT 65.825 111.275 67.795 111.370 ;
        RECT 58.160 111.260 67.795 111.275 ;
        RECT 56.780 110.565 67.795 111.260 ;
        RECT 67.830 110.565 69.640 111.295 ;
        RECT 49.560 110.320 69.720 110.565 ;
        RECT 10.200 110.075 36.120 110.320 ;
        RECT 10.280 109.345 12.090 110.075 ;
        RECT 12.200 109.345 14.010 110.075 ;
        RECT 15.005 109.420 16.915 110.075 ;
        RECT 20.765 109.420 22.675 110.075 ;
        RECT 23.645 109.420 25.555 110.075 ;
        RECT 15.005 109.400 16.880 109.420 ;
        RECT 20.800 109.400 22.675 109.420 ;
        RECT 23.680 109.400 25.555 109.420 ;
        RECT 25.640 109.345 27.450 110.075 ;
        RECT 27.485 109.080 29.775 110.075 ;
        RECT 29.960 109.345 31.770 110.075 ;
        RECT 31.805 109.420 33.715 110.075 ;
        RECT 31.840 109.400 33.715 109.420 ;
        RECT 33.800 109.345 35.610 110.075 ;
        RECT 36.145 109.045 36.575 110.130 ;
        RECT 36.600 110.075 62.040 110.320 ;
        RECT 37.085 109.080 39.075 110.075 ;
        RECT 44.780 109.380 55.795 110.075 ;
        RECT 46.160 109.365 55.795 109.380 ;
        RECT 46.160 109.080 51.470 109.365 ;
        RECT 53.825 109.270 55.795 109.365 ;
        RECT 55.880 109.345 57.690 110.075 ;
        RECT 59.165 109.400 62.020 110.075 ;
        RECT 54.815 109.080 55.795 109.270 ;
        RECT 62.065 109.045 62.495 110.130 ;
        RECT 62.520 110.075 69.720 110.320 ;
        RECT 62.600 109.345 64.410 110.075 ;
        RECT 64.925 109.400 67.780 110.075 ;
        RECT 67.830 109.345 69.640 110.075 ;
      LAYER nwell ;
        RECT 50.080 108.670 51.160 108.765 ;
        RECT 46.150 108.660 51.160 108.670 ;
        RECT 10.010 105.320 69.910 108.660 ;
        RECT 37.400 105.310 42.410 105.320 ;
        RECT 50.950 105.310 55.960 105.320 ;
        RECT 37.400 105.215 38.480 105.310 ;
        RECT 54.880 105.215 55.960 105.310 ;
      LAYER pwell ;
        RECT 10.280 103.905 12.090 104.635 ;
        RECT 12.125 103.905 21.715 104.580 ;
        RECT 10.200 103.660 23.160 103.905 ;
        RECT 23.185 103.850 23.615 104.935 ;
        RECT 23.725 103.905 27.410 104.965 ;
        RECT 27.525 103.905 30.835 104.900 ;
        RECT 32.765 104.710 33.745 104.900 ;
        RECT 32.765 104.615 34.735 104.710 ;
        RECT 37.090 104.615 42.400 104.900 ;
        RECT 32.765 104.600 42.400 104.615 ;
        RECT 30.880 104.560 32.755 104.580 ;
        RECT 30.845 103.905 32.755 104.560 ;
        RECT 32.765 103.905 43.780 104.600 ;
        RECT 43.880 103.905 45.690 104.635 ;
        RECT 46.685 103.905 48.675 104.900 ;
        RECT 23.640 103.660 49.080 103.905 ;
        RECT 49.105 103.850 49.535 104.935 ;
        RECT 50.960 104.615 56.270 104.900 ;
        RECT 59.615 104.710 60.595 104.900 ;
        RECT 58.625 104.615 60.595 104.710 ;
        RECT 50.960 104.600 60.595 104.615 ;
        RECT 49.580 103.905 60.595 104.600 ;
        RECT 62.045 103.905 64.900 104.580 ;
        RECT 64.925 103.905 67.780 104.580 ;
        RECT 67.830 103.905 69.640 104.635 ;
        RECT 49.560 103.660 69.720 103.905 ;
        RECT 10.200 103.415 36.120 103.660 ;
        RECT 10.280 102.685 12.090 103.415 ;
        RECT 13.565 102.605 21.715 103.415 ;
        RECT 13.565 102.485 17.120 102.605 ;
        RECT 18.200 102.490 21.715 102.605 ;
        RECT 13.565 102.420 16.645 102.485 ;
        RECT 20.770 102.420 21.715 102.490 ;
        RECT 16.025 102.230 16.645 102.420 ;
        RECT 22.350 102.290 24.480 103.415 ;
        RECT 24.605 102.605 32.755 103.415 ;
        RECT 32.840 102.685 34.650 103.415 ;
        RECT 24.605 102.485 28.160 102.605 ;
        RECT 29.240 102.490 32.755 102.605 ;
        RECT 24.605 102.420 27.685 102.485 ;
        RECT 31.810 102.420 32.755 102.490 ;
        RECT 22.350 102.210 23.295 102.290 ;
        RECT 27.065 102.230 27.685 102.420 ;
        RECT 36.145 102.385 36.575 103.470 ;
        RECT 36.600 103.415 62.040 103.660 ;
        RECT 40.520 102.685 42.330 103.415 ;
        RECT 43.340 102.720 54.355 103.415 ;
        RECT 59.165 102.740 62.020 103.415 ;
        RECT 44.720 102.705 54.355 102.720 ;
        RECT 44.720 102.420 50.030 102.705 ;
        RECT 52.385 102.610 54.355 102.705 ;
        RECT 53.375 102.420 54.355 102.610 ;
        RECT 62.065 102.385 62.495 103.470 ;
        RECT 62.520 103.415 69.720 103.660 ;
        RECT 63.005 102.420 64.915 103.415 ;
        RECT 64.925 102.740 67.780 103.415 ;
        RECT 67.830 102.685 69.640 103.415 ;
      LAYER nwell ;
        RECT 48.640 102.010 49.720 102.105 ;
        RECT 44.710 102.000 49.720 102.010 ;
        RECT 10.010 98.660 69.910 102.000 ;
        RECT 36.440 98.650 41.450 98.660 ;
        RECT 58.150 98.650 63.160 98.660 ;
        RECT 36.440 98.555 37.520 98.650 ;
        RECT 62.080 98.555 63.160 98.650 ;
      LAYER pwell ;
        RECT 10.280 97.245 12.090 97.975 ;
        RECT 12.200 97.245 14.010 97.975 ;
        RECT 15.520 97.900 17.395 97.920 ;
        RECT 15.485 97.245 17.395 97.900 ;
        RECT 18.845 97.245 23.145 98.240 ;
        RECT 10.200 97.000 23.160 97.245 ;
        RECT 23.185 97.190 23.615 98.275 ;
        RECT 23.720 97.245 25.530 97.975 ;
        RECT 25.600 97.900 27.475 97.920 ;
        RECT 25.565 97.245 27.475 97.900 ;
        RECT 27.550 97.245 31.235 98.305 ;
        RECT 31.805 98.050 32.785 98.240 ;
        RECT 31.805 97.955 33.775 98.050 ;
        RECT 36.130 97.955 41.440 98.240 ;
        RECT 31.805 97.940 41.440 97.955 ;
        RECT 31.805 97.245 42.820 97.940 ;
        RECT 46.760 97.245 48.570 97.975 ;
        RECT 23.640 97.000 49.080 97.245 ;
        RECT 49.105 97.190 49.535 98.275 ;
        RECT 58.160 97.955 63.470 98.240 ;
        RECT 66.815 98.050 67.795 98.240 ;
        RECT 65.825 97.955 67.795 98.050 ;
        RECT 58.160 97.940 67.795 97.955 ;
        RECT 50.045 97.245 52.900 97.920 ;
        RECT 53.885 97.245 56.740 97.920 ;
        RECT 56.780 97.245 67.795 97.940 ;
        RECT 67.830 97.245 69.640 97.975 ;
        RECT 49.560 97.000 69.720 97.245 ;
        RECT 10.200 96.755 36.120 97.000 ;
        RECT 10.280 96.025 12.090 96.755 ;
        RECT 23.720 96.025 25.530 96.755 ;
        RECT 27.005 96.080 28.915 96.755 ;
        RECT 28.925 95.760 30.835 96.755 ;
        RECT 30.845 96.100 32.755 96.755 ;
        RECT 30.880 96.080 32.755 96.100 ;
        RECT 32.765 95.760 34.755 96.755 ;
        RECT 36.145 95.725 36.575 96.810 ;
        RECT 36.600 96.755 62.040 97.000 ;
        RECT 38.060 96.060 49.075 96.755 ;
        RECT 39.440 96.045 49.075 96.060 ;
        RECT 39.440 95.760 44.750 96.045 ;
        RECT 47.105 95.950 49.075 96.045 ;
        RECT 48.095 95.760 49.075 95.950 ;
        RECT 49.085 96.060 60.100 96.755 ;
        RECT 49.085 96.045 58.720 96.060 ;
        RECT 49.085 95.950 51.055 96.045 ;
        RECT 49.085 95.760 50.065 95.950 ;
        RECT 53.410 95.760 58.720 96.045 ;
        RECT 60.200 96.025 62.010 96.755 ;
        RECT 62.065 95.725 62.495 96.810 ;
        RECT 62.520 96.755 69.720 97.000 ;
        RECT 62.600 96.025 64.410 96.755 ;
        RECT 64.925 96.080 67.780 96.755 ;
        RECT 67.830 96.025 69.640 96.755 ;
      LAYER nwell ;
        RECT 43.360 95.350 44.440 95.445 ;
        RECT 39.430 95.340 44.440 95.350 ;
        RECT 53.720 95.350 54.800 95.445 ;
        RECT 53.720 95.340 58.730 95.350 ;
        RECT 10.010 92.000 69.910 95.340 ;
        RECT 30.200 91.990 35.210 92.000 ;
        RECT 41.240 91.990 46.250 92.000 ;
        RECT 58.150 91.990 63.160 92.000 ;
        RECT 30.200 91.895 31.280 91.990 ;
        RECT 41.240 91.895 42.320 91.990 ;
        RECT 62.080 91.895 63.160 91.990 ;
      LAYER pwell ;
        RECT 10.280 90.585 12.090 91.315 ;
        RECT 19.880 90.585 21.690 91.315 ;
        RECT 10.200 90.340 23.160 90.585 ;
        RECT 23.185 90.530 23.615 91.615 ;
        RECT 25.565 91.390 26.545 91.580 ;
        RECT 25.565 91.295 27.535 91.390 ;
        RECT 29.890 91.295 35.200 91.580 ;
        RECT 25.565 91.280 35.200 91.295 ;
        RECT 36.605 91.390 37.585 91.580 ;
        RECT 36.605 91.295 38.575 91.390 ;
        RECT 40.930 91.295 46.240 91.580 ;
        RECT 36.605 91.280 46.240 91.295 ;
        RECT 23.645 90.585 25.555 91.260 ;
        RECT 25.565 90.585 36.580 91.280 ;
        RECT 36.605 90.585 47.620 91.280 ;
        RECT 23.640 90.340 49.080 90.585 ;
        RECT 49.105 90.530 49.535 91.615 ;
        RECT 58.160 91.295 63.470 91.580 ;
        RECT 66.815 91.390 67.795 91.580 ;
        RECT 65.825 91.295 67.795 91.390 ;
        RECT 58.160 91.280 67.795 91.295 ;
        RECT 51.005 90.585 53.860 91.260 ;
        RECT 53.885 90.585 56.740 91.260 ;
        RECT 56.780 90.585 67.795 91.280 ;
        RECT 67.830 90.585 69.640 91.315 ;
        RECT 49.560 90.340 69.720 90.585 ;
        RECT 10.200 90.095 36.120 90.340 ;
        RECT 10.280 89.365 12.090 90.095 ;
        RECT 25.100 89.400 36.115 90.095 ;
        RECT 26.480 89.385 36.115 89.400 ;
        RECT 26.480 89.100 31.790 89.385 ;
        RECT 34.145 89.290 36.115 89.385 ;
        RECT 35.135 89.100 36.115 89.290 ;
        RECT 36.145 89.065 36.575 90.150 ;
        RECT 36.600 90.095 62.040 90.340 ;
        RECT 36.605 89.100 38.515 90.095 ;
        RECT 39.965 89.420 42.820 90.095 ;
        RECT 42.845 89.420 45.700 90.095 ;
        RECT 45.740 89.400 56.755 90.095 ;
        RECT 56.765 89.440 58.675 90.095 ;
        RECT 56.800 89.420 58.675 89.440 ;
        RECT 59.165 89.420 62.020 90.095 ;
        RECT 47.120 89.385 56.755 89.400 ;
        RECT 47.120 89.100 52.430 89.385 ;
        RECT 54.785 89.290 56.755 89.385 ;
        RECT 55.775 89.100 56.755 89.290 ;
        RECT 62.065 89.065 62.495 90.150 ;
        RECT 62.520 90.095 69.720 90.340 ;
        RECT 62.600 89.365 64.410 90.095 ;
        RECT 64.925 89.420 67.780 90.095 ;
        RECT 67.830 89.365 69.640 90.095 ;
      LAYER nwell ;
        RECT 30.400 88.690 31.480 88.785 ;
        RECT 51.040 88.690 52.120 88.785 ;
        RECT 26.470 88.680 31.480 88.690 ;
        RECT 47.110 88.680 52.120 88.690 ;
        RECT 10.010 85.340 69.910 88.680 ;
      LAYER pwell ;
        RECT 112.850 87.695 115.210 93.345 ;
      LAYER nwell ;
        RECT 115.260 87.650 117.720 93.395 ;
      LAYER pwell ;
        RECT 117.770 87.700 120.130 93.350 ;
      LAYER nwell ;
        RECT 120.180 87.650 124.570 93.400 ;
      LAYER pwell ;
        RECT 124.620 87.700 128.910 93.350 ;
        RECT 129.205 93.115 129.450 93.210 ;
        RECT 129.205 88.910 130.445 93.115 ;
        RECT 129.205 88.795 129.450 88.910 ;
      LAYER nwell ;
        RECT 115.260 87.645 124.570 87.650 ;
        RECT 41.240 85.330 46.250 85.340 ;
        RECT 54.200 85.330 59.210 85.340 ;
        RECT 41.240 85.235 42.320 85.330 ;
        RECT 54.200 85.235 55.280 85.330 ;
      LAYER pwell ;
        RECT 10.280 83.925 12.090 84.655 ;
        RECT 12.620 83.925 15.475 84.600 ;
        RECT 10.200 83.680 23.160 83.925 ;
        RECT 23.185 83.870 23.615 84.955 ;
        RECT 23.720 83.925 25.530 84.655 ;
        RECT 26.525 84.580 28.400 84.600 ;
        RECT 26.525 83.925 28.435 84.580 ;
        RECT 32.360 83.925 34.170 84.655 ;
        RECT 34.205 84.580 36.080 84.600 ;
        RECT 34.205 83.925 36.115 84.580 ;
        RECT 23.640 83.680 36.120 83.925 ;
        RECT 36.145 83.870 36.575 84.955 ;
        RECT 36.605 84.730 37.585 84.920 ;
        RECT 36.605 84.635 38.575 84.730 ;
        RECT 40.930 84.635 46.240 84.920 ;
        RECT 36.605 84.620 46.240 84.635 ;
        RECT 36.605 83.925 47.620 84.620 ;
        RECT 36.600 83.680 49.080 83.925 ;
        RECT 49.105 83.870 49.535 84.955 ;
        RECT 49.565 84.730 50.545 84.920 ;
        RECT 49.565 84.635 51.535 84.730 ;
        RECT 53.890 84.635 59.200 84.920 ;
        RECT 49.565 84.620 59.200 84.635 ;
        RECT 49.565 83.925 60.580 84.620 ;
        RECT 49.560 83.680 62.040 83.925 ;
        RECT 62.065 83.870 62.495 84.955 ;
        RECT 62.560 84.580 64.435 84.600 ;
        RECT 62.525 83.925 64.435 84.580 ;
        RECT 64.925 83.925 67.780 84.600 ;
        RECT 67.830 83.925 69.640 84.655 ;
        RECT 62.520 83.680 69.720 83.925 ;
      LAYER nwell ;
        RECT 112.800 83.290 124.570 87.645 ;
      LAYER pwell ;
        RECT 129.205 84.590 130.445 88.795 ;
        RECT 129.205 84.570 129.450 84.590 ;
        RECT 129.395 84.115 130.480 84.545 ;
        RECT 129.205 84.085 129.450 84.090 ;
      LAYER nwell ;
        RECT 112.800 83.285 120.180 83.290 ;
        RECT 112.800 77.535 115.260 83.285 ;
      LAYER pwell ;
        RECT 115.310 77.585 117.670 83.235 ;
      LAYER nwell ;
        RECT 117.720 77.540 120.180 83.285 ;
      LAYER pwell ;
        RECT 129.205 81.695 130.445 84.085 ;
        RECT 129.205 81.675 129.450 81.695 ;
        RECT 129.205 80.625 130.445 81.675 ;
        RECT 129.205 80.250 129.450 80.625 ;
        RECT 129.395 79.795 130.480 80.225 ;
        RECT 129.205 79.755 129.450 79.770 ;
        RECT 129.205 78.705 130.445 79.755 ;
        RECT 129.205 78.280 129.450 78.705 ;
        RECT 129.205 76.910 130.445 78.280 ;
        RECT 129.205 76.875 129.450 76.910 ;
        RECT 129.205 75.825 130.445 76.875 ;
      LAYER nwell ;
        RECT 130.865 76.700 134.205 93.400 ;
      LAYER pwell ;
        RECT 135.620 93.115 135.865 93.210 ;
        RECT 134.625 88.910 135.865 93.115 ;
        RECT 135.620 88.795 135.865 88.910 ;
        RECT 134.625 84.590 135.865 88.795 ;
        RECT 136.860 87.695 139.220 93.345 ;
      LAYER nwell ;
        RECT 139.270 87.650 141.730 93.395 ;
      LAYER pwell ;
        RECT 141.780 87.700 144.140 93.350 ;
      LAYER nwell ;
        RECT 144.190 87.650 148.580 93.400 ;
      LAYER pwell ;
        RECT 148.630 87.700 152.920 93.350 ;
        RECT 153.215 93.115 153.460 93.210 ;
        RECT 153.215 88.910 154.455 93.115 ;
        RECT 153.215 88.795 153.460 88.910 ;
      LAYER nwell ;
        RECT 139.270 87.645 148.580 87.650 ;
      LAYER pwell ;
        RECT 135.620 84.570 135.865 84.590 ;
        RECT 134.590 84.115 135.675 84.545 ;
        RECT 135.620 84.085 135.865 84.090 ;
        RECT 134.625 81.695 135.865 84.085 ;
        RECT 135.620 81.675 135.865 81.695 ;
        RECT 134.625 80.625 135.865 81.675 ;
        RECT 135.620 80.250 135.865 80.625 ;
      LAYER nwell ;
        RECT 136.810 83.290 148.580 87.645 ;
      LAYER pwell ;
        RECT 153.215 84.590 154.455 88.795 ;
        RECT 153.215 84.570 153.460 84.590 ;
        RECT 153.405 84.115 154.490 84.545 ;
        RECT 153.215 84.085 153.460 84.090 ;
      LAYER nwell ;
        RECT 136.810 83.285 144.190 83.290 ;
      LAYER pwell ;
        RECT 134.590 79.795 135.675 80.225 ;
        RECT 135.620 79.755 135.865 79.770 ;
        RECT 134.625 78.705 135.865 79.755 ;
        RECT 135.620 78.310 135.865 78.705 ;
        RECT 134.625 76.940 135.865 78.310 ;
      LAYER nwell ;
        RECT 136.810 77.535 139.270 83.285 ;
      LAYER pwell ;
        RECT 139.320 77.585 141.680 83.235 ;
      LAYER nwell ;
        RECT 141.730 77.540 144.190 83.285 ;
      LAYER pwell ;
        RECT 153.215 81.695 154.455 84.085 ;
        RECT 153.215 81.675 153.460 81.695 ;
        RECT 153.215 80.625 154.455 81.675 ;
        RECT 153.215 80.250 153.460 80.625 ;
        RECT 153.405 79.795 154.490 80.225 ;
        RECT 153.215 79.755 153.460 79.770 ;
        RECT 153.215 78.705 154.455 79.755 ;
        RECT 153.215 78.280 153.460 78.705 ;
        RECT 135.620 76.890 135.865 76.940 ;
        RECT 153.215 76.910 154.455 78.280 ;
        RECT 153.215 76.875 153.460 76.910 ;
        RECT 129.205 75.450 129.450 75.825 ;
      LAYER nwell ;
        RECT 130.865 75.260 132.725 76.700 ;
      LAYER pwell ;
        RECT 153.215 75.825 154.455 76.875 ;
      LAYER nwell ;
        RECT 154.875 76.700 158.215 93.400 ;
      LAYER pwell ;
        RECT 159.630 93.115 159.875 93.210 ;
        RECT 158.635 88.910 159.875 93.115 ;
        RECT 159.630 88.795 159.875 88.910 ;
        RECT 158.635 84.590 159.875 88.795 ;
        RECT 160.870 87.695 163.230 93.345 ;
      LAYER nwell ;
        RECT 163.280 87.650 165.740 93.395 ;
      LAYER pwell ;
        RECT 165.790 87.700 168.150 93.350 ;
      LAYER nwell ;
        RECT 168.200 87.650 172.590 93.400 ;
      LAYER pwell ;
        RECT 172.640 87.700 176.930 93.350 ;
        RECT 177.225 93.115 177.470 93.210 ;
        RECT 177.225 88.910 178.465 93.115 ;
        RECT 177.225 88.795 177.470 88.910 ;
      LAYER nwell ;
        RECT 163.280 87.645 172.590 87.650 ;
      LAYER pwell ;
        RECT 159.630 84.570 159.875 84.590 ;
        RECT 158.600 84.115 159.685 84.545 ;
        RECT 159.630 84.085 159.875 84.090 ;
        RECT 158.635 81.695 159.875 84.085 ;
        RECT 159.630 81.675 159.875 81.695 ;
        RECT 158.635 80.625 159.875 81.675 ;
        RECT 159.630 80.250 159.875 80.625 ;
      LAYER nwell ;
        RECT 160.820 83.290 172.590 87.645 ;
      LAYER pwell ;
        RECT 177.225 84.590 178.465 88.795 ;
        RECT 177.225 84.570 177.470 84.590 ;
        RECT 177.415 84.115 178.500 84.545 ;
        RECT 177.225 84.085 177.470 84.090 ;
      LAYER nwell ;
        RECT 160.820 83.285 168.200 83.290 ;
      LAYER pwell ;
        RECT 158.600 79.795 159.685 80.225 ;
        RECT 159.630 79.755 159.875 79.770 ;
        RECT 158.635 78.705 159.875 79.755 ;
        RECT 159.630 78.310 159.875 78.705 ;
        RECT 158.635 76.940 159.875 78.310 ;
      LAYER nwell ;
        RECT 160.820 77.535 163.280 83.285 ;
      LAYER pwell ;
        RECT 163.330 77.585 165.690 83.235 ;
      LAYER nwell ;
        RECT 165.740 77.540 168.200 83.285 ;
      LAYER pwell ;
        RECT 177.225 81.695 178.465 84.085 ;
        RECT 177.225 81.675 177.470 81.695 ;
        RECT 177.225 80.625 178.465 81.675 ;
        RECT 177.225 80.250 177.470 80.625 ;
        RECT 177.415 79.795 178.500 80.225 ;
        RECT 177.225 79.755 177.470 79.770 ;
        RECT 177.225 78.705 178.465 79.755 ;
        RECT 177.225 78.280 177.470 78.705 ;
        RECT 159.630 76.890 159.875 76.940 ;
        RECT 177.225 76.910 178.465 78.280 ;
        RECT 177.225 76.875 177.470 76.910 ;
        RECT 153.215 75.450 153.460 75.825 ;
      LAYER nwell ;
        RECT 154.875 75.260 156.735 76.700 ;
      LAYER pwell ;
        RECT 177.225 75.825 178.465 76.875 ;
      LAYER nwell ;
        RECT 178.885 76.700 182.225 93.400 ;
      LAYER pwell ;
        RECT 183.640 93.115 183.885 93.210 ;
        RECT 182.645 88.910 183.885 93.115 ;
        RECT 183.640 88.795 183.885 88.910 ;
        RECT 182.645 84.590 183.885 88.795 ;
        RECT 184.880 87.695 187.240 93.345 ;
      LAYER nwell ;
        RECT 187.290 87.650 189.750 93.395 ;
      LAYER pwell ;
        RECT 189.800 87.700 192.160 93.350 ;
      LAYER nwell ;
        RECT 192.210 87.650 196.600 93.400 ;
      LAYER pwell ;
        RECT 196.650 87.700 200.940 93.350 ;
        RECT 201.235 93.115 201.480 93.210 ;
        RECT 201.235 88.910 202.475 93.115 ;
        RECT 201.235 88.795 201.480 88.910 ;
      LAYER nwell ;
        RECT 187.290 87.645 196.600 87.650 ;
      LAYER pwell ;
        RECT 183.640 84.570 183.885 84.590 ;
        RECT 182.610 84.115 183.695 84.545 ;
        RECT 183.640 84.085 183.885 84.090 ;
        RECT 182.645 81.695 183.885 84.085 ;
        RECT 183.640 81.675 183.885 81.695 ;
        RECT 182.645 80.625 183.885 81.675 ;
        RECT 183.640 80.250 183.885 80.625 ;
      LAYER nwell ;
        RECT 184.830 83.290 196.600 87.645 ;
      LAYER pwell ;
        RECT 201.235 84.590 202.475 88.795 ;
        RECT 201.235 84.570 201.480 84.590 ;
        RECT 201.425 84.115 202.510 84.545 ;
        RECT 201.235 84.085 201.480 84.090 ;
      LAYER nwell ;
        RECT 184.830 83.285 192.210 83.290 ;
      LAYER pwell ;
        RECT 182.610 79.795 183.695 80.225 ;
        RECT 183.640 79.755 183.885 79.770 ;
        RECT 182.645 78.705 183.885 79.755 ;
        RECT 183.640 78.310 183.885 78.705 ;
        RECT 182.645 76.940 183.885 78.310 ;
      LAYER nwell ;
        RECT 184.830 77.535 187.290 83.285 ;
      LAYER pwell ;
        RECT 187.340 77.585 189.700 83.235 ;
      LAYER nwell ;
        RECT 189.750 77.540 192.210 83.285 ;
      LAYER pwell ;
        RECT 201.235 81.695 202.475 84.085 ;
        RECT 201.235 81.675 201.480 81.695 ;
        RECT 201.235 80.625 202.475 81.675 ;
        RECT 201.235 80.250 201.480 80.625 ;
        RECT 201.425 79.795 202.510 80.225 ;
        RECT 201.235 79.755 201.480 79.770 ;
        RECT 201.235 78.705 202.475 79.755 ;
        RECT 201.235 78.280 201.480 78.705 ;
        RECT 183.640 76.890 183.885 76.940 ;
        RECT 201.235 76.910 202.475 78.280 ;
        RECT 201.235 76.875 201.480 76.910 ;
        RECT 177.225 75.450 177.470 75.825 ;
      LAYER nwell ;
        RECT 178.885 75.260 180.745 76.700 ;
      LAYER pwell ;
        RECT 201.235 75.825 202.475 76.875 ;
      LAYER nwell ;
        RECT 202.895 76.700 206.235 93.400 ;
      LAYER pwell ;
        RECT 207.650 93.115 207.895 93.210 ;
        RECT 206.655 88.910 207.895 93.115 ;
        RECT 207.650 88.795 207.895 88.910 ;
        RECT 206.655 84.590 207.895 88.795 ;
        RECT 208.890 87.695 211.250 93.345 ;
      LAYER nwell ;
        RECT 211.300 87.650 213.760 93.395 ;
      LAYER pwell ;
        RECT 213.810 87.700 216.170 93.350 ;
      LAYER nwell ;
        RECT 216.220 87.650 220.610 93.400 ;
      LAYER pwell ;
        RECT 220.660 87.700 224.950 93.350 ;
        RECT 225.245 93.115 225.490 93.210 ;
        RECT 225.245 88.910 226.485 93.115 ;
        RECT 225.245 88.795 225.490 88.910 ;
      LAYER nwell ;
        RECT 211.300 87.645 220.610 87.650 ;
      LAYER pwell ;
        RECT 207.650 84.570 207.895 84.590 ;
        RECT 206.620 84.115 207.705 84.545 ;
        RECT 207.650 84.085 207.895 84.090 ;
        RECT 206.655 81.695 207.895 84.085 ;
        RECT 207.650 81.675 207.895 81.695 ;
        RECT 206.655 80.625 207.895 81.675 ;
        RECT 207.650 80.250 207.895 80.625 ;
      LAYER nwell ;
        RECT 208.840 83.290 220.610 87.645 ;
      LAYER pwell ;
        RECT 225.245 84.590 226.485 88.795 ;
        RECT 225.245 84.570 225.490 84.590 ;
        RECT 225.435 84.115 226.520 84.545 ;
        RECT 225.245 84.085 225.490 84.090 ;
      LAYER nwell ;
        RECT 208.840 83.285 216.220 83.290 ;
      LAYER pwell ;
        RECT 206.620 79.795 207.705 80.225 ;
        RECT 207.650 79.755 207.895 79.770 ;
        RECT 206.655 78.705 207.895 79.755 ;
        RECT 207.650 78.310 207.895 78.705 ;
        RECT 206.655 76.940 207.895 78.310 ;
      LAYER nwell ;
        RECT 208.840 77.535 211.300 83.285 ;
      LAYER pwell ;
        RECT 211.350 77.585 213.710 83.235 ;
      LAYER nwell ;
        RECT 213.760 77.540 216.220 83.285 ;
      LAYER pwell ;
        RECT 225.245 81.695 226.485 84.085 ;
        RECT 225.245 81.675 225.490 81.695 ;
        RECT 225.245 80.625 226.485 81.675 ;
        RECT 225.245 80.250 225.490 80.625 ;
        RECT 225.435 79.795 226.520 80.225 ;
        RECT 225.245 79.755 225.490 79.770 ;
        RECT 225.245 78.705 226.485 79.755 ;
        RECT 225.245 78.280 225.490 78.705 ;
        RECT 207.650 76.890 207.895 76.940 ;
        RECT 225.245 76.910 226.485 78.280 ;
        RECT 225.245 76.875 225.490 76.910 ;
        RECT 201.235 75.450 201.480 75.825 ;
      LAYER nwell ;
        RECT 202.895 75.260 204.755 76.700 ;
      LAYER pwell ;
        RECT 225.245 75.825 226.485 76.875 ;
      LAYER nwell ;
        RECT 226.905 76.700 230.245 93.400 ;
      LAYER pwell ;
        RECT 231.660 93.115 231.905 93.210 ;
        RECT 230.665 88.910 231.905 93.115 ;
        RECT 231.660 88.795 231.905 88.910 ;
        RECT 230.665 84.590 231.905 88.795 ;
        RECT 232.905 87.695 235.265 93.345 ;
      LAYER nwell ;
        RECT 235.315 87.650 237.775 93.395 ;
      LAYER pwell ;
        RECT 237.825 87.700 240.185 93.350 ;
      LAYER nwell ;
        RECT 240.235 87.650 244.625 93.400 ;
      LAYER pwell ;
        RECT 244.675 87.700 248.965 93.350 ;
        RECT 249.260 93.115 249.505 93.210 ;
        RECT 249.260 88.910 250.500 93.115 ;
        RECT 249.260 88.795 249.505 88.910 ;
      LAYER nwell ;
        RECT 235.315 87.645 244.625 87.650 ;
      LAYER pwell ;
        RECT 231.660 84.570 231.905 84.590 ;
        RECT 230.630 84.115 231.715 84.545 ;
        RECT 231.660 84.085 231.905 84.090 ;
        RECT 230.665 81.695 231.905 84.085 ;
        RECT 231.660 81.675 231.905 81.695 ;
        RECT 230.665 80.625 231.905 81.675 ;
        RECT 231.660 80.250 231.905 80.625 ;
      LAYER nwell ;
        RECT 232.855 83.290 244.625 87.645 ;
      LAYER pwell ;
        RECT 249.260 84.590 250.500 88.795 ;
        RECT 249.260 84.570 249.505 84.590 ;
        RECT 249.450 84.115 250.535 84.545 ;
        RECT 249.260 84.085 249.505 84.090 ;
      LAYER nwell ;
        RECT 232.855 83.285 240.235 83.290 ;
      LAYER pwell ;
        RECT 230.630 79.795 231.715 80.225 ;
        RECT 231.660 79.755 231.905 79.770 ;
        RECT 230.665 78.705 231.905 79.755 ;
        RECT 231.660 78.310 231.905 78.705 ;
        RECT 230.665 76.940 231.905 78.310 ;
      LAYER nwell ;
        RECT 232.855 77.535 235.315 83.285 ;
      LAYER pwell ;
        RECT 235.365 77.585 237.725 83.235 ;
      LAYER nwell ;
        RECT 237.775 77.540 240.235 83.285 ;
      LAYER pwell ;
        RECT 249.260 81.695 250.500 84.085 ;
        RECT 249.260 81.675 249.505 81.695 ;
        RECT 249.260 80.625 250.500 81.675 ;
        RECT 249.260 80.250 249.505 80.625 ;
        RECT 249.450 79.795 250.535 80.225 ;
        RECT 249.260 79.755 249.505 79.770 ;
        RECT 249.260 78.705 250.500 79.755 ;
        RECT 249.260 78.280 249.505 78.705 ;
        RECT 231.660 76.890 231.905 76.940 ;
        RECT 249.260 76.910 250.500 78.280 ;
        RECT 249.260 76.875 249.505 76.910 ;
        RECT 225.245 75.450 225.490 75.825 ;
      LAYER nwell ;
        RECT 226.905 75.260 228.765 76.700 ;
      LAYER pwell ;
        RECT 249.260 75.825 250.500 76.875 ;
      LAYER nwell ;
        RECT 250.920 76.700 254.260 93.400 ;
      LAYER pwell ;
        RECT 255.675 93.115 255.920 93.210 ;
        RECT 254.680 88.910 255.920 93.115 ;
        RECT 255.675 88.795 255.920 88.910 ;
        RECT 254.680 84.590 255.920 88.795 ;
        RECT 256.960 87.695 259.320 93.345 ;
      LAYER nwell ;
        RECT 259.370 87.650 261.830 93.395 ;
      LAYER pwell ;
        RECT 261.880 87.700 264.240 93.350 ;
      LAYER nwell ;
        RECT 264.290 87.650 268.680 93.400 ;
      LAYER pwell ;
        RECT 268.730 87.700 273.020 93.350 ;
        RECT 273.315 93.115 273.560 93.210 ;
        RECT 273.315 88.910 274.555 93.115 ;
        RECT 273.315 88.795 273.560 88.910 ;
      LAYER nwell ;
        RECT 259.370 87.645 268.680 87.650 ;
      LAYER pwell ;
        RECT 255.675 84.570 255.920 84.590 ;
        RECT 254.645 84.115 255.730 84.545 ;
        RECT 255.675 84.085 255.920 84.090 ;
        RECT 254.680 81.695 255.920 84.085 ;
        RECT 255.675 81.675 255.920 81.695 ;
        RECT 254.680 80.625 255.920 81.675 ;
        RECT 255.675 80.250 255.920 80.625 ;
      LAYER nwell ;
        RECT 256.910 83.290 268.680 87.645 ;
      LAYER pwell ;
        RECT 273.315 84.590 274.555 88.795 ;
        RECT 273.315 84.570 273.560 84.590 ;
        RECT 273.505 84.115 274.590 84.545 ;
        RECT 273.315 84.085 273.560 84.090 ;
      LAYER nwell ;
        RECT 256.910 83.285 264.290 83.290 ;
      LAYER pwell ;
        RECT 254.645 79.795 255.730 80.225 ;
        RECT 255.675 79.755 255.920 79.770 ;
        RECT 254.680 78.705 255.920 79.755 ;
        RECT 255.675 78.310 255.920 78.705 ;
        RECT 254.680 76.940 255.920 78.310 ;
      LAYER nwell ;
        RECT 256.910 77.535 259.370 83.285 ;
      LAYER pwell ;
        RECT 259.420 77.585 261.780 83.235 ;
      LAYER nwell ;
        RECT 261.830 77.540 264.290 83.285 ;
      LAYER pwell ;
        RECT 273.315 81.695 274.555 84.085 ;
        RECT 273.315 81.675 273.560 81.695 ;
        RECT 273.315 80.625 274.555 81.675 ;
        RECT 273.315 80.250 273.560 80.625 ;
        RECT 273.505 79.795 274.590 80.225 ;
        RECT 273.315 79.755 273.560 79.770 ;
        RECT 273.315 78.705 274.555 79.755 ;
        RECT 273.315 78.280 273.560 78.705 ;
        RECT 255.675 76.890 255.920 76.940 ;
        RECT 273.315 76.910 274.555 78.280 ;
        RECT 273.315 76.875 273.560 76.910 ;
        RECT 249.260 75.450 249.505 75.825 ;
      LAYER nwell ;
        RECT 250.920 75.260 252.780 76.700 ;
      LAYER pwell ;
        RECT 273.315 75.825 274.555 76.875 ;
      LAYER nwell ;
        RECT 274.975 76.700 278.315 93.400 ;
      LAYER pwell ;
        RECT 279.730 93.115 279.975 93.210 ;
        RECT 278.735 88.910 279.975 93.115 ;
        RECT 279.730 88.795 279.975 88.910 ;
        RECT 278.735 84.590 279.975 88.795 ;
        RECT 280.920 87.695 283.280 93.345 ;
      LAYER nwell ;
        RECT 283.330 87.650 285.790 93.395 ;
      LAYER pwell ;
        RECT 285.840 87.700 288.200 93.350 ;
      LAYER nwell ;
        RECT 288.250 87.650 292.640 93.400 ;
      LAYER pwell ;
        RECT 292.690 87.700 296.980 93.350 ;
        RECT 297.275 93.115 297.520 93.210 ;
        RECT 297.275 88.910 298.515 93.115 ;
        RECT 297.275 88.795 297.520 88.910 ;
      LAYER nwell ;
        RECT 283.330 87.645 292.640 87.650 ;
      LAYER pwell ;
        RECT 279.730 84.570 279.975 84.590 ;
        RECT 278.700 84.115 279.785 84.545 ;
        RECT 279.730 84.085 279.975 84.090 ;
        RECT 278.735 81.695 279.975 84.085 ;
        RECT 279.730 81.675 279.975 81.695 ;
        RECT 278.735 80.625 279.975 81.675 ;
        RECT 279.730 80.250 279.975 80.625 ;
      LAYER nwell ;
        RECT 280.870 83.290 292.640 87.645 ;
      LAYER pwell ;
        RECT 297.275 84.590 298.515 88.795 ;
        RECT 297.275 84.570 297.520 84.590 ;
        RECT 297.465 84.115 298.550 84.545 ;
        RECT 297.275 84.085 297.520 84.090 ;
      LAYER nwell ;
        RECT 280.870 83.285 288.250 83.290 ;
      LAYER pwell ;
        RECT 278.700 79.795 279.785 80.225 ;
        RECT 279.730 79.755 279.975 79.770 ;
        RECT 278.735 78.705 279.975 79.755 ;
        RECT 279.730 78.310 279.975 78.705 ;
        RECT 278.735 76.940 279.975 78.310 ;
      LAYER nwell ;
        RECT 280.870 77.535 283.330 83.285 ;
      LAYER pwell ;
        RECT 283.380 77.585 285.740 83.235 ;
      LAYER nwell ;
        RECT 285.790 77.540 288.250 83.285 ;
      LAYER pwell ;
        RECT 297.275 81.695 298.515 84.085 ;
        RECT 297.275 81.675 297.520 81.695 ;
        RECT 297.275 80.625 298.515 81.675 ;
        RECT 297.275 80.250 297.520 80.625 ;
        RECT 297.465 79.795 298.550 80.225 ;
        RECT 297.275 79.755 297.520 79.770 ;
        RECT 297.275 78.705 298.515 79.755 ;
        RECT 297.275 78.280 297.520 78.705 ;
        RECT 279.730 76.890 279.975 76.940 ;
        RECT 297.275 76.910 298.515 78.280 ;
        RECT 297.275 76.875 297.520 76.910 ;
        RECT 273.315 75.450 273.560 75.825 ;
      LAYER nwell ;
        RECT 274.975 75.260 276.835 76.700 ;
      LAYER pwell ;
        RECT 297.275 75.825 298.515 76.875 ;
      LAYER nwell ;
        RECT 298.935 76.700 302.275 93.400 ;
      LAYER pwell ;
        RECT 303.690 93.115 303.935 93.210 ;
        RECT 302.695 88.910 303.935 93.115 ;
        RECT 303.690 88.795 303.935 88.910 ;
        RECT 302.695 84.590 303.935 88.795 ;
        RECT 304.930 87.695 307.290 93.345 ;
      LAYER nwell ;
        RECT 307.340 87.650 309.800 93.395 ;
      LAYER pwell ;
        RECT 309.850 87.700 312.210 93.350 ;
      LAYER nwell ;
        RECT 312.260 87.650 316.650 93.400 ;
      LAYER pwell ;
        RECT 316.700 87.700 320.990 93.350 ;
        RECT 321.285 93.115 321.530 93.210 ;
        RECT 321.285 88.910 322.525 93.115 ;
        RECT 321.285 88.795 321.530 88.910 ;
      LAYER nwell ;
        RECT 307.340 87.645 316.650 87.650 ;
      LAYER pwell ;
        RECT 303.690 84.570 303.935 84.590 ;
        RECT 302.660 84.115 303.745 84.545 ;
        RECT 303.690 84.085 303.935 84.090 ;
        RECT 302.695 81.695 303.935 84.085 ;
        RECT 303.690 81.675 303.935 81.695 ;
        RECT 302.695 80.625 303.935 81.675 ;
        RECT 303.690 80.250 303.935 80.625 ;
      LAYER nwell ;
        RECT 304.880 83.290 316.650 87.645 ;
      LAYER pwell ;
        RECT 321.285 84.590 322.525 88.795 ;
        RECT 321.285 84.570 321.530 84.590 ;
        RECT 321.475 84.115 322.560 84.545 ;
        RECT 321.285 84.085 321.530 84.090 ;
      LAYER nwell ;
        RECT 304.880 83.285 312.260 83.290 ;
      LAYER pwell ;
        RECT 302.660 79.795 303.745 80.225 ;
        RECT 303.690 79.755 303.935 79.770 ;
        RECT 302.695 78.705 303.935 79.755 ;
        RECT 303.690 78.310 303.935 78.705 ;
        RECT 302.695 76.940 303.935 78.310 ;
      LAYER nwell ;
        RECT 304.880 77.535 307.340 83.285 ;
      LAYER pwell ;
        RECT 307.390 77.585 309.750 83.235 ;
      LAYER nwell ;
        RECT 309.800 77.540 312.260 83.285 ;
      LAYER pwell ;
        RECT 321.285 81.695 322.525 84.085 ;
        RECT 321.285 81.675 321.530 81.695 ;
        RECT 321.285 80.625 322.525 81.675 ;
        RECT 321.285 80.250 321.530 80.625 ;
        RECT 321.475 79.795 322.560 80.225 ;
        RECT 321.285 79.755 321.530 79.770 ;
        RECT 321.285 78.705 322.525 79.755 ;
        RECT 321.285 78.280 321.530 78.705 ;
        RECT 303.690 76.890 303.935 76.940 ;
        RECT 321.285 76.910 322.525 78.280 ;
        RECT 321.285 76.875 321.530 76.910 ;
        RECT 297.275 75.450 297.520 75.825 ;
      LAYER nwell ;
        RECT 298.935 75.260 300.795 76.700 ;
      LAYER pwell ;
        RECT 321.285 75.825 322.525 76.875 ;
      LAYER nwell ;
        RECT 322.945 76.700 326.285 93.400 ;
      LAYER pwell ;
        RECT 327.700 93.115 327.945 93.210 ;
        RECT 326.705 88.910 327.945 93.115 ;
        RECT 327.700 88.795 327.945 88.910 ;
        RECT 326.705 84.590 327.945 88.795 ;
        RECT 327.700 84.570 327.945 84.590 ;
        RECT 326.670 84.115 327.755 84.545 ;
        RECT 327.700 84.085 327.945 84.090 ;
        RECT 326.705 81.695 327.945 84.085 ;
        RECT 327.700 81.675 327.945 81.695 ;
        RECT 326.705 80.625 327.945 81.675 ;
        RECT 327.700 80.250 327.945 80.625 ;
        RECT 326.670 79.795 327.755 80.225 ;
        RECT 327.700 79.755 327.945 79.770 ;
        RECT 326.705 78.705 327.945 79.755 ;
        RECT 327.700 78.310 327.945 78.705 ;
        RECT 326.705 76.940 327.945 78.310 ;
        RECT 327.700 76.890 327.945 76.940 ;
        RECT 321.285 75.450 321.530 75.825 ;
      LAYER nwell ;
        RECT 322.945 75.260 324.805 76.700 ;
        RECT 80.365 59.845 82.225 67.425 ;
      LAYER pwell ;
        RECT 83.640 67.165 83.885 67.235 ;
        RECT 82.580 63.480 83.885 67.165 ;
        RECT 83.640 63.395 83.885 63.480 ;
        RECT 82.610 62.940 83.695 63.370 ;
        RECT 83.640 62.865 83.885 62.915 ;
        RECT 82.645 61.495 83.885 62.865 ;
        RECT 83.640 61.425 83.885 61.495 ;
        RECT 82.645 60.055 83.885 61.425 ;
        RECT 83.640 60.035 83.885 60.055 ;
        RECT 75.130 56.450 76.390 57.880 ;
        RECT 75.240 56.000 76.280 56.430 ;
      LAYER nwell ;
        RECT 76.690 55.430 84.420 57.930 ;
      LAYER pwell ;
        RECT 84.720 56.450 85.980 57.880 ;
        RECT 84.830 56.000 85.870 56.430 ;
        RECT 75.385 52.845 75.630 52.965 ;
        RECT 75.385 51.660 76.755 52.845 ;
        RECT 75.385 50.715 76.835 51.660 ;
        RECT 75.385 50.565 75.630 50.715 ;
      LAYER nwell ;
        RECT 77.045 50.375 84.065 53.155 ;
      LAYER pwell ;
        RECT 85.480 52.845 85.725 52.965 ;
        RECT 84.355 51.660 85.725 52.845 ;
        RECT 84.275 50.715 85.725 51.660 ;
        RECT 85.480 50.565 85.725 50.715 ;
        RECT 74.295 49.795 75.675 50.225 ;
        RECT 74.355 45.355 75.615 49.775 ;
        RECT 74.295 44.905 75.675 45.335 ;
      LAYER nwell ;
        RECT 75.825 44.755 85.285 50.375 ;
      LAYER pwell ;
        RECT 85.435 49.795 86.815 50.225 ;
        RECT 85.495 45.355 86.755 49.775 ;
        RECT 85.435 44.905 86.815 45.335 ;
      LAYER nwell ;
        RECT 44.420 37.645 55.840 39.505 ;
        RECT 105.280 37.645 116.700 39.505 ;
      LAYER pwell ;
        RECT 44.635 36.175 45.065 37.260 ;
        RECT 45.095 36.230 55.630 37.225 ;
        RECT 105.490 36.230 116.025 37.225 ;
        RECT 45.090 35.985 55.650 36.230 ;
        RECT 105.470 35.985 116.030 36.230 ;
        RECT 116.055 36.175 116.485 37.260 ;
        RECT 50.190 30.640 53.780 34.140 ;
        RECT 50.190 30.450 55.360 30.640 ;
        RECT 51.770 19.690 55.360 30.450 ;
        RECT 58.580 28.605 80.270 33.775 ;
        RECT 80.850 28.605 102.540 33.775 ;
        RECT 107.340 30.640 110.930 34.140 ;
        RECT 105.760 30.450 110.930 30.640 ;
        RECT 105.760 19.690 109.350 30.450 ;
        RECT 51.770 18.380 53.780 19.690 ;
        RECT 50.190 16.190 53.780 18.380 ;
      LAYER nwell ;
        RECT 62.545 18.005 75.405 19.435 ;
        RECT 50.140 13.550 52.250 16.140 ;
        RECT 62.545 8.005 63.975 18.005 ;
        RECT 67.250 10.300 70.940 16.140 ;
        RECT 73.975 8.005 75.405 18.005 ;
        RECT 62.545 6.575 75.405 8.005 ;
        RECT 85.720 17.970 98.520 19.400 ;
        RECT 85.720 8.030 87.150 17.970 ;
        RECT 90.180 10.300 93.870 16.140 ;
        RECT 97.090 8.030 98.520 17.970 ;
      LAYER pwell ;
        RECT 107.340 18.380 109.350 19.690 ;
        RECT 107.340 16.190 110.930 18.380 ;
      LAYER nwell ;
        RECT 108.870 13.550 110.980 16.140 ;
        RECT 85.720 6.600 98.520 8.030 ;
      LAYER li1 ;
        RECT 129.120 151.365 129.290 151.850 ;
        RECT 129.120 151.035 130.335 151.365 ;
        RECT 130.505 151.035 130.985 151.725 ;
        RECT 132.450 151.365 132.620 151.850 ;
        RECT 131.155 151.035 132.620 151.365 ;
        RECT 129.120 150.280 129.290 151.035 ;
        RECT 129.555 150.535 132.185 150.865 ;
        RECT 130.490 150.305 130.690 150.535 ;
        RECT 132.450 150.305 132.620 151.035 ;
        RECT 153.130 151.365 153.300 151.850 ;
        RECT 153.130 151.035 154.345 151.365 ;
        RECT 154.515 151.035 154.995 151.725 ;
        RECT 156.460 151.365 156.630 151.850 ;
        RECT 155.165 151.035 156.630 151.365 ;
        RECT 129.120 149.950 130.215 150.280 ;
        RECT 130.385 149.975 130.755 150.305 ;
        RECT 131.025 149.975 134.045 150.305 ;
        RECT 134.315 149.975 134.685 150.305 ;
        RECT 112.980 149.415 115.080 149.585 ;
        RECT 10.200 143.535 69.720 143.705 ;
        RECT 10.370 142.035 10.940 143.535 ;
        RECT 11.650 142.815 11.980 143.535 ;
        RECT 12.685 142.810 13.045 143.270 ;
        RECT 13.215 142.810 13.465 143.535 ;
        RECT 13.635 142.830 13.975 143.270 ;
        RECT 14.155 142.830 14.405 143.535 ;
        RECT 10.295 140.375 10.625 141.690 ;
        RECT 11.345 140.375 11.915 142.370 ;
        RECT 12.685 141.300 12.855 142.810 ;
        RECT 13.025 141.470 13.435 142.610 ;
        RECT 13.635 141.800 13.805 142.830 ;
        RECT 14.605 142.810 14.980 143.140 ;
        RECT 15.150 142.810 15.480 143.535 ;
        RECT 13.975 141.990 14.305 142.660 ;
        RECT 13.635 141.470 13.965 141.800 ;
        RECT 14.135 141.300 14.305 141.990 ;
        RECT 12.685 141.130 14.305 141.300 ;
        RECT 14.605 142.040 14.775 142.810 ;
        RECT 15.650 142.640 15.980 143.270 ;
        RECT 16.160 142.810 16.330 143.535 ;
        RECT 16.510 142.640 16.840 143.270 ;
        RECT 17.020 142.810 17.270 143.535 ;
        RECT 14.945 142.210 15.345 142.540 ;
        RECT 15.650 142.470 16.865 142.640 ;
        RECT 15.515 142.040 16.525 142.270 ;
        RECT 14.605 141.870 16.525 142.040 ;
        RECT 12.685 140.640 12.985 141.130 ;
        RECT 13.185 140.375 13.515 140.960 ;
        RECT 14.085 140.375 14.415 140.960 ;
        RECT 14.605 140.640 14.985 141.870 ;
        RECT 16.695 141.700 16.865 142.470 ;
        RECT 17.995 142.610 18.325 143.170 ;
        RECT 18.505 142.780 18.835 143.535 ;
        RECT 17.995 142.440 18.795 142.610 ;
        RECT 19.005 142.440 19.335 143.270 ;
        RECT 19.515 142.490 19.765 143.535 ;
        RECT 20.365 142.810 20.740 143.140 ;
        RECT 20.910 142.810 21.240 143.535 ;
        RECT 18.005 141.840 18.455 142.270 ;
        RECT 15.155 140.375 15.405 141.700 ;
        RECT 15.605 141.530 16.865 141.700 ;
        RECT 15.605 140.640 15.935 141.530 ;
        RECT 16.135 140.375 16.385 141.360 ;
        RECT 16.585 140.640 16.865 141.530 ;
        RECT 17.035 140.375 17.285 141.800 ;
        RECT 17.995 141.300 18.350 141.670 ;
        RECT 18.625 141.300 18.795 142.440 ;
        RECT 18.965 141.470 19.335 142.440 ;
        RECT 19.505 141.990 20.175 142.320 ;
        RECT 20.365 142.040 20.535 142.810 ;
        RECT 21.410 142.640 21.740 143.270 ;
        RECT 21.920 142.810 22.090 143.535 ;
        RECT 22.270 142.640 22.600 143.270 ;
        RECT 22.780 142.810 23.030 143.535 ;
        RECT 20.705 142.210 21.105 142.540 ;
        RECT 21.410 142.470 22.625 142.640 ;
        RECT 23.250 142.515 23.550 143.535 ;
        RECT 23.755 142.490 24.005 143.535 ;
        RECT 24.185 142.490 24.515 143.270 ;
        RECT 21.275 142.040 22.285 142.270 ;
        RECT 19.505 141.300 19.675 141.990 ;
        RECT 20.365 141.870 22.285 142.040 ;
        RECT 17.995 141.130 19.675 141.300 ;
        RECT 17.995 140.740 18.350 141.130 ;
        RECT 18.555 140.375 18.885 140.960 ;
        RECT 19.860 140.885 20.165 141.800 ;
        RECT 19.455 140.375 20.165 140.885 ;
        RECT 20.365 140.640 20.745 141.870 ;
        RECT 22.455 141.700 22.625 142.470 ;
        RECT 20.915 140.375 21.165 141.700 ;
        RECT 21.365 141.530 22.625 141.700 ;
        RECT 21.365 140.640 21.695 141.530 ;
        RECT 21.895 140.375 22.145 141.360 ;
        RECT 22.345 140.640 22.625 141.530 ;
        RECT 22.795 140.375 23.045 141.800 ;
        RECT 23.250 140.375 23.550 141.415 ;
        RECT 23.755 140.375 24.085 141.800 ;
        RECT 24.255 141.735 24.515 142.490 ;
        RECT 24.745 142.235 25.075 143.270 ;
        RECT 25.255 142.775 25.505 143.535 ;
        RECT 25.735 142.605 26.065 143.235 ;
        RECT 26.605 142.775 26.935 143.535 ;
        RECT 27.260 143.195 29.200 143.365 ;
        RECT 29.370 143.225 29.765 143.535 ;
        RECT 27.260 142.605 27.430 143.195 ;
        RECT 29.030 143.055 29.200 143.195 ;
        RECT 30.245 143.120 32.170 143.290 ;
        RECT 30.245 143.055 30.415 143.120 ;
        RECT 27.600 142.775 28.360 143.025 ;
        RECT 25.490 142.435 27.090 142.605 ;
        RECT 24.745 141.905 25.295 142.235 ;
        RECT 24.255 140.640 24.955 141.735 ;
        RECT 25.125 140.715 25.295 141.905 ;
        RECT 25.490 141.765 25.660 142.435 ;
        RECT 26.760 142.275 27.090 142.435 ;
        RECT 27.260 142.275 27.990 142.605 ;
        RECT 25.830 142.105 26.160 142.265 ;
        RECT 25.830 141.935 27.215 142.105 ;
        RECT 25.490 141.595 26.165 141.765 ;
        RECT 25.495 140.375 25.825 141.425 ;
        RECT 25.995 141.175 26.165 141.595 ;
        RECT 26.335 141.365 26.875 141.700 ;
        RECT 25.995 140.715 26.360 141.175 ;
        RECT 26.545 140.375 26.875 141.175 ;
        RECT 27.045 141.145 27.215 141.935 ;
        RECT 27.385 141.315 27.715 142.275 ;
        RECT 28.190 142.105 28.360 142.775 ;
        RECT 28.030 141.935 28.360 142.105 ;
        RECT 28.530 142.715 28.860 142.955 ;
        RECT 29.030 142.885 30.415 143.055 ;
        RECT 28.530 142.545 30.415 142.715 ;
        RECT 28.530 142.490 28.860 142.545 ;
        RECT 28.030 141.145 28.200 141.935 ;
        RECT 28.530 141.755 28.700 142.490 ;
        RECT 29.030 142.045 30.065 142.375 ;
        RECT 27.045 140.815 28.200 141.145 ;
        RECT 28.370 140.865 28.700 141.755 ;
        RECT 28.870 140.375 29.200 141.875 ;
        RECT 29.395 141.470 29.725 141.825 ;
        RECT 29.895 141.300 30.065 142.045 ;
        RECT 30.235 141.495 30.415 142.545 ;
        RECT 30.585 142.570 31.055 142.950 ;
        RECT 29.430 141.220 30.065 141.300 ;
        RECT 30.585 141.220 30.755 142.570 ;
        RECT 31.225 142.400 31.475 142.950 ;
        RECT 30.925 142.230 31.475 142.400 ;
        RECT 31.645 142.820 32.170 143.120 ;
        RECT 32.340 142.820 32.670 143.535 ;
        RECT 30.925 141.560 31.095 142.230 ;
        RECT 31.645 142.060 31.815 142.820 ;
        RECT 32.840 142.650 33.225 143.270 ;
        RECT 33.400 142.790 33.650 143.535 ;
        RECT 34.220 142.960 34.550 143.250 ;
        RECT 33.825 142.790 34.550 142.960 ;
        RECT 31.985 142.480 33.225 142.650 ;
        RECT 31.985 142.070 32.235 142.480 ;
        RECT 31.265 141.900 31.815 142.060 ;
        RECT 32.405 141.980 32.885 142.310 ;
        RECT 31.265 141.730 32.165 141.900 ;
        RECT 32.405 141.840 32.635 141.980 ;
        RECT 33.055 141.810 33.225 142.480 ;
        RECT 30.925 141.390 31.670 141.560 ;
        RECT 31.915 141.450 32.165 141.730 ;
        RECT 32.815 141.480 33.225 141.810 ;
        RECT 33.395 141.480 33.655 142.490 ;
        RECT 31.420 141.280 31.670 141.390 ;
        RECT 33.825 141.310 33.995 142.790 ;
        RECT 34.165 141.450 34.555 142.620 ;
        RECT 36.210 142.515 36.510 143.535 ;
        RECT 37.645 142.810 38.020 143.140 ;
        RECT 38.190 142.810 38.520 143.535 ;
        RECT 37.645 142.040 37.815 142.810 ;
        RECT 38.690 142.640 39.020 143.270 ;
        RECT 39.200 142.810 39.370 143.535 ;
        RECT 39.550 142.640 39.880 143.270 ;
        RECT 40.060 142.810 40.310 143.535 ;
        RECT 40.525 142.810 40.900 143.140 ;
        RECT 41.070 142.810 41.400 143.535 ;
        RECT 37.985 142.210 38.385 142.540 ;
        RECT 38.690 142.470 39.905 142.640 ;
        RECT 38.555 142.040 39.565 142.270 ;
        RECT 37.645 141.870 39.565 142.040 ;
        RECT 33.005 141.280 33.995 141.310 ;
        RECT 29.430 141.050 31.220 141.220 ;
        RECT 30.890 140.895 31.220 141.050 ;
        RECT 31.420 141.140 33.995 141.280 ;
        RECT 31.420 141.110 33.175 141.140 ;
        RECT 31.420 140.895 31.670 141.110 ;
        RECT 33.795 141.100 33.995 141.140 ;
        RECT 29.965 140.375 30.295 140.880 ;
        RECT 32.365 140.375 32.695 140.940 ;
        RECT 33.345 140.375 33.595 140.970 ;
        RECT 33.795 140.640 34.125 141.100 ;
        RECT 34.325 140.375 34.575 141.100 ;
        RECT 36.210 140.375 36.510 141.415 ;
        RECT 37.645 140.640 38.025 141.870 ;
        RECT 39.735 141.700 39.905 142.470 ;
        RECT 40.525 142.040 40.695 142.810 ;
        RECT 41.570 142.640 41.900 143.270 ;
        RECT 42.080 142.810 42.250 143.535 ;
        RECT 42.430 142.640 42.760 143.270 ;
        RECT 42.940 142.810 43.190 143.535 ;
        RECT 43.405 142.810 43.780 143.140 ;
        RECT 43.950 142.810 44.280 143.535 ;
        RECT 40.865 142.210 41.265 142.540 ;
        RECT 41.570 142.470 42.785 142.640 ;
        RECT 41.435 142.040 42.445 142.270 ;
        RECT 40.525 141.870 42.445 142.040 ;
        RECT 38.195 140.375 38.445 141.700 ;
        RECT 38.645 141.530 39.905 141.700 ;
        RECT 38.645 140.640 38.975 141.530 ;
        RECT 39.175 140.375 39.425 141.360 ;
        RECT 39.625 140.640 39.905 141.530 ;
        RECT 40.075 140.375 40.325 141.800 ;
        RECT 40.525 140.640 40.905 141.870 ;
        RECT 42.615 141.700 42.785 142.470 ;
        RECT 43.405 142.040 43.575 142.810 ;
        RECT 44.450 142.640 44.780 143.270 ;
        RECT 44.960 142.810 45.130 143.535 ;
        RECT 45.310 142.640 45.640 143.270 ;
        RECT 45.820 142.810 46.070 143.535 ;
        RECT 46.330 142.810 46.580 143.535 ;
        RECT 46.760 142.640 47.090 143.270 ;
        RECT 47.270 142.810 47.440 143.535 ;
        RECT 47.620 142.640 47.950 143.270 ;
        RECT 48.120 142.810 48.450 143.535 ;
        RECT 48.620 142.810 48.995 143.140 ;
        RECT 43.745 142.210 44.145 142.540 ;
        RECT 44.450 142.470 45.665 142.640 ;
        RECT 44.315 142.040 45.325 142.270 ;
        RECT 43.405 141.870 45.325 142.040 ;
        RECT 41.075 140.375 41.325 141.700 ;
        RECT 41.525 141.530 42.785 141.700 ;
        RECT 41.525 140.640 41.855 141.530 ;
        RECT 42.055 140.375 42.305 141.360 ;
        RECT 42.505 140.640 42.785 141.530 ;
        RECT 42.955 140.375 43.205 141.800 ;
        RECT 43.405 140.640 43.785 141.870 ;
        RECT 45.495 141.700 45.665 142.470 ;
        RECT 46.735 142.470 47.950 142.640 ;
        RECT 43.955 140.375 44.205 141.700 ;
        RECT 44.405 141.530 45.665 141.700 ;
        RECT 44.405 140.640 44.735 141.530 ;
        RECT 44.935 140.375 45.185 141.360 ;
        RECT 45.385 140.640 45.665 141.530 ;
        RECT 45.835 140.375 46.085 141.800 ;
        RECT 46.315 140.375 46.565 141.800 ;
        RECT 46.735 141.700 46.905 142.470 ;
        RECT 47.075 142.040 48.085 142.270 ;
        RECT 48.255 142.210 48.655 142.540 ;
        RECT 48.825 142.040 48.995 142.810 ;
        RECT 49.170 142.515 49.470 143.535 ;
        RECT 49.645 142.810 50.020 143.140 ;
        RECT 50.190 142.810 50.520 143.535 ;
        RECT 47.075 141.870 48.995 142.040 ;
        RECT 46.735 141.530 47.995 141.700 ;
        RECT 46.735 140.640 47.015 141.530 ;
        RECT 47.215 140.375 47.465 141.360 ;
        RECT 47.665 140.640 47.995 141.530 ;
        RECT 48.195 140.375 48.445 141.700 ;
        RECT 48.615 140.640 48.995 141.870 ;
        RECT 49.645 142.040 49.815 142.810 ;
        RECT 50.690 142.640 51.020 143.270 ;
        RECT 51.200 142.810 51.370 143.535 ;
        RECT 51.550 142.640 51.880 143.270 ;
        RECT 52.060 142.810 52.310 143.535 ;
        RECT 49.985 142.210 50.385 142.540 ;
        RECT 50.690 142.470 51.905 142.640 ;
        RECT 50.555 142.040 51.565 142.270 ;
        RECT 49.645 141.870 51.565 142.040 ;
        RECT 49.170 140.375 49.470 141.415 ;
        RECT 49.645 140.640 50.025 141.870 ;
        RECT 51.735 141.700 51.905 142.470 ;
        RECT 52.610 142.035 53.180 143.535 ;
        RECT 53.890 142.815 54.220 143.535 ;
        RECT 54.925 142.810 55.300 143.140 ;
        RECT 55.470 142.810 55.800 143.535 ;
        RECT 50.195 140.375 50.445 141.700 ;
        RECT 50.645 141.530 51.905 141.700 ;
        RECT 50.645 140.640 50.975 141.530 ;
        RECT 51.175 140.375 51.425 141.360 ;
        RECT 51.625 140.640 51.905 141.530 ;
        RECT 52.075 140.375 52.325 141.800 ;
        RECT 52.535 140.375 52.865 141.690 ;
        RECT 53.585 140.375 54.155 142.370 ;
        RECT 54.925 142.040 55.095 142.810 ;
        RECT 55.970 142.640 56.300 143.270 ;
        RECT 56.480 142.810 56.650 143.535 ;
        RECT 56.830 142.640 57.160 143.270 ;
        RECT 57.340 142.810 57.590 143.535 ;
        RECT 59.290 142.810 59.540 143.535 ;
        RECT 59.720 142.640 60.050 143.270 ;
        RECT 60.230 142.810 60.400 143.535 ;
        RECT 60.580 142.640 60.910 143.270 ;
        RECT 61.080 142.810 61.410 143.535 ;
        RECT 61.580 142.810 61.955 143.140 ;
        RECT 55.265 142.210 55.665 142.540 ;
        RECT 55.970 142.470 57.185 142.640 ;
        RECT 55.835 142.040 56.845 142.270 ;
        RECT 54.925 141.870 56.845 142.040 ;
        RECT 54.925 140.640 55.305 141.870 ;
        RECT 57.015 141.700 57.185 142.470 ;
        RECT 59.695 142.470 60.910 142.640 ;
        RECT 55.475 140.375 55.725 141.700 ;
        RECT 55.925 141.530 57.185 141.700 ;
        RECT 55.925 140.640 56.255 141.530 ;
        RECT 56.455 140.375 56.705 141.360 ;
        RECT 56.905 140.640 57.185 141.530 ;
        RECT 57.355 140.375 57.605 141.800 ;
        RECT 59.275 140.375 59.525 141.800 ;
        RECT 59.695 141.700 59.865 142.470 ;
        RECT 60.035 142.040 61.045 142.270 ;
        RECT 61.215 142.210 61.615 142.540 ;
        RECT 61.785 142.040 61.955 142.810 ;
        RECT 62.130 142.515 62.430 143.535 ;
        RECT 62.605 142.810 62.980 143.140 ;
        RECT 63.150 142.810 63.480 143.535 ;
        RECT 60.035 141.870 61.955 142.040 ;
        RECT 59.695 141.530 60.955 141.700 ;
        RECT 59.695 140.640 59.975 141.530 ;
        RECT 60.175 140.375 60.425 141.360 ;
        RECT 60.625 140.640 60.955 141.530 ;
        RECT 61.155 140.375 61.405 141.700 ;
        RECT 61.575 140.640 61.955 141.870 ;
        RECT 62.605 142.040 62.775 142.810 ;
        RECT 63.650 142.640 63.980 143.270 ;
        RECT 64.160 142.810 64.330 143.535 ;
        RECT 64.510 142.640 64.840 143.270 ;
        RECT 65.020 142.810 65.270 143.535 ;
        RECT 65.515 142.830 65.845 143.270 ;
        RECT 66.015 142.940 66.705 143.535 ;
        RECT 62.945 142.210 63.345 142.540 ;
        RECT 63.650 142.470 64.865 142.640 ;
        RECT 63.515 142.040 64.525 142.270 ;
        RECT 62.605 141.870 64.525 142.040 ;
        RECT 62.130 140.375 62.430 141.415 ;
        RECT 62.605 140.640 62.985 141.870 ;
        RECT 64.695 141.700 64.865 142.470 ;
        RECT 65.515 141.800 65.755 142.830 ;
        RECT 66.875 142.660 67.205 143.270 ;
        RECT 67.940 142.815 68.270 143.535 ;
        RECT 65.925 142.490 67.205 142.660 ;
        RECT 65.925 141.990 66.315 142.490 ;
        RECT 63.155 140.375 63.405 141.700 ;
        RECT 63.605 141.530 64.865 141.700 ;
        RECT 63.605 140.640 63.935 141.530 ;
        RECT 64.135 140.375 64.385 141.360 ;
        RECT 64.585 140.640 64.865 141.530 ;
        RECT 65.035 140.375 65.285 141.800 ;
        RECT 65.515 140.640 65.975 141.800 ;
        RECT 66.145 141.670 66.315 141.990 ;
        RECT 66.485 141.840 67.195 142.320 ;
        RECT 66.145 141.500 66.975 141.670 ;
        RECT 66.145 140.375 66.475 141.330 ;
        RECT 66.645 140.640 66.975 141.500 ;
        RECT 68.005 140.375 68.575 142.370 ;
        RECT 68.980 142.035 69.550 143.535 ;
        RECT 69.295 140.375 69.625 141.690 ;
        RECT 10.200 140.205 69.720 140.375 ;
        RECT 10.295 138.890 10.625 140.205 ;
        RECT 10.370 137.045 10.940 138.545 ;
        RECT 11.345 138.210 11.915 140.205 ;
        RECT 12.235 138.780 12.565 140.205 ;
        RECT 12.735 138.845 13.435 139.940 ;
        RECT 12.735 138.090 12.995 138.845 ;
        RECT 13.605 138.675 13.775 139.865 ;
        RECT 13.975 139.155 14.305 140.205 ;
        RECT 14.475 139.405 14.840 139.865 ;
        RECT 15.025 139.405 15.355 140.205 ;
        RECT 15.525 139.435 16.680 139.765 ;
        RECT 14.475 138.985 14.645 139.405 ;
        RECT 11.650 137.045 11.980 137.765 ;
        RECT 12.235 137.045 12.485 138.090 ;
        RECT 12.665 137.310 12.995 138.090 ;
        RECT 13.225 138.345 13.775 138.675 ;
        RECT 13.970 138.815 14.645 138.985 ;
        RECT 14.815 138.880 15.355 139.215 ;
        RECT 13.225 137.310 13.555 138.345 ;
        RECT 13.970 138.145 14.140 138.815 ;
        RECT 15.525 138.645 15.695 139.435 ;
        RECT 14.310 138.475 15.695 138.645 ;
        RECT 14.310 138.315 14.640 138.475 ;
        RECT 15.865 138.305 16.195 139.265 ;
        RECT 16.510 138.645 16.680 139.435 ;
        RECT 16.850 138.825 17.180 139.715 ;
        RECT 16.510 138.475 16.840 138.645 ;
        RECT 15.240 138.145 15.570 138.305 ;
        RECT 13.970 137.975 15.570 138.145 ;
        RECT 15.740 137.975 16.470 138.305 ;
        RECT 13.735 137.045 13.985 137.805 ;
        RECT 14.215 137.345 14.545 137.975 ;
        RECT 15.085 137.045 15.415 137.805 ;
        RECT 15.740 137.385 15.910 137.975 ;
        RECT 16.670 137.805 16.840 138.475 ;
        RECT 16.080 137.555 16.840 137.805 ;
        RECT 17.010 138.090 17.180 138.825 ;
        RECT 17.350 138.705 17.680 140.205 ;
        RECT 18.445 139.700 18.775 140.205 ;
        RECT 19.370 139.530 19.700 139.685 ;
        RECT 17.910 139.360 19.700 139.530 ;
        RECT 19.900 139.470 20.150 139.685 ;
        RECT 20.845 139.640 21.175 140.205 ;
        RECT 21.825 139.610 22.075 140.205 ;
        RECT 22.275 139.480 22.605 139.940 ;
        RECT 22.805 139.480 23.055 140.205 ;
        RECT 19.900 139.440 21.655 139.470 ;
        RECT 22.275 139.440 22.475 139.480 ;
        RECT 17.910 139.280 18.545 139.360 ;
        RECT 17.875 138.755 18.205 139.110 ;
        RECT 18.375 138.535 18.545 139.280 ;
        RECT 17.510 138.205 18.545 138.535 ;
        RECT 17.010 138.035 17.340 138.090 ;
        RECT 18.715 138.035 18.895 139.085 ;
        RECT 17.010 137.865 18.895 138.035 ;
        RECT 19.065 138.010 19.235 139.360 ;
        RECT 19.900 139.300 22.475 139.440 ;
        RECT 19.900 139.190 20.150 139.300 ;
        RECT 21.485 139.270 22.475 139.300 ;
        RECT 19.405 139.020 20.150 139.190 ;
        RECT 19.405 138.350 19.575 139.020 ;
        RECT 20.395 138.850 20.645 139.130 ;
        RECT 19.745 138.680 20.645 138.850 ;
        RECT 21.295 138.770 21.705 139.100 ;
        RECT 19.745 138.520 20.295 138.680 ;
        RECT 19.405 138.180 19.955 138.350 ;
        RECT 17.010 137.625 17.340 137.865 ;
        RECT 17.510 137.525 18.895 137.695 ;
        RECT 19.065 137.630 19.535 138.010 ;
        RECT 19.705 137.630 19.955 138.180 ;
        RECT 20.125 137.760 20.295 138.520 ;
        RECT 20.885 138.600 21.115 138.740 ;
        RECT 20.465 138.100 20.715 138.510 ;
        RECT 20.885 138.270 21.365 138.600 ;
        RECT 21.535 138.100 21.705 138.770 ;
        RECT 20.465 137.930 21.705 138.100 ;
        RECT 21.875 138.090 22.135 139.100 ;
        RECT 17.510 137.385 17.680 137.525 ;
        RECT 15.740 137.215 17.680 137.385 ;
        RECT 18.725 137.460 18.895 137.525 ;
        RECT 20.125 137.460 20.650 137.760 ;
        RECT 17.850 137.045 18.245 137.355 ;
        RECT 18.725 137.290 20.650 137.460 ;
        RECT 20.820 137.045 21.150 137.760 ;
        RECT 21.320 137.310 21.705 137.930 ;
        RECT 22.305 137.790 22.475 139.270 ;
        RECT 23.250 139.165 23.550 140.205 ;
        RECT 23.755 139.695 24.465 140.205 ;
        RECT 22.645 137.960 23.035 139.130 ;
        RECT 23.755 138.780 24.060 139.695 ;
        RECT 25.035 139.620 25.365 140.205 ;
        RECT 25.570 139.450 25.925 139.840 ;
        RECT 24.245 139.280 25.925 139.450 ;
        RECT 24.245 138.590 24.415 139.280 ;
        RECT 23.745 138.260 24.415 138.590 ;
        RECT 24.585 138.140 24.955 139.110 ;
        RECT 25.125 138.140 25.295 139.280 ;
        RECT 25.570 138.910 25.925 139.280 ;
        RECT 25.465 138.310 25.915 138.740 ;
        RECT 26.125 138.710 26.505 139.940 ;
        RECT 26.675 138.880 26.925 140.205 ;
        RECT 27.125 139.050 27.455 139.940 ;
        RECT 27.655 139.220 27.905 140.205 ;
        RECT 28.105 139.050 28.385 139.940 ;
        RECT 27.125 138.880 28.385 139.050 ;
        RECT 26.125 138.540 28.045 138.710 ;
        RECT 21.880 137.045 22.130 137.790 ;
        RECT 22.305 137.620 23.030 137.790 ;
        RECT 22.700 137.330 23.030 137.620 ;
        RECT 23.250 137.045 23.550 138.065 ;
        RECT 24.155 137.045 24.405 138.090 ;
        RECT 24.585 137.310 24.915 138.140 ;
        RECT 25.125 137.970 25.925 138.140 ;
        RECT 25.085 137.045 25.415 137.800 ;
        RECT 25.595 137.410 25.925 137.970 ;
        RECT 26.125 137.770 26.295 138.540 ;
        RECT 26.465 138.040 26.865 138.370 ;
        RECT 27.035 138.310 28.045 138.540 ;
        RECT 28.215 138.110 28.385 138.880 ;
        RECT 28.555 138.780 28.805 140.205 ;
        RECT 29.015 138.890 29.345 140.205 ;
        RECT 27.170 137.940 28.385 138.110 ;
        RECT 26.125 137.440 26.500 137.770 ;
        RECT 26.670 137.045 27.000 137.770 ;
        RECT 27.170 137.310 27.500 137.940 ;
        RECT 27.680 137.045 27.850 137.770 ;
        RECT 28.030 137.310 28.360 137.940 ;
        RECT 28.540 137.045 28.790 137.770 ;
        RECT 29.090 137.045 29.660 138.545 ;
        RECT 30.065 138.210 30.635 140.205 ;
        RECT 31.425 139.620 31.755 140.205 ;
        RECT 32.325 139.620 32.655 140.205 ;
        RECT 32.855 139.450 33.155 139.940 ;
        RECT 33.345 139.480 33.595 140.205 ;
        RECT 33.795 139.480 34.125 139.940 ;
        RECT 34.325 139.610 34.575 140.205 ;
        RECT 35.225 139.640 35.555 140.205 ;
        RECT 37.625 139.700 37.955 140.205 ;
        RECT 31.535 139.280 33.155 139.450 ;
        RECT 31.535 138.590 31.705 139.280 ;
        RECT 31.875 138.780 32.205 139.110 ;
        RECT 31.535 137.920 31.865 138.590 ;
        RECT 30.370 137.045 30.700 137.765 ;
        RECT 32.035 137.750 32.205 138.780 ;
        RECT 32.405 137.970 32.815 139.110 ;
        RECT 32.985 137.770 33.155 139.280 ;
        RECT 33.925 139.440 34.125 139.480 ;
        RECT 36.250 139.470 36.500 139.685 ;
        RECT 34.745 139.440 36.500 139.470 ;
        RECT 33.925 139.300 36.500 139.440 ;
        RECT 36.700 139.530 37.030 139.685 ;
        RECT 36.700 139.360 38.490 139.530 ;
        RECT 33.925 139.270 34.915 139.300 ;
        RECT 33.365 137.960 33.755 139.130 ;
        RECT 33.925 137.790 34.095 139.270 ;
        RECT 36.250 139.190 36.500 139.300 ;
        RECT 34.265 138.090 34.525 139.100 ;
        RECT 34.695 138.770 35.105 139.100 ;
        RECT 35.755 138.850 36.005 139.130 ;
        RECT 36.250 139.020 36.995 139.190 ;
        RECT 34.695 138.100 34.865 138.770 ;
        RECT 35.285 138.600 35.515 138.740 ;
        RECT 35.755 138.680 36.655 138.850 ;
        RECT 35.035 138.270 35.515 138.600 ;
        RECT 36.105 138.520 36.655 138.680 ;
        RECT 35.685 138.100 35.935 138.510 ;
        RECT 34.695 137.930 35.935 138.100 ;
        RECT 31.435 137.045 31.685 137.750 ;
        RECT 31.865 137.310 32.205 137.750 ;
        RECT 32.375 137.045 32.625 137.770 ;
        RECT 32.795 137.310 33.155 137.770 ;
        RECT 33.370 137.620 34.095 137.790 ;
        RECT 33.370 137.330 33.700 137.620 ;
        RECT 34.270 137.045 34.520 137.790 ;
        RECT 34.695 137.310 35.080 137.930 ;
        RECT 36.105 137.760 36.275 138.520 ;
        RECT 36.825 138.350 36.995 139.020 ;
        RECT 35.250 137.045 35.580 137.760 ;
        RECT 35.750 137.460 36.275 137.760 ;
        RECT 36.445 138.180 36.995 138.350 ;
        RECT 36.445 137.630 36.695 138.180 ;
        RECT 37.165 138.010 37.335 139.360 ;
        RECT 37.855 139.280 38.490 139.360 ;
        RECT 36.865 137.630 37.335 138.010 ;
        RECT 37.505 138.035 37.685 139.085 ;
        RECT 37.855 138.535 38.025 139.280 ;
        RECT 38.195 138.755 38.525 139.110 ;
        RECT 38.720 138.705 39.050 140.205 ;
        RECT 39.220 138.825 39.550 139.715 ;
        RECT 39.720 139.435 40.875 139.765 ;
        RECT 37.855 138.205 38.890 138.535 ;
        RECT 39.220 138.090 39.390 138.825 ;
        RECT 39.720 138.645 39.890 139.435 ;
        RECT 39.060 138.035 39.390 138.090 ;
        RECT 37.505 137.865 39.390 138.035 ;
        RECT 37.505 137.525 38.890 137.695 ;
        RECT 39.060 137.625 39.390 137.865 ;
        RECT 39.560 138.475 39.890 138.645 ;
        RECT 39.560 137.805 39.730 138.475 ;
        RECT 40.205 138.305 40.535 139.265 ;
        RECT 40.705 138.645 40.875 139.435 ;
        RECT 41.045 139.405 41.375 140.205 ;
        RECT 41.560 139.405 41.925 139.865 ;
        RECT 41.045 138.880 41.585 139.215 ;
        RECT 41.755 138.985 41.925 139.405 ;
        RECT 42.095 139.155 42.425 140.205 ;
        RECT 41.755 138.815 42.430 138.985 ;
        RECT 40.705 138.475 42.090 138.645 ;
        RECT 41.760 138.315 42.090 138.475 ;
        RECT 39.930 137.975 40.660 138.305 ;
        RECT 40.830 138.145 41.160 138.305 ;
        RECT 42.260 138.145 42.430 138.815 ;
        RECT 42.625 138.675 42.795 139.865 ;
        RECT 42.965 138.845 43.665 139.940 ;
        RECT 42.625 138.345 43.175 138.675 ;
        RECT 40.830 137.975 42.430 138.145 ;
        RECT 39.560 137.555 40.320 137.805 ;
        RECT 37.505 137.460 37.675 137.525 ;
        RECT 35.750 137.290 37.675 137.460 ;
        RECT 38.720 137.385 38.890 137.525 ;
        RECT 40.490 137.385 40.660 137.975 ;
        RECT 38.155 137.045 38.550 137.355 ;
        RECT 38.720 137.215 40.660 137.385 ;
        RECT 40.985 137.045 41.315 137.805 ;
        RECT 41.855 137.345 42.185 137.975 ;
        RECT 42.415 137.045 42.665 137.805 ;
        RECT 42.845 137.310 43.175 138.345 ;
        RECT 43.405 138.090 43.665 138.845 ;
        RECT 43.835 138.780 44.165 140.205 ;
        RECT 44.365 139.450 44.665 139.940 ;
        RECT 44.865 139.620 45.195 140.205 ;
        RECT 45.765 139.620 46.095 140.205 ;
        RECT 44.365 139.280 45.985 139.450 ;
        RECT 43.405 137.310 43.735 138.090 ;
        RECT 43.915 137.045 44.165 138.090 ;
        RECT 44.365 137.770 44.535 139.280 ;
        RECT 44.705 137.970 45.115 139.110 ;
        RECT 45.315 138.780 45.645 139.110 ;
        RECT 44.365 137.310 44.725 137.770 ;
        RECT 44.895 137.045 45.145 137.770 ;
        RECT 45.315 137.750 45.485 138.780 ;
        RECT 45.815 138.590 45.985 139.280 ;
        RECT 46.315 138.780 46.565 140.205 ;
        RECT 46.735 139.050 47.015 139.940 ;
        RECT 47.215 139.220 47.465 140.205 ;
        RECT 47.665 139.050 47.995 139.940 ;
        RECT 46.735 138.880 47.995 139.050 ;
        RECT 48.195 138.880 48.445 140.205 ;
        RECT 45.655 137.920 45.985 138.590 ;
        RECT 46.735 138.110 46.905 138.880 ;
        RECT 48.615 138.710 48.995 139.940 ;
        RECT 49.170 139.165 49.470 140.205 ;
        RECT 49.665 139.480 49.915 140.205 ;
        RECT 50.115 139.480 50.445 139.940 ;
        RECT 50.645 139.610 50.895 140.205 ;
        RECT 51.545 139.640 51.875 140.205 ;
        RECT 53.945 139.700 54.275 140.205 ;
        RECT 50.245 139.440 50.445 139.480 ;
        RECT 52.570 139.470 52.820 139.685 ;
        RECT 51.065 139.440 52.820 139.470 ;
        RECT 50.245 139.300 52.820 139.440 ;
        RECT 53.020 139.530 53.350 139.685 ;
        RECT 53.020 139.360 54.810 139.530 ;
        RECT 50.245 139.270 51.235 139.300 ;
        RECT 47.075 138.540 48.995 138.710 ;
        RECT 47.075 138.310 48.085 138.540 ;
        RECT 46.735 137.940 47.950 138.110 ;
        RECT 48.255 138.040 48.655 138.370 ;
        RECT 45.315 137.310 45.655 137.750 ;
        RECT 45.835 137.045 46.085 137.750 ;
        RECT 46.330 137.045 46.580 137.770 ;
        RECT 46.760 137.310 47.090 137.940 ;
        RECT 47.270 137.045 47.440 137.770 ;
        RECT 47.620 137.310 47.950 137.940 ;
        RECT 48.825 137.770 48.995 138.540 ;
        RECT 48.120 137.045 48.450 137.770 ;
        RECT 48.620 137.440 48.995 137.770 ;
        RECT 49.170 137.045 49.470 138.065 ;
        RECT 49.685 137.960 50.075 139.130 ;
        RECT 50.245 137.790 50.415 139.270 ;
        RECT 52.570 139.190 52.820 139.300 ;
        RECT 50.585 138.090 50.845 139.100 ;
        RECT 51.015 138.770 51.425 139.100 ;
        RECT 52.075 138.850 52.325 139.130 ;
        RECT 52.570 139.020 53.315 139.190 ;
        RECT 51.015 138.100 51.185 138.770 ;
        RECT 51.605 138.600 51.835 138.740 ;
        RECT 52.075 138.680 52.975 138.850 ;
        RECT 51.355 138.270 51.835 138.600 ;
        RECT 52.425 138.520 52.975 138.680 ;
        RECT 52.005 138.100 52.255 138.510 ;
        RECT 51.015 137.930 52.255 138.100 ;
        RECT 49.690 137.620 50.415 137.790 ;
        RECT 49.690 137.330 50.020 137.620 ;
        RECT 50.590 137.045 50.840 137.790 ;
        RECT 51.015 137.310 51.400 137.930 ;
        RECT 52.425 137.760 52.595 138.520 ;
        RECT 53.145 138.350 53.315 139.020 ;
        RECT 51.570 137.045 51.900 137.760 ;
        RECT 52.070 137.460 52.595 137.760 ;
        RECT 52.765 138.180 53.315 138.350 ;
        RECT 52.765 137.630 53.015 138.180 ;
        RECT 53.485 138.010 53.655 139.360 ;
        RECT 54.175 139.280 54.810 139.360 ;
        RECT 53.185 137.630 53.655 138.010 ;
        RECT 53.825 138.035 54.005 139.085 ;
        RECT 54.175 138.535 54.345 139.280 ;
        RECT 54.515 138.755 54.845 139.110 ;
        RECT 55.040 138.705 55.370 140.205 ;
        RECT 55.540 138.825 55.870 139.715 ;
        RECT 56.040 139.435 57.195 139.765 ;
        RECT 54.175 138.205 55.210 138.535 ;
        RECT 55.540 138.090 55.710 138.825 ;
        RECT 56.040 138.645 56.210 139.435 ;
        RECT 55.380 138.035 55.710 138.090 ;
        RECT 53.825 137.865 55.710 138.035 ;
        RECT 53.825 137.525 55.210 137.695 ;
        RECT 55.380 137.625 55.710 137.865 ;
        RECT 55.880 138.475 56.210 138.645 ;
        RECT 55.880 137.805 56.050 138.475 ;
        RECT 56.525 138.305 56.855 139.265 ;
        RECT 57.025 138.645 57.195 139.435 ;
        RECT 57.365 139.405 57.695 140.205 ;
        RECT 57.880 139.405 58.245 139.865 ;
        RECT 57.365 138.880 57.905 139.215 ;
        RECT 58.075 138.985 58.245 139.405 ;
        RECT 58.415 139.155 58.745 140.205 ;
        RECT 58.075 138.815 58.750 138.985 ;
        RECT 57.025 138.475 58.410 138.645 ;
        RECT 58.080 138.315 58.410 138.475 ;
        RECT 56.250 137.975 56.980 138.305 ;
        RECT 57.150 138.145 57.480 138.305 ;
        RECT 58.580 138.145 58.750 138.815 ;
        RECT 58.945 138.675 59.115 139.865 ;
        RECT 59.285 138.845 59.985 139.940 ;
        RECT 58.945 138.345 59.495 138.675 ;
        RECT 57.150 137.975 58.750 138.145 ;
        RECT 55.880 137.555 56.640 137.805 ;
        RECT 53.825 137.460 53.995 137.525 ;
        RECT 52.070 137.290 53.995 137.460 ;
        RECT 55.040 137.385 55.210 137.525 ;
        RECT 56.810 137.385 56.980 137.975 ;
        RECT 54.475 137.045 54.870 137.355 ;
        RECT 55.040 137.215 56.980 137.385 ;
        RECT 57.305 137.045 57.635 137.805 ;
        RECT 58.175 137.345 58.505 137.975 ;
        RECT 58.735 137.045 58.985 137.805 ;
        RECT 59.165 137.310 59.495 138.345 ;
        RECT 59.725 138.090 59.985 138.845 ;
        RECT 60.155 138.780 60.485 140.205 ;
        RECT 62.155 138.780 62.405 140.205 ;
        RECT 62.575 139.050 62.855 139.940 ;
        RECT 63.055 139.220 63.305 140.205 ;
        RECT 63.505 139.050 63.835 139.940 ;
        RECT 62.575 138.880 63.835 139.050 ;
        RECT 64.035 138.880 64.285 140.205 ;
        RECT 62.575 138.110 62.745 138.880 ;
        RECT 64.455 138.710 64.835 139.940 ;
        RECT 65.035 138.780 65.285 140.205 ;
        RECT 65.455 139.050 65.735 139.940 ;
        RECT 65.935 139.220 66.185 140.205 ;
        RECT 66.385 139.050 66.715 139.940 ;
        RECT 65.455 138.880 66.715 139.050 ;
        RECT 66.915 138.880 67.165 140.205 ;
        RECT 62.915 138.540 64.835 138.710 ;
        RECT 62.915 138.310 63.925 138.540 ;
        RECT 59.725 137.310 60.055 138.090 ;
        RECT 60.235 137.045 60.485 138.090 ;
        RECT 62.575 137.940 63.790 138.110 ;
        RECT 64.095 138.040 64.495 138.370 ;
        RECT 62.170 137.045 62.420 137.770 ;
        RECT 62.600 137.310 62.930 137.940 ;
        RECT 63.110 137.045 63.280 137.770 ;
        RECT 63.460 137.310 63.790 137.940 ;
        RECT 64.665 137.770 64.835 138.540 ;
        RECT 65.455 138.110 65.625 138.880 ;
        RECT 67.335 138.710 67.715 139.940 ;
        RECT 65.795 138.540 67.715 138.710 ;
        RECT 65.795 138.310 66.805 138.540 ;
        RECT 65.455 137.940 66.670 138.110 ;
        RECT 66.975 138.040 67.375 138.370 ;
        RECT 63.960 137.045 64.290 137.770 ;
        RECT 64.460 137.440 64.835 137.770 ;
        RECT 65.050 137.045 65.300 137.770 ;
        RECT 65.480 137.310 65.810 137.940 ;
        RECT 65.990 137.045 66.160 137.770 ;
        RECT 66.340 137.310 66.670 137.940 ;
        RECT 67.545 137.770 67.715 138.540 ;
        RECT 68.005 138.210 68.575 140.205 ;
        RECT 69.295 138.890 69.625 140.205 ;
        RECT 112.980 140.005 113.150 149.415 ;
        RECT 113.780 148.905 114.280 149.075 ;
        RECT 113.550 147.150 113.720 148.690 ;
        RECT 114.340 147.150 114.510 148.690 ;
        RECT 113.780 146.765 114.280 146.935 ;
        RECT 113.550 145.010 113.720 146.550 ;
        RECT 114.340 145.010 114.510 146.550 ;
        RECT 113.780 144.625 114.280 144.795 ;
        RECT 113.550 142.870 113.720 144.410 ;
        RECT 114.340 142.870 114.510 144.410 ;
        RECT 113.780 142.485 114.280 142.655 ;
        RECT 113.550 140.730 113.720 142.270 ;
        RECT 114.340 140.730 114.510 142.270 ;
        RECT 113.780 140.345 114.280 140.515 ;
        RECT 114.910 140.005 115.080 149.415 ;
        RECT 115.440 149.415 117.540 149.585 ;
        RECT 115.440 144.365 115.610 149.415 ;
        RECT 116.240 148.905 116.740 149.075 ;
        RECT 116.010 148.195 116.180 148.735 ;
        RECT 116.800 148.195 116.970 148.735 ;
        RECT 116.240 147.855 116.740 148.025 ;
        RECT 116.010 147.145 116.180 147.685 ;
        RECT 116.800 147.145 116.970 147.685 ;
        RECT 116.240 146.805 116.740 146.975 ;
        RECT 116.010 146.095 116.180 146.635 ;
        RECT 116.800 146.095 116.970 146.635 ;
        RECT 116.240 145.755 116.740 145.925 ;
        RECT 116.010 145.045 116.180 145.585 ;
        RECT 116.800 145.045 116.970 145.585 ;
        RECT 116.240 144.705 116.740 144.875 ;
        RECT 117.370 144.365 117.540 149.415 ;
        RECT 115.440 144.195 117.540 144.365 ;
        RECT 117.900 149.410 120.000 149.580 ;
        RECT 112.980 139.835 115.080 140.005 ;
        RECT 115.440 143.665 117.540 143.835 ;
        RECT 112.980 139.305 115.080 139.475 ;
        RECT 66.840 137.045 67.170 137.770 ;
        RECT 67.340 137.440 67.715 137.770 ;
        RECT 67.940 137.045 68.270 137.765 ;
        RECT 68.980 137.045 69.550 138.545 ;
        RECT 10.200 136.875 69.720 137.045 ;
        RECT 10.370 135.375 10.940 136.875 ;
        RECT 11.650 136.155 11.980 136.875 ;
        RECT 12.235 136.000 12.565 136.610 ;
        RECT 12.735 136.280 13.425 136.875 ;
        RECT 13.595 136.170 13.925 136.610 ;
        RECT 12.235 135.830 13.515 136.000 ;
        RECT 10.295 133.715 10.625 135.030 ;
        RECT 11.345 133.715 11.915 135.710 ;
        RECT 12.245 135.180 12.955 135.660 ;
        RECT 13.125 135.330 13.515 135.830 ;
        RECT 13.125 135.010 13.295 135.330 ;
        RECT 13.685 135.140 13.925 136.170 ;
        RECT 14.155 135.830 14.405 136.875 ;
        RECT 14.585 135.830 14.915 136.610 ;
        RECT 12.465 134.840 13.295 135.010 ;
        RECT 12.465 133.980 12.795 134.840 ;
        RECT 12.965 133.715 13.295 134.670 ;
        RECT 13.465 133.980 13.925 135.140 ;
        RECT 14.155 133.715 14.485 135.140 ;
        RECT 14.655 135.075 14.915 135.830 ;
        RECT 15.145 135.575 15.475 136.610 ;
        RECT 15.655 136.115 15.905 136.875 ;
        RECT 16.135 135.945 16.465 136.575 ;
        RECT 17.005 136.115 17.335 136.875 ;
        RECT 17.660 136.535 19.600 136.705 ;
        RECT 19.770 136.565 20.165 136.875 ;
        RECT 17.660 135.945 17.830 136.535 ;
        RECT 19.430 136.395 19.600 136.535 ;
        RECT 20.645 136.460 22.570 136.630 ;
        RECT 20.645 136.395 20.815 136.460 ;
        RECT 18.000 136.115 18.760 136.365 ;
        RECT 15.890 135.775 17.490 135.945 ;
        RECT 15.145 135.245 15.695 135.575 ;
        RECT 14.655 133.980 15.355 135.075 ;
        RECT 15.525 134.055 15.695 135.245 ;
        RECT 15.890 135.105 16.060 135.775 ;
        RECT 17.160 135.615 17.490 135.775 ;
        RECT 17.660 135.615 18.390 135.945 ;
        RECT 16.230 135.445 16.560 135.605 ;
        RECT 16.230 135.275 17.615 135.445 ;
        RECT 15.890 134.935 16.565 135.105 ;
        RECT 15.895 133.715 16.225 134.765 ;
        RECT 16.395 134.515 16.565 134.935 ;
        RECT 16.735 134.705 17.275 135.040 ;
        RECT 16.395 134.055 16.760 134.515 ;
        RECT 16.945 133.715 17.275 134.515 ;
        RECT 17.445 134.485 17.615 135.275 ;
        RECT 17.785 134.655 18.115 135.615 ;
        RECT 18.590 135.445 18.760 136.115 ;
        RECT 18.430 135.275 18.760 135.445 ;
        RECT 18.930 136.055 19.260 136.295 ;
        RECT 19.430 136.225 20.815 136.395 ;
        RECT 18.930 135.885 20.815 136.055 ;
        RECT 18.930 135.830 19.260 135.885 ;
        RECT 18.430 134.485 18.600 135.275 ;
        RECT 18.930 135.095 19.100 135.830 ;
        RECT 19.430 135.385 20.465 135.715 ;
        RECT 17.445 134.155 18.600 134.485 ;
        RECT 18.770 134.205 19.100 135.095 ;
        RECT 19.270 133.715 19.600 135.215 ;
        RECT 19.795 134.810 20.125 135.165 ;
        RECT 20.295 134.640 20.465 135.385 ;
        RECT 20.635 134.835 20.815 135.885 ;
        RECT 20.985 135.910 21.455 136.290 ;
        RECT 19.830 134.560 20.465 134.640 ;
        RECT 20.985 134.560 21.155 135.910 ;
        RECT 21.625 135.740 21.875 136.290 ;
        RECT 21.325 135.570 21.875 135.740 ;
        RECT 22.045 136.160 22.570 136.460 ;
        RECT 22.740 136.160 23.070 136.875 ;
        RECT 21.325 134.900 21.495 135.570 ;
        RECT 22.045 135.400 22.215 136.160 ;
        RECT 23.240 135.990 23.625 136.610 ;
        RECT 23.800 136.130 24.050 136.875 ;
        RECT 24.620 136.300 24.950 136.590 ;
        RECT 24.225 136.130 24.950 136.300 ;
        RECT 25.210 136.300 25.540 136.590 ;
        RECT 25.210 136.130 25.935 136.300 ;
        RECT 26.110 136.130 26.360 136.875 ;
        RECT 22.385 135.820 23.625 135.990 ;
        RECT 22.385 135.410 22.635 135.820 ;
        RECT 21.665 135.240 22.215 135.400 ;
        RECT 22.805 135.320 23.285 135.650 ;
        RECT 21.665 135.070 22.565 135.240 ;
        RECT 22.805 135.180 23.035 135.320 ;
        RECT 23.455 135.150 23.625 135.820 ;
        RECT 21.325 134.730 22.070 134.900 ;
        RECT 22.315 134.790 22.565 135.070 ;
        RECT 23.215 134.820 23.625 135.150 ;
        RECT 23.795 134.820 24.055 135.830 ;
        RECT 21.820 134.620 22.070 134.730 ;
        RECT 24.225 134.650 24.395 136.130 ;
        RECT 24.565 134.790 24.955 135.960 ;
        RECT 25.205 134.790 25.595 135.960 ;
        RECT 23.405 134.620 24.395 134.650 ;
        RECT 19.830 134.390 21.620 134.560 ;
        RECT 21.290 134.235 21.620 134.390 ;
        RECT 21.820 134.480 24.395 134.620 ;
        RECT 21.820 134.450 23.575 134.480 ;
        RECT 21.820 134.235 22.070 134.450 ;
        RECT 24.195 134.440 24.395 134.480 ;
        RECT 25.765 134.650 25.935 136.130 ;
        RECT 26.535 135.990 26.920 136.610 ;
        RECT 27.090 136.160 27.420 136.875 ;
        RECT 27.590 136.460 29.515 136.630 ;
        RECT 29.995 136.565 30.390 136.875 ;
        RECT 27.590 136.160 28.115 136.460 ;
        RECT 29.345 136.395 29.515 136.460 ;
        RECT 30.560 136.535 32.500 136.705 ;
        RECT 30.560 136.395 30.730 136.535 ;
        RECT 26.105 134.820 26.365 135.830 ;
        RECT 26.535 135.820 27.775 135.990 ;
        RECT 26.535 135.150 26.705 135.820 ;
        RECT 26.875 135.320 27.355 135.650 ;
        RECT 27.525 135.410 27.775 135.820 ;
        RECT 27.125 135.180 27.355 135.320 ;
        RECT 27.945 135.400 28.115 136.160 ;
        RECT 28.285 135.740 28.535 136.290 ;
        RECT 28.705 135.910 29.175 136.290 ;
        RECT 29.345 136.225 30.730 136.395 ;
        RECT 30.900 136.055 31.230 136.295 ;
        RECT 28.285 135.570 28.835 135.740 ;
        RECT 27.945 135.240 28.495 135.400 ;
        RECT 26.535 134.820 26.945 135.150 ;
        RECT 27.595 135.070 28.495 135.240 ;
        RECT 27.595 134.790 27.845 135.070 ;
        RECT 28.665 134.900 28.835 135.570 ;
        RECT 28.090 134.730 28.835 134.900 ;
        RECT 25.765 134.620 26.755 134.650 ;
        RECT 28.090 134.620 28.340 134.730 ;
        RECT 25.765 134.480 28.340 134.620 ;
        RECT 29.005 134.560 29.175 135.910 ;
        RECT 29.345 135.885 31.230 136.055 ;
        RECT 29.345 134.835 29.525 135.885 ;
        RECT 30.900 135.830 31.230 135.885 ;
        RECT 29.695 135.385 30.730 135.715 ;
        RECT 29.695 134.640 29.865 135.385 ;
        RECT 30.035 134.810 30.365 135.165 ;
        RECT 29.695 134.560 30.330 134.640 ;
        RECT 25.765 134.440 25.965 134.480 ;
        RECT 26.585 134.450 28.340 134.480 ;
        RECT 20.365 133.715 20.695 134.220 ;
        RECT 22.765 133.715 23.095 134.280 ;
        RECT 23.745 133.715 23.995 134.310 ;
        RECT 24.195 133.980 24.525 134.440 ;
        RECT 24.725 133.715 24.975 134.440 ;
        RECT 25.185 133.715 25.435 134.440 ;
        RECT 25.635 133.980 25.965 134.440 ;
        RECT 26.165 133.715 26.415 134.310 ;
        RECT 27.065 133.715 27.395 134.280 ;
        RECT 28.090 134.235 28.340 134.450 ;
        RECT 28.540 134.390 30.330 134.560 ;
        RECT 28.540 134.235 28.870 134.390 ;
        RECT 29.465 133.715 29.795 134.220 ;
        RECT 30.560 133.715 30.890 135.215 ;
        RECT 31.060 135.095 31.230 135.830 ;
        RECT 31.400 136.115 32.160 136.365 ;
        RECT 31.400 135.445 31.570 136.115 ;
        RECT 32.330 135.945 32.500 136.535 ;
        RECT 32.825 136.115 33.155 136.875 ;
        RECT 33.695 135.945 34.025 136.575 ;
        RECT 34.255 136.115 34.505 136.875 ;
        RECT 31.770 135.615 32.500 135.945 ;
        RECT 32.670 135.775 34.270 135.945 ;
        RECT 32.670 135.615 33.000 135.775 ;
        RECT 31.400 135.275 31.730 135.445 ;
        RECT 31.060 134.205 31.390 135.095 ;
        RECT 31.560 134.485 31.730 135.275 ;
        RECT 32.045 134.655 32.375 135.615 ;
        RECT 33.600 135.445 33.930 135.605 ;
        RECT 32.545 135.275 33.930 135.445 ;
        RECT 32.545 134.485 32.715 135.275 ;
        RECT 34.100 135.105 34.270 135.775 ;
        RECT 34.685 135.575 35.015 136.610 ;
        RECT 32.885 134.705 33.425 135.040 ;
        RECT 33.595 134.935 34.270 135.105 ;
        RECT 34.465 135.245 35.015 135.575 ;
        RECT 35.245 135.830 35.575 136.610 ;
        RECT 35.755 135.830 36.005 136.875 ;
        RECT 36.210 135.855 36.510 136.875 ;
        RECT 44.395 135.830 44.645 136.875 ;
        RECT 44.825 135.830 45.155 136.610 ;
        RECT 33.595 134.515 33.765 134.935 ;
        RECT 31.560 134.155 32.715 134.485 ;
        RECT 32.885 133.715 33.215 134.515 ;
        RECT 33.400 134.055 33.765 134.515 ;
        RECT 33.935 133.715 34.265 134.765 ;
        RECT 34.465 134.055 34.635 135.245 ;
        RECT 35.245 135.075 35.505 135.830 ;
        RECT 34.805 133.980 35.505 135.075 ;
        RECT 35.675 133.715 36.005 135.140 ;
        RECT 36.210 133.715 36.510 134.755 ;
        RECT 44.395 133.715 44.725 135.140 ;
        RECT 44.895 135.075 45.155 135.830 ;
        RECT 45.385 135.575 45.715 136.610 ;
        RECT 45.895 136.115 46.145 136.875 ;
        RECT 46.375 135.945 46.705 136.575 ;
        RECT 47.245 136.115 47.575 136.875 ;
        RECT 47.900 136.535 49.840 136.705 ;
        RECT 50.010 136.565 50.405 136.875 ;
        RECT 47.900 135.945 48.070 136.535 ;
        RECT 49.670 136.395 49.840 136.535 ;
        RECT 50.885 136.460 52.810 136.630 ;
        RECT 50.885 136.395 51.055 136.460 ;
        RECT 48.240 136.115 49.000 136.365 ;
        RECT 46.130 135.775 47.730 135.945 ;
        RECT 45.385 135.245 45.935 135.575 ;
        RECT 44.895 133.980 45.595 135.075 ;
        RECT 45.765 134.055 45.935 135.245 ;
        RECT 46.130 135.105 46.300 135.775 ;
        RECT 47.400 135.615 47.730 135.775 ;
        RECT 47.900 135.615 48.630 135.945 ;
        RECT 46.470 135.445 46.800 135.605 ;
        RECT 46.470 135.275 47.855 135.445 ;
        RECT 46.130 134.935 46.805 135.105 ;
        RECT 46.135 133.715 46.465 134.765 ;
        RECT 46.635 134.515 46.805 134.935 ;
        RECT 46.975 134.705 47.515 135.040 ;
        RECT 46.635 134.055 47.000 134.515 ;
        RECT 47.185 133.715 47.515 134.515 ;
        RECT 47.685 134.485 47.855 135.275 ;
        RECT 48.025 134.655 48.355 135.615 ;
        RECT 48.830 135.445 49.000 136.115 ;
        RECT 48.670 135.275 49.000 135.445 ;
        RECT 49.170 136.055 49.500 136.295 ;
        RECT 49.670 136.225 51.055 136.395 ;
        RECT 49.170 135.885 51.055 136.055 ;
        RECT 49.170 135.830 49.500 135.885 ;
        RECT 48.670 134.485 48.840 135.275 ;
        RECT 49.170 135.095 49.340 135.830 ;
        RECT 49.670 135.385 50.705 135.715 ;
        RECT 47.685 134.155 48.840 134.485 ;
        RECT 49.010 134.205 49.340 135.095 ;
        RECT 49.510 133.715 49.840 135.215 ;
        RECT 50.035 134.810 50.365 135.165 ;
        RECT 50.535 134.640 50.705 135.385 ;
        RECT 50.875 134.835 51.055 135.885 ;
        RECT 51.225 135.910 51.695 136.290 ;
        RECT 50.070 134.560 50.705 134.640 ;
        RECT 51.225 134.560 51.395 135.910 ;
        RECT 51.865 135.740 52.115 136.290 ;
        RECT 51.565 135.570 52.115 135.740 ;
        RECT 52.285 136.160 52.810 136.460 ;
        RECT 52.980 136.160 53.310 136.875 ;
        RECT 51.565 134.900 51.735 135.570 ;
        RECT 52.285 135.400 52.455 136.160 ;
        RECT 53.480 135.990 53.865 136.610 ;
        RECT 54.040 136.130 54.290 136.875 ;
        RECT 54.860 136.300 55.190 136.590 ;
        RECT 54.465 136.130 55.190 136.300 ;
        RECT 56.410 136.150 56.660 136.875 ;
        RECT 52.625 135.820 53.865 135.990 ;
        RECT 52.625 135.410 52.875 135.820 ;
        RECT 51.905 135.240 52.455 135.400 ;
        RECT 53.045 135.320 53.525 135.650 ;
        RECT 51.905 135.070 52.805 135.240 ;
        RECT 53.045 135.180 53.275 135.320 ;
        RECT 53.695 135.150 53.865 135.820 ;
        RECT 51.565 134.730 52.310 134.900 ;
        RECT 52.555 134.790 52.805 135.070 ;
        RECT 53.455 134.820 53.865 135.150 ;
        RECT 54.035 134.820 54.295 135.830 ;
        RECT 52.060 134.620 52.310 134.730 ;
        RECT 54.465 134.650 54.635 136.130 ;
        RECT 56.840 135.980 57.170 136.610 ;
        RECT 57.350 136.150 57.520 136.875 ;
        RECT 57.700 135.980 58.030 136.610 ;
        RECT 58.200 136.150 58.530 136.875 ;
        RECT 58.700 136.150 59.075 136.480 ;
        RECT 59.290 136.150 59.540 136.875 ;
        RECT 54.805 134.790 55.195 135.960 ;
        RECT 56.815 135.810 58.030 135.980 ;
        RECT 53.645 134.620 54.635 134.650 ;
        RECT 50.070 134.390 51.860 134.560 ;
        RECT 51.530 134.235 51.860 134.390 ;
        RECT 52.060 134.480 54.635 134.620 ;
        RECT 52.060 134.450 53.815 134.480 ;
        RECT 52.060 134.235 52.310 134.450 ;
        RECT 54.435 134.440 54.635 134.480 ;
        RECT 50.605 133.715 50.935 134.220 ;
        RECT 53.005 133.715 53.335 134.280 ;
        RECT 53.985 133.715 54.235 134.310 ;
        RECT 54.435 133.980 54.765 134.440 ;
        RECT 54.965 133.715 55.215 134.440 ;
        RECT 56.395 133.715 56.645 135.140 ;
        RECT 56.815 135.040 56.985 135.810 ;
        RECT 57.155 135.380 58.165 135.610 ;
        RECT 58.335 135.550 58.735 135.880 ;
        RECT 58.905 135.380 59.075 136.150 ;
        RECT 59.720 135.980 60.050 136.610 ;
        RECT 60.230 136.150 60.400 136.875 ;
        RECT 60.580 135.980 60.910 136.610 ;
        RECT 61.080 136.150 61.410 136.875 ;
        RECT 61.580 136.150 61.955 136.480 ;
        RECT 57.155 135.210 59.075 135.380 ;
        RECT 56.815 134.870 58.075 135.040 ;
        RECT 56.815 133.980 57.095 134.870 ;
        RECT 57.295 133.715 57.545 134.700 ;
        RECT 57.745 133.980 58.075 134.870 ;
        RECT 58.275 133.715 58.525 135.040 ;
        RECT 58.695 133.980 59.075 135.210 ;
        RECT 59.695 135.810 60.910 135.980 ;
        RECT 59.275 133.715 59.525 135.140 ;
        RECT 59.695 135.040 59.865 135.810 ;
        RECT 60.035 135.380 61.045 135.610 ;
        RECT 61.215 135.550 61.615 135.880 ;
        RECT 61.785 135.380 61.955 136.150 ;
        RECT 62.130 135.855 62.430 136.875 ;
        RECT 62.625 136.290 63.355 136.705 ;
        RECT 60.035 135.210 61.955 135.380 ;
        RECT 59.695 134.870 60.955 135.040 ;
        RECT 59.695 133.980 59.975 134.870 ;
        RECT 60.175 133.715 60.425 134.700 ;
        RECT 60.625 133.980 60.955 134.870 ;
        RECT 61.155 133.715 61.405 135.040 ;
        RECT 61.575 133.980 61.955 135.210 ;
        RECT 62.780 135.110 63.110 136.120 ;
        RECT 63.860 135.950 64.190 136.875 ;
        RECT 64.360 135.780 64.835 136.490 ;
        RECT 63.595 135.280 63.925 135.780 ;
        RECT 64.100 135.280 64.495 135.610 ;
        RECT 64.100 135.110 64.270 135.280 ;
        RECT 64.665 135.110 64.835 135.780 ;
        RECT 62.780 134.940 64.270 135.110 ;
        RECT 62.130 133.715 62.430 134.755 ;
        RECT 62.870 133.715 63.205 134.770 ;
        RECT 63.375 133.960 63.705 134.940 ;
        RECT 63.910 133.715 64.240 134.770 ;
        RECT 64.440 133.980 64.835 135.110 ;
        RECT 65.005 136.150 65.380 136.480 ;
        RECT 65.550 136.150 65.880 136.875 ;
        RECT 65.005 135.380 65.175 136.150 ;
        RECT 66.050 135.980 66.380 136.610 ;
        RECT 66.560 136.150 66.730 136.875 ;
        RECT 66.910 135.980 67.240 136.610 ;
        RECT 67.420 136.150 67.670 136.875 ;
        RECT 67.940 136.155 68.270 136.875 ;
        RECT 65.345 135.550 65.745 135.880 ;
        RECT 66.050 135.810 67.265 135.980 ;
        RECT 65.915 135.380 66.925 135.610 ;
        RECT 65.005 135.210 66.925 135.380 ;
        RECT 65.005 133.980 65.385 135.210 ;
        RECT 67.095 135.040 67.265 135.810 ;
        RECT 65.555 133.715 65.805 135.040 ;
        RECT 66.005 134.870 67.265 135.040 ;
        RECT 66.005 133.980 66.335 134.870 ;
        RECT 66.535 133.715 66.785 134.700 ;
        RECT 66.985 133.980 67.265 134.870 ;
        RECT 67.435 133.715 67.685 135.140 ;
        RECT 68.005 133.715 68.575 135.710 ;
        RECT 68.980 135.375 69.550 136.875 ;
        RECT 69.295 133.715 69.625 135.030 ;
        RECT 112.980 134.255 113.150 139.305 ;
        RECT 113.780 138.795 114.280 138.965 ;
        RECT 113.550 138.085 113.720 138.625 ;
        RECT 114.340 138.085 114.510 138.625 ;
        RECT 113.780 137.745 114.280 137.915 ;
        RECT 113.550 137.035 113.720 137.575 ;
        RECT 114.340 137.035 114.510 137.575 ;
        RECT 113.780 136.695 114.280 136.865 ;
        RECT 113.550 135.985 113.720 136.525 ;
        RECT 114.340 135.985 114.510 136.525 ;
        RECT 113.780 135.645 114.280 135.815 ;
        RECT 113.550 134.935 113.720 135.475 ;
        RECT 114.340 134.935 114.510 135.475 ;
        RECT 113.780 134.595 114.280 134.765 ;
        RECT 114.910 134.255 115.080 139.305 ;
        RECT 112.980 134.085 115.080 134.255 ;
        RECT 115.440 134.255 115.610 143.665 ;
        RECT 116.240 143.155 116.740 143.325 ;
        RECT 116.010 141.400 116.180 142.940 ;
        RECT 116.800 141.400 116.970 142.940 ;
        RECT 116.240 141.015 116.740 141.185 ;
        RECT 116.010 139.260 116.180 140.800 ;
        RECT 116.800 139.260 116.970 140.800 ;
        RECT 116.240 138.875 116.740 139.045 ;
        RECT 116.010 137.120 116.180 138.660 ;
        RECT 116.800 137.120 116.970 138.660 ;
        RECT 116.240 136.735 116.740 136.905 ;
        RECT 116.010 134.980 116.180 136.520 ;
        RECT 116.800 134.980 116.970 136.520 ;
        RECT 116.240 134.595 116.740 134.765 ;
        RECT 117.370 134.255 117.540 143.665 ;
        RECT 117.900 140.000 118.070 149.410 ;
        RECT 118.700 148.900 119.200 149.070 ;
        RECT 118.470 147.145 118.640 148.685 ;
        RECT 119.260 147.145 119.430 148.685 ;
        RECT 118.700 146.760 119.200 146.930 ;
        RECT 118.470 145.005 118.640 146.545 ;
        RECT 119.260 145.005 119.430 146.545 ;
        RECT 118.700 144.620 119.200 144.790 ;
        RECT 118.470 142.865 118.640 144.405 ;
        RECT 119.260 142.865 119.430 144.405 ;
        RECT 118.700 142.480 119.200 142.650 ;
        RECT 118.470 140.725 118.640 142.265 ;
        RECT 119.260 140.725 119.430 142.265 ;
        RECT 118.700 140.340 119.200 140.510 ;
        RECT 119.830 140.000 120.000 149.410 ;
        RECT 129.120 148.485 129.290 149.950 ;
        RECT 130.385 149.745 132.185 149.805 ;
        RECT 130.045 149.575 132.185 149.745 ;
        RECT 130.045 149.460 130.215 149.575 ;
        RECT 129.555 149.130 130.215 149.460 ;
        RECT 132.450 149.405 132.620 149.975 ;
        RECT 134.855 149.920 135.515 150.250 ;
        RECT 134.855 149.805 135.025 149.920 ;
        RECT 132.885 149.635 135.025 149.805 ;
        RECT 132.885 149.575 134.685 149.635 ;
        RECT 135.780 149.430 135.950 150.410 ;
        RECT 153.130 150.280 153.300 151.035 ;
        RECT 153.565 150.535 156.195 150.865 ;
        RECT 154.500 150.305 154.700 150.535 ;
        RECT 156.460 150.305 156.630 151.035 ;
        RECT 177.140 151.365 177.310 151.850 ;
        RECT 177.140 151.035 178.355 151.365 ;
        RECT 178.525 151.035 179.005 151.725 ;
        RECT 180.470 151.365 180.640 151.850 ;
        RECT 179.175 151.035 180.640 151.365 ;
        RECT 153.130 149.950 154.225 150.280 ;
        RECT 154.395 149.975 154.765 150.305 ;
        RECT 155.035 149.975 158.055 150.305 ;
        RECT 158.325 149.975 158.695 150.305 ;
        RECT 130.385 149.075 130.755 149.405 ;
        RECT 131.025 149.075 134.045 149.405 ;
        RECT 134.315 149.075 134.685 149.405 ;
        RECT 134.855 149.100 135.950 149.430 ;
        RECT 129.120 148.155 130.335 148.485 ;
        RECT 130.505 148.155 130.985 148.845 ;
        RECT 132.450 148.485 132.620 149.075 ;
        RECT 131.155 148.155 133.915 148.485 ;
        RECT 134.085 148.155 134.565 148.845 ;
        RECT 135.780 148.485 135.950 149.100 ;
        RECT 134.735 148.155 135.950 148.485 ;
        RECT 129.120 147.440 129.290 148.155 ;
        RECT 129.555 147.655 132.185 147.985 ;
        RECT 129.120 147.140 130.310 147.440 ;
        RECT 129.120 146.565 129.290 147.140 ;
        RECT 130.570 146.925 130.770 147.655 ;
        RECT 132.450 147.440 132.620 148.155 ;
        RECT 132.885 147.655 135.515 147.985 ;
        RECT 131.410 147.140 133.660 147.440 ;
        RECT 129.120 146.235 130.335 146.565 ;
        RECT 130.505 146.235 130.985 146.925 ;
        RECT 132.450 146.565 132.620 147.140 ;
        RECT 134.300 146.925 134.500 147.655 ;
        RECT 135.780 147.440 135.950 148.155 ;
        RECT 134.760 147.140 135.950 147.440 ;
        RECT 131.155 146.235 133.915 146.565 ;
        RECT 134.085 146.235 134.565 146.925 ;
        RECT 135.780 146.565 135.950 147.140 ;
        RECT 134.735 146.235 135.950 146.565 ;
        RECT 129.120 145.495 129.290 146.235 ;
        RECT 129.555 145.735 132.185 146.065 ;
        RECT 129.120 145.165 130.335 145.495 ;
        RECT 130.620 145.485 130.820 145.735 ;
        RECT 129.120 144.565 129.290 145.165 ;
        RECT 129.555 144.745 130.385 144.995 ;
        RECT 129.120 144.235 130.045 144.565 ;
        RECT 117.900 139.830 120.000 140.000 ;
        RECT 120.360 143.660 124.390 143.830 ;
        RECT 115.440 134.085 117.540 134.255 ;
        RECT 117.900 139.300 120.000 139.470 ;
        RECT 117.900 134.250 118.070 139.300 ;
        RECT 118.700 138.790 119.200 138.960 ;
        RECT 118.470 138.080 118.640 138.620 ;
        RECT 119.260 138.080 119.430 138.620 ;
        RECT 118.700 137.740 119.200 137.910 ;
        RECT 118.470 137.030 118.640 137.570 ;
        RECT 119.260 137.030 119.430 137.570 ;
        RECT 118.700 136.690 119.200 136.860 ;
        RECT 118.470 135.980 118.640 136.520 ;
        RECT 119.260 135.980 119.430 136.520 ;
        RECT 118.700 135.640 119.200 135.810 ;
        RECT 118.470 134.930 118.640 135.470 ;
        RECT 119.260 134.930 119.430 135.470 ;
        RECT 118.700 134.590 119.200 134.760 ;
        RECT 119.830 134.250 120.000 139.300 ;
        RECT 117.900 134.080 120.000 134.250 ;
        RECT 120.360 134.250 120.530 143.660 ;
        RECT 121.160 143.150 121.660 143.320 ;
        RECT 120.930 141.395 121.100 142.935 ;
        RECT 121.720 141.395 121.890 142.935 ;
        RECT 121.160 141.010 121.660 141.180 ;
        RECT 120.930 139.255 121.100 140.795 ;
        RECT 121.720 139.255 121.890 140.795 ;
        RECT 121.160 138.870 121.660 139.040 ;
        RECT 120.930 137.115 121.100 138.655 ;
        RECT 121.720 137.115 121.890 138.655 ;
        RECT 121.160 136.730 121.660 136.900 ;
        RECT 120.930 134.975 121.100 136.515 ;
        RECT 121.720 134.975 121.890 136.515 ;
        RECT 121.160 134.590 121.660 134.760 ;
        RECT 122.290 134.250 122.460 143.660 ;
        RECT 123.090 143.150 123.590 143.320 ;
        RECT 122.860 141.395 123.030 142.935 ;
        RECT 123.650 141.395 123.820 142.935 ;
        RECT 123.090 141.010 123.590 141.180 ;
        RECT 122.860 139.255 123.030 140.795 ;
        RECT 123.650 139.255 123.820 140.795 ;
        RECT 123.090 138.870 123.590 139.040 ;
        RECT 122.860 137.115 123.030 138.655 ;
        RECT 123.650 137.115 123.820 138.655 ;
        RECT 123.090 136.730 123.590 136.900 ;
        RECT 122.860 134.975 123.030 136.515 ;
        RECT 123.650 134.975 123.820 136.515 ;
        RECT 123.090 134.590 123.590 134.760 ;
        RECT 124.220 134.250 124.390 143.660 ;
        RECT 129.120 143.655 129.290 144.235 ;
        RECT 130.215 144.005 130.385 144.745 ;
        RECT 129.555 143.835 130.385 144.005 ;
        RECT 129.120 143.325 130.045 143.655 ;
        RECT 130.215 143.565 130.385 143.835 ;
        RECT 130.555 143.810 130.985 145.485 ;
        RECT 132.450 145.460 132.620 146.235 ;
        RECT 132.885 145.735 135.515 146.065 ;
        RECT 134.250 145.485 134.450 145.735 ;
        RECT 135.780 145.495 135.950 146.235 ;
        RECT 131.155 145.210 133.915 145.460 ;
        RECT 131.155 144.680 132.185 145.010 ;
        RECT 131.155 144.110 131.325 144.680 ;
        RECT 132.450 144.480 132.620 145.210 ;
        RECT 132.885 144.680 133.915 145.010 ;
        RECT 131.495 144.310 133.575 144.480 ;
        RECT 131.155 143.780 132.185 144.110 ;
        RECT 131.155 143.565 131.325 143.780 ;
        RECT 132.450 143.580 132.620 144.310 ;
        RECT 133.745 144.110 133.915 144.680 ;
        RECT 132.885 143.780 133.915 144.110 ;
        RECT 134.085 143.810 134.515 145.485 ;
        RECT 134.735 145.165 135.950 145.495 ;
        RECT 134.685 144.745 135.515 144.995 ;
        RECT 134.685 144.005 134.855 144.745 ;
        RECT 135.780 144.565 135.950 145.165 ;
        RECT 135.025 144.235 135.950 144.565 ;
        RECT 134.685 143.835 135.515 144.005 ;
        RECT 130.215 143.335 131.325 143.565 ;
        RECT 129.120 143.120 129.290 143.325 ;
        RECT 129.120 142.820 130.310 143.120 ;
        RECT 129.120 142.600 129.290 142.820 ;
        RECT 129.120 142.350 130.335 142.600 ;
        RECT 129.120 141.740 129.290 142.350 ;
        RECT 130.620 142.170 130.820 143.335 ;
        RECT 131.495 143.330 133.575 143.580 ;
        RECT 133.745 143.565 133.915 143.780 ;
        RECT 134.685 143.565 134.855 143.835 ;
        RECT 135.780 143.655 135.950 144.235 ;
        RECT 133.745 143.335 134.855 143.565 ;
        RECT 132.450 143.120 132.620 143.330 ;
        RECT 131.410 142.820 133.660 143.120 ;
        RECT 132.450 142.615 132.620 142.820 ;
        RECT 131.025 142.365 134.045 142.615 ;
        RECT 129.555 141.920 130.385 142.170 ;
        RECT 129.120 141.410 130.045 141.740 ;
        RECT 129.120 140.880 129.290 141.410 ;
        RECT 130.215 141.230 130.385 141.920 ;
        RECT 129.555 141.060 130.385 141.230 ;
        RECT 129.120 140.550 130.045 140.880 ;
        RECT 129.120 139.880 129.290 140.550 ;
        RECT 130.215 140.380 130.385 141.060 ;
        RECT 130.555 140.480 130.985 142.170 ;
        RECT 131.155 141.915 132.185 142.165 ;
        RECT 131.155 141.215 131.325 141.915 ;
        RECT 132.450 141.715 132.620 142.365 ;
        RECT 134.255 142.170 134.455 143.335 ;
        RECT 135.025 143.325 135.950 143.655 ;
        RECT 135.780 143.120 135.950 143.325 ;
        RECT 134.760 142.820 135.950 143.120 ;
        RECT 135.780 142.600 135.950 142.820 ;
        RECT 134.735 142.350 135.950 142.600 ;
        RECT 132.885 141.915 133.915 142.165 ;
        RECT 131.495 141.385 133.575 141.715 ;
        RECT 131.155 140.885 132.185 141.215 ;
        RECT 129.555 140.310 130.385 140.380 ;
        RECT 129.555 140.235 130.515 140.310 ;
        RECT 131.155 140.235 131.325 140.885 ;
        RECT 132.450 140.685 132.620 141.385 ;
        RECT 133.745 141.215 133.915 141.915 ;
        RECT 132.885 140.885 133.915 141.215 ;
        RECT 131.495 140.435 133.575 140.685 ;
        RECT 129.555 140.065 132.185 140.235 ;
        RECT 129.555 140.050 130.825 140.065 ;
        RECT 129.120 139.550 130.175 139.880 ;
        RECT 120.360 134.080 124.390 134.250 ;
        RECT 124.750 139.300 128.780 139.470 ;
        RECT 124.750 134.250 124.920 139.300 ;
        RECT 125.550 138.790 126.050 138.960 ;
        RECT 125.320 138.080 125.490 138.620 ;
        RECT 126.110 138.080 126.280 138.620 ;
        RECT 125.550 137.740 126.050 137.910 ;
        RECT 125.320 137.030 125.490 137.570 ;
        RECT 126.110 137.030 126.280 137.570 ;
        RECT 125.550 136.690 126.050 136.860 ;
        RECT 125.320 135.980 125.490 136.520 ;
        RECT 126.110 135.980 126.280 136.520 ;
        RECT 125.550 135.640 126.050 135.810 ;
        RECT 125.320 134.930 125.490 135.470 ;
        RECT 126.110 134.930 126.280 135.470 ;
        RECT 125.550 134.590 126.050 134.760 ;
        RECT 126.680 134.250 126.850 139.300 ;
        RECT 127.480 138.790 127.980 138.960 ;
        RECT 127.250 138.080 127.420 138.620 ;
        RECT 128.040 138.080 128.210 138.620 ;
        RECT 127.480 137.740 127.980 137.910 ;
        RECT 127.250 137.030 127.420 137.570 ;
        RECT 128.040 137.030 128.210 137.570 ;
        RECT 127.480 136.690 127.980 136.860 ;
        RECT 127.250 135.980 127.420 136.520 ;
        RECT 128.040 135.980 128.210 136.520 ;
        RECT 127.480 135.640 127.980 135.810 ;
        RECT 127.250 134.930 127.420 135.470 ;
        RECT 128.040 134.930 128.210 135.470 ;
        RECT 127.480 134.590 127.980 134.760 ;
        RECT 128.610 134.250 128.780 139.300 ;
        RECT 124.750 134.080 128.780 134.250 ;
        RECT 129.120 138.950 129.290 139.550 ;
        RECT 130.345 139.380 130.825 140.050 ;
        RECT 132.450 139.865 132.620 140.435 ;
        RECT 133.745 140.235 133.915 140.885 ;
        RECT 134.085 140.480 134.515 142.170 ;
        RECT 134.685 141.920 135.515 142.170 ;
        RECT 134.685 141.230 134.855 141.920 ;
        RECT 135.780 141.740 135.950 142.350 ;
        RECT 135.025 141.410 135.950 141.740 ;
        RECT 134.685 141.060 135.515 141.230 ;
        RECT 134.685 140.380 134.855 141.060 ;
        RECT 135.780 140.880 135.950 141.410 ;
        RECT 135.025 140.550 135.950 140.880 ;
        RECT 134.685 140.310 135.515 140.380 ;
        RECT 134.555 140.235 135.515 140.310 ;
        RECT 132.885 140.065 135.515 140.235 ;
        RECT 134.245 140.050 135.515 140.065 ;
        RECT 131.025 139.535 134.045 139.865 ;
        RECT 129.555 139.365 130.825 139.380 ;
        RECT 129.555 139.120 132.185 139.365 ;
        RECT 130.345 139.035 132.185 139.120 ;
        RECT 129.120 138.620 130.175 138.950 ;
        RECT 129.120 138.280 129.290 138.620 ;
        RECT 130.345 138.535 130.825 139.035 ;
        RECT 132.450 138.865 132.620 139.535 ;
        RECT 134.245 139.380 134.725 140.050 ;
        RECT 135.780 139.880 135.950 140.550 ;
        RECT 134.895 139.550 135.950 139.880 ;
        RECT 136.990 149.415 139.090 149.585 ;
        RECT 136.990 140.005 137.160 149.415 ;
        RECT 137.790 148.905 138.290 149.075 ;
        RECT 137.560 147.150 137.730 148.690 ;
        RECT 138.350 147.150 138.520 148.690 ;
        RECT 137.790 146.765 138.290 146.935 ;
        RECT 137.560 145.010 137.730 146.550 ;
        RECT 138.350 145.010 138.520 146.550 ;
        RECT 137.790 144.625 138.290 144.795 ;
        RECT 137.560 142.870 137.730 144.410 ;
        RECT 138.350 142.870 138.520 144.410 ;
        RECT 137.790 142.485 138.290 142.655 ;
        RECT 137.560 140.730 137.730 142.270 ;
        RECT 138.350 140.730 138.520 142.270 ;
        RECT 137.790 140.345 138.290 140.515 ;
        RECT 138.920 140.005 139.090 149.415 ;
        RECT 139.450 149.415 141.550 149.585 ;
        RECT 139.450 144.365 139.620 149.415 ;
        RECT 140.250 148.905 140.750 149.075 ;
        RECT 140.020 148.195 140.190 148.735 ;
        RECT 140.810 148.195 140.980 148.735 ;
        RECT 140.250 147.855 140.750 148.025 ;
        RECT 140.020 147.145 140.190 147.685 ;
        RECT 140.810 147.145 140.980 147.685 ;
        RECT 140.250 146.805 140.750 146.975 ;
        RECT 140.020 146.095 140.190 146.635 ;
        RECT 140.810 146.095 140.980 146.635 ;
        RECT 140.250 145.755 140.750 145.925 ;
        RECT 140.020 145.045 140.190 145.585 ;
        RECT 140.810 145.045 140.980 145.585 ;
        RECT 140.250 144.705 140.750 144.875 ;
        RECT 141.380 144.365 141.550 149.415 ;
        RECT 139.450 144.195 141.550 144.365 ;
        RECT 141.910 149.410 144.010 149.580 ;
        RECT 136.990 139.835 139.090 140.005 ;
        RECT 139.450 143.665 141.550 143.835 ;
        RECT 134.245 139.365 135.515 139.380 ;
        RECT 132.885 139.120 135.515 139.365 ;
        RECT 132.885 139.035 134.725 139.120 ;
        RECT 131.025 138.535 134.045 138.865 ;
        RECT 134.245 138.535 134.725 139.035 ;
        RECT 135.780 138.950 135.950 139.550 ;
        RECT 134.895 138.620 135.950 138.950 ;
        RECT 129.120 138.030 130.335 138.280 ;
        RECT 129.120 137.420 129.290 138.030 ;
        RECT 130.620 137.850 130.820 138.535 ;
        RECT 132.450 138.295 132.620 138.535 ;
        RECT 131.025 138.045 134.045 138.295 ;
        RECT 129.555 137.600 130.385 137.850 ;
        RECT 129.120 137.090 130.045 137.420 ;
        RECT 129.120 136.560 129.290 137.090 ;
        RECT 130.215 136.910 130.385 137.600 ;
        RECT 129.555 136.740 130.385 136.910 ;
        RECT 129.120 136.230 130.045 136.560 ;
        RECT 129.120 135.560 129.290 136.230 ;
        RECT 130.215 136.060 130.385 136.740 ;
        RECT 130.555 136.160 130.985 137.850 ;
        RECT 131.155 137.595 132.185 137.845 ;
        RECT 131.155 136.895 131.325 137.595 ;
        RECT 132.450 137.395 132.620 138.045 ;
        RECT 134.250 137.850 134.450 138.535 ;
        RECT 135.780 138.280 135.950 138.620 ;
        RECT 134.735 138.030 135.950 138.280 ;
        RECT 132.885 137.595 133.915 137.845 ;
        RECT 131.495 137.065 133.575 137.395 ;
        RECT 131.155 136.565 132.185 136.895 ;
        RECT 129.555 135.990 130.385 136.060 ;
        RECT 129.555 135.915 130.515 135.990 ;
        RECT 131.155 135.915 131.325 136.565 ;
        RECT 132.450 136.365 132.620 137.065 ;
        RECT 133.745 136.895 133.915 137.595 ;
        RECT 132.885 136.565 133.915 136.895 ;
        RECT 131.495 136.115 133.575 136.365 ;
        RECT 129.555 135.745 132.185 135.915 ;
        RECT 129.555 135.730 130.825 135.745 ;
        RECT 129.120 135.230 130.175 135.560 ;
        RECT 129.120 134.630 129.290 135.230 ;
        RECT 130.345 135.060 130.825 135.730 ;
        RECT 132.450 135.545 132.620 136.115 ;
        RECT 133.745 135.915 133.915 136.565 ;
        RECT 134.085 136.160 134.515 137.850 ;
        RECT 134.685 137.600 135.515 137.850 ;
        RECT 134.685 136.910 134.855 137.600 ;
        RECT 135.780 137.420 135.950 138.030 ;
        RECT 135.025 137.090 135.950 137.420 ;
        RECT 134.685 136.740 135.515 136.910 ;
        RECT 134.685 136.060 134.855 136.740 ;
        RECT 135.780 136.560 135.950 137.090 ;
        RECT 135.025 136.230 135.950 136.560 ;
        RECT 134.685 135.990 135.515 136.060 ;
        RECT 134.555 135.915 135.515 135.990 ;
        RECT 132.885 135.745 135.515 135.915 ;
        RECT 134.245 135.730 135.515 135.745 ;
        RECT 131.025 135.215 134.045 135.545 ;
        RECT 129.555 135.045 130.825 135.060 ;
        RECT 129.555 134.800 132.185 135.045 ;
        RECT 130.345 134.715 132.185 134.800 ;
        RECT 129.120 134.300 130.175 134.630 ;
        RECT 129.120 134.090 129.290 134.300 ;
        RECT 130.345 134.215 130.825 134.715 ;
        RECT 132.450 134.545 132.620 135.215 ;
        RECT 134.245 135.060 134.725 135.730 ;
        RECT 135.780 135.560 135.950 136.230 ;
        RECT 134.895 135.230 135.950 135.560 ;
        RECT 134.245 135.045 135.515 135.060 ;
        RECT 132.885 134.800 135.515 135.045 ;
        RECT 132.885 134.715 134.725 134.800 ;
        RECT 131.025 134.215 134.045 134.545 ;
        RECT 134.245 134.215 134.725 134.715 ;
        RECT 135.780 134.630 135.950 135.230 ;
        RECT 134.895 134.300 135.950 134.630 ;
        RECT 132.450 134.090 132.620 134.215 ;
        RECT 135.780 134.090 135.950 134.300 ;
        RECT 136.990 139.305 139.090 139.475 ;
        RECT 136.990 134.255 137.160 139.305 ;
        RECT 137.790 138.795 138.290 138.965 ;
        RECT 137.560 138.085 137.730 138.625 ;
        RECT 138.350 138.085 138.520 138.625 ;
        RECT 137.790 137.745 138.290 137.915 ;
        RECT 137.560 137.035 137.730 137.575 ;
        RECT 138.350 137.035 138.520 137.575 ;
        RECT 137.790 136.695 138.290 136.865 ;
        RECT 137.560 135.985 137.730 136.525 ;
        RECT 138.350 135.985 138.520 136.525 ;
        RECT 137.790 135.645 138.290 135.815 ;
        RECT 137.560 134.935 137.730 135.475 ;
        RECT 138.350 134.935 138.520 135.475 ;
        RECT 137.790 134.595 138.290 134.765 ;
        RECT 138.920 134.255 139.090 139.305 ;
        RECT 136.990 134.085 139.090 134.255 ;
        RECT 139.450 134.255 139.620 143.665 ;
        RECT 140.250 143.155 140.750 143.325 ;
        RECT 140.020 141.400 140.190 142.940 ;
        RECT 140.810 141.400 140.980 142.940 ;
        RECT 140.250 141.015 140.750 141.185 ;
        RECT 140.020 139.260 140.190 140.800 ;
        RECT 140.810 139.260 140.980 140.800 ;
        RECT 140.250 138.875 140.750 139.045 ;
        RECT 140.020 137.120 140.190 138.660 ;
        RECT 140.810 137.120 140.980 138.660 ;
        RECT 140.250 136.735 140.750 136.905 ;
        RECT 140.020 134.980 140.190 136.520 ;
        RECT 140.810 134.980 140.980 136.520 ;
        RECT 140.250 134.595 140.750 134.765 ;
        RECT 141.380 134.255 141.550 143.665 ;
        RECT 141.910 140.000 142.080 149.410 ;
        RECT 142.710 148.900 143.210 149.070 ;
        RECT 142.480 147.145 142.650 148.685 ;
        RECT 143.270 147.145 143.440 148.685 ;
        RECT 142.710 146.760 143.210 146.930 ;
        RECT 142.480 145.005 142.650 146.545 ;
        RECT 143.270 145.005 143.440 146.545 ;
        RECT 142.710 144.620 143.210 144.790 ;
        RECT 142.480 142.865 142.650 144.405 ;
        RECT 143.270 142.865 143.440 144.405 ;
        RECT 142.710 142.480 143.210 142.650 ;
        RECT 142.480 140.725 142.650 142.265 ;
        RECT 143.270 140.725 143.440 142.265 ;
        RECT 142.710 140.340 143.210 140.510 ;
        RECT 143.840 140.000 144.010 149.410 ;
        RECT 153.130 148.485 153.300 149.950 ;
        RECT 154.395 149.745 156.195 149.805 ;
        RECT 154.055 149.575 156.195 149.745 ;
        RECT 154.055 149.460 154.225 149.575 ;
        RECT 153.565 149.130 154.225 149.460 ;
        RECT 156.460 149.405 156.630 149.975 ;
        RECT 158.865 149.920 159.525 150.250 ;
        RECT 158.865 149.805 159.035 149.920 ;
        RECT 156.895 149.635 159.035 149.805 ;
        RECT 156.895 149.575 158.695 149.635 ;
        RECT 159.790 149.430 159.960 150.410 ;
        RECT 177.140 150.280 177.310 151.035 ;
        RECT 177.575 150.535 180.205 150.865 ;
        RECT 178.510 150.305 178.710 150.535 ;
        RECT 180.470 150.305 180.640 151.035 ;
        RECT 201.150 151.365 201.320 151.850 ;
        RECT 201.150 151.035 202.365 151.365 ;
        RECT 202.535 151.035 203.015 151.725 ;
        RECT 204.480 151.365 204.650 151.850 ;
        RECT 203.185 151.035 204.650 151.365 ;
        RECT 177.140 149.950 178.235 150.280 ;
        RECT 178.405 149.975 178.775 150.305 ;
        RECT 179.045 149.975 182.065 150.305 ;
        RECT 182.335 149.975 182.705 150.305 ;
        RECT 154.395 149.075 154.765 149.405 ;
        RECT 155.035 149.075 158.055 149.405 ;
        RECT 158.325 149.075 158.695 149.405 ;
        RECT 158.865 149.100 159.960 149.430 ;
        RECT 153.130 148.155 154.345 148.485 ;
        RECT 154.515 148.155 154.995 148.845 ;
        RECT 156.460 148.485 156.630 149.075 ;
        RECT 155.165 148.155 157.925 148.485 ;
        RECT 158.095 148.155 158.575 148.845 ;
        RECT 159.790 148.485 159.960 149.100 ;
        RECT 158.745 148.155 159.960 148.485 ;
        RECT 153.130 147.440 153.300 148.155 ;
        RECT 153.565 147.655 156.195 147.985 ;
        RECT 153.130 147.140 154.320 147.440 ;
        RECT 153.130 146.565 153.300 147.140 ;
        RECT 154.580 146.925 154.780 147.655 ;
        RECT 156.460 147.440 156.630 148.155 ;
        RECT 156.895 147.655 159.525 147.985 ;
        RECT 155.420 147.140 157.670 147.440 ;
        RECT 153.130 146.235 154.345 146.565 ;
        RECT 154.515 146.235 154.995 146.925 ;
        RECT 156.460 146.565 156.630 147.140 ;
        RECT 158.310 146.925 158.510 147.655 ;
        RECT 159.790 147.440 159.960 148.155 ;
        RECT 158.770 147.140 159.960 147.440 ;
        RECT 155.165 146.235 157.925 146.565 ;
        RECT 158.095 146.235 158.575 146.925 ;
        RECT 159.790 146.565 159.960 147.140 ;
        RECT 158.745 146.235 159.960 146.565 ;
        RECT 153.130 145.495 153.300 146.235 ;
        RECT 153.565 145.735 156.195 146.065 ;
        RECT 153.130 145.165 154.345 145.495 ;
        RECT 154.630 145.485 154.830 145.735 ;
        RECT 153.130 144.565 153.300 145.165 ;
        RECT 153.565 144.745 154.395 144.995 ;
        RECT 153.130 144.235 154.055 144.565 ;
        RECT 141.910 139.830 144.010 140.000 ;
        RECT 144.370 143.660 148.400 143.830 ;
        RECT 139.450 134.085 141.550 134.255 ;
        RECT 141.910 139.300 144.010 139.470 ;
        RECT 141.910 134.250 142.080 139.300 ;
        RECT 142.710 138.790 143.210 138.960 ;
        RECT 142.480 138.080 142.650 138.620 ;
        RECT 143.270 138.080 143.440 138.620 ;
        RECT 142.710 137.740 143.210 137.910 ;
        RECT 142.480 137.030 142.650 137.570 ;
        RECT 143.270 137.030 143.440 137.570 ;
        RECT 142.710 136.690 143.210 136.860 ;
        RECT 142.480 135.980 142.650 136.520 ;
        RECT 143.270 135.980 143.440 136.520 ;
        RECT 142.710 135.640 143.210 135.810 ;
        RECT 142.480 134.930 142.650 135.470 ;
        RECT 143.270 134.930 143.440 135.470 ;
        RECT 142.710 134.590 143.210 134.760 ;
        RECT 143.840 134.250 144.010 139.300 ;
        RECT 141.910 134.080 144.010 134.250 ;
        RECT 144.370 134.250 144.540 143.660 ;
        RECT 145.170 143.150 145.670 143.320 ;
        RECT 144.940 141.395 145.110 142.935 ;
        RECT 145.730 141.395 145.900 142.935 ;
        RECT 145.170 141.010 145.670 141.180 ;
        RECT 144.940 139.255 145.110 140.795 ;
        RECT 145.730 139.255 145.900 140.795 ;
        RECT 145.170 138.870 145.670 139.040 ;
        RECT 144.940 137.115 145.110 138.655 ;
        RECT 145.730 137.115 145.900 138.655 ;
        RECT 145.170 136.730 145.670 136.900 ;
        RECT 144.940 134.975 145.110 136.515 ;
        RECT 145.730 134.975 145.900 136.515 ;
        RECT 145.170 134.590 145.670 134.760 ;
        RECT 146.300 134.250 146.470 143.660 ;
        RECT 147.100 143.150 147.600 143.320 ;
        RECT 146.870 141.395 147.040 142.935 ;
        RECT 147.660 141.395 147.830 142.935 ;
        RECT 147.100 141.010 147.600 141.180 ;
        RECT 146.870 139.255 147.040 140.795 ;
        RECT 147.660 139.255 147.830 140.795 ;
        RECT 147.100 138.870 147.600 139.040 ;
        RECT 146.870 137.115 147.040 138.655 ;
        RECT 147.660 137.115 147.830 138.655 ;
        RECT 147.100 136.730 147.600 136.900 ;
        RECT 146.870 134.975 147.040 136.515 ;
        RECT 147.660 134.975 147.830 136.515 ;
        RECT 147.100 134.590 147.600 134.760 ;
        RECT 148.230 134.250 148.400 143.660 ;
        RECT 153.130 143.655 153.300 144.235 ;
        RECT 154.225 144.005 154.395 144.745 ;
        RECT 153.565 143.835 154.395 144.005 ;
        RECT 153.130 143.325 154.055 143.655 ;
        RECT 154.225 143.565 154.395 143.835 ;
        RECT 154.565 143.810 154.995 145.485 ;
        RECT 156.460 145.460 156.630 146.235 ;
        RECT 156.895 145.735 159.525 146.065 ;
        RECT 158.260 145.485 158.460 145.735 ;
        RECT 159.790 145.495 159.960 146.235 ;
        RECT 155.165 145.210 157.925 145.460 ;
        RECT 155.165 144.680 156.195 145.010 ;
        RECT 155.165 144.110 155.335 144.680 ;
        RECT 156.460 144.480 156.630 145.210 ;
        RECT 156.895 144.680 157.925 145.010 ;
        RECT 155.505 144.310 157.585 144.480 ;
        RECT 155.165 143.780 156.195 144.110 ;
        RECT 155.165 143.565 155.335 143.780 ;
        RECT 156.460 143.580 156.630 144.310 ;
        RECT 157.755 144.110 157.925 144.680 ;
        RECT 156.895 143.780 157.925 144.110 ;
        RECT 158.095 143.810 158.525 145.485 ;
        RECT 158.745 145.165 159.960 145.495 ;
        RECT 158.695 144.745 159.525 144.995 ;
        RECT 158.695 144.005 158.865 144.745 ;
        RECT 159.790 144.565 159.960 145.165 ;
        RECT 159.035 144.235 159.960 144.565 ;
        RECT 158.695 143.835 159.525 144.005 ;
        RECT 154.225 143.335 155.335 143.565 ;
        RECT 153.130 143.120 153.300 143.325 ;
        RECT 153.130 142.820 154.320 143.120 ;
        RECT 153.130 142.600 153.300 142.820 ;
        RECT 153.130 142.350 154.345 142.600 ;
        RECT 153.130 141.740 153.300 142.350 ;
        RECT 154.630 142.170 154.830 143.335 ;
        RECT 155.505 143.330 157.585 143.580 ;
        RECT 157.755 143.565 157.925 143.780 ;
        RECT 158.695 143.565 158.865 143.835 ;
        RECT 159.790 143.655 159.960 144.235 ;
        RECT 157.755 143.335 158.865 143.565 ;
        RECT 156.460 143.120 156.630 143.330 ;
        RECT 155.420 142.820 157.670 143.120 ;
        RECT 156.460 142.615 156.630 142.820 ;
        RECT 155.035 142.365 158.055 142.615 ;
        RECT 153.565 141.920 154.395 142.170 ;
        RECT 153.130 141.410 154.055 141.740 ;
        RECT 153.130 140.880 153.300 141.410 ;
        RECT 154.225 141.230 154.395 141.920 ;
        RECT 153.565 141.060 154.395 141.230 ;
        RECT 153.130 140.550 154.055 140.880 ;
        RECT 153.130 139.880 153.300 140.550 ;
        RECT 154.225 140.380 154.395 141.060 ;
        RECT 154.565 140.480 154.995 142.170 ;
        RECT 155.165 141.915 156.195 142.165 ;
        RECT 155.165 141.215 155.335 141.915 ;
        RECT 156.460 141.715 156.630 142.365 ;
        RECT 158.265 142.170 158.465 143.335 ;
        RECT 159.035 143.325 159.960 143.655 ;
        RECT 159.790 143.120 159.960 143.325 ;
        RECT 158.770 142.820 159.960 143.120 ;
        RECT 159.790 142.600 159.960 142.820 ;
        RECT 158.745 142.350 159.960 142.600 ;
        RECT 156.895 141.915 157.925 142.165 ;
        RECT 155.505 141.385 157.585 141.715 ;
        RECT 155.165 140.885 156.195 141.215 ;
        RECT 153.565 140.310 154.395 140.380 ;
        RECT 153.565 140.235 154.525 140.310 ;
        RECT 155.165 140.235 155.335 140.885 ;
        RECT 156.460 140.685 156.630 141.385 ;
        RECT 157.755 141.215 157.925 141.915 ;
        RECT 156.895 140.885 157.925 141.215 ;
        RECT 155.505 140.435 157.585 140.685 ;
        RECT 153.565 140.065 156.195 140.235 ;
        RECT 153.565 140.050 154.835 140.065 ;
        RECT 153.130 139.550 154.185 139.880 ;
        RECT 144.370 134.080 148.400 134.250 ;
        RECT 148.760 139.300 152.790 139.470 ;
        RECT 148.760 134.250 148.930 139.300 ;
        RECT 149.560 138.790 150.060 138.960 ;
        RECT 149.330 138.080 149.500 138.620 ;
        RECT 150.120 138.080 150.290 138.620 ;
        RECT 149.560 137.740 150.060 137.910 ;
        RECT 149.330 137.030 149.500 137.570 ;
        RECT 150.120 137.030 150.290 137.570 ;
        RECT 149.560 136.690 150.060 136.860 ;
        RECT 149.330 135.980 149.500 136.520 ;
        RECT 150.120 135.980 150.290 136.520 ;
        RECT 149.560 135.640 150.060 135.810 ;
        RECT 149.330 134.930 149.500 135.470 ;
        RECT 150.120 134.930 150.290 135.470 ;
        RECT 149.560 134.590 150.060 134.760 ;
        RECT 150.690 134.250 150.860 139.300 ;
        RECT 151.490 138.790 151.990 138.960 ;
        RECT 151.260 138.080 151.430 138.620 ;
        RECT 152.050 138.080 152.220 138.620 ;
        RECT 151.490 137.740 151.990 137.910 ;
        RECT 151.260 137.030 151.430 137.570 ;
        RECT 152.050 137.030 152.220 137.570 ;
        RECT 151.490 136.690 151.990 136.860 ;
        RECT 151.260 135.980 151.430 136.520 ;
        RECT 152.050 135.980 152.220 136.520 ;
        RECT 151.490 135.640 151.990 135.810 ;
        RECT 151.260 134.930 151.430 135.470 ;
        RECT 152.050 134.930 152.220 135.470 ;
        RECT 151.490 134.590 151.990 134.760 ;
        RECT 152.620 134.250 152.790 139.300 ;
        RECT 148.760 134.080 152.790 134.250 ;
        RECT 153.130 138.950 153.300 139.550 ;
        RECT 154.355 139.380 154.835 140.050 ;
        RECT 156.460 139.865 156.630 140.435 ;
        RECT 157.755 140.235 157.925 140.885 ;
        RECT 158.095 140.480 158.525 142.170 ;
        RECT 158.695 141.920 159.525 142.170 ;
        RECT 158.695 141.230 158.865 141.920 ;
        RECT 159.790 141.740 159.960 142.350 ;
        RECT 159.035 141.410 159.960 141.740 ;
        RECT 158.695 141.060 159.525 141.230 ;
        RECT 158.695 140.380 158.865 141.060 ;
        RECT 159.790 140.880 159.960 141.410 ;
        RECT 159.035 140.550 159.960 140.880 ;
        RECT 158.695 140.310 159.525 140.380 ;
        RECT 158.565 140.235 159.525 140.310 ;
        RECT 156.895 140.065 159.525 140.235 ;
        RECT 158.255 140.050 159.525 140.065 ;
        RECT 155.035 139.535 158.055 139.865 ;
        RECT 153.565 139.365 154.835 139.380 ;
        RECT 153.565 139.120 156.195 139.365 ;
        RECT 154.355 139.035 156.195 139.120 ;
        RECT 153.130 138.620 154.185 138.950 ;
        RECT 153.130 138.280 153.300 138.620 ;
        RECT 154.355 138.535 154.835 139.035 ;
        RECT 156.460 138.865 156.630 139.535 ;
        RECT 158.255 139.380 158.735 140.050 ;
        RECT 159.790 139.880 159.960 140.550 ;
        RECT 158.905 139.550 159.960 139.880 ;
        RECT 161.000 149.415 163.100 149.585 ;
        RECT 161.000 140.005 161.170 149.415 ;
        RECT 161.800 148.905 162.300 149.075 ;
        RECT 161.570 147.150 161.740 148.690 ;
        RECT 162.360 147.150 162.530 148.690 ;
        RECT 161.800 146.765 162.300 146.935 ;
        RECT 161.570 145.010 161.740 146.550 ;
        RECT 162.360 145.010 162.530 146.550 ;
        RECT 161.800 144.625 162.300 144.795 ;
        RECT 161.570 142.870 161.740 144.410 ;
        RECT 162.360 142.870 162.530 144.410 ;
        RECT 161.800 142.485 162.300 142.655 ;
        RECT 161.570 140.730 161.740 142.270 ;
        RECT 162.360 140.730 162.530 142.270 ;
        RECT 161.800 140.345 162.300 140.515 ;
        RECT 162.930 140.005 163.100 149.415 ;
        RECT 163.460 149.415 165.560 149.585 ;
        RECT 163.460 144.365 163.630 149.415 ;
        RECT 164.260 148.905 164.760 149.075 ;
        RECT 164.030 148.195 164.200 148.735 ;
        RECT 164.820 148.195 164.990 148.735 ;
        RECT 164.260 147.855 164.760 148.025 ;
        RECT 164.030 147.145 164.200 147.685 ;
        RECT 164.820 147.145 164.990 147.685 ;
        RECT 164.260 146.805 164.760 146.975 ;
        RECT 164.030 146.095 164.200 146.635 ;
        RECT 164.820 146.095 164.990 146.635 ;
        RECT 164.260 145.755 164.760 145.925 ;
        RECT 164.030 145.045 164.200 145.585 ;
        RECT 164.820 145.045 164.990 145.585 ;
        RECT 164.260 144.705 164.760 144.875 ;
        RECT 165.390 144.365 165.560 149.415 ;
        RECT 163.460 144.195 165.560 144.365 ;
        RECT 165.920 149.410 168.020 149.580 ;
        RECT 161.000 139.835 163.100 140.005 ;
        RECT 163.460 143.665 165.560 143.835 ;
        RECT 158.255 139.365 159.525 139.380 ;
        RECT 156.895 139.120 159.525 139.365 ;
        RECT 156.895 139.035 158.735 139.120 ;
        RECT 155.035 138.535 158.055 138.865 ;
        RECT 158.255 138.535 158.735 139.035 ;
        RECT 159.790 138.950 159.960 139.550 ;
        RECT 158.905 138.620 159.960 138.950 ;
        RECT 153.130 138.030 154.345 138.280 ;
        RECT 153.130 137.420 153.300 138.030 ;
        RECT 154.630 137.850 154.830 138.535 ;
        RECT 156.460 138.295 156.630 138.535 ;
        RECT 155.035 138.045 158.055 138.295 ;
        RECT 153.565 137.600 154.395 137.850 ;
        RECT 153.130 137.090 154.055 137.420 ;
        RECT 153.130 136.560 153.300 137.090 ;
        RECT 154.225 136.910 154.395 137.600 ;
        RECT 153.565 136.740 154.395 136.910 ;
        RECT 153.130 136.230 154.055 136.560 ;
        RECT 153.130 135.560 153.300 136.230 ;
        RECT 154.225 136.060 154.395 136.740 ;
        RECT 154.565 136.160 154.995 137.850 ;
        RECT 155.165 137.595 156.195 137.845 ;
        RECT 155.165 136.895 155.335 137.595 ;
        RECT 156.460 137.395 156.630 138.045 ;
        RECT 158.260 137.850 158.460 138.535 ;
        RECT 159.790 138.280 159.960 138.620 ;
        RECT 158.745 138.030 159.960 138.280 ;
        RECT 156.895 137.595 157.925 137.845 ;
        RECT 155.505 137.065 157.585 137.395 ;
        RECT 155.165 136.565 156.195 136.895 ;
        RECT 153.565 135.990 154.395 136.060 ;
        RECT 153.565 135.915 154.525 135.990 ;
        RECT 155.165 135.915 155.335 136.565 ;
        RECT 156.460 136.365 156.630 137.065 ;
        RECT 157.755 136.895 157.925 137.595 ;
        RECT 156.895 136.565 157.925 136.895 ;
        RECT 155.505 136.115 157.585 136.365 ;
        RECT 153.565 135.745 156.195 135.915 ;
        RECT 153.565 135.730 154.835 135.745 ;
        RECT 153.130 135.230 154.185 135.560 ;
        RECT 153.130 134.630 153.300 135.230 ;
        RECT 154.355 135.060 154.835 135.730 ;
        RECT 156.460 135.545 156.630 136.115 ;
        RECT 157.755 135.915 157.925 136.565 ;
        RECT 158.095 136.160 158.525 137.850 ;
        RECT 158.695 137.600 159.525 137.850 ;
        RECT 158.695 136.910 158.865 137.600 ;
        RECT 159.790 137.420 159.960 138.030 ;
        RECT 159.035 137.090 159.960 137.420 ;
        RECT 158.695 136.740 159.525 136.910 ;
        RECT 158.695 136.060 158.865 136.740 ;
        RECT 159.790 136.560 159.960 137.090 ;
        RECT 159.035 136.230 159.960 136.560 ;
        RECT 158.695 135.990 159.525 136.060 ;
        RECT 158.565 135.915 159.525 135.990 ;
        RECT 156.895 135.745 159.525 135.915 ;
        RECT 158.255 135.730 159.525 135.745 ;
        RECT 155.035 135.215 158.055 135.545 ;
        RECT 153.565 135.045 154.835 135.060 ;
        RECT 153.565 134.800 156.195 135.045 ;
        RECT 154.355 134.715 156.195 134.800 ;
        RECT 153.130 134.300 154.185 134.630 ;
        RECT 153.130 134.090 153.300 134.300 ;
        RECT 154.355 134.215 154.835 134.715 ;
        RECT 156.460 134.545 156.630 135.215 ;
        RECT 158.255 135.060 158.735 135.730 ;
        RECT 159.790 135.560 159.960 136.230 ;
        RECT 158.905 135.230 159.960 135.560 ;
        RECT 158.255 135.045 159.525 135.060 ;
        RECT 156.895 134.800 159.525 135.045 ;
        RECT 156.895 134.715 158.735 134.800 ;
        RECT 155.035 134.215 158.055 134.545 ;
        RECT 158.255 134.215 158.735 134.715 ;
        RECT 159.790 134.630 159.960 135.230 ;
        RECT 158.905 134.300 159.960 134.630 ;
        RECT 156.460 134.090 156.630 134.215 ;
        RECT 159.790 134.090 159.960 134.300 ;
        RECT 161.000 139.305 163.100 139.475 ;
        RECT 161.000 134.255 161.170 139.305 ;
        RECT 161.800 138.795 162.300 138.965 ;
        RECT 161.570 138.085 161.740 138.625 ;
        RECT 162.360 138.085 162.530 138.625 ;
        RECT 161.800 137.745 162.300 137.915 ;
        RECT 161.570 137.035 161.740 137.575 ;
        RECT 162.360 137.035 162.530 137.575 ;
        RECT 161.800 136.695 162.300 136.865 ;
        RECT 161.570 135.985 161.740 136.525 ;
        RECT 162.360 135.985 162.530 136.525 ;
        RECT 161.800 135.645 162.300 135.815 ;
        RECT 161.570 134.935 161.740 135.475 ;
        RECT 162.360 134.935 162.530 135.475 ;
        RECT 161.800 134.595 162.300 134.765 ;
        RECT 162.930 134.255 163.100 139.305 ;
        RECT 161.000 134.085 163.100 134.255 ;
        RECT 163.460 134.255 163.630 143.665 ;
        RECT 164.260 143.155 164.760 143.325 ;
        RECT 164.030 141.400 164.200 142.940 ;
        RECT 164.820 141.400 164.990 142.940 ;
        RECT 164.260 141.015 164.760 141.185 ;
        RECT 164.030 139.260 164.200 140.800 ;
        RECT 164.820 139.260 164.990 140.800 ;
        RECT 164.260 138.875 164.760 139.045 ;
        RECT 164.030 137.120 164.200 138.660 ;
        RECT 164.820 137.120 164.990 138.660 ;
        RECT 164.260 136.735 164.760 136.905 ;
        RECT 164.030 134.980 164.200 136.520 ;
        RECT 164.820 134.980 164.990 136.520 ;
        RECT 164.260 134.595 164.760 134.765 ;
        RECT 165.390 134.255 165.560 143.665 ;
        RECT 165.920 140.000 166.090 149.410 ;
        RECT 166.720 148.900 167.220 149.070 ;
        RECT 166.490 147.145 166.660 148.685 ;
        RECT 167.280 147.145 167.450 148.685 ;
        RECT 166.720 146.760 167.220 146.930 ;
        RECT 166.490 145.005 166.660 146.545 ;
        RECT 167.280 145.005 167.450 146.545 ;
        RECT 166.720 144.620 167.220 144.790 ;
        RECT 166.490 142.865 166.660 144.405 ;
        RECT 167.280 142.865 167.450 144.405 ;
        RECT 166.720 142.480 167.220 142.650 ;
        RECT 166.490 140.725 166.660 142.265 ;
        RECT 167.280 140.725 167.450 142.265 ;
        RECT 166.720 140.340 167.220 140.510 ;
        RECT 167.850 140.000 168.020 149.410 ;
        RECT 177.140 148.485 177.310 149.950 ;
        RECT 178.405 149.745 180.205 149.805 ;
        RECT 178.065 149.575 180.205 149.745 ;
        RECT 178.065 149.460 178.235 149.575 ;
        RECT 177.575 149.130 178.235 149.460 ;
        RECT 180.470 149.405 180.640 149.975 ;
        RECT 182.875 149.920 183.535 150.250 ;
        RECT 182.875 149.805 183.045 149.920 ;
        RECT 180.905 149.635 183.045 149.805 ;
        RECT 180.905 149.575 182.705 149.635 ;
        RECT 183.800 149.430 183.970 150.410 ;
        RECT 201.150 150.280 201.320 151.035 ;
        RECT 201.585 150.535 204.215 150.865 ;
        RECT 202.520 150.305 202.720 150.535 ;
        RECT 204.480 150.305 204.650 151.035 ;
        RECT 225.160 151.365 225.330 151.850 ;
        RECT 225.160 151.035 226.375 151.365 ;
        RECT 226.545 151.035 227.025 151.725 ;
        RECT 228.490 151.365 228.660 151.850 ;
        RECT 227.195 151.035 228.660 151.365 ;
        RECT 201.150 149.950 202.245 150.280 ;
        RECT 202.415 149.975 202.785 150.305 ;
        RECT 203.055 149.975 206.075 150.305 ;
        RECT 206.345 149.975 206.715 150.305 ;
        RECT 178.405 149.075 178.775 149.405 ;
        RECT 179.045 149.075 182.065 149.405 ;
        RECT 182.335 149.075 182.705 149.405 ;
        RECT 182.875 149.100 183.970 149.430 ;
        RECT 177.140 148.155 178.355 148.485 ;
        RECT 178.525 148.155 179.005 148.845 ;
        RECT 180.470 148.485 180.640 149.075 ;
        RECT 179.175 148.155 181.935 148.485 ;
        RECT 182.105 148.155 182.585 148.845 ;
        RECT 183.800 148.485 183.970 149.100 ;
        RECT 182.755 148.155 183.970 148.485 ;
        RECT 177.140 147.440 177.310 148.155 ;
        RECT 177.575 147.655 180.205 147.985 ;
        RECT 177.140 147.140 178.330 147.440 ;
        RECT 177.140 146.565 177.310 147.140 ;
        RECT 178.590 146.925 178.790 147.655 ;
        RECT 180.470 147.440 180.640 148.155 ;
        RECT 180.905 147.655 183.535 147.985 ;
        RECT 179.430 147.140 181.680 147.440 ;
        RECT 177.140 146.235 178.355 146.565 ;
        RECT 178.525 146.235 179.005 146.925 ;
        RECT 180.470 146.565 180.640 147.140 ;
        RECT 182.320 146.925 182.520 147.655 ;
        RECT 183.800 147.440 183.970 148.155 ;
        RECT 182.780 147.140 183.970 147.440 ;
        RECT 179.175 146.235 181.935 146.565 ;
        RECT 182.105 146.235 182.585 146.925 ;
        RECT 183.800 146.565 183.970 147.140 ;
        RECT 182.755 146.235 183.970 146.565 ;
        RECT 177.140 145.495 177.310 146.235 ;
        RECT 177.575 145.735 180.205 146.065 ;
        RECT 177.140 145.165 178.355 145.495 ;
        RECT 178.640 145.485 178.840 145.735 ;
        RECT 177.140 144.565 177.310 145.165 ;
        RECT 177.575 144.745 178.405 144.995 ;
        RECT 177.140 144.235 178.065 144.565 ;
        RECT 165.920 139.830 168.020 140.000 ;
        RECT 168.380 143.660 172.410 143.830 ;
        RECT 163.460 134.085 165.560 134.255 ;
        RECT 165.920 139.300 168.020 139.470 ;
        RECT 165.920 134.250 166.090 139.300 ;
        RECT 166.720 138.790 167.220 138.960 ;
        RECT 166.490 138.080 166.660 138.620 ;
        RECT 167.280 138.080 167.450 138.620 ;
        RECT 166.720 137.740 167.220 137.910 ;
        RECT 166.490 137.030 166.660 137.570 ;
        RECT 167.280 137.030 167.450 137.570 ;
        RECT 166.720 136.690 167.220 136.860 ;
        RECT 166.490 135.980 166.660 136.520 ;
        RECT 167.280 135.980 167.450 136.520 ;
        RECT 166.720 135.640 167.220 135.810 ;
        RECT 166.490 134.930 166.660 135.470 ;
        RECT 167.280 134.930 167.450 135.470 ;
        RECT 166.720 134.590 167.220 134.760 ;
        RECT 167.850 134.250 168.020 139.300 ;
        RECT 165.920 134.080 168.020 134.250 ;
        RECT 168.380 134.250 168.550 143.660 ;
        RECT 169.180 143.150 169.680 143.320 ;
        RECT 168.950 141.395 169.120 142.935 ;
        RECT 169.740 141.395 169.910 142.935 ;
        RECT 169.180 141.010 169.680 141.180 ;
        RECT 168.950 139.255 169.120 140.795 ;
        RECT 169.740 139.255 169.910 140.795 ;
        RECT 169.180 138.870 169.680 139.040 ;
        RECT 168.950 137.115 169.120 138.655 ;
        RECT 169.740 137.115 169.910 138.655 ;
        RECT 169.180 136.730 169.680 136.900 ;
        RECT 168.950 134.975 169.120 136.515 ;
        RECT 169.740 134.975 169.910 136.515 ;
        RECT 169.180 134.590 169.680 134.760 ;
        RECT 170.310 134.250 170.480 143.660 ;
        RECT 171.110 143.150 171.610 143.320 ;
        RECT 170.880 141.395 171.050 142.935 ;
        RECT 171.670 141.395 171.840 142.935 ;
        RECT 171.110 141.010 171.610 141.180 ;
        RECT 170.880 139.255 171.050 140.795 ;
        RECT 171.670 139.255 171.840 140.795 ;
        RECT 171.110 138.870 171.610 139.040 ;
        RECT 170.880 137.115 171.050 138.655 ;
        RECT 171.670 137.115 171.840 138.655 ;
        RECT 171.110 136.730 171.610 136.900 ;
        RECT 170.880 134.975 171.050 136.515 ;
        RECT 171.670 134.975 171.840 136.515 ;
        RECT 171.110 134.590 171.610 134.760 ;
        RECT 172.240 134.250 172.410 143.660 ;
        RECT 177.140 143.655 177.310 144.235 ;
        RECT 178.235 144.005 178.405 144.745 ;
        RECT 177.575 143.835 178.405 144.005 ;
        RECT 177.140 143.325 178.065 143.655 ;
        RECT 178.235 143.565 178.405 143.835 ;
        RECT 178.575 143.810 179.005 145.485 ;
        RECT 180.470 145.460 180.640 146.235 ;
        RECT 180.905 145.735 183.535 146.065 ;
        RECT 182.270 145.485 182.470 145.735 ;
        RECT 183.800 145.495 183.970 146.235 ;
        RECT 179.175 145.210 181.935 145.460 ;
        RECT 179.175 144.680 180.205 145.010 ;
        RECT 179.175 144.110 179.345 144.680 ;
        RECT 180.470 144.480 180.640 145.210 ;
        RECT 180.905 144.680 181.935 145.010 ;
        RECT 179.515 144.310 181.595 144.480 ;
        RECT 179.175 143.780 180.205 144.110 ;
        RECT 179.175 143.565 179.345 143.780 ;
        RECT 180.470 143.580 180.640 144.310 ;
        RECT 181.765 144.110 181.935 144.680 ;
        RECT 180.905 143.780 181.935 144.110 ;
        RECT 182.105 143.810 182.535 145.485 ;
        RECT 182.755 145.165 183.970 145.495 ;
        RECT 182.705 144.745 183.535 144.995 ;
        RECT 182.705 144.005 182.875 144.745 ;
        RECT 183.800 144.565 183.970 145.165 ;
        RECT 183.045 144.235 183.970 144.565 ;
        RECT 182.705 143.835 183.535 144.005 ;
        RECT 178.235 143.335 179.345 143.565 ;
        RECT 177.140 143.120 177.310 143.325 ;
        RECT 177.140 142.820 178.330 143.120 ;
        RECT 177.140 142.600 177.310 142.820 ;
        RECT 177.140 142.350 178.355 142.600 ;
        RECT 177.140 141.740 177.310 142.350 ;
        RECT 178.640 142.170 178.840 143.335 ;
        RECT 179.515 143.330 181.595 143.580 ;
        RECT 181.765 143.565 181.935 143.780 ;
        RECT 182.705 143.565 182.875 143.835 ;
        RECT 183.800 143.655 183.970 144.235 ;
        RECT 181.765 143.335 182.875 143.565 ;
        RECT 180.470 143.120 180.640 143.330 ;
        RECT 179.430 142.820 181.680 143.120 ;
        RECT 180.470 142.615 180.640 142.820 ;
        RECT 179.045 142.365 182.065 142.615 ;
        RECT 177.575 141.920 178.405 142.170 ;
        RECT 177.140 141.410 178.065 141.740 ;
        RECT 177.140 140.880 177.310 141.410 ;
        RECT 178.235 141.230 178.405 141.920 ;
        RECT 177.575 141.060 178.405 141.230 ;
        RECT 177.140 140.550 178.065 140.880 ;
        RECT 177.140 139.880 177.310 140.550 ;
        RECT 178.235 140.380 178.405 141.060 ;
        RECT 178.575 140.480 179.005 142.170 ;
        RECT 179.175 141.915 180.205 142.165 ;
        RECT 179.175 141.215 179.345 141.915 ;
        RECT 180.470 141.715 180.640 142.365 ;
        RECT 182.275 142.170 182.475 143.335 ;
        RECT 183.045 143.325 183.970 143.655 ;
        RECT 183.800 143.120 183.970 143.325 ;
        RECT 182.780 142.820 183.970 143.120 ;
        RECT 183.800 142.600 183.970 142.820 ;
        RECT 182.755 142.350 183.970 142.600 ;
        RECT 180.905 141.915 181.935 142.165 ;
        RECT 179.515 141.385 181.595 141.715 ;
        RECT 179.175 140.885 180.205 141.215 ;
        RECT 177.575 140.310 178.405 140.380 ;
        RECT 177.575 140.235 178.535 140.310 ;
        RECT 179.175 140.235 179.345 140.885 ;
        RECT 180.470 140.685 180.640 141.385 ;
        RECT 181.765 141.215 181.935 141.915 ;
        RECT 180.905 140.885 181.935 141.215 ;
        RECT 179.515 140.435 181.595 140.685 ;
        RECT 177.575 140.065 180.205 140.235 ;
        RECT 177.575 140.050 178.845 140.065 ;
        RECT 177.140 139.550 178.195 139.880 ;
        RECT 168.380 134.080 172.410 134.250 ;
        RECT 172.770 139.300 176.800 139.470 ;
        RECT 172.770 134.250 172.940 139.300 ;
        RECT 173.570 138.790 174.070 138.960 ;
        RECT 173.340 138.080 173.510 138.620 ;
        RECT 174.130 138.080 174.300 138.620 ;
        RECT 173.570 137.740 174.070 137.910 ;
        RECT 173.340 137.030 173.510 137.570 ;
        RECT 174.130 137.030 174.300 137.570 ;
        RECT 173.570 136.690 174.070 136.860 ;
        RECT 173.340 135.980 173.510 136.520 ;
        RECT 174.130 135.980 174.300 136.520 ;
        RECT 173.570 135.640 174.070 135.810 ;
        RECT 173.340 134.930 173.510 135.470 ;
        RECT 174.130 134.930 174.300 135.470 ;
        RECT 173.570 134.590 174.070 134.760 ;
        RECT 174.700 134.250 174.870 139.300 ;
        RECT 175.500 138.790 176.000 138.960 ;
        RECT 175.270 138.080 175.440 138.620 ;
        RECT 176.060 138.080 176.230 138.620 ;
        RECT 175.500 137.740 176.000 137.910 ;
        RECT 175.270 137.030 175.440 137.570 ;
        RECT 176.060 137.030 176.230 137.570 ;
        RECT 175.500 136.690 176.000 136.860 ;
        RECT 175.270 135.980 175.440 136.520 ;
        RECT 176.060 135.980 176.230 136.520 ;
        RECT 175.500 135.640 176.000 135.810 ;
        RECT 175.270 134.930 175.440 135.470 ;
        RECT 176.060 134.930 176.230 135.470 ;
        RECT 175.500 134.590 176.000 134.760 ;
        RECT 176.630 134.250 176.800 139.300 ;
        RECT 172.770 134.080 176.800 134.250 ;
        RECT 177.140 138.950 177.310 139.550 ;
        RECT 178.365 139.380 178.845 140.050 ;
        RECT 180.470 139.865 180.640 140.435 ;
        RECT 181.765 140.235 181.935 140.885 ;
        RECT 182.105 140.480 182.535 142.170 ;
        RECT 182.705 141.920 183.535 142.170 ;
        RECT 182.705 141.230 182.875 141.920 ;
        RECT 183.800 141.740 183.970 142.350 ;
        RECT 183.045 141.410 183.970 141.740 ;
        RECT 182.705 141.060 183.535 141.230 ;
        RECT 182.705 140.380 182.875 141.060 ;
        RECT 183.800 140.880 183.970 141.410 ;
        RECT 183.045 140.550 183.970 140.880 ;
        RECT 182.705 140.310 183.535 140.380 ;
        RECT 182.575 140.235 183.535 140.310 ;
        RECT 180.905 140.065 183.535 140.235 ;
        RECT 182.265 140.050 183.535 140.065 ;
        RECT 179.045 139.535 182.065 139.865 ;
        RECT 177.575 139.365 178.845 139.380 ;
        RECT 177.575 139.120 180.205 139.365 ;
        RECT 178.365 139.035 180.205 139.120 ;
        RECT 177.140 138.620 178.195 138.950 ;
        RECT 177.140 138.280 177.310 138.620 ;
        RECT 178.365 138.535 178.845 139.035 ;
        RECT 180.470 138.865 180.640 139.535 ;
        RECT 182.265 139.380 182.745 140.050 ;
        RECT 183.800 139.880 183.970 140.550 ;
        RECT 182.915 139.550 183.970 139.880 ;
        RECT 185.010 149.415 187.110 149.585 ;
        RECT 185.010 140.005 185.180 149.415 ;
        RECT 185.810 148.905 186.310 149.075 ;
        RECT 185.580 147.150 185.750 148.690 ;
        RECT 186.370 147.150 186.540 148.690 ;
        RECT 185.810 146.765 186.310 146.935 ;
        RECT 185.580 145.010 185.750 146.550 ;
        RECT 186.370 145.010 186.540 146.550 ;
        RECT 185.810 144.625 186.310 144.795 ;
        RECT 185.580 142.870 185.750 144.410 ;
        RECT 186.370 142.870 186.540 144.410 ;
        RECT 185.810 142.485 186.310 142.655 ;
        RECT 185.580 140.730 185.750 142.270 ;
        RECT 186.370 140.730 186.540 142.270 ;
        RECT 185.810 140.345 186.310 140.515 ;
        RECT 186.940 140.005 187.110 149.415 ;
        RECT 187.470 149.415 189.570 149.585 ;
        RECT 187.470 144.365 187.640 149.415 ;
        RECT 188.270 148.905 188.770 149.075 ;
        RECT 188.040 148.195 188.210 148.735 ;
        RECT 188.830 148.195 189.000 148.735 ;
        RECT 188.270 147.855 188.770 148.025 ;
        RECT 188.040 147.145 188.210 147.685 ;
        RECT 188.830 147.145 189.000 147.685 ;
        RECT 188.270 146.805 188.770 146.975 ;
        RECT 188.040 146.095 188.210 146.635 ;
        RECT 188.830 146.095 189.000 146.635 ;
        RECT 188.270 145.755 188.770 145.925 ;
        RECT 188.040 145.045 188.210 145.585 ;
        RECT 188.830 145.045 189.000 145.585 ;
        RECT 188.270 144.705 188.770 144.875 ;
        RECT 189.400 144.365 189.570 149.415 ;
        RECT 187.470 144.195 189.570 144.365 ;
        RECT 189.930 149.410 192.030 149.580 ;
        RECT 185.010 139.835 187.110 140.005 ;
        RECT 187.470 143.665 189.570 143.835 ;
        RECT 182.265 139.365 183.535 139.380 ;
        RECT 180.905 139.120 183.535 139.365 ;
        RECT 180.905 139.035 182.745 139.120 ;
        RECT 179.045 138.535 182.065 138.865 ;
        RECT 182.265 138.535 182.745 139.035 ;
        RECT 183.800 138.950 183.970 139.550 ;
        RECT 182.915 138.620 183.970 138.950 ;
        RECT 177.140 138.030 178.355 138.280 ;
        RECT 177.140 137.420 177.310 138.030 ;
        RECT 178.640 137.850 178.840 138.535 ;
        RECT 180.470 138.295 180.640 138.535 ;
        RECT 179.045 138.045 182.065 138.295 ;
        RECT 177.575 137.600 178.405 137.850 ;
        RECT 177.140 137.090 178.065 137.420 ;
        RECT 177.140 136.560 177.310 137.090 ;
        RECT 178.235 136.910 178.405 137.600 ;
        RECT 177.575 136.740 178.405 136.910 ;
        RECT 177.140 136.230 178.065 136.560 ;
        RECT 177.140 135.560 177.310 136.230 ;
        RECT 178.235 136.060 178.405 136.740 ;
        RECT 178.575 136.160 179.005 137.850 ;
        RECT 179.175 137.595 180.205 137.845 ;
        RECT 179.175 136.895 179.345 137.595 ;
        RECT 180.470 137.395 180.640 138.045 ;
        RECT 182.270 137.850 182.470 138.535 ;
        RECT 183.800 138.280 183.970 138.620 ;
        RECT 182.755 138.030 183.970 138.280 ;
        RECT 180.905 137.595 181.935 137.845 ;
        RECT 179.515 137.065 181.595 137.395 ;
        RECT 179.175 136.565 180.205 136.895 ;
        RECT 177.575 135.990 178.405 136.060 ;
        RECT 177.575 135.915 178.535 135.990 ;
        RECT 179.175 135.915 179.345 136.565 ;
        RECT 180.470 136.365 180.640 137.065 ;
        RECT 181.765 136.895 181.935 137.595 ;
        RECT 180.905 136.565 181.935 136.895 ;
        RECT 179.515 136.115 181.595 136.365 ;
        RECT 177.575 135.745 180.205 135.915 ;
        RECT 177.575 135.730 178.845 135.745 ;
        RECT 177.140 135.230 178.195 135.560 ;
        RECT 177.140 134.630 177.310 135.230 ;
        RECT 178.365 135.060 178.845 135.730 ;
        RECT 180.470 135.545 180.640 136.115 ;
        RECT 181.765 135.915 181.935 136.565 ;
        RECT 182.105 136.160 182.535 137.850 ;
        RECT 182.705 137.600 183.535 137.850 ;
        RECT 182.705 136.910 182.875 137.600 ;
        RECT 183.800 137.420 183.970 138.030 ;
        RECT 183.045 137.090 183.970 137.420 ;
        RECT 182.705 136.740 183.535 136.910 ;
        RECT 182.705 136.060 182.875 136.740 ;
        RECT 183.800 136.560 183.970 137.090 ;
        RECT 183.045 136.230 183.970 136.560 ;
        RECT 182.705 135.990 183.535 136.060 ;
        RECT 182.575 135.915 183.535 135.990 ;
        RECT 180.905 135.745 183.535 135.915 ;
        RECT 182.265 135.730 183.535 135.745 ;
        RECT 179.045 135.215 182.065 135.545 ;
        RECT 177.575 135.045 178.845 135.060 ;
        RECT 177.575 134.800 180.205 135.045 ;
        RECT 178.365 134.715 180.205 134.800 ;
        RECT 177.140 134.300 178.195 134.630 ;
        RECT 177.140 134.090 177.310 134.300 ;
        RECT 178.365 134.215 178.845 134.715 ;
        RECT 180.470 134.545 180.640 135.215 ;
        RECT 182.265 135.060 182.745 135.730 ;
        RECT 183.800 135.560 183.970 136.230 ;
        RECT 182.915 135.230 183.970 135.560 ;
        RECT 182.265 135.045 183.535 135.060 ;
        RECT 180.905 134.800 183.535 135.045 ;
        RECT 180.905 134.715 182.745 134.800 ;
        RECT 179.045 134.215 182.065 134.545 ;
        RECT 182.265 134.215 182.745 134.715 ;
        RECT 183.800 134.630 183.970 135.230 ;
        RECT 182.915 134.300 183.970 134.630 ;
        RECT 180.470 134.090 180.640 134.215 ;
        RECT 183.800 134.090 183.970 134.300 ;
        RECT 185.010 139.305 187.110 139.475 ;
        RECT 185.010 134.255 185.180 139.305 ;
        RECT 185.810 138.795 186.310 138.965 ;
        RECT 185.580 138.085 185.750 138.625 ;
        RECT 186.370 138.085 186.540 138.625 ;
        RECT 185.810 137.745 186.310 137.915 ;
        RECT 185.580 137.035 185.750 137.575 ;
        RECT 186.370 137.035 186.540 137.575 ;
        RECT 185.810 136.695 186.310 136.865 ;
        RECT 185.580 135.985 185.750 136.525 ;
        RECT 186.370 135.985 186.540 136.525 ;
        RECT 185.810 135.645 186.310 135.815 ;
        RECT 185.580 134.935 185.750 135.475 ;
        RECT 186.370 134.935 186.540 135.475 ;
        RECT 185.810 134.595 186.310 134.765 ;
        RECT 186.940 134.255 187.110 139.305 ;
        RECT 185.010 134.085 187.110 134.255 ;
        RECT 187.470 134.255 187.640 143.665 ;
        RECT 188.270 143.155 188.770 143.325 ;
        RECT 188.040 141.400 188.210 142.940 ;
        RECT 188.830 141.400 189.000 142.940 ;
        RECT 188.270 141.015 188.770 141.185 ;
        RECT 188.040 139.260 188.210 140.800 ;
        RECT 188.830 139.260 189.000 140.800 ;
        RECT 188.270 138.875 188.770 139.045 ;
        RECT 188.040 137.120 188.210 138.660 ;
        RECT 188.830 137.120 189.000 138.660 ;
        RECT 188.270 136.735 188.770 136.905 ;
        RECT 188.040 134.980 188.210 136.520 ;
        RECT 188.830 134.980 189.000 136.520 ;
        RECT 188.270 134.595 188.770 134.765 ;
        RECT 189.400 134.255 189.570 143.665 ;
        RECT 189.930 140.000 190.100 149.410 ;
        RECT 190.730 148.900 191.230 149.070 ;
        RECT 190.500 147.145 190.670 148.685 ;
        RECT 191.290 147.145 191.460 148.685 ;
        RECT 190.730 146.760 191.230 146.930 ;
        RECT 190.500 145.005 190.670 146.545 ;
        RECT 191.290 145.005 191.460 146.545 ;
        RECT 190.730 144.620 191.230 144.790 ;
        RECT 190.500 142.865 190.670 144.405 ;
        RECT 191.290 142.865 191.460 144.405 ;
        RECT 190.730 142.480 191.230 142.650 ;
        RECT 190.500 140.725 190.670 142.265 ;
        RECT 191.290 140.725 191.460 142.265 ;
        RECT 190.730 140.340 191.230 140.510 ;
        RECT 191.860 140.000 192.030 149.410 ;
        RECT 201.150 148.485 201.320 149.950 ;
        RECT 202.415 149.745 204.215 149.805 ;
        RECT 202.075 149.575 204.215 149.745 ;
        RECT 202.075 149.460 202.245 149.575 ;
        RECT 201.585 149.130 202.245 149.460 ;
        RECT 204.480 149.405 204.650 149.975 ;
        RECT 206.885 149.920 207.545 150.250 ;
        RECT 206.885 149.805 207.055 149.920 ;
        RECT 204.915 149.635 207.055 149.805 ;
        RECT 204.915 149.575 206.715 149.635 ;
        RECT 207.810 149.430 207.980 150.410 ;
        RECT 225.160 150.280 225.330 151.035 ;
        RECT 225.595 150.535 228.225 150.865 ;
        RECT 226.530 150.305 226.730 150.535 ;
        RECT 228.490 150.305 228.660 151.035 ;
        RECT 249.175 151.365 249.345 151.850 ;
        RECT 249.175 151.035 250.390 151.365 ;
        RECT 250.560 151.035 251.040 151.725 ;
        RECT 252.505 151.365 252.675 151.850 ;
        RECT 251.210 151.035 252.675 151.365 ;
        RECT 225.160 149.950 226.255 150.280 ;
        RECT 226.425 149.975 226.795 150.305 ;
        RECT 227.065 149.975 230.085 150.305 ;
        RECT 230.355 149.975 230.725 150.305 ;
        RECT 202.415 149.075 202.785 149.405 ;
        RECT 203.055 149.075 206.075 149.405 ;
        RECT 206.345 149.075 206.715 149.405 ;
        RECT 206.885 149.100 207.980 149.430 ;
        RECT 201.150 148.155 202.365 148.485 ;
        RECT 202.535 148.155 203.015 148.845 ;
        RECT 204.480 148.485 204.650 149.075 ;
        RECT 203.185 148.155 205.945 148.485 ;
        RECT 206.115 148.155 206.595 148.845 ;
        RECT 207.810 148.485 207.980 149.100 ;
        RECT 206.765 148.155 207.980 148.485 ;
        RECT 201.150 147.440 201.320 148.155 ;
        RECT 201.585 147.655 204.215 147.985 ;
        RECT 201.150 147.140 202.340 147.440 ;
        RECT 201.150 146.565 201.320 147.140 ;
        RECT 202.600 146.925 202.800 147.655 ;
        RECT 204.480 147.440 204.650 148.155 ;
        RECT 204.915 147.655 207.545 147.985 ;
        RECT 203.440 147.140 205.690 147.440 ;
        RECT 201.150 146.235 202.365 146.565 ;
        RECT 202.535 146.235 203.015 146.925 ;
        RECT 204.480 146.565 204.650 147.140 ;
        RECT 206.330 146.925 206.530 147.655 ;
        RECT 207.810 147.440 207.980 148.155 ;
        RECT 206.790 147.140 207.980 147.440 ;
        RECT 203.185 146.235 205.945 146.565 ;
        RECT 206.115 146.235 206.595 146.925 ;
        RECT 207.810 146.565 207.980 147.140 ;
        RECT 206.765 146.235 207.980 146.565 ;
        RECT 201.150 145.495 201.320 146.235 ;
        RECT 201.585 145.735 204.215 146.065 ;
        RECT 201.150 145.165 202.365 145.495 ;
        RECT 202.650 145.485 202.850 145.735 ;
        RECT 201.150 144.565 201.320 145.165 ;
        RECT 201.585 144.745 202.415 144.995 ;
        RECT 201.150 144.235 202.075 144.565 ;
        RECT 189.930 139.830 192.030 140.000 ;
        RECT 192.390 143.660 196.420 143.830 ;
        RECT 187.470 134.085 189.570 134.255 ;
        RECT 189.930 139.300 192.030 139.470 ;
        RECT 189.930 134.250 190.100 139.300 ;
        RECT 190.730 138.790 191.230 138.960 ;
        RECT 190.500 138.080 190.670 138.620 ;
        RECT 191.290 138.080 191.460 138.620 ;
        RECT 190.730 137.740 191.230 137.910 ;
        RECT 190.500 137.030 190.670 137.570 ;
        RECT 191.290 137.030 191.460 137.570 ;
        RECT 190.730 136.690 191.230 136.860 ;
        RECT 190.500 135.980 190.670 136.520 ;
        RECT 191.290 135.980 191.460 136.520 ;
        RECT 190.730 135.640 191.230 135.810 ;
        RECT 190.500 134.930 190.670 135.470 ;
        RECT 191.290 134.930 191.460 135.470 ;
        RECT 190.730 134.590 191.230 134.760 ;
        RECT 191.860 134.250 192.030 139.300 ;
        RECT 189.930 134.080 192.030 134.250 ;
        RECT 192.390 134.250 192.560 143.660 ;
        RECT 193.190 143.150 193.690 143.320 ;
        RECT 192.960 141.395 193.130 142.935 ;
        RECT 193.750 141.395 193.920 142.935 ;
        RECT 193.190 141.010 193.690 141.180 ;
        RECT 192.960 139.255 193.130 140.795 ;
        RECT 193.750 139.255 193.920 140.795 ;
        RECT 193.190 138.870 193.690 139.040 ;
        RECT 192.960 137.115 193.130 138.655 ;
        RECT 193.750 137.115 193.920 138.655 ;
        RECT 193.190 136.730 193.690 136.900 ;
        RECT 192.960 134.975 193.130 136.515 ;
        RECT 193.750 134.975 193.920 136.515 ;
        RECT 193.190 134.590 193.690 134.760 ;
        RECT 194.320 134.250 194.490 143.660 ;
        RECT 195.120 143.150 195.620 143.320 ;
        RECT 194.890 141.395 195.060 142.935 ;
        RECT 195.680 141.395 195.850 142.935 ;
        RECT 195.120 141.010 195.620 141.180 ;
        RECT 194.890 139.255 195.060 140.795 ;
        RECT 195.680 139.255 195.850 140.795 ;
        RECT 195.120 138.870 195.620 139.040 ;
        RECT 194.890 137.115 195.060 138.655 ;
        RECT 195.680 137.115 195.850 138.655 ;
        RECT 195.120 136.730 195.620 136.900 ;
        RECT 194.890 134.975 195.060 136.515 ;
        RECT 195.680 134.975 195.850 136.515 ;
        RECT 195.120 134.590 195.620 134.760 ;
        RECT 196.250 134.250 196.420 143.660 ;
        RECT 201.150 143.655 201.320 144.235 ;
        RECT 202.245 144.005 202.415 144.745 ;
        RECT 201.585 143.835 202.415 144.005 ;
        RECT 201.150 143.325 202.075 143.655 ;
        RECT 202.245 143.565 202.415 143.835 ;
        RECT 202.585 143.810 203.015 145.485 ;
        RECT 204.480 145.460 204.650 146.235 ;
        RECT 204.915 145.735 207.545 146.065 ;
        RECT 206.280 145.485 206.480 145.735 ;
        RECT 207.810 145.495 207.980 146.235 ;
        RECT 203.185 145.210 205.945 145.460 ;
        RECT 203.185 144.680 204.215 145.010 ;
        RECT 203.185 144.110 203.355 144.680 ;
        RECT 204.480 144.480 204.650 145.210 ;
        RECT 204.915 144.680 205.945 145.010 ;
        RECT 203.525 144.310 205.605 144.480 ;
        RECT 203.185 143.780 204.215 144.110 ;
        RECT 203.185 143.565 203.355 143.780 ;
        RECT 204.480 143.580 204.650 144.310 ;
        RECT 205.775 144.110 205.945 144.680 ;
        RECT 204.915 143.780 205.945 144.110 ;
        RECT 206.115 143.810 206.545 145.485 ;
        RECT 206.765 145.165 207.980 145.495 ;
        RECT 206.715 144.745 207.545 144.995 ;
        RECT 206.715 144.005 206.885 144.745 ;
        RECT 207.810 144.565 207.980 145.165 ;
        RECT 207.055 144.235 207.980 144.565 ;
        RECT 206.715 143.835 207.545 144.005 ;
        RECT 202.245 143.335 203.355 143.565 ;
        RECT 201.150 143.120 201.320 143.325 ;
        RECT 201.150 142.820 202.340 143.120 ;
        RECT 201.150 142.600 201.320 142.820 ;
        RECT 201.150 142.350 202.365 142.600 ;
        RECT 201.150 141.740 201.320 142.350 ;
        RECT 202.650 142.170 202.850 143.335 ;
        RECT 203.525 143.330 205.605 143.580 ;
        RECT 205.775 143.565 205.945 143.780 ;
        RECT 206.715 143.565 206.885 143.835 ;
        RECT 207.810 143.655 207.980 144.235 ;
        RECT 205.775 143.335 206.885 143.565 ;
        RECT 204.480 143.120 204.650 143.330 ;
        RECT 203.440 142.820 205.690 143.120 ;
        RECT 204.480 142.615 204.650 142.820 ;
        RECT 203.055 142.365 206.075 142.615 ;
        RECT 201.585 141.920 202.415 142.170 ;
        RECT 201.150 141.410 202.075 141.740 ;
        RECT 201.150 140.880 201.320 141.410 ;
        RECT 202.245 141.230 202.415 141.920 ;
        RECT 201.585 141.060 202.415 141.230 ;
        RECT 201.150 140.550 202.075 140.880 ;
        RECT 201.150 139.880 201.320 140.550 ;
        RECT 202.245 140.380 202.415 141.060 ;
        RECT 202.585 140.480 203.015 142.170 ;
        RECT 203.185 141.915 204.215 142.165 ;
        RECT 203.185 141.215 203.355 141.915 ;
        RECT 204.480 141.715 204.650 142.365 ;
        RECT 206.285 142.170 206.485 143.335 ;
        RECT 207.055 143.325 207.980 143.655 ;
        RECT 207.810 143.120 207.980 143.325 ;
        RECT 206.790 142.820 207.980 143.120 ;
        RECT 207.810 142.600 207.980 142.820 ;
        RECT 206.765 142.350 207.980 142.600 ;
        RECT 204.915 141.915 205.945 142.165 ;
        RECT 203.525 141.385 205.605 141.715 ;
        RECT 203.185 140.885 204.215 141.215 ;
        RECT 201.585 140.310 202.415 140.380 ;
        RECT 201.585 140.235 202.545 140.310 ;
        RECT 203.185 140.235 203.355 140.885 ;
        RECT 204.480 140.685 204.650 141.385 ;
        RECT 205.775 141.215 205.945 141.915 ;
        RECT 204.915 140.885 205.945 141.215 ;
        RECT 203.525 140.435 205.605 140.685 ;
        RECT 201.585 140.065 204.215 140.235 ;
        RECT 201.585 140.050 202.855 140.065 ;
        RECT 201.150 139.550 202.205 139.880 ;
        RECT 192.390 134.080 196.420 134.250 ;
        RECT 196.780 139.300 200.810 139.470 ;
        RECT 196.780 134.250 196.950 139.300 ;
        RECT 197.580 138.790 198.080 138.960 ;
        RECT 197.350 138.080 197.520 138.620 ;
        RECT 198.140 138.080 198.310 138.620 ;
        RECT 197.580 137.740 198.080 137.910 ;
        RECT 197.350 137.030 197.520 137.570 ;
        RECT 198.140 137.030 198.310 137.570 ;
        RECT 197.580 136.690 198.080 136.860 ;
        RECT 197.350 135.980 197.520 136.520 ;
        RECT 198.140 135.980 198.310 136.520 ;
        RECT 197.580 135.640 198.080 135.810 ;
        RECT 197.350 134.930 197.520 135.470 ;
        RECT 198.140 134.930 198.310 135.470 ;
        RECT 197.580 134.590 198.080 134.760 ;
        RECT 198.710 134.250 198.880 139.300 ;
        RECT 199.510 138.790 200.010 138.960 ;
        RECT 199.280 138.080 199.450 138.620 ;
        RECT 200.070 138.080 200.240 138.620 ;
        RECT 199.510 137.740 200.010 137.910 ;
        RECT 199.280 137.030 199.450 137.570 ;
        RECT 200.070 137.030 200.240 137.570 ;
        RECT 199.510 136.690 200.010 136.860 ;
        RECT 199.280 135.980 199.450 136.520 ;
        RECT 200.070 135.980 200.240 136.520 ;
        RECT 199.510 135.640 200.010 135.810 ;
        RECT 199.280 134.930 199.450 135.470 ;
        RECT 200.070 134.930 200.240 135.470 ;
        RECT 199.510 134.590 200.010 134.760 ;
        RECT 200.640 134.250 200.810 139.300 ;
        RECT 196.780 134.080 200.810 134.250 ;
        RECT 201.150 138.950 201.320 139.550 ;
        RECT 202.375 139.380 202.855 140.050 ;
        RECT 204.480 139.865 204.650 140.435 ;
        RECT 205.775 140.235 205.945 140.885 ;
        RECT 206.115 140.480 206.545 142.170 ;
        RECT 206.715 141.920 207.545 142.170 ;
        RECT 206.715 141.230 206.885 141.920 ;
        RECT 207.810 141.740 207.980 142.350 ;
        RECT 207.055 141.410 207.980 141.740 ;
        RECT 206.715 141.060 207.545 141.230 ;
        RECT 206.715 140.380 206.885 141.060 ;
        RECT 207.810 140.880 207.980 141.410 ;
        RECT 207.055 140.550 207.980 140.880 ;
        RECT 206.715 140.310 207.545 140.380 ;
        RECT 206.585 140.235 207.545 140.310 ;
        RECT 204.915 140.065 207.545 140.235 ;
        RECT 206.275 140.050 207.545 140.065 ;
        RECT 203.055 139.535 206.075 139.865 ;
        RECT 201.585 139.365 202.855 139.380 ;
        RECT 201.585 139.120 204.215 139.365 ;
        RECT 202.375 139.035 204.215 139.120 ;
        RECT 201.150 138.620 202.205 138.950 ;
        RECT 201.150 138.280 201.320 138.620 ;
        RECT 202.375 138.535 202.855 139.035 ;
        RECT 204.480 138.865 204.650 139.535 ;
        RECT 206.275 139.380 206.755 140.050 ;
        RECT 207.810 139.880 207.980 140.550 ;
        RECT 206.925 139.550 207.980 139.880 ;
        RECT 209.020 149.415 211.120 149.585 ;
        RECT 209.020 140.005 209.190 149.415 ;
        RECT 209.820 148.905 210.320 149.075 ;
        RECT 209.590 147.150 209.760 148.690 ;
        RECT 210.380 147.150 210.550 148.690 ;
        RECT 209.820 146.765 210.320 146.935 ;
        RECT 209.590 145.010 209.760 146.550 ;
        RECT 210.380 145.010 210.550 146.550 ;
        RECT 209.820 144.625 210.320 144.795 ;
        RECT 209.590 142.870 209.760 144.410 ;
        RECT 210.380 142.870 210.550 144.410 ;
        RECT 209.820 142.485 210.320 142.655 ;
        RECT 209.590 140.730 209.760 142.270 ;
        RECT 210.380 140.730 210.550 142.270 ;
        RECT 209.820 140.345 210.320 140.515 ;
        RECT 210.950 140.005 211.120 149.415 ;
        RECT 211.480 149.415 213.580 149.585 ;
        RECT 211.480 144.365 211.650 149.415 ;
        RECT 212.280 148.905 212.780 149.075 ;
        RECT 212.050 148.195 212.220 148.735 ;
        RECT 212.840 148.195 213.010 148.735 ;
        RECT 212.280 147.855 212.780 148.025 ;
        RECT 212.050 147.145 212.220 147.685 ;
        RECT 212.840 147.145 213.010 147.685 ;
        RECT 212.280 146.805 212.780 146.975 ;
        RECT 212.050 146.095 212.220 146.635 ;
        RECT 212.840 146.095 213.010 146.635 ;
        RECT 212.280 145.755 212.780 145.925 ;
        RECT 212.050 145.045 212.220 145.585 ;
        RECT 212.840 145.045 213.010 145.585 ;
        RECT 212.280 144.705 212.780 144.875 ;
        RECT 213.410 144.365 213.580 149.415 ;
        RECT 211.480 144.195 213.580 144.365 ;
        RECT 213.940 149.410 216.040 149.580 ;
        RECT 209.020 139.835 211.120 140.005 ;
        RECT 211.480 143.665 213.580 143.835 ;
        RECT 206.275 139.365 207.545 139.380 ;
        RECT 204.915 139.120 207.545 139.365 ;
        RECT 204.915 139.035 206.755 139.120 ;
        RECT 203.055 138.535 206.075 138.865 ;
        RECT 206.275 138.535 206.755 139.035 ;
        RECT 207.810 138.950 207.980 139.550 ;
        RECT 206.925 138.620 207.980 138.950 ;
        RECT 201.150 138.030 202.365 138.280 ;
        RECT 201.150 137.420 201.320 138.030 ;
        RECT 202.650 137.850 202.850 138.535 ;
        RECT 204.480 138.295 204.650 138.535 ;
        RECT 203.055 138.045 206.075 138.295 ;
        RECT 201.585 137.600 202.415 137.850 ;
        RECT 201.150 137.090 202.075 137.420 ;
        RECT 201.150 136.560 201.320 137.090 ;
        RECT 202.245 136.910 202.415 137.600 ;
        RECT 201.585 136.740 202.415 136.910 ;
        RECT 201.150 136.230 202.075 136.560 ;
        RECT 201.150 135.560 201.320 136.230 ;
        RECT 202.245 136.060 202.415 136.740 ;
        RECT 202.585 136.160 203.015 137.850 ;
        RECT 203.185 137.595 204.215 137.845 ;
        RECT 203.185 136.895 203.355 137.595 ;
        RECT 204.480 137.395 204.650 138.045 ;
        RECT 206.280 137.850 206.480 138.535 ;
        RECT 207.810 138.280 207.980 138.620 ;
        RECT 206.765 138.030 207.980 138.280 ;
        RECT 204.915 137.595 205.945 137.845 ;
        RECT 203.525 137.065 205.605 137.395 ;
        RECT 203.185 136.565 204.215 136.895 ;
        RECT 201.585 135.990 202.415 136.060 ;
        RECT 201.585 135.915 202.545 135.990 ;
        RECT 203.185 135.915 203.355 136.565 ;
        RECT 204.480 136.365 204.650 137.065 ;
        RECT 205.775 136.895 205.945 137.595 ;
        RECT 204.915 136.565 205.945 136.895 ;
        RECT 203.525 136.115 205.605 136.365 ;
        RECT 201.585 135.745 204.215 135.915 ;
        RECT 201.585 135.730 202.855 135.745 ;
        RECT 201.150 135.230 202.205 135.560 ;
        RECT 201.150 134.630 201.320 135.230 ;
        RECT 202.375 135.060 202.855 135.730 ;
        RECT 204.480 135.545 204.650 136.115 ;
        RECT 205.775 135.915 205.945 136.565 ;
        RECT 206.115 136.160 206.545 137.850 ;
        RECT 206.715 137.600 207.545 137.850 ;
        RECT 206.715 136.910 206.885 137.600 ;
        RECT 207.810 137.420 207.980 138.030 ;
        RECT 207.055 137.090 207.980 137.420 ;
        RECT 206.715 136.740 207.545 136.910 ;
        RECT 206.715 136.060 206.885 136.740 ;
        RECT 207.810 136.560 207.980 137.090 ;
        RECT 207.055 136.230 207.980 136.560 ;
        RECT 206.715 135.990 207.545 136.060 ;
        RECT 206.585 135.915 207.545 135.990 ;
        RECT 204.915 135.745 207.545 135.915 ;
        RECT 206.275 135.730 207.545 135.745 ;
        RECT 203.055 135.215 206.075 135.545 ;
        RECT 201.585 135.045 202.855 135.060 ;
        RECT 201.585 134.800 204.215 135.045 ;
        RECT 202.375 134.715 204.215 134.800 ;
        RECT 201.150 134.300 202.205 134.630 ;
        RECT 201.150 134.090 201.320 134.300 ;
        RECT 202.375 134.215 202.855 134.715 ;
        RECT 204.480 134.545 204.650 135.215 ;
        RECT 206.275 135.060 206.755 135.730 ;
        RECT 207.810 135.560 207.980 136.230 ;
        RECT 206.925 135.230 207.980 135.560 ;
        RECT 206.275 135.045 207.545 135.060 ;
        RECT 204.915 134.800 207.545 135.045 ;
        RECT 204.915 134.715 206.755 134.800 ;
        RECT 203.055 134.215 206.075 134.545 ;
        RECT 206.275 134.215 206.755 134.715 ;
        RECT 207.810 134.630 207.980 135.230 ;
        RECT 206.925 134.300 207.980 134.630 ;
        RECT 204.480 134.090 204.650 134.215 ;
        RECT 207.810 134.090 207.980 134.300 ;
        RECT 209.020 139.305 211.120 139.475 ;
        RECT 209.020 134.255 209.190 139.305 ;
        RECT 209.820 138.795 210.320 138.965 ;
        RECT 209.590 138.085 209.760 138.625 ;
        RECT 210.380 138.085 210.550 138.625 ;
        RECT 209.820 137.745 210.320 137.915 ;
        RECT 209.590 137.035 209.760 137.575 ;
        RECT 210.380 137.035 210.550 137.575 ;
        RECT 209.820 136.695 210.320 136.865 ;
        RECT 209.590 135.985 209.760 136.525 ;
        RECT 210.380 135.985 210.550 136.525 ;
        RECT 209.820 135.645 210.320 135.815 ;
        RECT 209.590 134.935 209.760 135.475 ;
        RECT 210.380 134.935 210.550 135.475 ;
        RECT 209.820 134.595 210.320 134.765 ;
        RECT 210.950 134.255 211.120 139.305 ;
        RECT 209.020 134.085 211.120 134.255 ;
        RECT 211.480 134.255 211.650 143.665 ;
        RECT 212.280 143.155 212.780 143.325 ;
        RECT 212.050 141.400 212.220 142.940 ;
        RECT 212.840 141.400 213.010 142.940 ;
        RECT 212.280 141.015 212.780 141.185 ;
        RECT 212.050 139.260 212.220 140.800 ;
        RECT 212.840 139.260 213.010 140.800 ;
        RECT 212.280 138.875 212.780 139.045 ;
        RECT 212.050 137.120 212.220 138.660 ;
        RECT 212.840 137.120 213.010 138.660 ;
        RECT 212.280 136.735 212.780 136.905 ;
        RECT 212.050 134.980 212.220 136.520 ;
        RECT 212.840 134.980 213.010 136.520 ;
        RECT 212.280 134.595 212.780 134.765 ;
        RECT 213.410 134.255 213.580 143.665 ;
        RECT 213.940 140.000 214.110 149.410 ;
        RECT 214.740 148.900 215.240 149.070 ;
        RECT 214.510 147.145 214.680 148.685 ;
        RECT 215.300 147.145 215.470 148.685 ;
        RECT 214.740 146.760 215.240 146.930 ;
        RECT 214.510 145.005 214.680 146.545 ;
        RECT 215.300 145.005 215.470 146.545 ;
        RECT 214.740 144.620 215.240 144.790 ;
        RECT 214.510 142.865 214.680 144.405 ;
        RECT 215.300 142.865 215.470 144.405 ;
        RECT 214.740 142.480 215.240 142.650 ;
        RECT 214.510 140.725 214.680 142.265 ;
        RECT 215.300 140.725 215.470 142.265 ;
        RECT 214.740 140.340 215.240 140.510 ;
        RECT 215.870 140.000 216.040 149.410 ;
        RECT 225.160 148.485 225.330 149.950 ;
        RECT 226.425 149.745 228.225 149.805 ;
        RECT 226.085 149.575 228.225 149.745 ;
        RECT 226.085 149.460 226.255 149.575 ;
        RECT 225.595 149.130 226.255 149.460 ;
        RECT 228.490 149.405 228.660 149.975 ;
        RECT 230.895 149.920 231.555 150.250 ;
        RECT 230.895 149.805 231.065 149.920 ;
        RECT 228.925 149.635 231.065 149.805 ;
        RECT 228.925 149.575 230.725 149.635 ;
        RECT 231.820 149.430 231.990 150.410 ;
        RECT 249.175 150.280 249.345 151.035 ;
        RECT 249.610 150.535 252.240 150.865 ;
        RECT 250.545 150.305 250.745 150.535 ;
        RECT 252.505 150.305 252.675 151.035 ;
        RECT 273.230 151.365 273.400 151.850 ;
        RECT 273.230 151.035 274.445 151.365 ;
        RECT 274.615 151.035 275.095 151.725 ;
        RECT 276.560 151.365 276.730 151.850 ;
        RECT 275.265 151.035 276.730 151.365 ;
        RECT 249.175 149.950 250.270 150.280 ;
        RECT 250.440 149.975 250.810 150.305 ;
        RECT 251.080 149.975 254.100 150.305 ;
        RECT 254.370 149.975 254.740 150.305 ;
        RECT 226.425 149.075 226.795 149.405 ;
        RECT 227.065 149.075 230.085 149.405 ;
        RECT 230.355 149.075 230.725 149.405 ;
        RECT 230.895 149.100 231.990 149.430 ;
        RECT 225.160 148.155 226.375 148.485 ;
        RECT 226.545 148.155 227.025 148.845 ;
        RECT 228.490 148.485 228.660 149.075 ;
        RECT 227.195 148.155 229.955 148.485 ;
        RECT 230.125 148.155 230.605 148.845 ;
        RECT 231.820 148.485 231.990 149.100 ;
        RECT 230.775 148.155 231.990 148.485 ;
        RECT 225.160 147.440 225.330 148.155 ;
        RECT 225.595 147.655 228.225 147.985 ;
        RECT 225.160 147.140 226.350 147.440 ;
        RECT 225.160 146.565 225.330 147.140 ;
        RECT 226.610 146.925 226.810 147.655 ;
        RECT 228.490 147.440 228.660 148.155 ;
        RECT 228.925 147.655 231.555 147.985 ;
        RECT 227.450 147.140 229.700 147.440 ;
        RECT 225.160 146.235 226.375 146.565 ;
        RECT 226.545 146.235 227.025 146.925 ;
        RECT 228.490 146.565 228.660 147.140 ;
        RECT 230.340 146.925 230.540 147.655 ;
        RECT 231.820 147.440 231.990 148.155 ;
        RECT 230.800 147.140 231.990 147.440 ;
        RECT 227.195 146.235 229.955 146.565 ;
        RECT 230.125 146.235 230.605 146.925 ;
        RECT 231.820 146.565 231.990 147.140 ;
        RECT 230.775 146.235 231.990 146.565 ;
        RECT 225.160 145.495 225.330 146.235 ;
        RECT 225.595 145.735 228.225 146.065 ;
        RECT 225.160 145.165 226.375 145.495 ;
        RECT 226.660 145.485 226.860 145.735 ;
        RECT 225.160 144.565 225.330 145.165 ;
        RECT 225.595 144.745 226.425 144.995 ;
        RECT 225.160 144.235 226.085 144.565 ;
        RECT 213.940 139.830 216.040 140.000 ;
        RECT 216.400 143.660 220.430 143.830 ;
        RECT 211.480 134.085 213.580 134.255 ;
        RECT 213.940 139.300 216.040 139.470 ;
        RECT 213.940 134.250 214.110 139.300 ;
        RECT 214.740 138.790 215.240 138.960 ;
        RECT 214.510 138.080 214.680 138.620 ;
        RECT 215.300 138.080 215.470 138.620 ;
        RECT 214.740 137.740 215.240 137.910 ;
        RECT 214.510 137.030 214.680 137.570 ;
        RECT 215.300 137.030 215.470 137.570 ;
        RECT 214.740 136.690 215.240 136.860 ;
        RECT 214.510 135.980 214.680 136.520 ;
        RECT 215.300 135.980 215.470 136.520 ;
        RECT 214.740 135.640 215.240 135.810 ;
        RECT 214.510 134.930 214.680 135.470 ;
        RECT 215.300 134.930 215.470 135.470 ;
        RECT 214.740 134.590 215.240 134.760 ;
        RECT 215.870 134.250 216.040 139.300 ;
        RECT 213.940 134.080 216.040 134.250 ;
        RECT 216.400 134.250 216.570 143.660 ;
        RECT 217.200 143.150 217.700 143.320 ;
        RECT 216.970 141.395 217.140 142.935 ;
        RECT 217.760 141.395 217.930 142.935 ;
        RECT 217.200 141.010 217.700 141.180 ;
        RECT 216.970 139.255 217.140 140.795 ;
        RECT 217.760 139.255 217.930 140.795 ;
        RECT 217.200 138.870 217.700 139.040 ;
        RECT 216.970 137.115 217.140 138.655 ;
        RECT 217.760 137.115 217.930 138.655 ;
        RECT 217.200 136.730 217.700 136.900 ;
        RECT 216.970 134.975 217.140 136.515 ;
        RECT 217.760 134.975 217.930 136.515 ;
        RECT 217.200 134.590 217.700 134.760 ;
        RECT 218.330 134.250 218.500 143.660 ;
        RECT 219.130 143.150 219.630 143.320 ;
        RECT 218.900 141.395 219.070 142.935 ;
        RECT 219.690 141.395 219.860 142.935 ;
        RECT 219.130 141.010 219.630 141.180 ;
        RECT 218.900 139.255 219.070 140.795 ;
        RECT 219.690 139.255 219.860 140.795 ;
        RECT 219.130 138.870 219.630 139.040 ;
        RECT 218.900 137.115 219.070 138.655 ;
        RECT 219.690 137.115 219.860 138.655 ;
        RECT 219.130 136.730 219.630 136.900 ;
        RECT 218.900 134.975 219.070 136.515 ;
        RECT 219.690 134.975 219.860 136.515 ;
        RECT 219.130 134.590 219.630 134.760 ;
        RECT 220.260 134.250 220.430 143.660 ;
        RECT 225.160 143.655 225.330 144.235 ;
        RECT 226.255 144.005 226.425 144.745 ;
        RECT 225.595 143.835 226.425 144.005 ;
        RECT 225.160 143.325 226.085 143.655 ;
        RECT 226.255 143.565 226.425 143.835 ;
        RECT 226.595 143.810 227.025 145.485 ;
        RECT 228.490 145.460 228.660 146.235 ;
        RECT 228.925 145.735 231.555 146.065 ;
        RECT 230.290 145.485 230.490 145.735 ;
        RECT 231.820 145.495 231.990 146.235 ;
        RECT 227.195 145.210 229.955 145.460 ;
        RECT 227.195 144.680 228.225 145.010 ;
        RECT 227.195 144.110 227.365 144.680 ;
        RECT 228.490 144.480 228.660 145.210 ;
        RECT 228.925 144.680 229.955 145.010 ;
        RECT 227.535 144.310 229.615 144.480 ;
        RECT 227.195 143.780 228.225 144.110 ;
        RECT 227.195 143.565 227.365 143.780 ;
        RECT 228.490 143.580 228.660 144.310 ;
        RECT 229.785 144.110 229.955 144.680 ;
        RECT 228.925 143.780 229.955 144.110 ;
        RECT 230.125 143.810 230.555 145.485 ;
        RECT 230.775 145.165 231.990 145.495 ;
        RECT 230.725 144.745 231.555 144.995 ;
        RECT 230.725 144.005 230.895 144.745 ;
        RECT 231.820 144.565 231.990 145.165 ;
        RECT 231.065 144.235 231.990 144.565 ;
        RECT 230.725 143.835 231.555 144.005 ;
        RECT 226.255 143.335 227.365 143.565 ;
        RECT 225.160 143.120 225.330 143.325 ;
        RECT 225.160 142.820 226.350 143.120 ;
        RECT 225.160 142.600 225.330 142.820 ;
        RECT 225.160 142.350 226.375 142.600 ;
        RECT 225.160 141.740 225.330 142.350 ;
        RECT 226.660 142.170 226.860 143.335 ;
        RECT 227.535 143.330 229.615 143.580 ;
        RECT 229.785 143.565 229.955 143.780 ;
        RECT 230.725 143.565 230.895 143.835 ;
        RECT 231.820 143.655 231.990 144.235 ;
        RECT 229.785 143.335 230.895 143.565 ;
        RECT 228.490 143.120 228.660 143.330 ;
        RECT 227.450 142.820 229.700 143.120 ;
        RECT 228.490 142.615 228.660 142.820 ;
        RECT 227.065 142.365 230.085 142.615 ;
        RECT 225.595 141.920 226.425 142.170 ;
        RECT 225.160 141.410 226.085 141.740 ;
        RECT 225.160 140.880 225.330 141.410 ;
        RECT 226.255 141.230 226.425 141.920 ;
        RECT 225.595 141.060 226.425 141.230 ;
        RECT 225.160 140.550 226.085 140.880 ;
        RECT 225.160 139.880 225.330 140.550 ;
        RECT 226.255 140.380 226.425 141.060 ;
        RECT 226.595 140.480 227.025 142.170 ;
        RECT 227.195 141.915 228.225 142.165 ;
        RECT 227.195 141.215 227.365 141.915 ;
        RECT 228.490 141.715 228.660 142.365 ;
        RECT 230.295 142.170 230.495 143.335 ;
        RECT 231.065 143.325 231.990 143.655 ;
        RECT 231.820 143.120 231.990 143.325 ;
        RECT 230.800 142.820 231.990 143.120 ;
        RECT 231.820 142.600 231.990 142.820 ;
        RECT 230.775 142.350 231.990 142.600 ;
        RECT 228.925 141.915 229.955 142.165 ;
        RECT 227.535 141.385 229.615 141.715 ;
        RECT 227.195 140.885 228.225 141.215 ;
        RECT 225.595 140.310 226.425 140.380 ;
        RECT 225.595 140.235 226.555 140.310 ;
        RECT 227.195 140.235 227.365 140.885 ;
        RECT 228.490 140.685 228.660 141.385 ;
        RECT 229.785 141.215 229.955 141.915 ;
        RECT 228.925 140.885 229.955 141.215 ;
        RECT 227.535 140.435 229.615 140.685 ;
        RECT 225.595 140.065 228.225 140.235 ;
        RECT 225.595 140.050 226.865 140.065 ;
        RECT 225.160 139.550 226.215 139.880 ;
        RECT 216.400 134.080 220.430 134.250 ;
        RECT 220.790 139.300 224.820 139.470 ;
        RECT 220.790 134.250 220.960 139.300 ;
        RECT 221.590 138.790 222.090 138.960 ;
        RECT 221.360 138.080 221.530 138.620 ;
        RECT 222.150 138.080 222.320 138.620 ;
        RECT 221.590 137.740 222.090 137.910 ;
        RECT 221.360 137.030 221.530 137.570 ;
        RECT 222.150 137.030 222.320 137.570 ;
        RECT 221.590 136.690 222.090 136.860 ;
        RECT 221.360 135.980 221.530 136.520 ;
        RECT 222.150 135.980 222.320 136.520 ;
        RECT 221.590 135.640 222.090 135.810 ;
        RECT 221.360 134.930 221.530 135.470 ;
        RECT 222.150 134.930 222.320 135.470 ;
        RECT 221.590 134.590 222.090 134.760 ;
        RECT 222.720 134.250 222.890 139.300 ;
        RECT 223.520 138.790 224.020 138.960 ;
        RECT 223.290 138.080 223.460 138.620 ;
        RECT 224.080 138.080 224.250 138.620 ;
        RECT 223.520 137.740 224.020 137.910 ;
        RECT 223.290 137.030 223.460 137.570 ;
        RECT 224.080 137.030 224.250 137.570 ;
        RECT 223.520 136.690 224.020 136.860 ;
        RECT 223.290 135.980 223.460 136.520 ;
        RECT 224.080 135.980 224.250 136.520 ;
        RECT 223.520 135.640 224.020 135.810 ;
        RECT 223.290 134.930 223.460 135.470 ;
        RECT 224.080 134.930 224.250 135.470 ;
        RECT 223.520 134.590 224.020 134.760 ;
        RECT 224.650 134.250 224.820 139.300 ;
        RECT 220.790 134.080 224.820 134.250 ;
        RECT 225.160 138.950 225.330 139.550 ;
        RECT 226.385 139.380 226.865 140.050 ;
        RECT 228.490 139.865 228.660 140.435 ;
        RECT 229.785 140.235 229.955 140.885 ;
        RECT 230.125 140.480 230.555 142.170 ;
        RECT 230.725 141.920 231.555 142.170 ;
        RECT 230.725 141.230 230.895 141.920 ;
        RECT 231.820 141.740 231.990 142.350 ;
        RECT 231.065 141.410 231.990 141.740 ;
        RECT 230.725 141.060 231.555 141.230 ;
        RECT 230.725 140.380 230.895 141.060 ;
        RECT 231.820 140.880 231.990 141.410 ;
        RECT 231.065 140.550 231.990 140.880 ;
        RECT 230.725 140.310 231.555 140.380 ;
        RECT 230.595 140.235 231.555 140.310 ;
        RECT 228.925 140.065 231.555 140.235 ;
        RECT 230.285 140.050 231.555 140.065 ;
        RECT 227.065 139.535 230.085 139.865 ;
        RECT 225.595 139.365 226.865 139.380 ;
        RECT 225.595 139.120 228.225 139.365 ;
        RECT 226.385 139.035 228.225 139.120 ;
        RECT 225.160 138.620 226.215 138.950 ;
        RECT 225.160 138.280 225.330 138.620 ;
        RECT 226.385 138.535 226.865 139.035 ;
        RECT 228.490 138.865 228.660 139.535 ;
        RECT 230.285 139.380 230.765 140.050 ;
        RECT 231.820 139.880 231.990 140.550 ;
        RECT 230.935 139.550 231.990 139.880 ;
        RECT 233.035 149.415 235.135 149.585 ;
        RECT 233.035 140.005 233.205 149.415 ;
        RECT 233.835 148.905 234.335 149.075 ;
        RECT 233.605 147.150 233.775 148.690 ;
        RECT 234.395 147.150 234.565 148.690 ;
        RECT 233.835 146.765 234.335 146.935 ;
        RECT 233.605 145.010 233.775 146.550 ;
        RECT 234.395 145.010 234.565 146.550 ;
        RECT 233.835 144.625 234.335 144.795 ;
        RECT 233.605 142.870 233.775 144.410 ;
        RECT 234.395 142.870 234.565 144.410 ;
        RECT 233.835 142.485 234.335 142.655 ;
        RECT 233.605 140.730 233.775 142.270 ;
        RECT 234.395 140.730 234.565 142.270 ;
        RECT 233.835 140.345 234.335 140.515 ;
        RECT 234.965 140.005 235.135 149.415 ;
        RECT 235.495 149.415 237.595 149.585 ;
        RECT 235.495 144.365 235.665 149.415 ;
        RECT 236.295 148.905 236.795 149.075 ;
        RECT 236.065 148.195 236.235 148.735 ;
        RECT 236.855 148.195 237.025 148.735 ;
        RECT 236.295 147.855 236.795 148.025 ;
        RECT 236.065 147.145 236.235 147.685 ;
        RECT 236.855 147.145 237.025 147.685 ;
        RECT 236.295 146.805 236.795 146.975 ;
        RECT 236.065 146.095 236.235 146.635 ;
        RECT 236.855 146.095 237.025 146.635 ;
        RECT 236.295 145.755 236.795 145.925 ;
        RECT 236.065 145.045 236.235 145.585 ;
        RECT 236.855 145.045 237.025 145.585 ;
        RECT 236.295 144.705 236.795 144.875 ;
        RECT 237.425 144.365 237.595 149.415 ;
        RECT 235.495 144.195 237.595 144.365 ;
        RECT 237.955 149.410 240.055 149.580 ;
        RECT 233.035 139.835 235.135 140.005 ;
        RECT 235.495 143.665 237.595 143.835 ;
        RECT 230.285 139.365 231.555 139.380 ;
        RECT 228.925 139.120 231.555 139.365 ;
        RECT 228.925 139.035 230.765 139.120 ;
        RECT 227.065 138.535 230.085 138.865 ;
        RECT 230.285 138.535 230.765 139.035 ;
        RECT 231.820 138.950 231.990 139.550 ;
        RECT 230.935 138.620 231.990 138.950 ;
        RECT 225.160 138.030 226.375 138.280 ;
        RECT 225.160 137.420 225.330 138.030 ;
        RECT 226.660 137.850 226.860 138.535 ;
        RECT 228.490 138.295 228.660 138.535 ;
        RECT 227.065 138.045 230.085 138.295 ;
        RECT 225.595 137.600 226.425 137.850 ;
        RECT 225.160 137.090 226.085 137.420 ;
        RECT 225.160 136.560 225.330 137.090 ;
        RECT 226.255 136.910 226.425 137.600 ;
        RECT 225.595 136.740 226.425 136.910 ;
        RECT 225.160 136.230 226.085 136.560 ;
        RECT 225.160 135.560 225.330 136.230 ;
        RECT 226.255 136.060 226.425 136.740 ;
        RECT 226.595 136.160 227.025 137.850 ;
        RECT 227.195 137.595 228.225 137.845 ;
        RECT 227.195 136.895 227.365 137.595 ;
        RECT 228.490 137.395 228.660 138.045 ;
        RECT 230.290 137.850 230.490 138.535 ;
        RECT 231.820 138.280 231.990 138.620 ;
        RECT 230.775 138.030 231.990 138.280 ;
        RECT 228.925 137.595 229.955 137.845 ;
        RECT 227.535 137.065 229.615 137.395 ;
        RECT 227.195 136.565 228.225 136.895 ;
        RECT 225.595 135.990 226.425 136.060 ;
        RECT 225.595 135.915 226.555 135.990 ;
        RECT 227.195 135.915 227.365 136.565 ;
        RECT 228.490 136.365 228.660 137.065 ;
        RECT 229.785 136.895 229.955 137.595 ;
        RECT 228.925 136.565 229.955 136.895 ;
        RECT 227.535 136.115 229.615 136.365 ;
        RECT 225.595 135.745 228.225 135.915 ;
        RECT 225.595 135.730 226.865 135.745 ;
        RECT 225.160 135.230 226.215 135.560 ;
        RECT 225.160 134.630 225.330 135.230 ;
        RECT 226.385 135.060 226.865 135.730 ;
        RECT 228.490 135.545 228.660 136.115 ;
        RECT 229.785 135.915 229.955 136.565 ;
        RECT 230.125 136.160 230.555 137.850 ;
        RECT 230.725 137.600 231.555 137.850 ;
        RECT 230.725 136.910 230.895 137.600 ;
        RECT 231.820 137.420 231.990 138.030 ;
        RECT 231.065 137.090 231.990 137.420 ;
        RECT 230.725 136.740 231.555 136.910 ;
        RECT 230.725 136.060 230.895 136.740 ;
        RECT 231.820 136.560 231.990 137.090 ;
        RECT 231.065 136.230 231.990 136.560 ;
        RECT 230.725 135.990 231.555 136.060 ;
        RECT 230.595 135.915 231.555 135.990 ;
        RECT 228.925 135.745 231.555 135.915 ;
        RECT 230.285 135.730 231.555 135.745 ;
        RECT 227.065 135.215 230.085 135.545 ;
        RECT 225.595 135.045 226.865 135.060 ;
        RECT 225.595 134.800 228.225 135.045 ;
        RECT 226.385 134.715 228.225 134.800 ;
        RECT 225.160 134.300 226.215 134.630 ;
        RECT 225.160 134.090 225.330 134.300 ;
        RECT 226.385 134.215 226.865 134.715 ;
        RECT 228.490 134.545 228.660 135.215 ;
        RECT 230.285 135.060 230.765 135.730 ;
        RECT 231.820 135.560 231.990 136.230 ;
        RECT 230.935 135.230 231.990 135.560 ;
        RECT 230.285 135.045 231.555 135.060 ;
        RECT 228.925 134.800 231.555 135.045 ;
        RECT 228.925 134.715 230.765 134.800 ;
        RECT 227.065 134.215 230.085 134.545 ;
        RECT 230.285 134.215 230.765 134.715 ;
        RECT 231.820 134.630 231.990 135.230 ;
        RECT 230.935 134.300 231.990 134.630 ;
        RECT 228.490 134.090 228.660 134.215 ;
        RECT 231.820 134.090 231.990 134.300 ;
        RECT 233.035 139.305 235.135 139.475 ;
        RECT 233.035 134.255 233.205 139.305 ;
        RECT 233.835 138.795 234.335 138.965 ;
        RECT 233.605 138.085 233.775 138.625 ;
        RECT 234.395 138.085 234.565 138.625 ;
        RECT 233.835 137.745 234.335 137.915 ;
        RECT 233.605 137.035 233.775 137.575 ;
        RECT 234.395 137.035 234.565 137.575 ;
        RECT 233.835 136.695 234.335 136.865 ;
        RECT 233.605 135.985 233.775 136.525 ;
        RECT 234.395 135.985 234.565 136.525 ;
        RECT 233.835 135.645 234.335 135.815 ;
        RECT 233.605 134.935 233.775 135.475 ;
        RECT 234.395 134.935 234.565 135.475 ;
        RECT 233.835 134.595 234.335 134.765 ;
        RECT 234.965 134.255 235.135 139.305 ;
        RECT 233.035 134.085 235.135 134.255 ;
        RECT 235.495 134.255 235.665 143.665 ;
        RECT 236.295 143.155 236.795 143.325 ;
        RECT 236.065 141.400 236.235 142.940 ;
        RECT 236.855 141.400 237.025 142.940 ;
        RECT 236.295 141.015 236.795 141.185 ;
        RECT 236.065 139.260 236.235 140.800 ;
        RECT 236.855 139.260 237.025 140.800 ;
        RECT 236.295 138.875 236.795 139.045 ;
        RECT 236.065 137.120 236.235 138.660 ;
        RECT 236.855 137.120 237.025 138.660 ;
        RECT 236.295 136.735 236.795 136.905 ;
        RECT 236.065 134.980 236.235 136.520 ;
        RECT 236.855 134.980 237.025 136.520 ;
        RECT 236.295 134.595 236.795 134.765 ;
        RECT 237.425 134.255 237.595 143.665 ;
        RECT 237.955 140.000 238.125 149.410 ;
        RECT 238.755 148.900 239.255 149.070 ;
        RECT 238.525 147.145 238.695 148.685 ;
        RECT 239.315 147.145 239.485 148.685 ;
        RECT 238.755 146.760 239.255 146.930 ;
        RECT 238.525 145.005 238.695 146.545 ;
        RECT 239.315 145.005 239.485 146.545 ;
        RECT 238.755 144.620 239.255 144.790 ;
        RECT 238.525 142.865 238.695 144.405 ;
        RECT 239.315 142.865 239.485 144.405 ;
        RECT 238.755 142.480 239.255 142.650 ;
        RECT 238.525 140.725 238.695 142.265 ;
        RECT 239.315 140.725 239.485 142.265 ;
        RECT 238.755 140.340 239.255 140.510 ;
        RECT 239.885 140.000 240.055 149.410 ;
        RECT 249.175 148.485 249.345 149.950 ;
        RECT 250.440 149.745 252.240 149.805 ;
        RECT 250.100 149.575 252.240 149.745 ;
        RECT 250.100 149.460 250.270 149.575 ;
        RECT 249.610 149.130 250.270 149.460 ;
        RECT 252.505 149.405 252.675 149.975 ;
        RECT 254.910 149.920 255.570 150.250 ;
        RECT 254.910 149.805 255.080 149.920 ;
        RECT 252.940 149.635 255.080 149.805 ;
        RECT 252.940 149.575 254.740 149.635 ;
        RECT 255.835 149.430 256.005 150.410 ;
        RECT 273.230 150.280 273.400 151.035 ;
        RECT 273.665 150.535 276.295 150.865 ;
        RECT 274.600 150.305 274.800 150.535 ;
        RECT 276.560 150.305 276.730 151.035 ;
        RECT 297.190 151.365 297.360 151.850 ;
        RECT 297.190 151.035 298.405 151.365 ;
        RECT 298.575 151.035 299.055 151.725 ;
        RECT 300.520 151.365 300.690 151.850 ;
        RECT 299.225 151.035 300.690 151.365 ;
        RECT 273.230 149.950 274.325 150.280 ;
        RECT 274.495 149.975 274.865 150.305 ;
        RECT 275.135 149.975 278.155 150.305 ;
        RECT 278.425 149.975 278.795 150.305 ;
        RECT 250.440 149.075 250.810 149.405 ;
        RECT 251.080 149.075 254.100 149.405 ;
        RECT 254.370 149.075 254.740 149.405 ;
        RECT 254.910 149.100 256.005 149.430 ;
        RECT 249.175 148.155 250.390 148.485 ;
        RECT 250.560 148.155 251.040 148.845 ;
        RECT 252.505 148.485 252.675 149.075 ;
        RECT 251.210 148.155 253.970 148.485 ;
        RECT 254.140 148.155 254.620 148.845 ;
        RECT 255.835 148.485 256.005 149.100 ;
        RECT 254.790 148.155 256.005 148.485 ;
        RECT 249.175 147.440 249.345 148.155 ;
        RECT 249.610 147.655 252.240 147.985 ;
        RECT 249.175 147.140 250.365 147.440 ;
        RECT 249.175 146.565 249.345 147.140 ;
        RECT 250.625 146.925 250.825 147.655 ;
        RECT 252.505 147.440 252.675 148.155 ;
        RECT 252.940 147.655 255.570 147.985 ;
        RECT 251.465 147.140 253.715 147.440 ;
        RECT 249.175 146.235 250.390 146.565 ;
        RECT 250.560 146.235 251.040 146.925 ;
        RECT 252.505 146.565 252.675 147.140 ;
        RECT 254.355 146.925 254.555 147.655 ;
        RECT 255.835 147.440 256.005 148.155 ;
        RECT 254.815 147.140 256.005 147.440 ;
        RECT 251.210 146.235 253.970 146.565 ;
        RECT 254.140 146.235 254.620 146.925 ;
        RECT 255.835 146.565 256.005 147.140 ;
        RECT 254.790 146.235 256.005 146.565 ;
        RECT 249.175 145.495 249.345 146.235 ;
        RECT 249.610 145.735 252.240 146.065 ;
        RECT 249.175 145.165 250.390 145.495 ;
        RECT 250.675 145.485 250.875 145.735 ;
        RECT 249.175 144.565 249.345 145.165 ;
        RECT 249.610 144.745 250.440 144.995 ;
        RECT 249.175 144.235 250.100 144.565 ;
        RECT 237.955 139.830 240.055 140.000 ;
        RECT 240.415 143.660 244.445 143.830 ;
        RECT 235.495 134.085 237.595 134.255 ;
        RECT 237.955 139.300 240.055 139.470 ;
        RECT 237.955 134.250 238.125 139.300 ;
        RECT 238.755 138.790 239.255 138.960 ;
        RECT 238.525 138.080 238.695 138.620 ;
        RECT 239.315 138.080 239.485 138.620 ;
        RECT 238.755 137.740 239.255 137.910 ;
        RECT 238.525 137.030 238.695 137.570 ;
        RECT 239.315 137.030 239.485 137.570 ;
        RECT 238.755 136.690 239.255 136.860 ;
        RECT 238.525 135.980 238.695 136.520 ;
        RECT 239.315 135.980 239.485 136.520 ;
        RECT 238.755 135.640 239.255 135.810 ;
        RECT 238.525 134.930 238.695 135.470 ;
        RECT 239.315 134.930 239.485 135.470 ;
        RECT 238.755 134.590 239.255 134.760 ;
        RECT 239.885 134.250 240.055 139.300 ;
        RECT 237.955 134.080 240.055 134.250 ;
        RECT 240.415 134.250 240.585 143.660 ;
        RECT 241.215 143.150 241.715 143.320 ;
        RECT 240.985 141.395 241.155 142.935 ;
        RECT 241.775 141.395 241.945 142.935 ;
        RECT 241.215 141.010 241.715 141.180 ;
        RECT 240.985 139.255 241.155 140.795 ;
        RECT 241.775 139.255 241.945 140.795 ;
        RECT 241.215 138.870 241.715 139.040 ;
        RECT 240.985 137.115 241.155 138.655 ;
        RECT 241.775 137.115 241.945 138.655 ;
        RECT 241.215 136.730 241.715 136.900 ;
        RECT 240.985 134.975 241.155 136.515 ;
        RECT 241.775 134.975 241.945 136.515 ;
        RECT 241.215 134.590 241.715 134.760 ;
        RECT 242.345 134.250 242.515 143.660 ;
        RECT 243.145 143.150 243.645 143.320 ;
        RECT 242.915 141.395 243.085 142.935 ;
        RECT 243.705 141.395 243.875 142.935 ;
        RECT 243.145 141.010 243.645 141.180 ;
        RECT 242.915 139.255 243.085 140.795 ;
        RECT 243.705 139.255 243.875 140.795 ;
        RECT 243.145 138.870 243.645 139.040 ;
        RECT 242.915 137.115 243.085 138.655 ;
        RECT 243.705 137.115 243.875 138.655 ;
        RECT 243.145 136.730 243.645 136.900 ;
        RECT 242.915 134.975 243.085 136.515 ;
        RECT 243.705 134.975 243.875 136.515 ;
        RECT 243.145 134.590 243.645 134.760 ;
        RECT 244.275 134.250 244.445 143.660 ;
        RECT 249.175 143.655 249.345 144.235 ;
        RECT 250.270 144.005 250.440 144.745 ;
        RECT 249.610 143.835 250.440 144.005 ;
        RECT 249.175 143.325 250.100 143.655 ;
        RECT 250.270 143.565 250.440 143.835 ;
        RECT 250.610 143.810 251.040 145.485 ;
        RECT 252.505 145.460 252.675 146.235 ;
        RECT 252.940 145.735 255.570 146.065 ;
        RECT 254.305 145.485 254.505 145.735 ;
        RECT 255.835 145.495 256.005 146.235 ;
        RECT 251.210 145.210 253.970 145.460 ;
        RECT 251.210 144.680 252.240 145.010 ;
        RECT 251.210 144.110 251.380 144.680 ;
        RECT 252.505 144.480 252.675 145.210 ;
        RECT 252.940 144.680 253.970 145.010 ;
        RECT 251.550 144.310 253.630 144.480 ;
        RECT 251.210 143.780 252.240 144.110 ;
        RECT 251.210 143.565 251.380 143.780 ;
        RECT 252.505 143.580 252.675 144.310 ;
        RECT 253.800 144.110 253.970 144.680 ;
        RECT 252.940 143.780 253.970 144.110 ;
        RECT 254.140 143.810 254.570 145.485 ;
        RECT 254.790 145.165 256.005 145.495 ;
        RECT 254.740 144.745 255.570 144.995 ;
        RECT 254.740 144.005 254.910 144.745 ;
        RECT 255.835 144.565 256.005 145.165 ;
        RECT 255.080 144.235 256.005 144.565 ;
        RECT 254.740 143.835 255.570 144.005 ;
        RECT 250.270 143.335 251.380 143.565 ;
        RECT 249.175 143.120 249.345 143.325 ;
        RECT 249.175 142.820 250.365 143.120 ;
        RECT 249.175 142.600 249.345 142.820 ;
        RECT 249.175 142.350 250.390 142.600 ;
        RECT 249.175 141.740 249.345 142.350 ;
        RECT 250.675 142.170 250.875 143.335 ;
        RECT 251.550 143.330 253.630 143.580 ;
        RECT 253.800 143.565 253.970 143.780 ;
        RECT 254.740 143.565 254.910 143.835 ;
        RECT 255.835 143.655 256.005 144.235 ;
        RECT 253.800 143.335 254.910 143.565 ;
        RECT 252.505 143.120 252.675 143.330 ;
        RECT 251.465 142.820 253.715 143.120 ;
        RECT 252.505 142.615 252.675 142.820 ;
        RECT 251.080 142.365 254.100 142.615 ;
        RECT 249.610 141.920 250.440 142.170 ;
        RECT 249.175 141.410 250.100 141.740 ;
        RECT 249.175 140.880 249.345 141.410 ;
        RECT 250.270 141.230 250.440 141.920 ;
        RECT 249.610 141.060 250.440 141.230 ;
        RECT 249.175 140.550 250.100 140.880 ;
        RECT 249.175 139.880 249.345 140.550 ;
        RECT 250.270 140.380 250.440 141.060 ;
        RECT 250.610 140.480 251.040 142.170 ;
        RECT 251.210 141.915 252.240 142.165 ;
        RECT 251.210 141.215 251.380 141.915 ;
        RECT 252.505 141.715 252.675 142.365 ;
        RECT 254.310 142.170 254.510 143.335 ;
        RECT 255.080 143.325 256.005 143.655 ;
        RECT 255.835 143.120 256.005 143.325 ;
        RECT 254.815 142.820 256.005 143.120 ;
        RECT 255.835 142.600 256.005 142.820 ;
        RECT 254.790 142.350 256.005 142.600 ;
        RECT 252.940 141.915 253.970 142.165 ;
        RECT 251.550 141.385 253.630 141.715 ;
        RECT 251.210 140.885 252.240 141.215 ;
        RECT 249.610 140.310 250.440 140.380 ;
        RECT 249.610 140.235 250.570 140.310 ;
        RECT 251.210 140.235 251.380 140.885 ;
        RECT 252.505 140.685 252.675 141.385 ;
        RECT 253.800 141.215 253.970 141.915 ;
        RECT 252.940 140.885 253.970 141.215 ;
        RECT 251.550 140.435 253.630 140.685 ;
        RECT 249.610 140.065 252.240 140.235 ;
        RECT 249.610 140.050 250.880 140.065 ;
        RECT 249.175 139.550 250.230 139.880 ;
        RECT 240.415 134.080 244.445 134.250 ;
        RECT 244.805 139.300 248.835 139.470 ;
        RECT 244.805 134.250 244.975 139.300 ;
        RECT 245.605 138.790 246.105 138.960 ;
        RECT 245.375 138.080 245.545 138.620 ;
        RECT 246.165 138.080 246.335 138.620 ;
        RECT 245.605 137.740 246.105 137.910 ;
        RECT 245.375 137.030 245.545 137.570 ;
        RECT 246.165 137.030 246.335 137.570 ;
        RECT 245.605 136.690 246.105 136.860 ;
        RECT 245.375 135.980 245.545 136.520 ;
        RECT 246.165 135.980 246.335 136.520 ;
        RECT 245.605 135.640 246.105 135.810 ;
        RECT 245.375 134.930 245.545 135.470 ;
        RECT 246.165 134.930 246.335 135.470 ;
        RECT 245.605 134.590 246.105 134.760 ;
        RECT 246.735 134.250 246.905 139.300 ;
        RECT 247.535 138.790 248.035 138.960 ;
        RECT 247.305 138.080 247.475 138.620 ;
        RECT 248.095 138.080 248.265 138.620 ;
        RECT 247.535 137.740 248.035 137.910 ;
        RECT 247.305 137.030 247.475 137.570 ;
        RECT 248.095 137.030 248.265 137.570 ;
        RECT 247.535 136.690 248.035 136.860 ;
        RECT 247.305 135.980 247.475 136.520 ;
        RECT 248.095 135.980 248.265 136.520 ;
        RECT 247.535 135.640 248.035 135.810 ;
        RECT 247.305 134.930 247.475 135.470 ;
        RECT 248.095 134.930 248.265 135.470 ;
        RECT 247.535 134.590 248.035 134.760 ;
        RECT 248.665 134.250 248.835 139.300 ;
        RECT 244.805 134.080 248.835 134.250 ;
        RECT 249.175 138.950 249.345 139.550 ;
        RECT 250.400 139.380 250.880 140.050 ;
        RECT 252.505 139.865 252.675 140.435 ;
        RECT 253.800 140.235 253.970 140.885 ;
        RECT 254.140 140.480 254.570 142.170 ;
        RECT 254.740 141.920 255.570 142.170 ;
        RECT 254.740 141.230 254.910 141.920 ;
        RECT 255.835 141.740 256.005 142.350 ;
        RECT 255.080 141.410 256.005 141.740 ;
        RECT 254.740 141.060 255.570 141.230 ;
        RECT 254.740 140.380 254.910 141.060 ;
        RECT 255.835 140.880 256.005 141.410 ;
        RECT 255.080 140.550 256.005 140.880 ;
        RECT 254.740 140.310 255.570 140.380 ;
        RECT 254.610 140.235 255.570 140.310 ;
        RECT 252.940 140.065 255.570 140.235 ;
        RECT 254.300 140.050 255.570 140.065 ;
        RECT 251.080 139.535 254.100 139.865 ;
        RECT 249.610 139.365 250.880 139.380 ;
        RECT 249.610 139.120 252.240 139.365 ;
        RECT 250.400 139.035 252.240 139.120 ;
        RECT 249.175 138.620 250.230 138.950 ;
        RECT 249.175 138.280 249.345 138.620 ;
        RECT 250.400 138.535 250.880 139.035 ;
        RECT 252.505 138.865 252.675 139.535 ;
        RECT 254.300 139.380 254.780 140.050 ;
        RECT 255.835 139.880 256.005 140.550 ;
        RECT 254.950 139.550 256.005 139.880 ;
        RECT 257.090 149.415 259.190 149.585 ;
        RECT 257.090 140.005 257.260 149.415 ;
        RECT 257.890 148.905 258.390 149.075 ;
        RECT 257.660 147.150 257.830 148.690 ;
        RECT 258.450 147.150 258.620 148.690 ;
        RECT 257.890 146.765 258.390 146.935 ;
        RECT 257.660 145.010 257.830 146.550 ;
        RECT 258.450 145.010 258.620 146.550 ;
        RECT 257.890 144.625 258.390 144.795 ;
        RECT 257.660 142.870 257.830 144.410 ;
        RECT 258.450 142.870 258.620 144.410 ;
        RECT 257.890 142.485 258.390 142.655 ;
        RECT 257.660 140.730 257.830 142.270 ;
        RECT 258.450 140.730 258.620 142.270 ;
        RECT 257.890 140.345 258.390 140.515 ;
        RECT 259.020 140.005 259.190 149.415 ;
        RECT 259.550 149.415 261.650 149.585 ;
        RECT 259.550 144.365 259.720 149.415 ;
        RECT 260.350 148.905 260.850 149.075 ;
        RECT 260.120 148.195 260.290 148.735 ;
        RECT 260.910 148.195 261.080 148.735 ;
        RECT 260.350 147.855 260.850 148.025 ;
        RECT 260.120 147.145 260.290 147.685 ;
        RECT 260.910 147.145 261.080 147.685 ;
        RECT 260.350 146.805 260.850 146.975 ;
        RECT 260.120 146.095 260.290 146.635 ;
        RECT 260.910 146.095 261.080 146.635 ;
        RECT 260.350 145.755 260.850 145.925 ;
        RECT 260.120 145.045 260.290 145.585 ;
        RECT 260.910 145.045 261.080 145.585 ;
        RECT 260.350 144.705 260.850 144.875 ;
        RECT 261.480 144.365 261.650 149.415 ;
        RECT 259.550 144.195 261.650 144.365 ;
        RECT 262.010 149.410 264.110 149.580 ;
        RECT 257.090 139.835 259.190 140.005 ;
        RECT 259.550 143.665 261.650 143.835 ;
        RECT 254.300 139.365 255.570 139.380 ;
        RECT 252.940 139.120 255.570 139.365 ;
        RECT 252.940 139.035 254.780 139.120 ;
        RECT 251.080 138.535 254.100 138.865 ;
        RECT 254.300 138.535 254.780 139.035 ;
        RECT 255.835 138.950 256.005 139.550 ;
        RECT 254.950 138.620 256.005 138.950 ;
        RECT 249.175 138.030 250.390 138.280 ;
        RECT 249.175 137.420 249.345 138.030 ;
        RECT 250.675 137.850 250.875 138.535 ;
        RECT 252.505 138.295 252.675 138.535 ;
        RECT 251.080 138.045 254.100 138.295 ;
        RECT 249.610 137.600 250.440 137.850 ;
        RECT 249.175 137.090 250.100 137.420 ;
        RECT 249.175 136.560 249.345 137.090 ;
        RECT 250.270 136.910 250.440 137.600 ;
        RECT 249.610 136.740 250.440 136.910 ;
        RECT 249.175 136.230 250.100 136.560 ;
        RECT 249.175 135.560 249.345 136.230 ;
        RECT 250.270 136.060 250.440 136.740 ;
        RECT 250.610 136.160 251.040 137.850 ;
        RECT 251.210 137.595 252.240 137.845 ;
        RECT 251.210 136.895 251.380 137.595 ;
        RECT 252.505 137.395 252.675 138.045 ;
        RECT 254.305 137.850 254.505 138.535 ;
        RECT 255.835 138.280 256.005 138.620 ;
        RECT 254.790 138.030 256.005 138.280 ;
        RECT 252.940 137.595 253.970 137.845 ;
        RECT 251.550 137.065 253.630 137.395 ;
        RECT 251.210 136.565 252.240 136.895 ;
        RECT 249.610 135.990 250.440 136.060 ;
        RECT 249.610 135.915 250.570 135.990 ;
        RECT 251.210 135.915 251.380 136.565 ;
        RECT 252.505 136.365 252.675 137.065 ;
        RECT 253.800 136.895 253.970 137.595 ;
        RECT 252.940 136.565 253.970 136.895 ;
        RECT 251.550 136.115 253.630 136.365 ;
        RECT 249.610 135.745 252.240 135.915 ;
        RECT 249.610 135.730 250.880 135.745 ;
        RECT 249.175 135.230 250.230 135.560 ;
        RECT 249.175 134.630 249.345 135.230 ;
        RECT 250.400 135.060 250.880 135.730 ;
        RECT 252.505 135.545 252.675 136.115 ;
        RECT 253.800 135.915 253.970 136.565 ;
        RECT 254.140 136.160 254.570 137.850 ;
        RECT 254.740 137.600 255.570 137.850 ;
        RECT 254.740 136.910 254.910 137.600 ;
        RECT 255.835 137.420 256.005 138.030 ;
        RECT 255.080 137.090 256.005 137.420 ;
        RECT 254.740 136.740 255.570 136.910 ;
        RECT 254.740 136.060 254.910 136.740 ;
        RECT 255.835 136.560 256.005 137.090 ;
        RECT 255.080 136.230 256.005 136.560 ;
        RECT 254.740 135.990 255.570 136.060 ;
        RECT 254.610 135.915 255.570 135.990 ;
        RECT 252.940 135.745 255.570 135.915 ;
        RECT 254.300 135.730 255.570 135.745 ;
        RECT 251.080 135.215 254.100 135.545 ;
        RECT 249.610 135.045 250.880 135.060 ;
        RECT 249.610 134.800 252.240 135.045 ;
        RECT 250.400 134.715 252.240 134.800 ;
        RECT 249.175 134.300 250.230 134.630 ;
        RECT 249.175 134.090 249.345 134.300 ;
        RECT 250.400 134.215 250.880 134.715 ;
        RECT 252.505 134.545 252.675 135.215 ;
        RECT 254.300 135.060 254.780 135.730 ;
        RECT 255.835 135.560 256.005 136.230 ;
        RECT 254.950 135.230 256.005 135.560 ;
        RECT 254.300 135.045 255.570 135.060 ;
        RECT 252.940 134.800 255.570 135.045 ;
        RECT 252.940 134.715 254.780 134.800 ;
        RECT 251.080 134.215 254.100 134.545 ;
        RECT 254.300 134.215 254.780 134.715 ;
        RECT 255.835 134.630 256.005 135.230 ;
        RECT 254.950 134.300 256.005 134.630 ;
        RECT 252.505 134.090 252.675 134.215 ;
        RECT 255.835 134.090 256.005 134.300 ;
        RECT 257.090 139.305 259.190 139.475 ;
        RECT 257.090 134.255 257.260 139.305 ;
        RECT 257.890 138.795 258.390 138.965 ;
        RECT 257.660 138.085 257.830 138.625 ;
        RECT 258.450 138.085 258.620 138.625 ;
        RECT 257.890 137.745 258.390 137.915 ;
        RECT 257.660 137.035 257.830 137.575 ;
        RECT 258.450 137.035 258.620 137.575 ;
        RECT 257.890 136.695 258.390 136.865 ;
        RECT 257.660 135.985 257.830 136.525 ;
        RECT 258.450 135.985 258.620 136.525 ;
        RECT 257.890 135.645 258.390 135.815 ;
        RECT 257.660 134.935 257.830 135.475 ;
        RECT 258.450 134.935 258.620 135.475 ;
        RECT 257.890 134.595 258.390 134.765 ;
        RECT 259.020 134.255 259.190 139.305 ;
        RECT 257.090 134.085 259.190 134.255 ;
        RECT 259.550 134.255 259.720 143.665 ;
        RECT 260.350 143.155 260.850 143.325 ;
        RECT 260.120 141.400 260.290 142.940 ;
        RECT 260.910 141.400 261.080 142.940 ;
        RECT 260.350 141.015 260.850 141.185 ;
        RECT 260.120 139.260 260.290 140.800 ;
        RECT 260.910 139.260 261.080 140.800 ;
        RECT 260.350 138.875 260.850 139.045 ;
        RECT 260.120 137.120 260.290 138.660 ;
        RECT 260.910 137.120 261.080 138.660 ;
        RECT 260.350 136.735 260.850 136.905 ;
        RECT 260.120 134.980 260.290 136.520 ;
        RECT 260.910 134.980 261.080 136.520 ;
        RECT 260.350 134.595 260.850 134.765 ;
        RECT 261.480 134.255 261.650 143.665 ;
        RECT 262.010 140.000 262.180 149.410 ;
        RECT 262.810 148.900 263.310 149.070 ;
        RECT 262.580 147.145 262.750 148.685 ;
        RECT 263.370 147.145 263.540 148.685 ;
        RECT 262.810 146.760 263.310 146.930 ;
        RECT 262.580 145.005 262.750 146.545 ;
        RECT 263.370 145.005 263.540 146.545 ;
        RECT 262.810 144.620 263.310 144.790 ;
        RECT 262.580 142.865 262.750 144.405 ;
        RECT 263.370 142.865 263.540 144.405 ;
        RECT 262.810 142.480 263.310 142.650 ;
        RECT 262.580 140.725 262.750 142.265 ;
        RECT 263.370 140.725 263.540 142.265 ;
        RECT 262.810 140.340 263.310 140.510 ;
        RECT 263.940 140.000 264.110 149.410 ;
        RECT 273.230 148.485 273.400 149.950 ;
        RECT 274.495 149.745 276.295 149.805 ;
        RECT 274.155 149.575 276.295 149.745 ;
        RECT 274.155 149.460 274.325 149.575 ;
        RECT 273.665 149.130 274.325 149.460 ;
        RECT 276.560 149.405 276.730 149.975 ;
        RECT 278.965 149.920 279.625 150.250 ;
        RECT 278.965 149.805 279.135 149.920 ;
        RECT 276.995 149.635 279.135 149.805 ;
        RECT 276.995 149.575 278.795 149.635 ;
        RECT 279.890 149.430 280.060 150.410 ;
        RECT 297.190 150.280 297.360 151.035 ;
        RECT 297.625 150.535 300.255 150.865 ;
        RECT 298.560 150.305 298.760 150.535 ;
        RECT 300.520 150.305 300.690 151.035 ;
        RECT 321.200 151.365 321.370 151.850 ;
        RECT 321.200 151.035 322.415 151.365 ;
        RECT 322.585 151.035 323.065 151.725 ;
        RECT 324.530 151.365 324.700 151.850 ;
        RECT 323.235 151.035 324.700 151.365 ;
        RECT 297.190 149.950 298.285 150.280 ;
        RECT 298.455 149.975 298.825 150.305 ;
        RECT 299.095 149.975 302.115 150.305 ;
        RECT 302.385 149.975 302.755 150.305 ;
        RECT 274.495 149.075 274.865 149.405 ;
        RECT 275.135 149.075 278.155 149.405 ;
        RECT 278.425 149.075 278.795 149.405 ;
        RECT 278.965 149.100 280.060 149.430 ;
        RECT 273.230 148.155 274.445 148.485 ;
        RECT 274.615 148.155 275.095 148.845 ;
        RECT 276.560 148.485 276.730 149.075 ;
        RECT 275.265 148.155 278.025 148.485 ;
        RECT 278.195 148.155 278.675 148.845 ;
        RECT 279.890 148.485 280.060 149.100 ;
        RECT 278.845 148.155 280.060 148.485 ;
        RECT 273.230 147.440 273.400 148.155 ;
        RECT 273.665 147.655 276.295 147.985 ;
        RECT 273.230 147.140 274.420 147.440 ;
        RECT 273.230 146.565 273.400 147.140 ;
        RECT 274.680 146.925 274.880 147.655 ;
        RECT 276.560 147.440 276.730 148.155 ;
        RECT 276.995 147.655 279.625 147.985 ;
        RECT 275.520 147.140 277.770 147.440 ;
        RECT 273.230 146.235 274.445 146.565 ;
        RECT 274.615 146.235 275.095 146.925 ;
        RECT 276.560 146.565 276.730 147.140 ;
        RECT 278.410 146.925 278.610 147.655 ;
        RECT 279.890 147.440 280.060 148.155 ;
        RECT 278.870 147.140 280.060 147.440 ;
        RECT 275.265 146.235 278.025 146.565 ;
        RECT 278.195 146.235 278.675 146.925 ;
        RECT 279.890 146.565 280.060 147.140 ;
        RECT 278.845 146.235 280.060 146.565 ;
        RECT 273.230 145.495 273.400 146.235 ;
        RECT 273.665 145.735 276.295 146.065 ;
        RECT 273.230 145.165 274.445 145.495 ;
        RECT 274.730 145.485 274.930 145.735 ;
        RECT 273.230 144.565 273.400 145.165 ;
        RECT 273.665 144.745 274.495 144.995 ;
        RECT 273.230 144.235 274.155 144.565 ;
        RECT 262.010 139.830 264.110 140.000 ;
        RECT 264.470 143.660 268.500 143.830 ;
        RECT 259.550 134.085 261.650 134.255 ;
        RECT 262.010 139.300 264.110 139.470 ;
        RECT 262.010 134.250 262.180 139.300 ;
        RECT 262.810 138.790 263.310 138.960 ;
        RECT 262.580 138.080 262.750 138.620 ;
        RECT 263.370 138.080 263.540 138.620 ;
        RECT 262.810 137.740 263.310 137.910 ;
        RECT 262.580 137.030 262.750 137.570 ;
        RECT 263.370 137.030 263.540 137.570 ;
        RECT 262.810 136.690 263.310 136.860 ;
        RECT 262.580 135.980 262.750 136.520 ;
        RECT 263.370 135.980 263.540 136.520 ;
        RECT 262.810 135.640 263.310 135.810 ;
        RECT 262.580 134.930 262.750 135.470 ;
        RECT 263.370 134.930 263.540 135.470 ;
        RECT 262.810 134.590 263.310 134.760 ;
        RECT 263.940 134.250 264.110 139.300 ;
        RECT 262.010 134.080 264.110 134.250 ;
        RECT 264.470 134.250 264.640 143.660 ;
        RECT 265.270 143.150 265.770 143.320 ;
        RECT 265.040 141.395 265.210 142.935 ;
        RECT 265.830 141.395 266.000 142.935 ;
        RECT 265.270 141.010 265.770 141.180 ;
        RECT 265.040 139.255 265.210 140.795 ;
        RECT 265.830 139.255 266.000 140.795 ;
        RECT 265.270 138.870 265.770 139.040 ;
        RECT 265.040 137.115 265.210 138.655 ;
        RECT 265.830 137.115 266.000 138.655 ;
        RECT 265.270 136.730 265.770 136.900 ;
        RECT 265.040 134.975 265.210 136.515 ;
        RECT 265.830 134.975 266.000 136.515 ;
        RECT 265.270 134.590 265.770 134.760 ;
        RECT 266.400 134.250 266.570 143.660 ;
        RECT 267.200 143.150 267.700 143.320 ;
        RECT 266.970 141.395 267.140 142.935 ;
        RECT 267.760 141.395 267.930 142.935 ;
        RECT 267.200 141.010 267.700 141.180 ;
        RECT 266.970 139.255 267.140 140.795 ;
        RECT 267.760 139.255 267.930 140.795 ;
        RECT 267.200 138.870 267.700 139.040 ;
        RECT 266.970 137.115 267.140 138.655 ;
        RECT 267.760 137.115 267.930 138.655 ;
        RECT 267.200 136.730 267.700 136.900 ;
        RECT 266.970 134.975 267.140 136.515 ;
        RECT 267.760 134.975 267.930 136.515 ;
        RECT 267.200 134.590 267.700 134.760 ;
        RECT 268.330 134.250 268.500 143.660 ;
        RECT 273.230 143.655 273.400 144.235 ;
        RECT 274.325 144.005 274.495 144.745 ;
        RECT 273.665 143.835 274.495 144.005 ;
        RECT 273.230 143.325 274.155 143.655 ;
        RECT 274.325 143.565 274.495 143.835 ;
        RECT 274.665 143.810 275.095 145.485 ;
        RECT 276.560 145.460 276.730 146.235 ;
        RECT 276.995 145.735 279.625 146.065 ;
        RECT 278.360 145.485 278.560 145.735 ;
        RECT 279.890 145.495 280.060 146.235 ;
        RECT 275.265 145.210 278.025 145.460 ;
        RECT 275.265 144.680 276.295 145.010 ;
        RECT 275.265 144.110 275.435 144.680 ;
        RECT 276.560 144.480 276.730 145.210 ;
        RECT 276.995 144.680 278.025 145.010 ;
        RECT 275.605 144.310 277.685 144.480 ;
        RECT 275.265 143.780 276.295 144.110 ;
        RECT 275.265 143.565 275.435 143.780 ;
        RECT 276.560 143.580 276.730 144.310 ;
        RECT 277.855 144.110 278.025 144.680 ;
        RECT 276.995 143.780 278.025 144.110 ;
        RECT 278.195 143.810 278.625 145.485 ;
        RECT 278.845 145.165 280.060 145.495 ;
        RECT 278.795 144.745 279.625 144.995 ;
        RECT 278.795 144.005 278.965 144.745 ;
        RECT 279.890 144.565 280.060 145.165 ;
        RECT 279.135 144.235 280.060 144.565 ;
        RECT 278.795 143.835 279.625 144.005 ;
        RECT 274.325 143.335 275.435 143.565 ;
        RECT 273.230 143.120 273.400 143.325 ;
        RECT 273.230 142.820 274.420 143.120 ;
        RECT 273.230 142.600 273.400 142.820 ;
        RECT 273.230 142.350 274.445 142.600 ;
        RECT 273.230 141.740 273.400 142.350 ;
        RECT 274.730 142.170 274.930 143.335 ;
        RECT 275.605 143.330 277.685 143.580 ;
        RECT 277.855 143.565 278.025 143.780 ;
        RECT 278.795 143.565 278.965 143.835 ;
        RECT 279.890 143.655 280.060 144.235 ;
        RECT 277.855 143.335 278.965 143.565 ;
        RECT 276.560 143.120 276.730 143.330 ;
        RECT 275.520 142.820 277.770 143.120 ;
        RECT 276.560 142.615 276.730 142.820 ;
        RECT 275.135 142.365 278.155 142.615 ;
        RECT 273.665 141.920 274.495 142.170 ;
        RECT 273.230 141.410 274.155 141.740 ;
        RECT 273.230 140.880 273.400 141.410 ;
        RECT 274.325 141.230 274.495 141.920 ;
        RECT 273.665 141.060 274.495 141.230 ;
        RECT 273.230 140.550 274.155 140.880 ;
        RECT 273.230 139.880 273.400 140.550 ;
        RECT 274.325 140.380 274.495 141.060 ;
        RECT 274.665 140.480 275.095 142.170 ;
        RECT 275.265 141.915 276.295 142.165 ;
        RECT 275.265 141.215 275.435 141.915 ;
        RECT 276.560 141.715 276.730 142.365 ;
        RECT 278.365 142.170 278.565 143.335 ;
        RECT 279.135 143.325 280.060 143.655 ;
        RECT 279.890 143.120 280.060 143.325 ;
        RECT 278.870 142.820 280.060 143.120 ;
        RECT 279.890 142.600 280.060 142.820 ;
        RECT 278.845 142.350 280.060 142.600 ;
        RECT 276.995 141.915 278.025 142.165 ;
        RECT 275.605 141.385 277.685 141.715 ;
        RECT 275.265 140.885 276.295 141.215 ;
        RECT 273.665 140.310 274.495 140.380 ;
        RECT 273.665 140.235 274.625 140.310 ;
        RECT 275.265 140.235 275.435 140.885 ;
        RECT 276.560 140.685 276.730 141.385 ;
        RECT 277.855 141.215 278.025 141.915 ;
        RECT 276.995 140.885 278.025 141.215 ;
        RECT 275.605 140.435 277.685 140.685 ;
        RECT 273.665 140.065 276.295 140.235 ;
        RECT 273.665 140.050 274.935 140.065 ;
        RECT 273.230 139.550 274.285 139.880 ;
        RECT 264.470 134.080 268.500 134.250 ;
        RECT 268.860 139.300 272.890 139.470 ;
        RECT 268.860 134.250 269.030 139.300 ;
        RECT 269.660 138.790 270.160 138.960 ;
        RECT 269.430 138.080 269.600 138.620 ;
        RECT 270.220 138.080 270.390 138.620 ;
        RECT 269.660 137.740 270.160 137.910 ;
        RECT 269.430 137.030 269.600 137.570 ;
        RECT 270.220 137.030 270.390 137.570 ;
        RECT 269.660 136.690 270.160 136.860 ;
        RECT 269.430 135.980 269.600 136.520 ;
        RECT 270.220 135.980 270.390 136.520 ;
        RECT 269.660 135.640 270.160 135.810 ;
        RECT 269.430 134.930 269.600 135.470 ;
        RECT 270.220 134.930 270.390 135.470 ;
        RECT 269.660 134.590 270.160 134.760 ;
        RECT 270.790 134.250 270.960 139.300 ;
        RECT 271.590 138.790 272.090 138.960 ;
        RECT 271.360 138.080 271.530 138.620 ;
        RECT 272.150 138.080 272.320 138.620 ;
        RECT 271.590 137.740 272.090 137.910 ;
        RECT 271.360 137.030 271.530 137.570 ;
        RECT 272.150 137.030 272.320 137.570 ;
        RECT 271.590 136.690 272.090 136.860 ;
        RECT 271.360 135.980 271.530 136.520 ;
        RECT 272.150 135.980 272.320 136.520 ;
        RECT 271.590 135.640 272.090 135.810 ;
        RECT 271.360 134.930 271.530 135.470 ;
        RECT 272.150 134.930 272.320 135.470 ;
        RECT 271.590 134.590 272.090 134.760 ;
        RECT 272.720 134.250 272.890 139.300 ;
        RECT 268.860 134.080 272.890 134.250 ;
        RECT 273.230 138.950 273.400 139.550 ;
        RECT 274.455 139.380 274.935 140.050 ;
        RECT 276.560 139.865 276.730 140.435 ;
        RECT 277.855 140.235 278.025 140.885 ;
        RECT 278.195 140.480 278.625 142.170 ;
        RECT 278.795 141.920 279.625 142.170 ;
        RECT 278.795 141.230 278.965 141.920 ;
        RECT 279.890 141.740 280.060 142.350 ;
        RECT 279.135 141.410 280.060 141.740 ;
        RECT 278.795 141.060 279.625 141.230 ;
        RECT 278.795 140.380 278.965 141.060 ;
        RECT 279.890 140.880 280.060 141.410 ;
        RECT 279.135 140.550 280.060 140.880 ;
        RECT 278.795 140.310 279.625 140.380 ;
        RECT 278.665 140.235 279.625 140.310 ;
        RECT 276.995 140.065 279.625 140.235 ;
        RECT 278.355 140.050 279.625 140.065 ;
        RECT 275.135 139.535 278.155 139.865 ;
        RECT 273.665 139.365 274.935 139.380 ;
        RECT 273.665 139.120 276.295 139.365 ;
        RECT 274.455 139.035 276.295 139.120 ;
        RECT 273.230 138.620 274.285 138.950 ;
        RECT 273.230 138.280 273.400 138.620 ;
        RECT 274.455 138.535 274.935 139.035 ;
        RECT 276.560 138.865 276.730 139.535 ;
        RECT 278.355 139.380 278.835 140.050 ;
        RECT 279.890 139.880 280.060 140.550 ;
        RECT 279.005 139.550 280.060 139.880 ;
        RECT 281.050 149.415 283.150 149.585 ;
        RECT 281.050 140.005 281.220 149.415 ;
        RECT 281.850 148.905 282.350 149.075 ;
        RECT 281.620 147.150 281.790 148.690 ;
        RECT 282.410 147.150 282.580 148.690 ;
        RECT 281.850 146.765 282.350 146.935 ;
        RECT 281.620 145.010 281.790 146.550 ;
        RECT 282.410 145.010 282.580 146.550 ;
        RECT 281.850 144.625 282.350 144.795 ;
        RECT 281.620 142.870 281.790 144.410 ;
        RECT 282.410 142.870 282.580 144.410 ;
        RECT 281.850 142.485 282.350 142.655 ;
        RECT 281.620 140.730 281.790 142.270 ;
        RECT 282.410 140.730 282.580 142.270 ;
        RECT 281.850 140.345 282.350 140.515 ;
        RECT 282.980 140.005 283.150 149.415 ;
        RECT 283.510 149.415 285.610 149.585 ;
        RECT 283.510 144.365 283.680 149.415 ;
        RECT 284.310 148.905 284.810 149.075 ;
        RECT 284.080 148.195 284.250 148.735 ;
        RECT 284.870 148.195 285.040 148.735 ;
        RECT 284.310 147.855 284.810 148.025 ;
        RECT 284.080 147.145 284.250 147.685 ;
        RECT 284.870 147.145 285.040 147.685 ;
        RECT 284.310 146.805 284.810 146.975 ;
        RECT 284.080 146.095 284.250 146.635 ;
        RECT 284.870 146.095 285.040 146.635 ;
        RECT 284.310 145.755 284.810 145.925 ;
        RECT 284.080 145.045 284.250 145.585 ;
        RECT 284.870 145.045 285.040 145.585 ;
        RECT 284.310 144.705 284.810 144.875 ;
        RECT 285.440 144.365 285.610 149.415 ;
        RECT 283.510 144.195 285.610 144.365 ;
        RECT 285.970 149.410 288.070 149.580 ;
        RECT 281.050 139.835 283.150 140.005 ;
        RECT 283.510 143.665 285.610 143.835 ;
        RECT 278.355 139.365 279.625 139.380 ;
        RECT 276.995 139.120 279.625 139.365 ;
        RECT 276.995 139.035 278.835 139.120 ;
        RECT 275.135 138.535 278.155 138.865 ;
        RECT 278.355 138.535 278.835 139.035 ;
        RECT 279.890 138.950 280.060 139.550 ;
        RECT 279.005 138.620 280.060 138.950 ;
        RECT 273.230 138.030 274.445 138.280 ;
        RECT 273.230 137.420 273.400 138.030 ;
        RECT 274.730 137.850 274.930 138.535 ;
        RECT 276.560 138.295 276.730 138.535 ;
        RECT 275.135 138.045 278.155 138.295 ;
        RECT 273.665 137.600 274.495 137.850 ;
        RECT 273.230 137.090 274.155 137.420 ;
        RECT 273.230 136.560 273.400 137.090 ;
        RECT 274.325 136.910 274.495 137.600 ;
        RECT 273.665 136.740 274.495 136.910 ;
        RECT 273.230 136.230 274.155 136.560 ;
        RECT 273.230 135.560 273.400 136.230 ;
        RECT 274.325 136.060 274.495 136.740 ;
        RECT 274.665 136.160 275.095 137.850 ;
        RECT 275.265 137.595 276.295 137.845 ;
        RECT 275.265 136.895 275.435 137.595 ;
        RECT 276.560 137.395 276.730 138.045 ;
        RECT 278.360 137.850 278.560 138.535 ;
        RECT 279.890 138.280 280.060 138.620 ;
        RECT 278.845 138.030 280.060 138.280 ;
        RECT 276.995 137.595 278.025 137.845 ;
        RECT 275.605 137.065 277.685 137.395 ;
        RECT 275.265 136.565 276.295 136.895 ;
        RECT 273.665 135.990 274.495 136.060 ;
        RECT 273.665 135.915 274.625 135.990 ;
        RECT 275.265 135.915 275.435 136.565 ;
        RECT 276.560 136.365 276.730 137.065 ;
        RECT 277.855 136.895 278.025 137.595 ;
        RECT 276.995 136.565 278.025 136.895 ;
        RECT 275.605 136.115 277.685 136.365 ;
        RECT 273.665 135.745 276.295 135.915 ;
        RECT 273.665 135.730 274.935 135.745 ;
        RECT 273.230 135.230 274.285 135.560 ;
        RECT 273.230 134.630 273.400 135.230 ;
        RECT 274.455 135.060 274.935 135.730 ;
        RECT 276.560 135.545 276.730 136.115 ;
        RECT 277.855 135.915 278.025 136.565 ;
        RECT 278.195 136.160 278.625 137.850 ;
        RECT 278.795 137.600 279.625 137.850 ;
        RECT 278.795 136.910 278.965 137.600 ;
        RECT 279.890 137.420 280.060 138.030 ;
        RECT 279.135 137.090 280.060 137.420 ;
        RECT 278.795 136.740 279.625 136.910 ;
        RECT 278.795 136.060 278.965 136.740 ;
        RECT 279.890 136.560 280.060 137.090 ;
        RECT 279.135 136.230 280.060 136.560 ;
        RECT 278.795 135.990 279.625 136.060 ;
        RECT 278.665 135.915 279.625 135.990 ;
        RECT 276.995 135.745 279.625 135.915 ;
        RECT 278.355 135.730 279.625 135.745 ;
        RECT 275.135 135.215 278.155 135.545 ;
        RECT 273.665 135.045 274.935 135.060 ;
        RECT 273.665 134.800 276.295 135.045 ;
        RECT 274.455 134.715 276.295 134.800 ;
        RECT 273.230 134.300 274.285 134.630 ;
        RECT 273.230 134.090 273.400 134.300 ;
        RECT 274.455 134.215 274.935 134.715 ;
        RECT 276.560 134.545 276.730 135.215 ;
        RECT 278.355 135.060 278.835 135.730 ;
        RECT 279.890 135.560 280.060 136.230 ;
        RECT 279.005 135.230 280.060 135.560 ;
        RECT 278.355 135.045 279.625 135.060 ;
        RECT 276.995 134.800 279.625 135.045 ;
        RECT 276.995 134.715 278.835 134.800 ;
        RECT 275.135 134.215 278.155 134.545 ;
        RECT 278.355 134.215 278.835 134.715 ;
        RECT 279.890 134.630 280.060 135.230 ;
        RECT 279.005 134.300 280.060 134.630 ;
        RECT 276.560 134.090 276.730 134.215 ;
        RECT 279.890 134.090 280.060 134.300 ;
        RECT 281.050 139.305 283.150 139.475 ;
        RECT 281.050 134.255 281.220 139.305 ;
        RECT 281.850 138.795 282.350 138.965 ;
        RECT 281.620 138.085 281.790 138.625 ;
        RECT 282.410 138.085 282.580 138.625 ;
        RECT 281.850 137.745 282.350 137.915 ;
        RECT 281.620 137.035 281.790 137.575 ;
        RECT 282.410 137.035 282.580 137.575 ;
        RECT 281.850 136.695 282.350 136.865 ;
        RECT 281.620 135.985 281.790 136.525 ;
        RECT 282.410 135.985 282.580 136.525 ;
        RECT 281.850 135.645 282.350 135.815 ;
        RECT 281.620 134.935 281.790 135.475 ;
        RECT 282.410 134.935 282.580 135.475 ;
        RECT 281.850 134.595 282.350 134.765 ;
        RECT 282.980 134.255 283.150 139.305 ;
        RECT 281.050 134.085 283.150 134.255 ;
        RECT 283.510 134.255 283.680 143.665 ;
        RECT 284.310 143.155 284.810 143.325 ;
        RECT 284.080 141.400 284.250 142.940 ;
        RECT 284.870 141.400 285.040 142.940 ;
        RECT 284.310 141.015 284.810 141.185 ;
        RECT 284.080 139.260 284.250 140.800 ;
        RECT 284.870 139.260 285.040 140.800 ;
        RECT 284.310 138.875 284.810 139.045 ;
        RECT 284.080 137.120 284.250 138.660 ;
        RECT 284.870 137.120 285.040 138.660 ;
        RECT 284.310 136.735 284.810 136.905 ;
        RECT 284.080 134.980 284.250 136.520 ;
        RECT 284.870 134.980 285.040 136.520 ;
        RECT 284.310 134.595 284.810 134.765 ;
        RECT 285.440 134.255 285.610 143.665 ;
        RECT 285.970 140.000 286.140 149.410 ;
        RECT 286.770 148.900 287.270 149.070 ;
        RECT 286.540 147.145 286.710 148.685 ;
        RECT 287.330 147.145 287.500 148.685 ;
        RECT 286.770 146.760 287.270 146.930 ;
        RECT 286.540 145.005 286.710 146.545 ;
        RECT 287.330 145.005 287.500 146.545 ;
        RECT 286.770 144.620 287.270 144.790 ;
        RECT 286.540 142.865 286.710 144.405 ;
        RECT 287.330 142.865 287.500 144.405 ;
        RECT 286.770 142.480 287.270 142.650 ;
        RECT 286.540 140.725 286.710 142.265 ;
        RECT 287.330 140.725 287.500 142.265 ;
        RECT 286.770 140.340 287.270 140.510 ;
        RECT 287.900 140.000 288.070 149.410 ;
        RECT 297.190 148.485 297.360 149.950 ;
        RECT 298.455 149.745 300.255 149.805 ;
        RECT 298.115 149.575 300.255 149.745 ;
        RECT 298.115 149.460 298.285 149.575 ;
        RECT 297.625 149.130 298.285 149.460 ;
        RECT 300.520 149.405 300.690 149.975 ;
        RECT 302.925 149.920 303.585 150.250 ;
        RECT 302.925 149.805 303.095 149.920 ;
        RECT 300.955 149.635 303.095 149.805 ;
        RECT 300.955 149.575 302.755 149.635 ;
        RECT 303.850 149.430 304.020 150.410 ;
        RECT 321.200 150.280 321.370 151.035 ;
        RECT 321.635 150.535 324.265 150.865 ;
        RECT 322.570 150.305 322.770 150.535 ;
        RECT 324.530 150.305 324.700 151.035 ;
        RECT 321.200 149.950 322.295 150.280 ;
        RECT 322.465 149.975 322.835 150.305 ;
        RECT 323.105 149.975 326.125 150.305 ;
        RECT 326.395 149.975 326.765 150.305 ;
        RECT 298.455 149.075 298.825 149.405 ;
        RECT 299.095 149.075 302.115 149.405 ;
        RECT 302.385 149.075 302.755 149.405 ;
        RECT 302.925 149.100 304.020 149.430 ;
        RECT 297.190 148.155 298.405 148.485 ;
        RECT 298.575 148.155 299.055 148.845 ;
        RECT 300.520 148.485 300.690 149.075 ;
        RECT 299.225 148.155 301.985 148.485 ;
        RECT 302.155 148.155 302.635 148.845 ;
        RECT 303.850 148.485 304.020 149.100 ;
        RECT 302.805 148.155 304.020 148.485 ;
        RECT 297.190 147.440 297.360 148.155 ;
        RECT 297.625 147.655 300.255 147.985 ;
        RECT 297.190 147.140 298.380 147.440 ;
        RECT 297.190 146.565 297.360 147.140 ;
        RECT 298.640 146.925 298.840 147.655 ;
        RECT 300.520 147.440 300.690 148.155 ;
        RECT 300.955 147.655 303.585 147.985 ;
        RECT 299.480 147.140 301.730 147.440 ;
        RECT 297.190 146.235 298.405 146.565 ;
        RECT 298.575 146.235 299.055 146.925 ;
        RECT 300.520 146.565 300.690 147.140 ;
        RECT 302.370 146.925 302.570 147.655 ;
        RECT 303.850 147.440 304.020 148.155 ;
        RECT 302.830 147.140 304.020 147.440 ;
        RECT 299.225 146.235 301.985 146.565 ;
        RECT 302.155 146.235 302.635 146.925 ;
        RECT 303.850 146.565 304.020 147.140 ;
        RECT 302.805 146.235 304.020 146.565 ;
        RECT 297.190 145.495 297.360 146.235 ;
        RECT 297.625 145.735 300.255 146.065 ;
        RECT 297.190 145.165 298.405 145.495 ;
        RECT 298.690 145.485 298.890 145.735 ;
        RECT 297.190 144.565 297.360 145.165 ;
        RECT 297.625 144.745 298.455 144.995 ;
        RECT 297.190 144.235 298.115 144.565 ;
        RECT 285.970 139.830 288.070 140.000 ;
        RECT 288.430 143.660 292.460 143.830 ;
        RECT 283.510 134.085 285.610 134.255 ;
        RECT 285.970 139.300 288.070 139.470 ;
        RECT 285.970 134.250 286.140 139.300 ;
        RECT 286.770 138.790 287.270 138.960 ;
        RECT 286.540 138.080 286.710 138.620 ;
        RECT 287.330 138.080 287.500 138.620 ;
        RECT 286.770 137.740 287.270 137.910 ;
        RECT 286.540 137.030 286.710 137.570 ;
        RECT 287.330 137.030 287.500 137.570 ;
        RECT 286.770 136.690 287.270 136.860 ;
        RECT 286.540 135.980 286.710 136.520 ;
        RECT 287.330 135.980 287.500 136.520 ;
        RECT 286.770 135.640 287.270 135.810 ;
        RECT 286.540 134.930 286.710 135.470 ;
        RECT 287.330 134.930 287.500 135.470 ;
        RECT 286.770 134.590 287.270 134.760 ;
        RECT 287.900 134.250 288.070 139.300 ;
        RECT 285.970 134.080 288.070 134.250 ;
        RECT 288.430 134.250 288.600 143.660 ;
        RECT 289.230 143.150 289.730 143.320 ;
        RECT 289.000 141.395 289.170 142.935 ;
        RECT 289.790 141.395 289.960 142.935 ;
        RECT 289.230 141.010 289.730 141.180 ;
        RECT 289.000 139.255 289.170 140.795 ;
        RECT 289.790 139.255 289.960 140.795 ;
        RECT 289.230 138.870 289.730 139.040 ;
        RECT 289.000 137.115 289.170 138.655 ;
        RECT 289.790 137.115 289.960 138.655 ;
        RECT 289.230 136.730 289.730 136.900 ;
        RECT 289.000 134.975 289.170 136.515 ;
        RECT 289.790 134.975 289.960 136.515 ;
        RECT 289.230 134.590 289.730 134.760 ;
        RECT 290.360 134.250 290.530 143.660 ;
        RECT 291.160 143.150 291.660 143.320 ;
        RECT 290.930 141.395 291.100 142.935 ;
        RECT 291.720 141.395 291.890 142.935 ;
        RECT 291.160 141.010 291.660 141.180 ;
        RECT 290.930 139.255 291.100 140.795 ;
        RECT 291.720 139.255 291.890 140.795 ;
        RECT 291.160 138.870 291.660 139.040 ;
        RECT 290.930 137.115 291.100 138.655 ;
        RECT 291.720 137.115 291.890 138.655 ;
        RECT 291.160 136.730 291.660 136.900 ;
        RECT 290.930 134.975 291.100 136.515 ;
        RECT 291.720 134.975 291.890 136.515 ;
        RECT 291.160 134.590 291.660 134.760 ;
        RECT 292.290 134.250 292.460 143.660 ;
        RECT 297.190 143.655 297.360 144.235 ;
        RECT 298.285 144.005 298.455 144.745 ;
        RECT 297.625 143.835 298.455 144.005 ;
        RECT 297.190 143.325 298.115 143.655 ;
        RECT 298.285 143.565 298.455 143.835 ;
        RECT 298.625 143.810 299.055 145.485 ;
        RECT 300.520 145.460 300.690 146.235 ;
        RECT 300.955 145.735 303.585 146.065 ;
        RECT 302.320 145.485 302.520 145.735 ;
        RECT 303.850 145.495 304.020 146.235 ;
        RECT 299.225 145.210 301.985 145.460 ;
        RECT 299.225 144.680 300.255 145.010 ;
        RECT 299.225 144.110 299.395 144.680 ;
        RECT 300.520 144.480 300.690 145.210 ;
        RECT 300.955 144.680 301.985 145.010 ;
        RECT 299.565 144.310 301.645 144.480 ;
        RECT 299.225 143.780 300.255 144.110 ;
        RECT 299.225 143.565 299.395 143.780 ;
        RECT 300.520 143.580 300.690 144.310 ;
        RECT 301.815 144.110 301.985 144.680 ;
        RECT 300.955 143.780 301.985 144.110 ;
        RECT 302.155 143.810 302.585 145.485 ;
        RECT 302.805 145.165 304.020 145.495 ;
        RECT 302.755 144.745 303.585 144.995 ;
        RECT 302.755 144.005 302.925 144.745 ;
        RECT 303.850 144.565 304.020 145.165 ;
        RECT 303.095 144.235 304.020 144.565 ;
        RECT 302.755 143.835 303.585 144.005 ;
        RECT 298.285 143.335 299.395 143.565 ;
        RECT 297.190 143.120 297.360 143.325 ;
        RECT 297.190 142.820 298.380 143.120 ;
        RECT 297.190 142.600 297.360 142.820 ;
        RECT 297.190 142.350 298.405 142.600 ;
        RECT 297.190 141.740 297.360 142.350 ;
        RECT 298.690 142.170 298.890 143.335 ;
        RECT 299.565 143.330 301.645 143.580 ;
        RECT 301.815 143.565 301.985 143.780 ;
        RECT 302.755 143.565 302.925 143.835 ;
        RECT 303.850 143.655 304.020 144.235 ;
        RECT 301.815 143.335 302.925 143.565 ;
        RECT 300.520 143.120 300.690 143.330 ;
        RECT 299.480 142.820 301.730 143.120 ;
        RECT 300.520 142.615 300.690 142.820 ;
        RECT 299.095 142.365 302.115 142.615 ;
        RECT 297.625 141.920 298.455 142.170 ;
        RECT 297.190 141.410 298.115 141.740 ;
        RECT 297.190 140.880 297.360 141.410 ;
        RECT 298.285 141.230 298.455 141.920 ;
        RECT 297.625 141.060 298.455 141.230 ;
        RECT 297.190 140.550 298.115 140.880 ;
        RECT 297.190 139.880 297.360 140.550 ;
        RECT 298.285 140.380 298.455 141.060 ;
        RECT 298.625 140.480 299.055 142.170 ;
        RECT 299.225 141.915 300.255 142.165 ;
        RECT 299.225 141.215 299.395 141.915 ;
        RECT 300.520 141.715 300.690 142.365 ;
        RECT 302.325 142.170 302.525 143.335 ;
        RECT 303.095 143.325 304.020 143.655 ;
        RECT 303.850 143.120 304.020 143.325 ;
        RECT 302.830 142.820 304.020 143.120 ;
        RECT 303.850 142.600 304.020 142.820 ;
        RECT 302.805 142.350 304.020 142.600 ;
        RECT 300.955 141.915 301.985 142.165 ;
        RECT 299.565 141.385 301.645 141.715 ;
        RECT 299.225 140.885 300.255 141.215 ;
        RECT 297.625 140.310 298.455 140.380 ;
        RECT 297.625 140.235 298.585 140.310 ;
        RECT 299.225 140.235 299.395 140.885 ;
        RECT 300.520 140.685 300.690 141.385 ;
        RECT 301.815 141.215 301.985 141.915 ;
        RECT 300.955 140.885 301.985 141.215 ;
        RECT 299.565 140.435 301.645 140.685 ;
        RECT 297.625 140.065 300.255 140.235 ;
        RECT 297.625 140.050 298.895 140.065 ;
        RECT 297.190 139.550 298.245 139.880 ;
        RECT 288.430 134.080 292.460 134.250 ;
        RECT 292.820 139.300 296.850 139.470 ;
        RECT 292.820 134.250 292.990 139.300 ;
        RECT 293.620 138.790 294.120 138.960 ;
        RECT 293.390 138.080 293.560 138.620 ;
        RECT 294.180 138.080 294.350 138.620 ;
        RECT 293.620 137.740 294.120 137.910 ;
        RECT 293.390 137.030 293.560 137.570 ;
        RECT 294.180 137.030 294.350 137.570 ;
        RECT 293.620 136.690 294.120 136.860 ;
        RECT 293.390 135.980 293.560 136.520 ;
        RECT 294.180 135.980 294.350 136.520 ;
        RECT 293.620 135.640 294.120 135.810 ;
        RECT 293.390 134.930 293.560 135.470 ;
        RECT 294.180 134.930 294.350 135.470 ;
        RECT 293.620 134.590 294.120 134.760 ;
        RECT 294.750 134.250 294.920 139.300 ;
        RECT 295.550 138.790 296.050 138.960 ;
        RECT 295.320 138.080 295.490 138.620 ;
        RECT 296.110 138.080 296.280 138.620 ;
        RECT 295.550 137.740 296.050 137.910 ;
        RECT 295.320 137.030 295.490 137.570 ;
        RECT 296.110 137.030 296.280 137.570 ;
        RECT 295.550 136.690 296.050 136.860 ;
        RECT 295.320 135.980 295.490 136.520 ;
        RECT 296.110 135.980 296.280 136.520 ;
        RECT 295.550 135.640 296.050 135.810 ;
        RECT 295.320 134.930 295.490 135.470 ;
        RECT 296.110 134.930 296.280 135.470 ;
        RECT 295.550 134.590 296.050 134.760 ;
        RECT 296.680 134.250 296.850 139.300 ;
        RECT 292.820 134.080 296.850 134.250 ;
        RECT 297.190 138.950 297.360 139.550 ;
        RECT 298.415 139.380 298.895 140.050 ;
        RECT 300.520 139.865 300.690 140.435 ;
        RECT 301.815 140.235 301.985 140.885 ;
        RECT 302.155 140.480 302.585 142.170 ;
        RECT 302.755 141.920 303.585 142.170 ;
        RECT 302.755 141.230 302.925 141.920 ;
        RECT 303.850 141.740 304.020 142.350 ;
        RECT 303.095 141.410 304.020 141.740 ;
        RECT 302.755 141.060 303.585 141.230 ;
        RECT 302.755 140.380 302.925 141.060 ;
        RECT 303.850 140.880 304.020 141.410 ;
        RECT 303.095 140.550 304.020 140.880 ;
        RECT 302.755 140.310 303.585 140.380 ;
        RECT 302.625 140.235 303.585 140.310 ;
        RECT 300.955 140.065 303.585 140.235 ;
        RECT 302.315 140.050 303.585 140.065 ;
        RECT 299.095 139.535 302.115 139.865 ;
        RECT 297.625 139.365 298.895 139.380 ;
        RECT 297.625 139.120 300.255 139.365 ;
        RECT 298.415 139.035 300.255 139.120 ;
        RECT 297.190 138.620 298.245 138.950 ;
        RECT 297.190 138.280 297.360 138.620 ;
        RECT 298.415 138.535 298.895 139.035 ;
        RECT 300.520 138.865 300.690 139.535 ;
        RECT 302.315 139.380 302.795 140.050 ;
        RECT 303.850 139.880 304.020 140.550 ;
        RECT 302.965 139.550 304.020 139.880 ;
        RECT 305.060 149.415 307.160 149.585 ;
        RECT 305.060 140.005 305.230 149.415 ;
        RECT 305.860 148.905 306.360 149.075 ;
        RECT 305.630 147.150 305.800 148.690 ;
        RECT 306.420 147.150 306.590 148.690 ;
        RECT 305.860 146.765 306.360 146.935 ;
        RECT 305.630 145.010 305.800 146.550 ;
        RECT 306.420 145.010 306.590 146.550 ;
        RECT 305.860 144.625 306.360 144.795 ;
        RECT 305.630 142.870 305.800 144.410 ;
        RECT 306.420 142.870 306.590 144.410 ;
        RECT 305.860 142.485 306.360 142.655 ;
        RECT 305.630 140.730 305.800 142.270 ;
        RECT 306.420 140.730 306.590 142.270 ;
        RECT 305.860 140.345 306.360 140.515 ;
        RECT 306.990 140.005 307.160 149.415 ;
        RECT 307.520 149.415 309.620 149.585 ;
        RECT 307.520 144.365 307.690 149.415 ;
        RECT 308.320 148.905 308.820 149.075 ;
        RECT 308.090 148.195 308.260 148.735 ;
        RECT 308.880 148.195 309.050 148.735 ;
        RECT 308.320 147.855 308.820 148.025 ;
        RECT 308.090 147.145 308.260 147.685 ;
        RECT 308.880 147.145 309.050 147.685 ;
        RECT 308.320 146.805 308.820 146.975 ;
        RECT 308.090 146.095 308.260 146.635 ;
        RECT 308.880 146.095 309.050 146.635 ;
        RECT 308.320 145.755 308.820 145.925 ;
        RECT 308.090 145.045 308.260 145.585 ;
        RECT 308.880 145.045 309.050 145.585 ;
        RECT 308.320 144.705 308.820 144.875 ;
        RECT 309.450 144.365 309.620 149.415 ;
        RECT 307.520 144.195 309.620 144.365 ;
        RECT 309.980 149.410 312.080 149.580 ;
        RECT 305.060 139.835 307.160 140.005 ;
        RECT 307.520 143.665 309.620 143.835 ;
        RECT 302.315 139.365 303.585 139.380 ;
        RECT 300.955 139.120 303.585 139.365 ;
        RECT 300.955 139.035 302.795 139.120 ;
        RECT 299.095 138.535 302.115 138.865 ;
        RECT 302.315 138.535 302.795 139.035 ;
        RECT 303.850 138.950 304.020 139.550 ;
        RECT 302.965 138.620 304.020 138.950 ;
        RECT 297.190 138.030 298.405 138.280 ;
        RECT 297.190 137.420 297.360 138.030 ;
        RECT 298.690 137.850 298.890 138.535 ;
        RECT 300.520 138.295 300.690 138.535 ;
        RECT 299.095 138.045 302.115 138.295 ;
        RECT 297.625 137.600 298.455 137.850 ;
        RECT 297.190 137.090 298.115 137.420 ;
        RECT 297.190 136.560 297.360 137.090 ;
        RECT 298.285 136.910 298.455 137.600 ;
        RECT 297.625 136.740 298.455 136.910 ;
        RECT 297.190 136.230 298.115 136.560 ;
        RECT 297.190 135.560 297.360 136.230 ;
        RECT 298.285 136.060 298.455 136.740 ;
        RECT 298.625 136.160 299.055 137.850 ;
        RECT 299.225 137.595 300.255 137.845 ;
        RECT 299.225 136.895 299.395 137.595 ;
        RECT 300.520 137.395 300.690 138.045 ;
        RECT 302.320 137.850 302.520 138.535 ;
        RECT 303.850 138.280 304.020 138.620 ;
        RECT 302.805 138.030 304.020 138.280 ;
        RECT 300.955 137.595 301.985 137.845 ;
        RECT 299.565 137.065 301.645 137.395 ;
        RECT 299.225 136.565 300.255 136.895 ;
        RECT 297.625 135.990 298.455 136.060 ;
        RECT 297.625 135.915 298.585 135.990 ;
        RECT 299.225 135.915 299.395 136.565 ;
        RECT 300.520 136.365 300.690 137.065 ;
        RECT 301.815 136.895 301.985 137.595 ;
        RECT 300.955 136.565 301.985 136.895 ;
        RECT 299.565 136.115 301.645 136.365 ;
        RECT 297.625 135.745 300.255 135.915 ;
        RECT 297.625 135.730 298.895 135.745 ;
        RECT 297.190 135.230 298.245 135.560 ;
        RECT 297.190 134.630 297.360 135.230 ;
        RECT 298.415 135.060 298.895 135.730 ;
        RECT 300.520 135.545 300.690 136.115 ;
        RECT 301.815 135.915 301.985 136.565 ;
        RECT 302.155 136.160 302.585 137.850 ;
        RECT 302.755 137.600 303.585 137.850 ;
        RECT 302.755 136.910 302.925 137.600 ;
        RECT 303.850 137.420 304.020 138.030 ;
        RECT 303.095 137.090 304.020 137.420 ;
        RECT 302.755 136.740 303.585 136.910 ;
        RECT 302.755 136.060 302.925 136.740 ;
        RECT 303.850 136.560 304.020 137.090 ;
        RECT 303.095 136.230 304.020 136.560 ;
        RECT 302.755 135.990 303.585 136.060 ;
        RECT 302.625 135.915 303.585 135.990 ;
        RECT 300.955 135.745 303.585 135.915 ;
        RECT 302.315 135.730 303.585 135.745 ;
        RECT 299.095 135.215 302.115 135.545 ;
        RECT 297.625 135.045 298.895 135.060 ;
        RECT 297.625 134.800 300.255 135.045 ;
        RECT 298.415 134.715 300.255 134.800 ;
        RECT 297.190 134.300 298.245 134.630 ;
        RECT 297.190 134.090 297.360 134.300 ;
        RECT 298.415 134.215 298.895 134.715 ;
        RECT 300.520 134.545 300.690 135.215 ;
        RECT 302.315 135.060 302.795 135.730 ;
        RECT 303.850 135.560 304.020 136.230 ;
        RECT 302.965 135.230 304.020 135.560 ;
        RECT 302.315 135.045 303.585 135.060 ;
        RECT 300.955 134.800 303.585 135.045 ;
        RECT 300.955 134.715 302.795 134.800 ;
        RECT 299.095 134.215 302.115 134.545 ;
        RECT 302.315 134.215 302.795 134.715 ;
        RECT 303.850 134.630 304.020 135.230 ;
        RECT 302.965 134.300 304.020 134.630 ;
        RECT 300.520 134.090 300.690 134.215 ;
        RECT 303.850 134.090 304.020 134.300 ;
        RECT 305.060 139.305 307.160 139.475 ;
        RECT 305.060 134.255 305.230 139.305 ;
        RECT 305.860 138.795 306.360 138.965 ;
        RECT 305.630 138.085 305.800 138.625 ;
        RECT 306.420 138.085 306.590 138.625 ;
        RECT 305.860 137.745 306.360 137.915 ;
        RECT 305.630 137.035 305.800 137.575 ;
        RECT 306.420 137.035 306.590 137.575 ;
        RECT 305.860 136.695 306.360 136.865 ;
        RECT 305.630 135.985 305.800 136.525 ;
        RECT 306.420 135.985 306.590 136.525 ;
        RECT 305.860 135.645 306.360 135.815 ;
        RECT 305.630 134.935 305.800 135.475 ;
        RECT 306.420 134.935 306.590 135.475 ;
        RECT 305.860 134.595 306.360 134.765 ;
        RECT 306.990 134.255 307.160 139.305 ;
        RECT 305.060 134.085 307.160 134.255 ;
        RECT 307.520 134.255 307.690 143.665 ;
        RECT 308.320 143.155 308.820 143.325 ;
        RECT 308.090 141.400 308.260 142.940 ;
        RECT 308.880 141.400 309.050 142.940 ;
        RECT 308.320 141.015 308.820 141.185 ;
        RECT 308.090 139.260 308.260 140.800 ;
        RECT 308.880 139.260 309.050 140.800 ;
        RECT 308.320 138.875 308.820 139.045 ;
        RECT 308.090 137.120 308.260 138.660 ;
        RECT 308.880 137.120 309.050 138.660 ;
        RECT 308.320 136.735 308.820 136.905 ;
        RECT 308.090 134.980 308.260 136.520 ;
        RECT 308.880 134.980 309.050 136.520 ;
        RECT 308.320 134.595 308.820 134.765 ;
        RECT 309.450 134.255 309.620 143.665 ;
        RECT 309.980 140.000 310.150 149.410 ;
        RECT 310.780 148.900 311.280 149.070 ;
        RECT 310.550 147.145 310.720 148.685 ;
        RECT 311.340 147.145 311.510 148.685 ;
        RECT 310.780 146.760 311.280 146.930 ;
        RECT 310.550 145.005 310.720 146.545 ;
        RECT 311.340 145.005 311.510 146.545 ;
        RECT 310.780 144.620 311.280 144.790 ;
        RECT 310.550 142.865 310.720 144.405 ;
        RECT 311.340 142.865 311.510 144.405 ;
        RECT 310.780 142.480 311.280 142.650 ;
        RECT 310.550 140.725 310.720 142.265 ;
        RECT 311.340 140.725 311.510 142.265 ;
        RECT 310.780 140.340 311.280 140.510 ;
        RECT 311.910 140.000 312.080 149.410 ;
        RECT 321.200 148.485 321.370 149.950 ;
        RECT 322.465 149.745 324.265 149.805 ;
        RECT 322.125 149.575 324.265 149.745 ;
        RECT 322.125 149.460 322.295 149.575 ;
        RECT 321.635 149.130 322.295 149.460 ;
        RECT 324.530 149.405 324.700 149.975 ;
        RECT 326.935 149.920 327.595 150.250 ;
        RECT 326.935 149.805 327.105 149.920 ;
        RECT 324.965 149.635 327.105 149.805 ;
        RECT 324.965 149.575 326.765 149.635 ;
        RECT 327.860 149.430 328.030 150.410 ;
        RECT 322.465 149.075 322.835 149.405 ;
        RECT 323.105 149.075 326.125 149.405 ;
        RECT 326.395 149.075 326.765 149.405 ;
        RECT 326.935 149.100 328.030 149.430 ;
        RECT 321.200 148.155 322.415 148.485 ;
        RECT 322.585 148.155 323.065 148.845 ;
        RECT 324.530 148.485 324.700 149.075 ;
        RECT 323.235 148.155 325.995 148.485 ;
        RECT 326.165 148.155 326.645 148.845 ;
        RECT 327.860 148.485 328.030 149.100 ;
        RECT 326.815 148.155 328.030 148.485 ;
        RECT 321.200 147.440 321.370 148.155 ;
        RECT 321.635 147.655 324.265 147.985 ;
        RECT 321.200 147.140 322.390 147.440 ;
        RECT 321.200 146.565 321.370 147.140 ;
        RECT 322.650 146.925 322.850 147.655 ;
        RECT 324.530 147.440 324.700 148.155 ;
        RECT 324.965 147.655 327.595 147.985 ;
        RECT 323.490 147.140 325.740 147.440 ;
        RECT 321.200 146.235 322.415 146.565 ;
        RECT 322.585 146.235 323.065 146.925 ;
        RECT 324.530 146.565 324.700 147.140 ;
        RECT 326.380 146.925 326.580 147.655 ;
        RECT 327.860 147.440 328.030 148.155 ;
        RECT 326.840 147.140 328.030 147.440 ;
        RECT 323.235 146.235 325.995 146.565 ;
        RECT 326.165 146.235 326.645 146.925 ;
        RECT 327.860 146.565 328.030 147.140 ;
        RECT 326.815 146.235 328.030 146.565 ;
        RECT 321.200 145.495 321.370 146.235 ;
        RECT 321.635 145.735 324.265 146.065 ;
        RECT 321.200 145.165 322.415 145.495 ;
        RECT 322.700 145.485 322.900 145.735 ;
        RECT 321.200 144.565 321.370 145.165 ;
        RECT 321.635 144.745 322.465 144.995 ;
        RECT 321.200 144.235 322.125 144.565 ;
        RECT 309.980 139.830 312.080 140.000 ;
        RECT 312.440 143.660 316.470 143.830 ;
        RECT 307.520 134.085 309.620 134.255 ;
        RECT 309.980 139.300 312.080 139.470 ;
        RECT 309.980 134.250 310.150 139.300 ;
        RECT 310.780 138.790 311.280 138.960 ;
        RECT 310.550 138.080 310.720 138.620 ;
        RECT 311.340 138.080 311.510 138.620 ;
        RECT 310.780 137.740 311.280 137.910 ;
        RECT 310.550 137.030 310.720 137.570 ;
        RECT 311.340 137.030 311.510 137.570 ;
        RECT 310.780 136.690 311.280 136.860 ;
        RECT 310.550 135.980 310.720 136.520 ;
        RECT 311.340 135.980 311.510 136.520 ;
        RECT 310.780 135.640 311.280 135.810 ;
        RECT 310.550 134.930 310.720 135.470 ;
        RECT 311.340 134.930 311.510 135.470 ;
        RECT 310.780 134.590 311.280 134.760 ;
        RECT 311.910 134.250 312.080 139.300 ;
        RECT 309.980 134.080 312.080 134.250 ;
        RECT 312.440 134.250 312.610 143.660 ;
        RECT 313.240 143.150 313.740 143.320 ;
        RECT 313.010 141.395 313.180 142.935 ;
        RECT 313.800 141.395 313.970 142.935 ;
        RECT 313.240 141.010 313.740 141.180 ;
        RECT 313.010 139.255 313.180 140.795 ;
        RECT 313.800 139.255 313.970 140.795 ;
        RECT 313.240 138.870 313.740 139.040 ;
        RECT 313.010 137.115 313.180 138.655 ;
        RECT 313.800 137.115 313.970 138.655 ;
        RECT 313.240 136.730 313.740 136.900 ;
        RECT 313.010 134.975 313.180 136.515 ;
        RECT 313.800 134.975 313.970 136.515 ;
        RECT 313.240 134.590 313.740 134.760 ;
        RECT 314.370 134.250 314.540 143.660 ;
        RECT 315.170 143.150 315.670 143.320 ;
        RECT 314.940 141.395 315.110 142.935 ;
        RECT 315.730 141.395 315.900 142.935 ;
        RECT 315.170 141.010 315.670 141.180 ;
        RECT 314.940 139.255 315.110 140.795 ;
        RECT 315.730 139.255 315.900 140.795 ;
        RECT 315.170 138.870 315.670 139.040 ;
        RECT 314.940 137.115 315.110 138.655 ;
        RECT 315.730 137.115 315.900 138.655 ;
        RECT 315.170 136.730 315.670 136.900 ;
        RECT 314.940 134.975 315.110 136.515 ;
        RECT 315.730 134.975 315.900 136.515 ;
        RECT 315.170 134.590 315.670 134.760 ;
        RECT 316.300 134.250 316.470 143.660 ;
        RECT 321.200 143.655 321.370 144.235 ;
        RECT 322.295 144.005 322.465 144.745 ;
        RECT 321.635 143.835 322.465 144.005 ;
        RECT 321.200 143.325 322.125 143.655 ;
        RECT 322.295 143.565 322.465 143.835 ;
        RECT 322.635 143.810 323.065 145.485 ;
        RECT 324.530 145.460 324.700 146.235 ;
        RECT 324.965 145.735 327.595 146.065 ;
        RECT 326.330 145.485 326.530 145.735 ;
        RECT 327.860 145.495 328.030 146.235 ;
        RECT 323.235 145.210 325.995 145.460 ;
        RECT 323.235 144.680 324.265 145.010 ;
        RECT 323.235 144.110 323.405 144.680 ;
        RECT 324.530 144.480 324.700 145.210 ;
        RECT 324.965 144.680 325.995 145.010 ;
        RECT 323.575 144.310 325.655 144.480 ;
        RECT 323.235 143.780 324.265 144.110 ;
        RECT 323.235 143.565 323.405 143.780 ;
        RECT 324.530 143.580 324.700 144.310 ;
        RECT 325.825 144.110 325.995 144.680 ;
        RECT 324.965 143.780 325.995 144.110 ;
        RECT 326.165 143.810 326.595 145.485 ;
        RECT 326.815 145.165 328.030 145.495 ;
        RECT 326.765 144.745 327.595 144.995 ;
        RECT 326.765 144.005 326.935 144.745 ;
        RECT 327.860 144.565 328.030 145.165 ;
        RECT 327.105 144.235 328.030 144.565 ;
        RECT 326.765 143.835 327.595 144.005 ;
        RECT 322.295 143.335 323.405 143.565 ;
        RECT 321.200 143.120 321.370 143.325 ;
        RECT 321.200 142.820 322.390 143.120 ;
        RECT 321.200 142.600 321.370 142.820 ;
        RECT 321.200 142.350 322.415 142.600 ;
        RECT 321.200 141.740 321.370 142.350 ;
        RECT 322.700 142.170 322.900 143.335 ;
        RECT 323.575 143.330 325.655 143.580 ;
        RECT 325.825 143.565 325.995 143.780 ;
        RECT 326.765 143.565 326.935 143.835 ;
        RECT 327.860 143.655 328.030 144.235 ;
        RECT 325.825 143.335 326.935 143.565 ;
        RECT 324.530 143.120 324.700 143.330 ;
        RECT 323.490 142.820 325.740 143.120 ;
        RECT 324.530 142.615 324.700 142.820 ;
        RECT 323.105 142.365 326.125 142.615 ;
        RECT 321.635 141.920 322.465 142.170 ;
        RECT 321.200 141.410 322.125 141.740 ;
        RECT 321.200 140.880 321.370 141.410 ;
        RECT 322.295 141.230 322.465 141.920 ;
        RECT 321.635 141.060 322.465 141.230 ;
        RECT 321.200 140.550 322.125 140.880 ;
        RECT 321.200 139.880 321.370 140.550 ;
        RECT 322.295 140.380 322.465 141.060 ;
        RECT 322.635 140.480 323.065 142.170 ;
        RECT 323.235 141.915 324.265 142.165 ;
        RECT 323.235 141.215 323.405 141.915 ;
        RECT 324.530 141.715 324.700 142.365 ;
        RECT 326.335 142.170 326.535 143.335 ;
        RECT 327.105 143.325 328.030 143.655 ;
        RECT 327.860 143.120 328.030 143.325 ;
        RECT 326.840 142.820 328.030 143.120 ;
        RECT 327.860 142.600 328.030 142.820 ;
        RECT 326.815 142.350 328.030 142.600 ;
        RECT 324.965 141.915 325.995 142.165 ;
        RECT 323.575 141.385 325.655 141.715 ;
        RECT 323.235 140.885 324.265 141.215 ;
        RECT 321.635 140.310 322.465 140.380 ;
        RECT 321.635 140.235 322.595 140.310 ;
        RECT 323.235 140.235 323.405 140.885 ;
        RECT 324.530 140.685 324.700 141.385 ;
        RECT 325.825 141.215 325.995 141.915 ;
        RECT 324.965 140.885 325.995 141.215 ;
        RECT 323.575 140.435 325.655 140.685 ;
        RECT 321.635 140.065 324.265 140.235 ;
        RECT 321.635 140.050 322.905 140.065 ;
        RECT 321.200 139.550 322.255 139.880 ;
        RECT 312.440 134.080 316.470 134.250 ;
        RECT 316.830 139.300 320.860 139.470 ;
        RECT 316.830 134.250 317.000 139.300 ;
        RECT 317.630 138.790 318.130 138.960 ;
        RECT 317.400 138.080 317.570 138.620 ;
        RECT 318.190 138.080 318.360 138.620 ;
        RECT 317.630 137.740 318.130 137.910 ;
        RECT 317.400 137.030 317.570 137.570 ;
        RECT 318.190 137.030 318.360 137.570 ;
        RECT 317.630 136.690 318.130 136.860 ;
        RECT 317.400 135.980 317.570 136.520 ;
        RECT 318.190 135.980 318.360 136.520 ;
        RECT 317.630 135.640 318.130 135.810 ;
        RECT 317.400 134.930 317.570 135.470 ;
        RECT 318.190 134.930 318.360 135.470 ;
        RECT 317.630 134.590 318.130 134.760 ;
        RECT 318.760 134.250 318.930 139.300 ;
        RECT 319.560 138.790 320.060 138.960 ;
        RECT 319.330 138.080 319.500 138.620 ;
        RECT 320.120 138.080 320.290 138.620 ;
        RECT 319.560 137.740 320.060 137.910 ;
        RECT 319.330 137.030 319.500 137.570 ;
        RECT 320.120 137.030 320.290 137.570 ;
        RECT 319.560 136.690 320.060 136.860 ;
        RECT 319.330 135.980 319.500 136.520 ;
        RECT 320.120 135.980 320.290 136.520 ;
        RECT 319.560 135.640 320.060 135.810 ;
        RECT 319.330 134.930 319.500 135.470 ;
        RECT 320.120 134.930 320.290 135.470 ;
        RECT 319.560 134.590 320.060 134.760 ;
        RECT 320.690 134.250 320.860 139.300 ;
        RECT 316.830 134.080 320.860 134.250 ;
        RECT 321.200 138.950 321.370 139.550 ;
        RECT 322.425 139.380 322.905 140.050 ;
        RECT 324.530 139.865 324.700 140.435 ;
        RECT 325.825 140.235 325.995 140.885 ;
        RECT 326.165 140.480 326.595 142.170 ;
        RECT 326.765 141.920 327.595 142.170 ;
        RECT 326.765 141.230 326.935 141.920 ;
        RECT 327.860 141.740 328.030 142.350 ;
        RECT 327.105 141.410 328.030 141.740 ;
        RECT 326.765 141.060 327.595 141.230 ;
        RECT 326.765 140.380 326.935 141.060 ;
        RECT 327.860 140.880 328.030 141.410 ;
        RECT 327.105 140.550 328.030 140.880 ;
        RECT 326.765 140.310 327.595 140.380 ;
        RECT 326.635 140.235 327.595 140.310 ;
        RECT 324.965 140.065 327.595 140.235 ;
        RECT 326.325 140.050 327.595 140.065 ;
        RECT 323.105 139.535 326.125 139.865 ;
        RECT 321.635 139.365 322.905 139.380 ;
        RECT 321.635 139.120 324.265 139.365 ;
        RECT 322.425 139.035 324.265 139.120 ;
        RECT 321.200 138.620 322.255 138.950 ;
        RECT 321.200 138.280 321.370 138.620 ;
        RECT 322.425 138.535 322.905 139.035 ;
        RECT 324.530 138.865 324.700 139.535 ;
        RECT 326.325 139.380 326.805 140.050 ;
        RECT 327.860 139.880 328.030 140.550 ;
        RECT 326.975 139.550 328.030 139.880 ;
        RECT 326.325 139.365 327.595 139.380 ;
        RECT 324.965 139.120 327.595 139.365 ;
        RECT 324.965 139.035 326.805 139.120 ;
        RECT 323.105 138.535 326.125 138.865 ;
        RECT 326.325 138.535 326.805 139.035 ;
        RECT 327.860 138.950 328.030 139.550 ;
        RECT 326.975 138.620 328.030 138.950 ;
        RECT 321.200 138.030 322.415 138.280 ;
        RECT 321.200 137.420 321.370 138.030 ;
        RECT 322.700 137.850 322.900 138.535 ;
        RECT 324.530 138.295 324.700 138.535 ;
        RECT 323.105 138.045 326.125 138.295 ;
        RECT 321.635 137.600 322.465 137.850 ;
        RECT 321.200 137.090 322.125 137.420 ;
        RECT 321.200 136.560 321.370 137.090 ;
        RECT 322.295 136.910 322.465 137.600 ;
        RECT 321.635 136.740 322.465 136.910 ;
        RECT 321.200 136.230 322.125 136.560 ;
        RECT 321.200 135.560 321.370 136.230 ;
        RECT 322.295 136.060 322.465 136.740 ;
        RECT 322.635 136.160 323.065 137.850 ;
        RECT 323.235 137.595 324.265 137.845 ;
        RECT 323.235 136.895 323.405 137.595 ;
        RECT 324.530 137.395 324.700 138.045 ;
        RECT 326.330 137.850 326.530 138.535 ;
        RECT 327.860 138.280 328.030 138.620 ;
        RECT 326.815 138.030 328.030 138.280 ;
        RECT 324.965 137.595 325.995 137.845 ;
        RECT 323.575 137.065 325.655 137.395 ;
        RECT 323.235 136.565 324.265 136.895 ;
        RECT 321.635 135.990 322.465 136.060 ;
        RECT 321.635 135.915 322.595 135.990 ;
        RECT 323.235 135.915 323.405 136.565 ;
        RECT 324.530 136.365 324.700 137.065 ;
        RECT 325.825 136.895 325.995 137.595 ;
        RECT 324.965 136.565 325.995 136.895 ;
        RECT 323.575 136.115 325.655 136.365 ;
        RECT 321.635 135.745 324.265 135.915 ;
        RECT 321.635 135.730 322.905 135.745 ;
        RECT 321.200 135.230 322.255 135.560 ;
        RECT 321.200 134.630 321.370 135.230 ;
        RECT 322.425 135.060 322.905 135.730 ;
        RECT 324.530 135.545 324.700 136.115 ;
        RECT 325.825 135.915 325.995 136.565 ;
        RECT 326.165 136.160 326.595 137.850 ;
        RECT 326.765 137.600 327.595 137.850 ;
        RECT 326.765 136.910 326.935 137.600 ;
        RECT 327.860 137.420 328.030 138.030 ;
        RECT 327.105 137.090 328.030 137.420 ;
        RECT 326.765 136.740 327.595 136.910 ;
        RECT 326.765 136.060 326.935 136.740 ;
        RECT 327.860 136.560 328.030 137.090 ;
        RECT 327.105 136.230 328.030 136.560 ;
        RECT 326.765 135.990 327.595 136.060 ;
        RECT 326.635 135.915 327.595 135.990 ;
        RECT 324.965 135.745 327.595 135.915 ;
        RECT 326.325 135.730 327.595 135.745 ;
        RECT 323.105 135.215 326.125 135.545 ;
        RECT 321.635 135.045 322.905 135.060 ;
        RECT 321.635 134.800 324.265 135.045 ;
        RECT 322.425 134.715 324.265 134.800 ;
        RECT 321.200 134.300 322.255 134.630 ;
        RECT 321.200 134.090 321.370 134.300 ;
        RECT 322.425 134.215 322.905 134.715 ;
        RECT 324.530 134.545 324.700 135.215 ;
        RECT 326.325 135.060 326.805 135.730 ;
        RECT 327.860 135.560 328.030 136.230 ;
        RECT 326.975 135.230 328.030 135.560 ;
        RECT 326.325 135.045 327.595 135.060 ;
        RECT 324.965 134.800 327.595 135.045 ;
        RECT 324.965 134.715 326.805 134.800 ;
        RECT 323.105 134.215 326.125 134.545 ;
        RECT 326.325 134.215 326.805 134.715 ;
        RECT 327.860 134.630 328.030 135.230 ;
        RECT 326.975 134.300 328.030 134.630 ;
        RECT 324.530 134.090 324.700 134.215 ;
        RECT 327.860 134.090 328.030 134.300 ;
        RECT 10.200 133.545 69.720 133.715 ;
        RECT 10.295 132.230 10.625 133.545 ;
        RECT 10.370 130.385 10.940 131.885 ;
        RECT 11.345 131.550 11.915 133.545 ;
        RECT 12.235 132.120 12.565 133.545 ;
        RECT 12.735 132.185 13.435 133.280 ;
        RECT 12.735 131.430 12.995 132.185 ;
        RECT 13.605 132.015 13.775 133.205 ;
        RECT 13.975 132.495 14.305 133.545 ;
        RECT 14.475 132.745 14.840 133.205 ;
        RECT 15.025 132.745 15.355 133.545 ;
        RECT 15.525 132.775 16.680 133.105 ;
        RECT 14.475 132.325 14.645 132.745 ;
        RECT 11.650 130.385 11.980 131.105 ;
        RECT 12.235 130.385 12.485 131.430 ;
        RECT 12.665 130.650 12.995 131.430 ;
        RECT 13.225 131.685 13.775 132.015 ;
        RECT 13.970 132.155 14.645 132.325 ;
        RECT 14.815 132.220 15.355 132.555 ;
        RECT 13.225 130.650 13.555 131.685 ;
        RECT 13.970 131.485 14.140 132.155 ;
        RECT 15.525 131.985 15.695 132.775 ;
        RECT 14.310 131.815 15.695 131.985 ;
        RECT 14.310 131.655 14.640 131.815 ;
        RECT 15.865 131.645 16.195 132.605 ;
        RECT 16.510 131.985 16.680 132.775 ;
        RECT 16.850 132.165 17.180 133.055 ;
        RECT 16.510 131.815 16.840 131.985 ;
        RECT 15.240 131.485 15.570 131.645 ;
        RECT 13.970 131.315 15.570 131.485 ;
        RECT 15.740 131.315 16.470 131.645 ;
        RECT 13.735 130.385 13.985 131.145 ;
        RECT 14.215 130.685 14.545 131.315 ;
        RECT 15.085 130.385 15.415 131.145 ;
        RECT 15.740 130.725 15.910 131.315 ;
        RECT 16.670 131.145 16.840 131.815 ;
        RECT 16.080 130.895 16.840 131.145 ;
        RECT 17.010 131.430 17.180 132.165 ;
        RECT 17.350 132.045 17.680 133.545 ;
        RECT 18.445 133.040 18.775 133.545 ;
        RECT 19.370 132.870 19.700 133.025 ;
        RECT 17.910 132.700 19.700 132.870 ;
        RECT 19.900 132.810 20.150 133.025 ;
        RECT 20.845 132.980 21.175 133.545 ;
        RECT 21.825 132.950 22.075 133.545 ;
        RECT 22.275 132.820 22.605 133.280 ;
        RECT 22.805 132.820 23.055 133.545 ;
        RECT 19.900 132.780 21.655 132.810 ;
        RECT 22.275 132.780 22.475 132.820 ;
        RECT 17.910 132.620 18.545 132.700 ;
        RECT 17.875 132.095 18.205 132.450 ;
        RECT 18.375 131.875 18.545 132.620 ;
        RECT 17.510 131.545 18.545 131.875 ;
        RECT 17.010 131.375 17.340 131.430 ;
        RECT 18.715 131.375 18.895 132.425 ;
        RECT 17.010 131.205 18.895 131.375 ;
        RECT 19.065 131.350 19.235 132.700 ;
        RECT 19.900 132.640 22.475 132.780 ;
        RECT 19.900 132.530 20.150 132.640 ;
        RECT 21.485 132.610 22.475 132.640 ;
        RECT 19.405 132.360 20.150 132.530 ;
        RECT 19.405 131.690 19.575 132.360 ;
        RECT 20.395 132.190 20.645 132.470 ;
        RECT 19.745 132.020 20.645 132.190 ;
        RECT 21.295 132.110 21.705 132.440 ;
        RECT 19.745 131.860 20.295 132.020 ;
        RECT 19.405 131.520 19.955 131.690 ;
        RECT 17.010 130.965 17.340 131.205 ;
        RECT 17.510 130.865 18.895 131.035 ;
        RECT 19.065 130.970 19.535 131.350 ;
        RECT 19.705 130.970 19.955 131.520 ;
        RECT 20.125 131.100 20.295 131.860 ;
        RECT 20.885 131.940 21.115 132.080 ;
        RECT 20.465 131.440 20.715 131.850 ;
        RECT 20.885 131.610 21.365 131.940 ;
        RECT 21.535 131.440 21.705 132.110 ;
        RECT 20.465 131.270 21.705 131.440 ;
        RECT 21.875 131.430 22.135 132.440 ;
        RECT 17.510 130.725 17.680 130.865 ;
        RECT 15.740 130.555 17.680 130.725 ;
        RECT 18.725 130.800 18.895 130.865 ;
        RECT 20.125 130.800 20.650 131.100 ;
        RECT 17.850 130.385 18.245 130.695 ;
        RECT 18.725 130.630 20.650 130.800 ;
        RECT 20.820 130.385 21.150 131.100 ;
        RECT 21.320 130.650 21.705 131.270 ;
        RECT 22.305 131.130 22.475 132.610 ;
        RECT 23.250 132.505 23.550 133.545 ;
        RECT 22.645 131.300 23.035 132.470 ;
        RECT 35.255 132.230 35.585 133.545 ;
        RECT 21.880 130.385 22.130 131.130 ;
        RECT 22.305 130.960 23.030 131.130 ;
        RECT 22.700 130.670 23.030 130.960 ;
        RECT 23.250 130.385 23.550 131.405 ;
        RECT 35.330 130.385 35.900 131.885 ;
        RECT 36.305 131.550 36.875 133.545 ;
        RECT 38.155 132.120 38.485 133.545 ;
        RECT 38.655 132.185 39.355 133.280 ;
        RECT 38.655 131.430 38.915 132.185 ;
        RECT 39.525 132.015 39.695 133.205 ;
        RECT 39.895 132.495 40.225 133.545 ;
        RECT 40.395 132.745 40.760 133.205 ;
        RECT 40.945 132.745 41.275 133.545 ;
        RECT 41.445 132.775 42.600 133.105 ;
        RECT 40.395 132.325 40.565 132.745 ;
        RECT 36.610 130.385 36.940 131.105 ;
        RECT 38.155 130.385 38.405 131.430 ;
        RECT 38.585 130.650 38.915 131.430 ;
        RECT 39.145 131.685 39.695 132.015 ;
        RECT 39.890 132.155 40.565 132.325 ;
        RECT 40.735 132.220 41.275 132.555 ;
        RECT 39.145 130.650 39.475 131.685 ;
        RECT 39.890 131.485 40.060 132.155 ;
        RECT 41.445 131.985 41.615 132.775 ;
        RECT 40.230 131.815 41.615 131.985 ;
        RECT 40.230 131.655 40.560 131.815 ;
        RECT 41.785 131.645 42.115 132.605 ;
        RECT 42.430 131.985 42.600 132.775 ;
        RECT 42.770 132.165 43.100 133.055 ;
        RECT 42.430 131.815 42.760 131.985 ;
        RECT 41.160 131.485 41.490 131.645 ;
        RECT 39.890 131.315 41.490 131.485 ;
        RECT 41.660 131.315 42.390 131.645 ;
        RECT 39.655 130.385 39.905 131.145 ;
        RECT 40.135 130.685 40.465 131.315 ;
        RECT 41.005 130.385 41.335 131.145 ;
        RECT 41.660 130.725 41.830 131.315 ;
        RECT 42.590 131.145 42.760 131.815 ;
        RECT 42.000 130.895 42.760 131.145 ;
        RECT 42.930 131.430 43.100 132.165 ;
        RECT 43.270 132.045 43.600 133.545 ;
        RECT 44.365 133.040 44.695 133.545 ;
        RECT 45.290 132.870 45.620 133.025 ;
        RECT 43.830 132.700 45.620 132.870 ;
        RECT 45.820 132.810 46.070 133.025 ;
        RECT 46.765 132.980 47.095 133.545 ;
        RECT 47.745 132.950 47.995 133.545 ;
        RECT 48.195 132.820 48.525 133.280 ;
        RECT 48.725 132.820 48.975 133.545 ;
        RECT 45.820 132.780 47.575 132.810 ;
        RECT 48.195 132.780 48.395 132.820 ;
        RECT 43.830 132.620 44.465 132.700 ;
        RECT 43.795 132.095 44.125 132.450 ;
        RECT 44.295 131.875 44.465 132.620 ;
        RECT 43.430 131.545 44.465 131.875 ;
        RECT 42.930 131.375 43.260 131.430 ;
        RECT 44.635 131.375 44.815 132.425 ;
        RECT 42.930 131.205 44.815 131.375 ;
        RECT 44.985 131.350 45.155 132.700 ;
        RECT 45.820 132.640 48.395 132.780 ;
        RECT 45.820 132.530 46.070 132.640 ;
        RECT 47.405 132.610 48.395 132.640 ;
        RECT 45.325 132.360 46.070 132.530 ;
        RECT 45.325 131.690 45.495 132.360 ;
        RECT 46.315 132.190 46.565 132.470 ;
        RECT 45.665 132.020 46.565 132.190 ;
        RECT 47.215 132.110 47.625 132.440 ;
        RECT 45.665 131.860 46.215 132.020 ;
        RECT 45.325 131.520 45.875 131.690 ;
        RECT 42.930 130.965 43.260 131.205 ;
        RECT 43.430 130.865 44.815 131.035 ;
        RECT 44.985 130.970 45.455 131.350 ;
        RECT 45.625 130.970 45.875 131.520 ;
        RECT 46.045 131.100 46.215 131.860 ;
        RECT 46.805 131.940 47.035 132.080 ;
        RECT 46.385 131.440 46.635 131.850 ;
        RECT 46.805 131.610 47.285 131.940 ;
        RECT 47.455 131.440 47.625 132.110 ;
        RECT 46.385 131.270 47.625 131.440 ;
        RECT 47.795 131.430 48.055 132.440 ;
        RECT 43.430 130.725 43.600 130.865 ;
        RECT 41.660 130.555 43.600 130.725 ;
        RECT 44.645 130.800 44.815 130.865 ;
        RECT 46.045 130.800 46.570 131.100 ;
        RECT 43.770 130.385 44.165 130.695 ;
        RECT 44.645 130.630 46.570 130.800 ;
        RECT 46.740 130.385 47.070 131.100 ;
        RECT 47.240 130.650 47.625 131.270 ;
        RECT 48.225 131.130 48.395 132.610 ;
        RECT 49.170 132.505 49.470 133.545 ;
        RECT 48.565 131.300 48.955 132.470 ;
        RECT 53.995 132.120 54.245 133.545 ;
        RECT 54.415 132.390 54.695 133.280 ;
        RECT 54.895 132.560 55.145 133.545 ;
        RECT 55.345 132.390 55.675 133.280 ;
        RECT 54.415 132.220 55.675 132.390 ;
        RECT 55.875 132.220 56.125 133.545 ;
        RECT 54.415 131.450 54.585 132.220 ;
        RECT 56.295 132.050 56.675 133.280 ;
        RECT 56.865 132.820 57.115 133.545 ;
        RECT 57.315 132.820 57.645 133.280 ;
        RECT 57.845 132.950 58.095 133.545 ;
        RECT 58.745 132.980 59.075 133.545 ;
        RECT 61.145 133.040 61.475 133.545 ;
        RECT 57.445 132.780 57.645 132.820 ;
        RECT 59.770 132.810 60.020 133.025 ;
        RECT 58.265 132.780 60.020 132.810 ;
        RECT 57.445 132.640 60.020 132.780 ;
        RECT 60.220 132.870 60.550 133.025 ;
        RECT 60.220 132.700 62.010 132.870 ;
        RECT 57.445 132.610 58.435 132.640 ;
        RECT 54.755 131.880 56.675 132.050 ;
        RECT 54.755 131.650 55.765 131.880 ;
        RECT 47.800 130.385 48.050 131.130 ;
        RECT 48.225 130.960 48.950 131.130 ;
        RECT 48.620 130.670 48.950 130.960 ;
        RECT 49.170 130.385 49.470 131.405 ;
        RECT 54.415 131.280 55.630 131.450 ;
        RECT 55.935 131.380 56.335 131.710 ;
        RECT 54.010 130.385 54.260 131.110 ;
        RECT 54.440 130.650 54.770 131.280 ;
        RECT 54.950 130.385 55.120 131.110 ;
        RECT 55.300 130.650 55.630 131.280 ;
        RECT 56.505 131.110 56.675 131.880 ;
        RECT 56.885 131.300 57.275 132.470 ;
        RECT 57.445 131.130 57.615 132.610 ;
        RECT 59.770 132.530 60.020 132.640 ;
        RECT 57.785 131.430 58.045 132.440 ;
        RECT 58.215 132.110 58.625 132.440 ;
        RECT 59.275 132.190 59.525 132.470 ;
        RECT 59.770 132.360 60.515 132.530 ;
        RECT 58.215 131.440 58.385 132.110 ;
        RECT 58.805 131.940 59.035 132.080 ;
        RECT 59.275 132.020 60.175 132.190 ;
        RECT 58.555 131.610 59.035 131.940 ;
        RECT 59.625 131.860 60.175 132.020 ;
        RECT 59.205 131.440 59.455 131.850 ;
        RECT 58.215 131.270 59.455 131.440 ;
        RECT 55.800 130.385 56.130 131.110 ;
        RECT 56.300 130.780 56.675 131.110 ;
        RECT 56.890 130.960 57.615 131.130 ;
        RECT 56.890 130.670 57.220 130.960 ;
        RECT 57.790 130.385 58.040 131.130 ;
        RECT 58.215 130.650 58.600 131.270 ;
        RECT 59.625 131.100 59.795 131.860 ;
        RECT 60.345 131.690 60.515 132.360 ;
        RECT 58.770 130.385 59.100 131.100 ;
        RECT 59.270 130.800 59.795 131.100 ;
        RECT 59.965 131.520 60.515 131.690 ;
        RECT 59.965 130.970 60.215 131.520 ;
        RECT 60.685 131.350 60.855 132.700 ;
        RECT 61.375 132.620 62.010 132.700 ;
        RECT 60.385 130.970 60.855 131.350 ;
        RECT 61.025 131.375 61.205 132.425 ;
        RECT 61.375 131.875 61.545 132.620 ;
        RECT 61.715 132.095 62.045 132.450 ;
        RECT 62.240 132.045 62.570 133.545 ;
        RECT 62.740 132.165 63.070 133.055 ;
        RECT 63.240 132.775 64.395 133.105 ;
        RECT 61.375 131.545 62.410 131.875 ;
        RECT 62.740 131.430 62.910 132.165 ;
        RECT 63.240 131.985 63.410 132.775 ;
        RECT 62.580 131.375 62.910 131.430 ;
        RECT 61.025 131.205 62.910 131.375 ;
        RECT 61.025 130.865 62.410 131.035 ;
        RECT 62.580 130.965 62.910 131.205 ;
        RECT 63.080 131.815 63.410 131.985 ;
        RECT 63.080 131.145 63.250 131.815 ;
        RECT 63.725 131.645 64.055 132.605 ;
        RECT 64.225 131.985 64.395 132.775 ;
        RECT 64.565 132.745 64.895 133.545 ;
        RECT 65.080 132.745 65.445 133.205 ;
        RECT 64.565 132.220 65.105 132.555 ;
        RECT 65.275 132.325 65.445 132.745 ;
        RECT 65.615 132.495 65.945 133.545 ;
        RECT 65.275 132.155 65.950 132.325 ;
        RECT 64.225 131.815 65.610 131.985 ;
        RECT 65.280 131.655 65.610 131.815 ;
        RECT 63.450 131.315 64.180 131.645 ;
        RECT 64.350 131.485 64.680 131.645 ;
        RECT 65.780 131.485 65.950 132.155 ;
        RECT 66.145 132.015 66.315 133.205 ;
        RECT 66.485 132.185 67.185 133.280 ;
        RECT 66.145 131.685 66.695 132.015 ;
        RECT 64.350 131.315 65.950 131.485 ;
        RECT 63.080 130.895 63.840 131.145 ;
        RECT 61.025 130.800 61.195 130.865 ;
        RECT 59.270 130.630 61.195 130.800 ;
        RECT 62.240 130.725 62.410 130.865 ;
        RECT 64.010 130.725 64.180 131.315 ;
        RECT 61.675 130.385 62.070 130.695 ;
        RECT 62.240 130.555 64.180 130.725 ;
        RECT 64.505 130.385 64.835 131.145 ;
        RECT 65.375 130.685 65.705 131.315 ;
        RECT 65.935 130.385 66.185 131.145 ;
        RECT 66.365 130.650 66.695 131.685 ;
        RECT 66.925 131.430 67.185 132.185 ;
        RECT 67.355 132.120 67.685 133.545 ;
        RECT 68.005 131.550 68.575 133.545 ;
        RECT 69.295 132.230 69.625 133.545 ;
        RECT 66.925 130.650 67.255 131.430 ;
        RECT 67.435 130.385 67.685 131.430 ;
        RECT 67.940 130.385 68.270 131.105 ;
        RECT 68.980 130.385 69.550 131.885 ;
        RECT 10.200 130.215 69.720 130.385 ;
        RECT 10.370 128.715 10.940 130.215 ;
        RECT 11.650 129.495 11.980 130.215 ;
        RECT 16.555 129.510 16.885 129.950 ;
        RECT 17.055 129.620 17.745 130.215 ;
        RECT 10.295 127.055 10.625 128.370 ;
        RECT 11.345 127.055 11.915 129.050 ;
        RECT 16.555 128.480 16.795 129.510 ;
        RECT 17.915 129.340 18.245 129.950 ;
        RECT 16.965 129.170 18.245 129.340 ;
        RECT 18.445 129.170 18.805 129.950 ;
        RECT 18.985 129.620 19.300 130.215 ;
        RECT 19.480 129.450 19.730 129.950 ;
        RECT 18.975 129.280 19.730 129.450 ;
        RECT 16.965 128.670 17.355 129.170 ;
        RECT 16.555 127.320 17.015 128.480 ;
        RECT 17.185 128.350 17.355 128.670 ;
        RECT 17.525 128.520 18.235 129.000 ;
        RECT 17.185 128.180 18.015 128.350 ;
        RECT 17.185 127.055 17.515 128.010 ;
        RECT 17.685 127.320 18.015 128.180 ;
        RECT 18.445 128.270 18.615 129.170 ;
        RECT 18.975 128.950 19.145 129.280 ;
        RECT 19.960 129.240 20.290 130.215 ;
        RECT 20.625 129.875 22.030 130.045 ;
        RECT 20.625 129.790 20.955 129.875 ;
        RECT 20.700 129.320 21.300 129.570 ;
        RECT 18.785 128.610 19.145 128.950 ;
        RECT 19.315 129.070 19.645 129.110 ;
        RECT 20.700 129.070 20.870 129.320 ;
        RECT 21.520 129.270 21.690 129.705 ;
        RECT 21.860 129.610 22.030 129.875 ;
        RECT 22.200 129.780 22.450 130.215 ;
        RECT 22.760 129.855 24.035 130.025 ;
        RECT 22.760 129.610 22.930 129.855 ;
        RECT 21.860 129.440 22.930 129.610 ;
        RECT 19.315 128.900 20.870 129.070 ;
        RECT 19.315 128.780 19.645 128.900 ;
        RECT 20.140 128.610 20.470 128.730 ;
        RECT 18.785 128.440 20.470 128.610 ;
        RECT 18.445 127.320 18.805 128.270 ;
        RECT 18.980 127.055 19.310 128.270 ;
        RECT 19.510 127.600 19.760 128.440 ;
        RECT 20.140 128.060 20.470 128.440 ;
        RECT 20.700 128.590 20.870 128.900 ;
        RECT 21.040 128.930 21.350 129.150 ;
        RECT 21.520 129.100 22.590 129.270 ;
        RECT 21.040 128.760 21.740 128.930 ;
        RECT 20.700 128.420 21.400 128.590 ;
        RECT 19.990 127.055 20.320 127.780 ;
        RECT 20.680 127.395 21.010 128.250 ;
        RECT 21.230 127.565 21.400 128.420 ;
        RECT 21.570 127.675 21.740 128.760 ;
        RECT 21.910 128.175 22.080 129.100 ;
        RECT 22.260 128.885 22.590 129.100 ;
        RECT 22.250 128.345 22.550 128.675 ;
        RECT 21.910 127.845 22.185 128.175 ;
        RECT 22.380 128.015 22.550 128.345 ;
        RECT 22.760 128.550 22.930 129.440 ;
        RECT 23.100 128.890 23.365 129.685 ;
        RECT 23.865 129.570 24.035 129.855 ;
        RECT 24.205 129.740 24.535 130.215 ;
        RECT 24.705 129.875 25.555 130.045 ;
        RECT 24.705 129.570 24.875 129.875 ;
        RECT 23.865 129.400 24.875 129.570 ;
        RECT 23.545 129.060 24.100 129.230 ;
        RECT 23.100 128.720 23.760 128.890 ;
        RECT 22.760 128.220 23.420 128.550 ;
        RECT 23.590 128.015 23.760 128.720 ;
        RECT 22.380 127.845 23.760 128.015 ;
        RECT 23.400 127.675 23.760 127.845 ;
        RECT 23.930 127.675 24.100 129.060 ;
        RECT 24.270 128.275 24.550 129.175 ;
        RECT 25.045 128.950 25.215 129.705 ;
        RECT 24.760 128.620 25.215 128.950 ;
        RECT 25.385 129.340 25.555 129.875 ;
        RECT 25.725 129.510 25.975 130.215 ;
        RECT 26.155 129.340 26.405 129.950 ;
        RECT 25.385 129.170 26.405 129.340 ;
        RECT 25.385 128.750 25.845 129.170 ;
        RECT 25.045 128.480 25.215 128.620 ;
        RECT 24.270 127.945 24.650 128.275 ;
        RECT 25.045 127.675 25.505 128.480 ;
        RECT 25.675 128.350 25.845 128.750 ;
        RECT 26.015 128.520 26.395 129.000 ;
        RECT 34.370 128.715 34.940 130.215 ;
        RECT 35.650 129.495 35.980 130.215 ;
        RECT 36.210 129.195 36.510 130.215 ;
        RECT 25.675 128.180 26.405 128.350 ;
        RECT 21.570 127.505 23.230 127.675 ;
        RECT 24.270 127.505 25.505 127.675 ;
        RECT 21.570 127.395 21.740 127.505 ;
        RECT 20.680 127.225 21.740 127.395 ;
        RECT 23.060 127.335 24.440 127.505 ;
        RECT 22.390 127.055 22.720 127.335 ;
        RECT 24.610 127.055 24.945 127.335 ;
        RECT 25.175 127.320 25.505 127.505 ;
        RECT 25.705 127.055 25.875 128.010 ;
        RECT 26.075 127.320 26.405 128.180 ;
        RECT 34.295 127.055 34.625 128.370 ;
        RECT 35.345 127.055 35.915 129.050 ;
        RECT 48.290 128.715 48.860 130.215 ;
        RECT 49.570 129.495 49.900 130.215 ;
        RECT 51.115 129.170 51.365 130.215 ;
        RECT 51.545 129.170 51.875 129.950 ;
        RECT 36.210 127.055 36.510 128.095 ;
        RECT 48.215 127.055 48.545 128.370 ;
        RECT 49.265 127.055 49.835 129.050 ;
        RECT 51.115 127.055 51.445 128.480 ;
        RECT 51.615 128.415 51.875 129.170 ;
        RECT 52.105 128.915 52.435 129.950 ;
        RECT 52.615 129.455 52.865 130.215 ;
        RECT 53.095 129.285 53.425 129.915 ;
        RECT 53.965 129.455 54.295 130.215 ;
        RECT 54.620 129.875 56.560 130.045 ;
        RECT 56.730 129.905 57.125 130.215 ;
        RECT 54.620 129.285 54.790 129.875 ;
        RECT 56.390 129.735 56.560 129.875 ;
        RECT 57.605 129.800 59.530 129.970 ;
        RECT 57.605 129.735 57.775 129.800 ;
        RECT 54.960 129.455 55.720 129.705 ;
        RECT 52.850 129.115 54.450 129.285 ;
        RECT 52.105 128.585 52.655 128.915 ;
        RECT 51.615 127.320 52.315 128.415 ;
        RECT 52.485 127.395 52.655 128.585 ;
        RECT 52.850 128.445 53.020 129.115 ;
        RECT 54.120 128.955 54.450 129.115 ;
        RECT 54.620 128.955 55.350 129.285 ;
        RECT 53.190 128.785 53.520 128.945 ;
        RECT 53.190 128.615 54.575 128.785 ;
        RECT 52.850 128.275 53.525 128.445 ;
        RECT 52.855 127.055 53.185 128.105 ;
        RECT 53.355 127.855 53.525 128.275 ;
        RECT 53.695 128.045 54.235 128.380 ;
        RECT 53.355 127.395 53.720 127.855 ;
        RECT 53.905 127.055 54.235 127.855 ;
        RECT 54.405 127.825 54.575 128.615 ;
        RECT 54.745 127.995 55.075 128.955 ;
        RECT 55.550 128.785 55.720 129.455 ;
        RECT 55.390 128.615 55.720 128.785 ;
        RECT 55.890 129.395 56.220 129.635 ;
        RECT 56.390 129.565 57.775 129.735 ;
        RECT 55.890 129.225 57.775 129.395 ;
        RECT 55.890 129.170 56.220 129.225 ;
        RECT 55.390 127.825 55.560 128.615 ;
        RECT 55.890 128.435 56.060 129.170 ;
        RECT 56.390 128.725 57.425 129.055 ;
        RECT 54.405 127.495 55.560 127.825 ;
        RECT 55.730 127.545 56.060 128.435 ;
        RECT 56.230 127.055 56.560 128.555 ;
        RECT 56.755 128.150 57.085 128.505 ;
        RECT 57.255 127.980 57.425 128.725 ;
        RECT 57.595 128.175 57.775 129.225 ;
        RECT 57.945 129.250 58.415 129.630 ;
        RECT 56.790 127.900 57.425 127.980 ;
        RECT 57.945 127.900 58.115 129.250 ;
        RECT 58.585 129.080 58.835 129.630 ;
        RECT 58.285 128.910 58.835 129.080 ;
        RECT 59.005 129.500 59.530 129.800 ;
        RECT 59.700 129.500 60.030 130.215 ;
        RECT 58.285 128.240 58.455 128.910 ;
        RECT 59.005 128.740 59.175 129.500 ;
        RECT 60.200 129.330 60.585 129.950 ;
        RECT 60.760 129.470 61.010 130.215 ;
        RECT 61.580 129.640 61.910 129.930 ;
        RECT 61.185 129.470 61.910 129.640 ;
        RECT 59.345 129.160 60.585 129.330 ;
        RECT 59.345 128.750 59.595 129.160 ;
        RECT 58.625 128.580 59.175 128.740 ;
        RECT 59.765 128.660 60.245 128.990 ;
        RECT 58.625 128.410 59.525 128.580 ;
        RECT 59.765 128.520 59.995 128.660 ;
        RECT 60.415 128.490 60.585 129.160 ;
        RECT 58.285 128.070 59.030 128.240 ;
        RECT 59.275 128.130 59.525 128.410 ;
        RECT 60.175 128.160 60.585 128.490 ;
        RECT 60.755 128.160 61.015 129.170 ;
        RECT 58.780 127.960 59.030 128.070 ;
        RECT 61.185 127.990 61.355 129.470 ;
        RECT 61.525 128.130 61.915 129.300 ;
        RECT 62.130 129.195 62.430 130.215 ;
        RECT 62.690 128.715 63.260 130.215 ;
        RECT 63.970 129.495 64.300 130.215 ;
        RECT 65.005 129.490 65.380 129.820 ;
        RECT 65.550 129.490 65.880 130.215 ;
        RECT 60.365 127.960 61.355 127.990 ;
        RECT 56.790 127.730 58.580 127.900 ;
        RECT 58.250 127.575 58.580 127.730 ;
        RECT 58.780 127.820 61.355 127.960 ;
        RECT 58.780 127.790 60.535 127.820 ;
        RECT 58.780 127.575 59.030 127.790 ;
        RECT 61.155 127.780 61.355 127.820 ;
        RECT 57.325 127.055 57.655 127.560 ;
        RECT 59.725 127.055 60.055 127.620 ;
        RECT 60.705 127.055 60.955 127.650 ;
        RECT 61.155 127.320 61.485 127.780 ;
        RECT 61.685 127.055 61.935 127.780 ;
        RECT 62.130 127.055 62.430 128.095 ;
        RECT 62.615 127.055 62.945 128.370 ;
        RECT 63.665 127.055 64.235 129.050 ;
        RECT 65.005 128.720 65.175 129.490 ;
        RECT 66.050 129.320 66.380 129.950 ;
        RECT 66.560 129.490 66.730 130.215 ;
        RECT 66.910 129.320 67.240 129.950 ;
        RECT 67.420 129.490 67.670 130.215 ;
        RECT 67.940 129.495 68.270 130.215 ;
        RECT 65.345 128.890 65.745 129.220 ;
        RECT 66.050 129.150 67.265 129.320 ;
        RECT 65.915 128.720 66.925 128.950 ;
        RECT 65.005 128.550 66.925 128.720 ;
        RECT 65.005 127.320 65.385 128.550 ;
        RECT 67.095 128.380 67.265 129.150 ;
        RECT 65.555 127.055 65.805 128.380 ;
        RECT 66.005 128.210 67.265 128.380 ;
        RECT 66.005 127.320 66.335 128.210 ;
        RECT 66.535 127.055 66.785 128.040 ;
        RECT 66.985 127.320 67.265 128.210 ;
        RECT 67.435 127.055 67.685 128.480 ;
        RECT 68.005 127.055 68.575 129.050 ;
        RECT 68.980 128.715 69.550 130.215 ;
        RECT 69.295 127.055 69.625 128.370 ;
        RECT 10.200 126.885 69.720 127.055 ;
        RECT 10.295 125.570 10.625 126.885 ;
        RECT 10.370 123.725 10.940 125.225 ;
        RECT 11.345 124.890 11.915 126.885 ;
        RECT 12.705 125.460 13.035 126.885 ;
        RECT 12.705 124.820 13.035 125.190 ;
        RECT 13.205 124.820 13.435 126.620 ;
        RECT 13.605 125.460 13.935 126.885 ;
        RECT 14.125 125.460 14.515 126.620 ;
        RECT 14.685 126.100 15.015 126.620 ;
        RECT 15.185 126.290 15.625 126.885 ;
        RECT 15.795 126.100 16.125 126.620 ;
        RECT 14.685 125.930 16.125 126.100 ;
        RECT 16.355 125.760 16.935 126.620 ;
        RECT 14.685 125.590 16.935 125.760 ;
        RECT 13.605 124.820 13.935 125.190 ;
        RECT 13.265 124.650 13.435 124.820 ;
        RECT 14.125 124.790 14.295 125.460 ;
        RECT 14.685 125.290 14.855 125.590 ;
        RECT 14.465 124.960 14.855 125.290 ;
        RECT 15.035 125.335 15.365 125.420 ;
        RECT 16.115 125.335 16.285 125.390 ;
        RECT 15.035 125.005 16.595 125.335 ;
        RECT 15.035 124.990 15.365 125.005 ;
        RECT 11.650 123.725 11.980 124.445 ;
        RECT 12.730 123.725 13.060 124.650 ;
        RECT 13.265 124.480 13.885 124.650 ;
        RECT 14.125 124.620 15.355 124.790 ;
        RECT 13.550 123.990 13.880 124.480 ;
        RECT 14.340 123.725 14.670 124.385 ;
        RECT 14.910 124.055 15.355 124.620 ;
        RECT 15.730 123.725 16.060 124.835 ;
        RECT 16.765 124.680 16.935 125.590 ;
        RECT 17.225 125.580 17.555 126.885 ;
        RECT 17.975 125.570 18.305 126.885 ;
        RECT 17.105 124.820 17.775 125.255 ;
        RECT 16.240 124.350 16.935 124.680 ;
        RECT 17.105 123.725 17.705 124.630 ;
        RECT 18.050 123.725 18.620 125.225 ;
        RECT 19.025 124.890 19.595 126.885 ;
        RECT 19.915 125.460 20.375 126.620 ;
        RECT 20.545 125.930 20.875 126.885 ;
        RECT 21.045 125.760 21.375 126.620 ;
        RECT 23.250 125.845 23.550 126.885 ;
        RECT 20.545 125.590 21.375 125.760 ;
        RECT 19.330 123.725 19.660 124.445 ;
        RECT 19.915 124.430 20.155 125.460 ;
        RECT 20.545 125.270 20.715 125.590 ;
        RECT 23.735 125.570 24.065 126.885 ;
        RECT 20.325 124.770 20.715 125.270 ;
        RECT 20.885 124.940 21.595 125.420 ;
        RECT 20.325 124.600 21.605 124.770 ;
        RECT 19.915 123.990 20.245 124.430 ;
        RECT 20.415 123.725 21.105 124.320 ;
        RECT 21.275 123.990 21.605 124.600 ;
        RECT 23.250 123.725 23.550 124.745 ;
        RECT 23.810 123.725 24.380 125.225 ;
        RECT 24.785 124.890 25.355 126.885 ;
        RECT 25.675 125.460 26.135 126.620 ;
        RECT 26.305 125.930 26.635 126.885 ;
        RECT 26.805 125.760 27.135 126.620 ;
        RECT 26.305 125.590 27.135 125.760 ;
        RECT 25.090 123.725 25.420 124.445 ;
        RECT 25.675 124.430 25.915 125.460 ;
        RECT 26.305 125.270 26.475 125.590 ;
        RECT 27.595 125.460 28.055 126.620 ;
        RECT 28.225 125.930 28.555 126.885 ;
        RECT 28.725 125.760 29.055 126.620 ;
        RECT 30.465 126.160 30.715 126.885 ;
        RECT 30.915 126.160 31.245 126.620 ;
        RECT 31.445 126.290 31.695 126.885 ;
        RECT 32.345 126.320 32.675 126.885 ;
        RECT 34.745 126.380 35.075 126.885 ;
        RECT 31.045 126.120 31.245 126.160 ;
        RECT 33.370 126.150 33.620 126.365 ;
        RECT 31.865 126.120 33.620 126.150 ;
        RECT 31.045 125.980 33.620 126.120 ;
        RECT 33.820 126.210 34.150 126.365 ;
        RECT 33.820 126.040 35.610 126.210 ;
        RECT 31.045 125.950 32.035 125.980 ;
        RECT 28.225 125.590 29.055 125.760 ;
        RECT 26.085 124.770 26.475 125.270 ;
        RECT 26.645 124.940 27.355 125.420 ;
        RECT 26.085 124.600 27.365 124.770 ;
        RECT 25.675 123.990 26.005 124.430 ;
        RECT 26.175 123.725 26.865 124.320 ;
        RECT 27.035 123.990 27.365 124.600 ;
        RECT 27.595 124.430 27.835 125.460 ;
        RECT 28.225 125.270 28.395 125.590 ;
        RECT 28.005 124.770 28.395 125.270 ;
        RECT 28.565 124.940 29.275 125.420 ;
        RECT 28.005 124.600 29.285 124.770 ;
        RECT 30.485 124.640 30.875 125.810 ;
        RECT 27.595 123.990 27.925 124.430 ;
        RECT 28.095 123.725 28.785 124.320 ;
        RECT 28.955 123.990 29.285 124.600 ;
        RECT 31.045 124.470 31.215 125.950 ;
        RECT 33.370 125.870 33.620 125.980 ;
        RECT 31.385 124.770 31.645 125.780 ;
        RECT 31.815 125.450 32.225 125.780 ;
        RECT 32.875 125.530 33.125 125.810 ;
        RECT 33.370 125.700 34.115 125.870 ;
        RECT 31.815 124.780 31.985 125.450 ;
        RECT 32.405 125.280 32.635 125.420 ;
        RECT 32.875 125.360 33.775 125.530 ;
        RECT 32.155 124.950 32.635 125.280 ;
        RECT 33.225 125.200 33.775 125.360 ;
        RECT 32.805 124.780 33.055 125.190 ;
        RECT 31.815 124.610 33.055 124.780 ;
        RECT 30.490 124.300 31.215 124.470 ;
        RECT 30.490 124.010 30.820 124.300 ;
        RECT 31.390 123.725 31.640 124.470 ;
        RECT 31.815 123.990 32.200 124.610 ;
        RECT 33.225 124.440 33.395 125.200 ;
        RECT 33.945 125.030 34.115 125.700 ;
        RECT 32.370 123.725 32.700 124.440 ;
        RECT 32.870 124.140 33.395 124.440 ;
        RECT 33.565 124.860 34.115 125.030 ;
        RECT 33.565 124.310 33.815 124.860 ;
        RECT 34.285 124.690 34.455 126.040 ;
        RECT 34.975 125.960 35.610 126.040 ;
        RECT 33.985 124.310 34.455 124.690 ;
        RECT 34.625 124.715 34.805 125.765 ;
        RECT 34.975 125.215 35.145 125.960 ;
        RECT 35.315 125.435 35.645 125.790 ;
        RECT 35.840 125.385 36.170 126.885 ;
        RECT 36.340 125.505 36.670 126.395 ;
        RECT 36.840 126.115 37.995 126.445 ;
        RECT 34.975 124.885 36.010 125.215 ;
        RECT 36.340 124.770 36.510 125.505 ;
        RECT 36.840 125.325 37.010 126.115 ;
        RECT 36.180 124.715 36.510 124.770 ;
        RECT 34.625 124.545 36.510 124.715 ;
        RECT 34.625 124.205 36.010 124.375 ;
        RECT 36.180 124.305 36.510 124.545 ;
        RECT 36.680 125.155 37.010 125.325 ;
        RECT 36.680 124.485 36.850 125.155 ;
        RECT 37.325 124.985 37.655 125.945 ;
        RECT 37.825 125.325 37.995 126.115 ;
        RECT 38.165 126.085 38.495 126.885 ;
        RECT 38.680 126.085 39.045 126.545 ;
        RECT 38.165 125.560 38.705 125.895 ;
        RECT 38.875 125.665 39.045 126.085 ;
        RECT 39.215 125.835 39.545 126.885 ;
        RECT 38.875 125.495 39.550 125.665 ;
        RECT 37.825 125.155 39.210 125.325 ;
        RECT 38.880 124.995 39.210 125.155 ;
        RECT 37.050 124.655 37.780 124.985 ;
        RECT 37.950 124.825 38.280 124.985 ;
        RECT 39.380 124.825 39.550 125.495 ;
        RECT 39.745 125.355 39.915 126.545 ;
        RECT 40.085 125.525 40.785 126.620 ;
        RECT 39.745 125.025 40.295 125.355 ;
        RECT 37.950 124.655 39.550 124.825 ;
        RECT 36.680 124.235 37.440 124.485 ;
        RECT 34.625 124.140 34.795 124.205 ;
        RECT 32.870 123.970 34.795 124.140 ;
        RECT 35.840 124.065 36.010 124.205 ;
        RECT 37.610 124.065 37.780 124.655 ;
        RECT 35.275 123.725 35.670 124.035 ;
        RECT 35.840 123.895 37.780 124.065 ;
        RECT 38.105 123.725 38.435 124.485 ;
        RECT 38.975 124.025 39.305 124.655 ;
        RECT 39.535 123.725 39.785 124.485 ;
        RECT 39.965 123.990 40.295 125.025 ;
        RECT 40.525 124.770 40.785 125.525 ;
        RECT 40.955 125.460 41.285 126.885 ;
        RECT 45.835 126.375 46.545 126.885 ;
        RECT 45.835 125.460 46.140 126.375 ;
        RECT 47.115 126.300 47.445 126.885 ;
        RECT 47.650 126.130 48.005 126.520 ;
        RECT 46.325 125.960 48.005 126.130 ;
        RECT 46.325 125.270 46.495 125.960 ;
        RECT 45.825 124.940 46.495 125.270 ;
        RECT 46.665 124.820 47.035 125.790 ;
        RECT 47.205 124.820 47.375 125.960 ;
        RECT 47.650 125.590 48.005 125.960 ;
        RECT 49.170 125.845 49.470 126.885 ;
        RECT 49.665 126.160 49.915 126.885 ;
        RECT 50.115 126.160 50.445 126.620 ;
        RECT 50.645 126.290 50.895 126.885 ;
        RECT 51.545 126.320 51.875 126.885 ;
        RECT 53.945 126.380 54.275 126.885 ;
        RECT 50.245 126.120 50.445 126.160 ;
        RECT 52.570 126.150 52.820 126.365 ;
        RECT 51.065 126.120 52.820 126.150 ;
        RECT 50.245 125.980 52.820 126.120 ;
        RECT 53.020 126.210 53.350 126.365 ;
        RECT 53.020 126.040 54.810 126.210 ;
        RECT 50.245 125.950 51.235 125.980 ;
        RECT 47.545 124.990 47.995 125.420 ;
        RECT 40.525 123.990 40.855 124.770 ;
        RECT 41.035 123.725 41.285 124.770 ;
        RECT 46.235 123.725 46.485 124.770 ;
        RECT 46.665 123.990 46.995 124.820 ;
        RECT 47.205 124.650 48.005 124.820 ;
        RECT 47.165 123.725 47.495 124.480 ;
        RECT 47.675 124.090 48.005 124.650 ;
        RECT 49.170 123.725 49.470 124.745 ;
        RECT 49.685 124.640 50.075 125.810 ;
        RECT 50.245 124.470 50.415 125.950 ;
        RECT 52.570 125.870 52.820 125.980 ;
        RECT 50.585 124.770 50.845 125.780 ;
        RECT 51.015 125.450 51.425 125.780 ;
        RECT 52.075 125.530 52.325 125.810 ;
        RECT 52.570 125.700 53.315 125.870 ;
        RECT 51.015 124.780 51.185 125.450 ;
        RECT 51.605 125.280 51.835 125.420 ;
        RECT 52.075 125.360 52.975 125.530 ;
        RECT 51.355 124.950 51.835 125.280 ;
        RECT 52.425 125.200 52.975 125.360 ;
        RECT 52.005 124.780 52.255 125.190 ;
        RECT 51.015 124.610 52.255 124.780 ;
        RECT 49.690 124.300 50.415 124.470 ;
        RECT 49.690 124.010 50.020 124.300 ;
        RECT 50.590 123.725 50.840 124.470 ;
        RECT 51.015 123.990 51.400 124.610 ;
        RECT 52.425 124.440 52.595 125.200 ;
        RECT 53.145 125.030 53.315 125.700 ;
        RECT 51.570 123.725 51.900 124.440 ;
        RECT 52.070 124.140 52.595 124.440 ;
        RECT 52.765 124.860 53.315 125.030 ;
        RECT 52.765 124.310 53.015 124.860 ;
        RECT 53.485 124.690 53.655 126.040 ;
        RECT 54.175 125.960 54.810 126.040 ;
        RECT 53.185 124.310 53.655 124.690 ;
        RECT 53.825 124.715 54.005 125.765 ;
        RECT 54.175 125.215 54.345 125.960 ;
        RECT 54.515 125.435 54.845 125.790 ;
        RECT 55.040 125.385 55.370 126.885 ;
        RECT 55.540 125.505 55.870 126.395 ;
        RECT 56.040 126.115 57.195 126.445 ;
        RECT 54.175 124.885 55.210 125.215 ;
        RECT 55.540 124.770 55.710 125.505 ;
        RECT 56.040 125.325 56.210 126.115 ;
        RECT 55.380 124.715 55.710 124.770 ;
        RECT 53.825 124.545 55.710 124.715 ;
        RECT 53.825 124.205 55.210 124.375 ;
        RECT 55.380 124.305 55.710 124.545 ;
        RECT 55.880 125.155 56.210 125.325 ;
        RECT 55.880 124.485 56.050 125.155 ;
        RECT 56.525 124.985 56.855 125.945 ;
        RECT 57.025 125.325 57.195 126.115 ;
        RECT 57.365 126.085 57.695 126.885 ;
        RECT 57.880 126.085 58.245 126.545 ;
        RECT 57.365 125.560 57.905 125.895 ;
        RECT 58.075 125.665 58.245 126.085 ;
        RECT 58.415 125.835 58.745 126.885 ;
        RECT 58.075 125.495 58.750 125.665 ;
        RECT 57.025 125.155 58.410 125.325 ;
        RECT 58.080 124.995 58.410 125.155 ;
        RECT 56.250 124.655 56.980 124.985 ;
        RECT 57.150 124.825 57.480 124.985 ;
        RECT 58.580 124.825 58.750 125.495 ;
        RECT 58.945 125.355 59.115 126.545 ;
        RECT 59.285 125.525 59.985 126.620 ;
        RECT 58.945 125.025 59.495 125.355 ;
        RECT 57.150 124.655 58.750 124.825 ;
        RECT 55.880 124.235 56.640 124.485 ;
        RECT 53.825 124.140 53.995 124.205 ;
        RECT 52.070 123.970 53.995 124.140 ;
        RECT 55.040 124.065 55.210 124.205 ;
        RECT 56.810 124.065 56.980 124.655 ;
        RECT 54.475 123.725 54.870 124.035 ;
        RECT 55.040 123.895 56.980 124.065 ;
        RECT 57.305 123.725 57.635 124.485 ;
        RECT 58.175 124.025 58.505 124.655 ;
        RECT 58.735 123.725 58.985 124.485 ;
        RECT 59.165 123.990 59.495 125.025 ;
        RECT 59.725 124.770 59.985 125.525 ;
        RECT 60.155 125.460 60.485 126.885 ;
        RECT 62.125 125.390 62.505 126.620 ;
        RECT 62.675 125.560 62.925 126.885 ;
        RECT 63.125 125.730 63.455 126.620 ;
        RECT 63.655 125.900 63.905 126.885 ;
        RECT 64.105 125.730 64.385 126.620 ;
        RECT 63.125 125.560 64.385 125.730 ;
        RECT 62.125 125.220 64.045 125.390 ;
        RECT 59.725 123.990 60.055 124.770 ;
        RECT 60.235 123.725 60.485 124.770 ;
        RECT 62.125 124.450 62.295 125.220 ;
        RECT 62.465 124.720 62.865 125.050 ;
        RECT 63.035 124.990 64.045 125.220 ;
        RECT 64.215 124.790 64.385 125.560 ;
        RECT 64.555 125.460 64.805 126.885 ;
        RECT 63.170 124.620 64.385 124.790 ;
        RECT 65.005 125.390 65.385 126.620 ;
        RECT 65.555 125.560 65.805 126.885 ;
        RECT 66.005 125.730 66.335 126.620 ;
        RECT 66.535 125.900 66.785 126.885 ;
        RECT 66.985 125.730 67.265 126.620 ;
        RECT 66.005 125.560 67.265 125.730 ;
        RECT 65.005 125.220 66.925 125.390 ;
        RECT 62.125 124.120 62.500 124.450 ;
        RECT 62.670 123.725 63.000 124.450 ;
        RECT 63.170 123.990 63.500 124.620 ;
        RECT 63.680 123.725 63.850 124.450 ;
        RECT 64.030 123.990 64.360 124.620 ;
        RECT 65.005 124.450 65.175 125.220 ;
        RECT 65.345 124.720 65.745 125.050 ;
        RECT 65.915 124.990 66.925 125.220 ;
        RECT 67.095 124.790 67.265 125.560 ;
        RECT 67.435 125.460 67.685 126.885 ;
        RECT 68.005 124.890 68.575 126.885 ;
        RECT 69.295 125.570 69.625 126.885 ;
        RECT 66.050 124.620 67.265 124.790 ;
        RECT 64.540 123.725 64.790 124.450 ;
        RECT 65.005 124.120 65.380 124.450 ;
        RECT 65.550 123.725 65.880 124.450 ;
        RECT 66.050 123.990 66.380 124.620 ;
        RECT 66.560 123.725 66.730 124.450 ;
        RECT 66.910 123.990 67.240 124.620 ;
        RECT 67.420 123.725 67.670 124.450 ;
        RECT 67.940 123.725 68.270 124.445 ;
        RECT 68.980 123.725 69.550 125.225 ;
        RECT 10.200 123.555 69.720 123.725 ;
        RECT 10.370 122.055 10.940 123.555 ;
        RECT 11.650 122.835 11.980 123.555 ;
        RECT 10.295 120.395 10.625 121.710 ;
        RECT 11.345 120.395 11.915 122.390 ;
        RECT 12.290 122.055 12.860 123.555 ;
        RECT 13.570 122.835 13.900 123.555 ;
        RECT 14.155 122.680 14.405 123.290 ;
        RECT 14.585 122.850 14.835 123.555 ;
        RECT 15.005 123.215 15.855 123.385 ;
        RECT 15.005 122.680 15.175 123.215 ;
        RECT 14.155 122.510 15.175 122.680 ;
        RECT 12.215 120.395 12.545 121.710 ;
        RECT 13.265 120.395 13.835 122.390 ;
        RECT 14.165 121.860 14.545 122.340 ;
        RECT 14.715 122.090 15.175 122.510 ;
        RECT 15.345 122.290 15.515 123.045 ;
        RECT 15.685 122.910 15.855 123.215 ;
        RECT 16.025 123.080 16.355 123.555 ;
        RECT 16.525 123.195 17.800 123.365 ;
        RECT 16.525 122.910 16.695 123.195 ;
        RECT 15.685 122.740 16.695 122.910 ;
        RECT 14.715 121.690 14.885 122.090 ;
        RECT 15.345 121.960 15.800 122.290 ;
        RECT 15.345 121.820 15.515 121.960 ;
        RECT 14.155 121.520 14.885 121.690 ;
        RECT 14.155 120.660 14.485 121.520 ;
        RECT 14.685 120.395 14.855 121.350 ;
        RECT 15.055 121.015 15.515 121.820 ;
        RECT 16.010 121.615 16.290 122.515 ;
        RECT 15.910 121.285 16.290 121.615 ;
        RECT 16.460 122.400 17.015 122.570 ;
        RECT 16.460 121.015 16.630 122.400 ;
        RECT 17.195 122.230 17.460 123.025 ;
        RECT 16.800 122.060 17.460 122.230 ;
        RECT 17.630 122.950 17.800 123.195 ;
        RECT 18.110 123.120 18.360 123.555 ;
        RECT 18.530 123.215 19.935 123.385 ;
        RECT 18.530 122.950 18.700 123.215 ;
        RECT 19.605 123.130 19.935 123.215 ;
        RECT 17.630 122.780 18.700 122.950 ;
        RECT 16.800 121.355 16.970 122.060 ;
        RECT 17.630 121.890 17.800 122.780 ;
        RECT 18.870 122.610 19.040 123.045 ;
        RECT 19.260 122.660 19.860 122.910 ;
        RECT 17.970 122.440 19.040 122.610 ;
        RECT 17.970 122.225 18.300 122.440 ;
        RECT 17.140 121.560 17.800 121.890 ;
        RECT 18.010 121.685 18.310 122.015 ;
        RECT 18.010 121.355 18.180 121.685 ;
        RECT 18.480 121.515 18.650 122.440 ;
        RECT 19.210 122.270 19.520 122.490 ;
        RECT 16.800 121.185 18.180 121.355 ;
        RECT 18.375 121.185 18.650 121.515 ;
        RECT 18.820 122.100 19.520 122.270 ;
        RECT 19.690 122.410 19.860 122.660 ;
        RECT 20.270 122.580 20.600 123.555 ;
        RECT 20.830 122.790 21.080 123.290 ;
        RECT 21.260 122.960 21.575 123.555 ;
        RECT 20.830 122.620 21.585 122.790 ;
        RECT 20.915 122.410 21.245 122.450 ;
        RECT 19.690 122.240 21.245 122.410 ;
        RECT 16.800 121.015 17.160 121.185 ;
        RECT 18.820 121.015 18.990 122.100 ;
        RECT 19.690 121.930 19.860 122.240 ;
        RECT 20.915 122.120 21.245 122.240 ;
        RECT 21.415 122.290 21.585 122.620 ;
        RECT 21.755 122.510 22.115 123.290 ;
        RECT 22.305 123.070 23.515 123.385 ;
        RECT 23.285 122.970 23.515 123.070 ;
        RECT 15.055 120.845 16.290 121.015 ;
        RECT 17.330 120.845 18.990 121.015 ;
        RECT 19.160 121.760 19.860 121.930 ;
        RECT 20.090 121.950 20.420 122.070 ;
        RECT 21.415 121.950 21.775 122.290 ;
        RECT 20.090 121.780 21.775 121.950 ;
        RECT 19.160 120.905 19.330 121.760 ;
        RECT 15.055 120.660 15.385 120.845 ;
        RECT 16.120 120.675 17.500 120.845 ;
        RECT 18.820 120.735 18.990 120.845 ;
        RECT 19.550 120.735 19.880 121.590 ;
        RECT 20.090 121.400 20.420 121.780 ;
        RECT 15.615 120.395 15.950 120.675 ;
        RECT 17.840 120.395 18.170 120.675 ;
        RECT 18.820 120.565 19.880 120.735 ;
        RECT 20.240 120.395 20.570 121.120 ;
        RECT 20.800 120.940 21.050 121.780 ;
        RECT 21.945 121.610 22.115 122.510 ;
        RECT 21.250 120.395 21.580 121.610 ;
        RECT 21.755 120.660 22.115 121.610 ;
        RECT 22.315 121.690 22.680 122.900 ;
        RECT 23.895 122.460 24.225 123.555 ;
        RECT 24.395 122.630 24.725 123.160 ;
        RECT 24.395 122.460 24.965 122.630 ;
        RECT 25.195 122.510 25.445 123.555 ;
        RECT 25.625 122.510 25.955 123.290 ;
        RECT 23.045 121.860 23.515 122.460 ;
        RECT 23.685 121.860 24.015 122.190 ;
        RECT 24.270 121.960 24.600 122.290 ;
        RECT 24.270 121.690 24.440 121.960 ;
        RECT 24.795 121.790 24.965 122.460 ;
        RECT 22.315 121.520 24.440 121.690 ;
        RECT 22.315 120.790 22.645 121.520 ;
        RECT 22.815 120.395 23.145 121.350 ;
        RECT 23.315 120.790 23.600 121.520 ;
        RECT 23.770 120.395 24.510 121.350 ;
        RECT 24.680 120.660 24.965 121.790 ;
        RECT 25.195 120.395 25.525 121.820 ;
        RECT 25.695 121.755 25.955 122.510 ;
        RECT 26.185 122.255 26.515 123.290 ;
        RECT 26.695 122.795 26.945 123.555 ;
        RECT 27.175 122.625 27.505 123.255 ;
        RECT 28.045 122.795 28.375 123.555 ;
        RECT 28.700 123.215 30.640 123.385 ;
        RECT 30.810 123.245 31.205 123.555 ;
        RECT 28.700 122.625 28.870 123.215 ;
        RECT 30.470 123.075 30.640 123.215 ;
        RECT 31.685 123.140 33.610 123.310 ;
        RECT 31.685 123.075 31.855 123.140 ;
        RECT 29.040 122.795 29.800 123.045 ;
        RECT 26.930 122.455 28.530 122.625 ;
        RECT 26.185 121.925 26.735 122.255 ;
        RECT 25.695 120.660 26.395 121.755 ;
        RECT 26.565 120.735 26.735 121.925 ;
        RECT 26.930 121.785 27.100 122.455 ;
        RECT 28.200 122.295 28.530 122.455 ;
        RECT 28.700 122.295 29.430 122.625 ;
        RECT 27.270 122.125 27.600 122.285 ;
        RECT 27.270 121.955 28.655 122.125 ;
        RECT 26.930 121.615 27.605 121.785 ;
        RECT 26.935 120.395 27.265 121.445 ;
        RECT 27.435 121.195 27.605 121.615 ;
        RECT 27.775 121.385 28.315 121.720 ;
        RECT 27.435 120.735 27.800 121.195 ;
        RECT 27.985 120.395 28.315 121.195 ;
        RECT 28.485 121.165 28.655 121.955 ;
        RECT 28.825 121.335 29.155 122.295 ;
        RECT 29.630 122.125 29.800 122.795 ;
        RECT 29.470 121.955 29.800 122.125 ;
        RECT 29.970 122.735 30.300 122.975 ;
        RECT 30.470 122.905 31.855 123.075 ;
        RECT 29.970 122.565 31.855 122.735 ;
        RECT 29.970 122.510 30.300 122.565 ;
        RECT 29.470 121.165 29.640 121.955 ;
        RECT 29.970 121.775 30.140 122.510 ;
        RECT 30.470 122.065 31.505 122.395 ;
        RECT 28.485 120.835 29.640 121.165 ;
        RECT 29.810 120.885 30.140 121.775 ;
        RECT 30.310 120.395 30.640 121.895 ;
        RECT 30.835 121.490 31.165 121.845 ;
        RECT 31.335 121.320 31.505 122.065 ;
        RECT 31.675 121.515 31.855 122.565 ;
        RECT 32.025 122.590 32.495 122.970 ;
        RECT 30.870 121.240 31.505 121.320 ;
        RECT 32.025 121.240 32.195 122.590 ;
        RECT 32.665 122.420 32.915 122.970 ;
        RECT 32.365 122.250 32.915 122.420 ;
        RECT 33.085 122.840 33.610 123.140 ;
        RECT 33.780 122.840 34.110 123.555 ;
        RECT 32.365 121.580 32.535 122.250 ;
        RECT 33.085 122.080 33.255 122.840 ;
        RECT 34.280 122.670 34.665 123.290 ;
        RECT 34.840 122.810 35.090 123.555 ;
        RECT 35.660 122.980 35.990 123.270 ;
        RECT 35.265 122.810 35.990 122.980 ;
        RECT 33.425 122.500 34.665 122.670 ;
        RECT 33.425 122.090 33.675 122.500 ;
        RECT 32.705 121.920 33.255 122.080 ;
        RECT 33.845 122.000 34.325 122.330 ;
        RECT 32.705 121.750 33.605 121.920 ;
        RECT 33.845 121.860 34.075 122.000 ;
        RECT 34.495 121.830 34.665 122.500 ;
        RECT 32.365 121.410 33.110 121.580 ;
        RECT 33.355 121.470 33.605 121.750 ;
        RECT 34.255 121.500 34.665 121.830 ;
        RECT 34.835 121.500 35.095 122.510 ;
        RECT 32.860 121.300 33.110 121.410 ;
        RECT 35.265 121.330 35.435 122.810 ;
        RECT 35.605 121.470 35.995 122.640 ;
        RECT 36.210 122.535 36.510 123.555 ;
        RECT 36.715 122.630 37.045 123.190 ;
        RECT 37.225 122.800 37.555 123.555 ;
        RECT 36.715 122.460 37.515 122.630 ;
        RECT 37.725 122.460 38.055 123.290 ;
        RECT 38.235 122.510 38.485 123.555 ;
        RECT 44.395 122.850 44.725 123.290 ;
        RECT 44.895 122.960 45.585 123.555 ;
        RECT 36.725 121.860 37.175 122.290 ;
        RECT 34.445 121.300 35.435 121.330 ;
        RECT 30.870 121.070 32.660 121.240 ;
        RECT 32.330 120.915 32.660 121.070 ;
        RECT 32.860 121.160 35.435 121.300 ;
        RECT 32.860 121.130 34.615 121.160 ;
        RECT 32.860 120.915 33.110 121.130 ;
        RECT 35.235 121.120 35.435 121.160 ;
        RECT 31.405 120.395 31.735 120.900 ;
        RECT 33.805 120.395 34.135 120.960 ;
        RECT 34.785 120.395 35.035 120.990 ;
        RECT 35.235 120.660 35.565 121.120 ;
        RECT 35.765 120.395 36.015 121.120 ;
        RECT 36.210 120.395 36.510 121.435 ;
        RECT 36.715 121.320 37.070 121.690 ;
        RECT 37.345 121.320 37.515 122.460 ;
        RECT 37.685 121.490 38.055 122.460 ;
        RECT 38.225 122.010 38.895 122.340 ;
        RECT 38.225 121.320 38.395 122.010 ;
        RECT 44.395 121.820 44.635 122.850 ;
        RECT 45.755 122.680 46.085 123.290 ;
        RECT 46.330 122.980 46.660 123.270 ;
        RECT 46.330 122.810 47.055 122.980 ;
        RECT 47.230 122.810 47.480 123.555 ;
        RECT 44.805 122.510 46.085 122.680 ;
        RECT 44.805 122.010 45.195 122.510 ;
        RECT 36.715 121.150 38.395 121.320 ;
        RECT 36.715 120.760 37.070 121.150 ;
        RECT 37.275 120.395 37.605 120.980 ;
        RECT 38.580 120.905 38.885 121.820 ;
        RECT 38.175 120.395 38.885 120.905 ;
        RECT 44.395 120.660 44.855 121.820 ;
        RECT 45.025 121.690 45.195 122.010 ;
        RECT 45.365 121.860 46.075 122.340 ;
        RECT 45.025 121.520 45.855 121.690 ;
        RECT 45.025 120.395 45.355 121.350 ;
        RECT 45.525 120.660 45.855 121.520 ;
        RECT 46.325 121.470 46.715 122.640 ;
        RECT 46.885 121.330 47.055 122.810 ;
        RECT 47.655 122.670 48.040 123.290 ;
        RECT 48.210 122.840 48.540 123.555 ;
        RECT 48.710 123.140 50.635 123.310 ;
        RECT 51.115 123.245 51.510 123.555 ;
        RECT 48.710 122.840 49.235 123.140 ;
        RECT 50.465 123.075 50.635 123.140 ;
        RECT 51.680 123.215 53.620 123.385 ;
        RECT 51.680 123.075 51.850 123.215 ;
        RECT 47.225 121.500 47.485 122.510 ;
        RECT 47.655 122.500 48.895 122.670 ;
        RECT 47.655 121.830 47.825 122.500 ;
        RECT 47.995 122.000 48.475 122.330 ;
        RECT 48.645 122.090 48.895 122.500 ;
        RECT 48.245 121.860 48.475 122.000 ;
        RECT 49.065 122.080 49.235 122.840 ;
        RECT 49.405 122.420 49.655 122.970 ;
        RECT 49.825 122.590 50.295 122.970 ;
        RECT 50.465 122.905 51.850 123.075 ;
        RECT 52.020 122.735 52.350 122.975 ;
        RECT 49.405 122.250 49.955 122.420 ;
        RECT 49.065 121.920 49.615 122.080 ;
        RECT 47.655 121.500 48.065 121.830 ;
        RECT 48.715 121.750 49.615 121.920 ;
        RECT 48.715 121.470 48.965 121.750 ;
        RECT 49.785 121.580 49.955 122.250 ;
        RECT 49.210 121.410 49.955 121.580 ;
        RECT 46.885 121.300 47.875 121.330 ;
        RECT 49.210 121.300 49.460 121.410 ;
        RECT 46.885 121.160 49.460 121.300 ;
        RECT 50.125 121.240 50.295 122.590 ;
        RECT 50.465 122.565 52.350 122.735 ;
        RECT 50.465 121.515 50.645 122.565 ;
        RECT 52.020 122.510 52.350 122.565 ;
        RECT 50.815 122.065 51.850 122.395 ;
        RECT 50.815 121.320 50.985 122.065 ;
        RECT 51.155 121.490 51.485 121.845 ;
        RECT 50.815 121.240 51.450 121.320 ;
        RECT 46.885 121.120 47.085 121.160 ;
        RECT 47.705 121.130 49.460 121.160 ;
        RECT 46.305 120.395 46.555 121.120 ;
        RECT 46.755 120.660 47.085 121.120 ;
        RECT 47.285 120.395 47.535 120.990 ;
        RECT 48.185 120.395 48.515 120.960 ;
        RECT 49.210 120.915 49.460 121.130 ;
        RECT 49.660 121.070 51.450 121.240 ;
        RECT 49.660 120.915 49.990 121.070 ;
        RECT 50.585 120.395 50.915 120.900 ;
        RECT 51.680 120.395 52.010 121.895 ;
        RECT 52.180 121.775 52.350 122.510 ;
        RECT 52.520 122.795 53.280 123.045 ;
        RECT 52.520 122.125 52.690 122.795 ;
        RECT 53.450 122.625 53.620 123.215 ;
        RECT 53.945 122.795 54.275 123.555 ;
        RECT 54.815 122.625 55.145 123.255 ;
        RECT 55.375 122.795 55.625 123.555 ;
        RECT 52.890 122.295 53.620 122.625 ;
        RECT 53.790 122.455 55.390 122.625 ;
        RECT 53.790 122.295 54.120 122.455 ;
        RECT 52.520 121.955 52.850 122.125 ;
        RECT 52.180 120.885 52.510 121.775 ;
        RECT 52.680 121.165 52.850 121.955 ;
        RECT 53.165 121.335 53.495 122.295 ;
        RECT 54.720 122.125 55.050 122.285 ;
        RECT 53.665 121.955 55.050 122.125 ;
        RECT 53.665 121.165 53.835 121.955 ;
        RECT 55.220 121.785 55.390 122.455 ;
        RECT 55.805 122.255 56.135 123.290 ;
        RECT 54.005 121.385 54.545 121.720 ;
        RECT 54.715 121.615 55.390 121.785 ;
        RECT 55.585 121.925 56.135 122.255 ;
        RECT 56.365 122.510 56.695 123.290 ;
        RECT 56.875 122.510 57.125 123.555 ;
        RECT 62.130 122.535 62.430 123.555 ;
        RECT 54.715 121.195 54.885 121.615 ;
        RECT 52.680 120.835 53.835 121.165 ;
        RECT 54.005 120.395 54.335 121.195 ;
        RECT 54.520 120.735 54.885 121.195 ;
        RECT 55.055 120.395 55.385 121.445 ;
        RECT 55.585 120.735 55.755 121.925 ;
        RECT 56.365 121.755 56.625 122.510 ;
        RECT 62.690 122.055 63.260 123.555 ;
        RECT 63.970 122.835 64.300 123.555 ;
        RECT 65.005 122.830 65.380 123.160 ;
        RECT 65.550 122.830 65.880 123.555 ;
        RECT 55.925 120.660 56.625 121.755 ;
        RECT 56.795 120.395 57.125 121.820 ;
        RECT 62.130 120.395 62.430 121.435 ;
        RECT 62.615 120.395 62.945 121.710 ;
        RECT 63.665 120.395 64.235 122.390 ;
        RECT 65.005 122.060 65.175 122.830 ;
        RECT 66.050 122.660 66.380 123.290 ;
        RECT 66.560 122.830 66.730 123.555 ;
        RECT 66.910 122.660 67.240 123.290 ;
        RECT 67.420 122.830 67.670 123.555 ;
        RECT 67.940 122.835 68.270 123.555 ;
        RECT 65.345 122.230 65.745 122.560 ;
        RECT 66.050 122.490 67.265 122.660 ;
        RECT 65.915 122.060 66.925 122.290 ;
        RECT 65.005 121.890 66.925 122.060 ;
        RECT 65.005 120.660 65.385 121.890 ;
        RECT 67.095 121.720 67.265 122.490 ;
        RECT 65.555 120.395 65.805 121.720 ;
        RECT 66.005 121.550 67.265 121.720 ;
        RECT 66.005 120.660 66.335 121.550 ;
        RECT 66.535 120.395 66.785 121.380 ;
        RECT 66.985 120.660 67.265 121.550 ;
        RECT 67.435 120.395 67.685 121.820 ;
        RECT 68.005 120.395 68.575 122.390 ;
        RECT 68.980 122.055 69.550 123.555 ;
        RECT 69.295 120.395 69.625 121.710 ;
        RECT 10.200 120.225 69.720 120.395 ;
        RECT 10.295 118.910 10.625 120.225 ;
        RECT 10.370 117.065 10.940 118.565 ;
        RECT 11.345 118.230 11.915 120.225 ;
        RECT 12.240 119.010 12.570 120.225 ;
        RECT 12.750 118.840 12.970 119.960 ;
        RECT 13.160 119.010 13.490 120.225 ;
        RECT 13.670 118.840 13.880 119.960 ;
        RECT 14.060 119.010 14.390 120.225 ;
        RECT 14.570 118.840 14.775 119.960 ;
        RECT 14.960 119.010 15.290 120.225 ;
        RECT 15.475 118.840 15.680 119.960 ;
        RECT 15.860 119.010 16.190 120.225 ;
        RECT 16.370 118.840 16.580 119.960 ;
        RECT 16.760 119.010 17.090 120.225 ;
        RECT 17.290 118.840 17.490 119.960 ;
        RECT 17.660 119.010 17.990 120.225 ;
        RECT 18.175 118.840 18.380 119.960 ;
        RECT 18.560 119.010 18.890 120.225 ;
        RECT 19.060 119.100 19.290 119.960 ;
        RECT 19.470 119.270 19.720 120.225 ;
        RECT 19.920 119.100 20.250 119.960 ;
        RECT 20.450 119.270 20.620 120.225 ;
        RECT 20.820 119.100 21.150 119.960 ;
        RECT 12.750 118.810 12.995 118.840 ;
        RECT 11.650 117.065 11.980 117.785 ;
        RECT 12.235 117.065 12.565 117.725 ;
        RECT 12.745 117.330 12.995 118.810 ;
        RECT 13.670 118.670 13.925 118.840 ;
        RECT 14.570 118.670 14.855 118.840 ;
        RECT 15.475 118.670 15.785 118.840 ;
        RECT 16.370 118.670 16.695 118.840 ;
        RECT 17.290 118.670 17.550 118.840 ;
        RECT 18.175 118.670 18.445 118.840 ;
        RECT 13.165 118.170 13.495 118.500 ;
        RECT 13.165 117.065 13.495 117.660 ;
        RECT 13.675 117.330 13.925 118.670 ;
        RECT 14.095 118.170 14.425 118.500 ;
        RECT 14.095 117.065 14.425 117.660 ;
        RECT 14.605 117.330 14.855 118.670 ;
        RECT 15.025 118.170 15.355 118.500 ;
        RECT 15.025 117.065 15.355 117.660 ;
        RECT 15.535 117.330 15.785 118.670 ;
        RECT 15.965 118.170 16.295 118.500 ;
        RECT 15.955 117.065 16.285 117.660 ;
        RECT 16.465 117.330 16.695 118.670 ;
        RECT 16.880 118.170 17.210 118.500 ;
        RECT 17.380 117.725 17.550 118.670 ;
        RECT 17.720 118.170 18.050 118.500 ;
        RECT 16.885 117.065 17.210 117.720 ;
        RECT 17.380 117.330 17.645 117.725 ;
        RECT 17.825 117.065 18.050 117.705 ;
        RECT 18.220 117.330 18.445 118.670 ;
        RECT 18.615 118.170 18.885 118.500 ;
        RECT 18.685 117.065 18.855 117.660 ;
        RECT 19.060 117.330 19.330 119.100 ;
        RECT 19.585 118.930 21.150 119.100 ;
        RECT 21.350 118.930 21.600 120.225 ;
        RECT 23.250 119.185 23.550 120.225 ;
        RECT 19.585 118.390 19.755 118.930 ;
        RECT 23.730 118.800 24.085 119.960 ;
        RECT 24.255 119.270 24.875 120.225 ;
        RECT 25.415 119.100 25.745 119.680 ;
        RECT 24.255 118.930 25.745 119.100 ;
        RECT 19.510 118.160 19.755 118.390 ;
        RECT 19.925 118.330 21.595 118.760 ;
        RECT 19.585 118.130 19.755 118.160 ;
        RECT 19.585 117.960 21.175 118.130 ;
        RECT 23.730 118.110 23.900 118.800 ;
        RECT 24.255 118.610 24.425 118.930 ;
        RECT 25.415 118.800 25.745 118.930 ;
        RECT 27.115 118.800 27.445 120.225 ;
        RECT 27.615 118.865 28.315 119.960 ;
        RECT 24.070 118.280 24.425 118.610 ;
        RECT 24.665 118.330 24.995 118.760 ;
        RECT 24.255 118.160 24.425 118.280 ;
        RECT 25.265 118.160 25.935 118.530 ;
        RECT 19.535 117.065 19.865 117.790 ;
        RECT 20.045 117.330 20.295 117.960 ;
        RECT 20.495 117.065 20.745 117.790 ;
        RECT 20.925 117.330 21.175 117.960 ;
        RECT 21.355 117.065 21.605 117.790 ;
        RECT 23.250 117.065 23.550 118.085 ;
        RECT 23.730 117.330 24.085 118.110 ;
        RECT 24.255 117.990 25.095 118.160 ;
        RECT 27.615 118.110 27.875 118.865 ;
        RECT 28.485 118.695 28.655 119.885 ;
        RECT 28.855 119.175 29.185 120.225 ;
        RECT 29.355 119.425 29.720 119.885 ;
        RECT 29.905 119.425 30.235 120.225 ;
        RECT 30.405 119.455 31.560 119.785 ;
        RECT 29.355 119.005 29.525 119.425 ;
        RECT 24.255 117.065 24.585 117.820 ;
        RECT 24.800 117.520 25.095 117.990 ;
        RECT 25.390 117.065 25.745 117.975 ;
        RECT 27.115 117.065 27.365 118.110 ;
        RECT 27.545 117.330 27.875 118.110 ;
        RECT 28.105 118.365 28.655 118.695 ;
        RECT 28.850 118.835 29.525 119.005 ;
        RECT 29.695 118.900 30.235 119.235 ;
        RECT 28.105 117.330 28.435 118.365 ;
        RECT 28.850 118.165 29.020 118.835 ;
        RECT 30.405 118.665 30.575 119.455 ;
        RECT 29.190 118.495 30.575 118.665 ;
        RECT 29.190 118.335 29.520 118.495 ;
        RECT 30.745 118.325 31.075 119.285 ;
        RECT 31.390 118.665 31.560 119.455 ;
        RECT 31.730 118.845 32.060 119.735 ;
        RECT 31.390 118.495 31.720 118.665 ;
        RECT 30.120 118.165 30.450 118.325 ;
        RECT 28.850 117.995 30.450 118.165 ;
        RECT 30.620 117.995 31.350 118.325 ;
        RECT 28.615 117.065 28.865 117.825 ;
        RECT 29.095 117.365 29.425 117.995 ;
        RECT 29.965 117.065 30.295 117.825 ;
        RECT 30.620 117.405 30.790 117.995 ;
        RECT 31.550 117.825 31.720 118.495 ;
        RECT 30.960 117.575 31.720 117.825 ;
        RECT 31.890 118.110 32.060 118.845 ;
        RECT 32.230 118.725 32.560 120.225 ;
        RECT 33.325 119.720 33.655 120.225 ;
        RECT 34.250 119.550 34.580 119.705 ;
        RECT 32.790 119.380 34.580 119.550 ;
        RECT 34.780 119.490 35.030 119.705 ;
        RECT 35.725 119.660 36.055 120.225 ;
        RECT 36.705 119.630 36.955 120.225 ;
        RECT 37.155 119.500 37.485 119.960 ;
        RECT 37.685 119.500 37.935 120.225 ;
        RECT 38.145 119.500 38.395 120.225 ;
        RECT 38.595 119.500 38.925 119.960 ;
        RECT 39.125 119.630 39.375 120.225 ;
        RECT 40.025 119.660 40.355 120.225 ;
        RECT 42.425 119.720 42.755 120.225 ;
        RECT 34.780 119.460 36.535 119.490 ;
        RECT 37.155 119.460 37.355 119.500 ;
        RECT 32.790 119.300 33.425 119.380 ;
        RECT 32.755 118.775 33.085 119.130 ;
        RECT 33.255 118.555 33.425 119.300 ;
        RECT 32.390 118.225 33.425 118.555 ;
        RECT 31.890 118.055 32.220 118.110 ;
        RECT 33.595 118.055 33.775 119.105 ;
        RECT 31.890 117.885 33.775 118.055 ;
        RECT 33.945 118.030 34.115 119.380 ;
        RECT 34.780 119.320 37.355 119.460 ;
        RECT 34.780 119.210 35.030 119.320 ;
        RECT 36.365 119.290 37.355 119.320 ;
        RECT 34.285 119.040 35.030 119.210 ;
        RECT 34.285 118.370 34.455 119.040 ;
        RECT 35.275 118.870 35.525 119.150 ;
        RECT 34.625 118.700 35.525 118.870 ;
        RECT 36.175 118.790 36.585 119.120 ;
        RECT 34.625 118.540 35.175 118.700 ;
        RECT 34.285 118.200 34.835 118.370 ;
        RECT 31.890 117.645 32.220 117.885 ;
        RECT 32.390 117.545 33.775 117.715 ;
        RECT 33.945 117.650 34.415 118.030 ;
        RECT 34.585 117.650 34.835 118.200 ;
        RECT 35.005 117.780 35.175 118.540 ;
        RECT 35.765 118.620 35.995 118.760 ;
        RECT 35.345 118.120 35.595 118.530 ;
        RECT 35.765 118.290 36.245 118.620 ;
        RECT 36.415 118.120 36.585 118.790 ;
        RECT 35.345 117.950 36.585 118.120 ;
        RECT 36.755 118.110 37.015 119.120 ;
        RECT 32.390 117.405 32.560 117.545 ;
        RECT 30.620 117.235 32.560 117.405 ;
        RECT 33.605 117.480 33.775 117.545 ;
        RECT 35.005 117.480 35.530 117.780 ;
        RECT 32.730 117.065 33.125 117.375 ;
        RECT 33.605 117.310 35.530 117.480 ;
        RECT 35.700 117.065 36.030 117.780 ;
        RECT 36.200 117.330 36.585 117.950 ;
        RECT 37.185 117.810 37.355 119.290 ;
        RECT 38.725 119.460 38.925 119.500 ;
        RECT 41.050 119.490 41.300 119.705 ;
        RECT 39.545 119.460 41.300 119.490 ;
        RECT 38.725 119.320 41.300 119.460 ;
        RECT 41.500 119.550 41.830 119.705 ;
        RECT 41.500 119.380 43.290 119.550 ;
        RECT 38.725 119.290 39.715 119.320 ;
        RECT 37.525 117.980 37.915 119.150 ;
        RECT 38.165 117.980 38.555 119.150 ;
        RECT 38.725 117.810 38.895 119.290 ;
        RECT 41.050 119.210 41.300 119.320 ;
        RECT 39.065 118.110 39.325 119.120 ;
        RECT 39.495 118.790 39.905 119.120 ;
        RECT 40.555 118.870 40.805 119.150 ;
        RECT 41.050 119.040 41.795 119.210 ;
        RECT 39.495 118.120 39.665 118.790 ;
        RECT 40.085 118.620 40.315 118.760 ;
        RECT 40.555 118.700 41.455 118.870 ;
        RECT 39.835 118.290 40.315 118.620 ;
        RECT 40.905 118.540 41.455 118.700 ;
        RECT 40.485 118.120 40.735 118.530 ;
        RECT 39.495 117.950 40.735 118.120 ;
        RECT 36.760 117.065 37.010 117.810 ;
        RECT 37.185 117.640 37.910 117.810 ;
        RECT 37.580 117.350 37.910 117.640 ;
        RECT 38.170 117.640 38.895 117.810 ;
        RECT 38.170 117.350 38.500 117.640 ;
        RECT 39.070 117.065 39.320 117.810 ;
        RECT 39.495 117.330 39.880 117.950 ;
        RECT 40.905 117.780 41.075 118.540 ;
        RECT 41.625 118.370 41.795 119.040 ;
        RECT 40.050 117.065 40.380 117.780 ;
        RECT 40.550 117.480 41.075 117.780 ;
        RECT 41.245 118.200 41.795 118.370 ;
        RECT 41.245 117.650 41.495 118.200 ;
        RECT 41.965 118.030 42.135 119.380 ;
        RECT 42.655 119.300 43.290 119.380 ;
        RECT 41.665 117.650 42.135 118.030 ;
        RECT 42.305 118.055 42.485 119.105 ;
        RECT 42.655 118.555 42.825 119.300 ;
        RECT 42.995 118.775 43.325 119.130 ;
        RECT 43.520 118.725 43.850 120.225 ;
        RECT 44.020 118.845 44.350 119.735 ;
        RECT 44.520 119.455 45.675 119.785 ;
        RECT 42.655 118.225 43.690 118.555 ;
        RECT 44.020 118.110 44.190 118.845 ;
        RECT 44.520 118.665 44.690 119.455 ;
        RECT 43.860 118.055 44.190 118.110 ;
        RECT 42.305 117.885 44.190 118.055 ;
        RECT 42.305 117.545 43.690 117.715 ;
        RECT 43.860 117.645 44.190 117.885 ;
        RECT 44.360 118.495 44.690 118.665 ;
        RECT 44.360 117.825 44.530 118.495 ;
        RECT 45.005 118.325 45.335 119.285 ;
        RECT 45.505 118.665 45.675 119.455 ;
        RECT 45.845 119.425 46.175 120.225 ;
        RECT 46.360 119.425 46.725 119.885 ;
        RECT 45.845 118.900 46.385 119.235 ;
        RECT 46.555 119.005 46.725 119.425 ;
        RECT 46.895 119.175 47.225 120.225 ;
        RECT 46.555 118.835 47.230 119.005 ;
        RECT 45.505 118.495 46.890 118.665 ;
        RECT 46.560 118.335 46.890 118.495 ;
        RECT 44.730 117.995 45.460 118.325 ;
        RECT 45.630 118.165 45.960 118.325 ;
        RECT 47.060 118.165 47.230 118.835 ;
        RECT 47.425 118.695 47.595 119.885 ;
        RECT 47.765 118.865 48.465 119.960 ;
        RECT 47.425 118.365 47.975 118.695 ;
        RECT 45.630 117.995 47.230 118.165 ;
        RECT 44.360 117.575 45.120 117.825 ;
        RECT 42.305 117.480 42.475 117.545 ;
        RECT 40.550 117.310 42.475 117.480 ;
        RECT 43.520 117.405 43.690 117.545 ;
        RECT 45.290 117.405 45.460 117.995 ;
        RECT 42.955 117.065 43.350 117.375 ;
        RECT 43.520 117.235 45.460 117.405 ;
        RECT 45.785 117.065 46.115 117.825 ;
        RECT 46.655 117.365 46.985 117.995 ;
        RECT 47.215 117.065 47.465 117.825 ;
        RECT 47.645 117.330 47.975 118.365 ;
        RECT 48.205 118.110 48.465 118.865 ;
        RECT 48.635 118.800 48.965 120.225 ;
        RECT 49.170 119.185 49.470 120.225 ;
        RECT 51.115 119.470 51.470 119.860 ;
        RECT 51.675 119.640 52.005 120.225 ;
        RECT 52.575 119.715 53.285 120.225 ;
        RECT 51.115 119.300 52.795 119.470 ;
        RECT 51.115 118.930 51.470 119.300 ;
        RECT 51.125 118.330 51.575 118.760 ;
        RECT 51.745 118.160 51.915 119.300 ;
        RECT 52.085 118.160 52.455 119.130 ;
        RECT 52.625 118.610 52.795 119.300 ;
        RECT 52.980 118.800 53.285 119.715 ;
        RECT 53.745 119.100 54.075 119.960 ;
        RECT 54.245 119.270 54.575 120.225 ;
        RECT 53.745 118.930 54.575 119.100 ;
        RECT 52.625 118.280 53.295 118.610 ;
        RECT 53.525 118.280 54.235 118.760 ;
        RECT 54.405 118.610 54.575 118.930 ;
        RECT 54.745 118.800 55.205 119.960 ;
        RECT 56.865 119.500 57.115 120.225 ;
        RECT 57.315 119.500 57.645 119.960 ;
        RECT 57.845 119.630 58.095 120.225 ;
        RECT 58.745 119.660 59.075 120.225 ;
        RECT 61.145 119.720 61.475 120.225 ;
        RECT 57.445 119.460 57.645 119.500 ;
        RECT 59.770 119.490 60.020 119.705 ;
        RECT 58.265 119.460 60.020 119.490 ;
        RECT 57.445 119.320 60.020 119.460 ;
        RECT 60.220 119.550 60.550 119.705 ;
        RECT 60.220 119.380 62.010 119.550 ;
        RECT 57.445 119.290 58.435 119.320 ;
        RECT 48.205 117.330 48.535 118.110 ;
        RECT 48.715 117.065 48.965 118.110 ;
        RECT 49.170 117.065 49.470 118.085 ;
        RECT 51.115 117.990 51.915 118.160 ;
        RECT 51.115 117.430 51.445 117.990 ;
        RECT 51.625 117.065 51.955 117.820 ;
        RECT 52.125 117.330 52.455 118.160 ;
        RECT 54.405 118.110 54.795 118.610 ;
        RECT 52.635 117.065 52.885 118.110 ;
        RECT 53.515 117.940 54.795 118.110 ;
        RECT 53.515 117.330 53.845 117.940 ;
        RECT 54.965 117.770 55.205 118.800 ;
        RECT 56.885 117.980 57.275 119.150 ;
        RECT 57.445 117.810 57.615 119.290 ;
        RECT 59.770 119.210 60.020 119.320 ;
        RECT 57.785 118.110 58.045 119.120 ;
        RECT 58.215 118.790 58.625 119.120 ;
        RECT 59.275 118.870 59.525 119.150 ;
        RECT 59.770 119.040 60.515 119.210 ;
        RECT 58.215 118.120 58.385 118.790 ;
        RECT 58.805 118.620 59.035 118.760 ;
        RECT 59.275 118.700 60.175 118.870 ;
        RECT 58.555 118.290 59.035 118.620 ;
        RECT 59.625 118.540 60.175 118.700 ;
        RECT 59.205 118.120 59.455 118.530 ;
        RECT 58.215 117.950 59.455 118.120 ;
        RECT 54.015 117.065 54.705 117.660 ;
        RECT 54.875 117.330 55.205 117.770 ;
        RECT 56.890 117.640 57.615 117.810 ;
        RECT 56.890 117.350 57.220 117.640 ;
        RECT 57.790 117.065 58.040 117.810 ;
        RECT 58.215 117.330 58.600 117.950 ;
        RECT 59.625 117.780 59.795 118.540 ;
        RECT 60.345 118.370 60.515 119.040 ;
        RECT 58.770 117.065 59.100 117.780 ;
        RECT 59.270 117.480 59.795 117.780 ;
        RECT 59.965 118.200 60.515 118.370 ;
        RECT 59.965 117.650 60.215 118.200 ;
        RECT 60.685 118.030 60.855 119.380 ;
        RECT 61.375 119.300 62.010 119.380 ;
        RECT 60.385 117.650 60.855 118.030 ;
        RECT 61.025 118.055 61.205 119.105 ;
        RECT 61.375 118.555 61.545 119.300 ;
        RECT 61.715 118.775 62.045 119.130 ;
        RECT 62.240 118.725 62.570 120.225 ;
        RECT 62.740 118.845 63.070 119.735 ;
        RECT 63.240 119.455 64.395 119.785 ;
        RECT 61.375 118.225 62.410 118.555 ;
        RECT 62.740 118.110 62.910 118.845 ;
        RECT 63.240 118.665 63.410 119.455 ;
        RECT 62.580 118.055 62.910 118.110 ;
        RECT 61.025 117.885 62.910 118.055 ;
        RECT 61.025 117.545 62.410 117.715 ;
        RECT 62.580 117.645 62.910 117.885 ;
        RECT 63.080 118.495 63.410 118.665 ;
        RECT 63.080 117.825 63.250 118.495 ;
        RECT 63.725 118.325 64.055 119.285 ;
        RECT 64.225 118.665 64.395 119.455 ;
        RECT 64.565 119.425 64.895 120.225 ;
        RECT 65.080 119.425 65.445 119.885 ;
        RECT 64.565 118.900 65.105 119.235 ;
        RECT 65.275 119.005 65.445 119.425 ;
        RECT 65.615 119.175 65.945 120.225 ;
        RECT 65.275 118.835 65.950 119.005 ;
        RECT 64.225 118.495 65.610 118.665 ;
        RECT 65.280 118.335 65.610 118.495 ;
        RECT 63.450 117.995 64.180 118.325 ;
        RECT 64.350 118.165 64.680 118.325 ;
        RECT 65.780 118.165 65.950 118.835 ;
        RECT 66.145 118.695 66.315 119.885 ;
        RECT 66.485 118.865 67.185 119.960 ;
        RECT 66.145 118.365 66.695 118.695 ;
        RECT 64.350 117.995 65.950 118.165 ;
        RECT 63.080 117.575 63.840 117.825 ;
        RECT 61.025 117.480 61.195 117.545 ;
        RECT 59.270 117.310 61.195 117.480 ;
        RECT 62.240 117.405 62.410 117.545 ;
        RECT 64.010 117.405 64.180 117.995 ;
        RECT 61.675 117.065 62.070 117.375 ;
        RECT 62.240 117.235 64.180 117.405 ;
        RECT 64.505 117.065 64.835 117.825 ;
        RECT 65.375 117.365 65.705 117.995 ;
        RECT 65.935 117.065 66.185 117.825 ;
        RECT 66.365 117.330 66.695 118.365 ;
        RECT 66.925 118.110 67.185 118.865 ;
        RECT 67.355 118.800 67.685 120.225 ;
        RECT 68.005 118.230 68.575 120.225 ;
        RECT 69.295 118.910 69.625 120.225 ;
        RECT 66.925 117.330 67.255 118.110 ;
        RECT 67.435 117.065 67.685 118.110 ;
        RECT 67.940 117.065 68.270 117.785 ;
        RECT 68.980 117.065 69.550 118.565 ;
        RECT 10.200 116.895 69.720 117.065 ;
        RECT 10.370 115.395 10.940 116.895 ;
        RECT 11.650 116.175 11.980 116.895 ;
        RECT 10.295 113.735 10.625 115.050 ;
        RECT 11.345 113.735 11.915 115.730 ;
        RECT 12.290 115.395 12.860 116.895 ;
        RECT 13.570 116.175 13.900 116.895 ;
        RECT 14.155 116.190 14.485 116.630 ;
        RECT 14.655 116.300 15.345 116.895 ;
        RECT 12.215 113.735 12.545 115.050 ;
        RECT 13.265 113.735 13.835 115.730 ;
        RECT 14.155 115.160 14.395 116.190 ;
        RECT 15.515 116.020 15.845 116.630 ;
        RECT 14.565 115.850 15.845 116.020 ;
        RECT 16.075 116.020 16.325 116.630 ;
        RECT 16.505 116.190 16.835 116.895 ;
        RECT 17.040 116.510 17.230 116.630 ;
        RECT 17.040 116.340 17.245 116.510 ;
        RECT 17.040 116.020 17.230 116.340 ;
        RECT 17.780 116.120 18.345 116.630 ;
        RECT 19.680 116.300 20.070 116.895 ;
        RECT 20.315 116.130 20.645 116.540 ;
        RECT 21.355 116.235 21.685 116.895 ;
        RECT 16.075 115.850 16.700 116.020 ;
        RECT 14.565 115.350 14.955 115.850 ;
        RECT 14.155 114.000 14.615 115.160 ;
        RECT 14.785 115.030 14.955 115.350 ;
        RECT 15.125 115.200 15.835 115.680 ;
        RECT 16.065 115.200 16.360 115.680 ;
        RECT 16.530 115.030 16.700 115.850 ;
        RECT 14.785 114.860 15.615 115.030 ;
        RECT 14.785 113.735 15.115 114.690 ;
        RECT 15.285 114.000 15.615 114.860 ;
        RECT 16.075 114.660 16.700 115.030 ;
        RECT 16.870 115.850 17.230 116.020 ;
        RECT 17.400 115.950 18.345 116.120 ;
        RECT 16.870 115.160 17.040 115.850 ;
        RECT 17.400 115.680 17.570 115.950 ;
        RECT 17.210 115.350 17.570 115.680 ;
        RECT 16.870 114.830 17.525 115.160 ;
        RECT 17.740 114.660 18.005 115.690 ;
        RECT 18.175 114.950 18.345 115.950 ;
        RECT 18.515 115.960 20.645 116.130 ;
        RECT 18.515 115.190 18.805 115.960 ;
        RECT 20.020 115.950 20.645 115.960 ;
        RECT 18.975 115.120 19.305 115.790 ;
        RECT 19.475 115.120 19.850 115.790 ;
        RECT 20.020 115.030 20.190 115.950 ;
        RECT 20.360 115.200 20.655 115.680 ;
        RECT 21.865 115.150 22.115 116.630 ;
        RECT 22.285 116.300 22.615 116.895 ;
        RECT 22.285 115.460 22.615 115.790 ;
        RECT 22.795 115.290 23.045 116.630 ;
        RECT 23.215 116.300 23.545 116.895 ;
        RECT 23.215 115.460 23.545 115.790 ;
        RECT 23.725 115.290 23.975 116.630 ;
        RECT 24.145 116.300 24.475 116.895 ;
        RECT 24.145 115.460 24.475 115.790 ;
        RECT 24.655 115.290 24.905 116.630 ;
        RECT 25.075 116.300 25.405 116.895 ;
        RECT 25.085 115.460 25.415 115.790 ;
        RECT 25.585 115.290 25.815 116.630 ;
        RECT 26.005 116.240 26.330 116.895 ;
        RECT 26.500 116.235 26.765 116.630 ;
        RECT 26.945 116.255 27.170 116.895 ;
        RECT 26.000 115.460 26.330 115.790 ;
        RECT 26.500 115.290 26.670 116.235 ;
        RECT 26.840 115.460 27.170 115.790 ;
        RECT 27.340 115.290 27.565 116.630 ;
        RECT 27.805 116.300 27.975 116.895 ;
        RECT 27.735 115.460 28.005 115.790 ;
        RECT 21.870 115.120 22.115 115.150 ;
        RECT 22.790 115.120 23.045 115.290 ;
        RECT 23.690 115.120 23.975 115.290 ;
        RECT 24.595 115.120 24.905 115.290 ;
        RECT 25.490 115.120 25.815 115.290 ;
        RECT 26.410 115.120 26.670 115.290 ;
        RECT 27.295 115.120 27.565 115.290 ;
        RECT 18.175 114.780 19.585 114.950 ;
        RECT 20.020 114.860 20.605 115.030 ;
        RECT 16.075 114.490 18.005 114.660 ;
        RECT 16.075 114.280 16.405 114.490 ;
        RECT 16.610 113.735 16.940 114.320 ;
        RECT 17.755 113.735 18.085 114.320 ;
        RECT 18.255 114.000 18.585 114.780 ;
        RECT 18.755 113.735 19.085 114.610 ;
        RECT 19.255 114.000 19.585 114.780 ;
        RECT 19.775 113.735 20.105 114.690 ;
        RECT 20.275 114.000 20.605 114.860 ;
        RECT 21.360 113.735 21.690 114.950 ;
        RECT 21.870 114.000 22.090 115.120 ;
        RECT 22.280 113.735 22.610 114.950 ;
        RECT 22.790 114.000 23.000 115.120 ;
        RECT 23.180 113.735 23.510 114.950 ;
        RECT 23.690 114.000 23.895 115.120 ;
        RECT 24.080 113.735 24.410 114.950 ;
        RECT 24.595 114.000 24.800 115.120 ;
        RECT 24.980 113.735 25.310 114.950 ;
        RECT 25.490 114.000 25.700 115.120 ;
        RECT 25.880 113.735 26.210 114.950 ;
        RECT 26.410 114.000 26.610 115.120 ;
        RECT 26.780 113.735 27.110 114.950 ;
        RECT 27.295 114.000 27.500 115.120 ;
        RECT 27.680 113.735 28.010 114.950 ;
        RECT 28.180 114.860 28.450 116.630 ;
        RECT 28.655 116.170 28.985 116.895 ;
        RECT 29.165 116.000 29.415 116.630 ;
        RECT 29.615 116.170 29.865 116.895 ;
        RECT 30.045 116.000 30.295 116.630 ;
        RECT 30.475 116.170 30.725 116.895 ;
        RECT 28.705 115.830 30.295 116.000 ;
        RECT 30.955 115.850 31.285 116.895 ;
        RECT 31.465 115.850 31.715 116.630 ;
        RECT 31.895 115.850 32.145 116.895 ;
        RECT 32.375 116.160 32.690 116.675 ;
        RECT 32.865 116.330 33.195 116.895 ;
        RECT 33.695 116.345 34.000 116.675 ;
        RECT 32.375 115.960 33.585 116.160 ;
        RECT 28.705 115.800 28.875 115.830 ;
        RECT 28.630 115.570 28.875 115.800 ;
        RECT 28.705 115.030 28.875 115.570 ;
        RECT 29.045 115.200 30.715 115.630 ;
        RECT 30.965 115.200 31.295 115.680 ;
        RECT 31.465 115.030 31.635 115.850 ;
        RECT 31.825 115.200 32.155 115.680 ;
        RECT 32.380 115.120 33.010 115.790 ;
        RECT 28.705 114.860 30.270 115.030 ;
        RECT 28.180 114.000 28.410 114.860 ;
        RECT 28.590 113.735 28.840 114.690 ;
        RECT 29.040 114.000 29.370 114.860 ;
        RECT 29.570 113.735 29.740 114.690 ;
        RECT 29.940 114.000 30.270 114.860 ;
        RECT 30.470 113.735 30.720 115.030 ;
        RECT 30.965 114.290 31.635 115.030 ;
        RECT 30.965 114.120 31.645 114.290 ;
        RECT 30.965 114.090 31.635 114.120 ;
        RECT 30.965 114.000 31.295 114.090 ;
        RECT 31.835 113.735 32.165 115.030 ;
        RECT 33.255 114.950 33.585 115.960 ;
        RECT 32.375 114.775 33.585 114.950 ;
        RECT 33.755 115.600 34.000 116.345 ;
        RECT 34.265 115.940 34.625 116.270 ;
        RECT 35.105 116.110 35.435 116.895 ;
        RECT 34.265 115.770 35.435 115.940 ;
        RECT 35.605 115.860 36.020 116.625 ;
        RECT 36.210 115.875 36.510 116.895 ;
        RECT 36.960 116.140 37.290 116.630 ;
        RECT 36.745 115.970 37.290 116.140 ;
        RECT 35.190 115.685 35.435 115.770 ;
        RECT 33.755 115.370 35.020 115.600 ;
        RECT 32.375 114.255 32.680 114.775 ;
        RECT 32.855 113.735 33.185 114.600 ;
        RECT 33.755 114.585 34.000 115.370 ;
        RECT 35.190 115.355 35.560 115.685 ;
        RECT 35.190 115.155 35.435 115.355 ;
        RECT 35.730 115.165 36.020 115.860 ;
        RECT 34.265 114.985 35.435 115.155 ;
        RECT 34.265 114.790 34.625 114.985 ;
        RECT 33.695 114.255 34.000 114.585 ;
        RECT 35.105 113.735 35.435 114.815 ;
        RECT 35.605 113.920 36.020 115.165 ;
        RECT 36.745 115.260 36.915 115.970 ;
        RECT 37.085 115.430 37.435 115.800 ;
        RECT 37.655 115.430 37.985 116.540 ;
        RECT 38.350 115.970 38.680 116.895 ;
        RECT 39.610 116.320 39.940 116.610 ;
        RECT 39.610 116.150 40.335 116.320 ;
        RECT 40.510 116.150 40.760 116.895 ;
        RECT 38.165 115.430 38.895 115.800 ;
        RECT 36.745 115.090 38.395 115.260 ;
        RECT 36.210 113.735 36.510 114.775 ;
        RECT 36.745 114.000 37.265 115.090 ;
        RECT 37.455 113.735 37.785 114.920 ;
        RECT 37.955 114.000 38.395 115.090 ;
        RECT 38.565 113.735 38.815 115.160 ;
        RECT 39.605 114.810 39.995 115.980 ;
        RECT 40.165 114.670 40.335 116.150 ;
        RECT 40.935 116.010 41.320 116.630 ;
        RECT 41.490 116.180 41.820 116.895 ;
        RECT 41.990 116.480 43.915 116.650 ;
        RECT 44.395 116.585 44.790 116.895 ;
        RECT 41.990 116.180 42.515 116.480 ;
        RECT 43.745 116.415 43.915 116.480 ;
        RECT 44.960 116.555 46.900 116.725 ;
        RECT 44.960 116.415 45.130 116.555 ;
        RECT 40.505 114.840 40.765 115.850 ;
        RECT 40.935 115.840 42.175 116.010 ;
        RECT 40.935 115.170 41.105 115.840 ;
        RECT 41.275 115.340 41.755 115.670 ;
        RECT 41.925 115.430 42.175 115.840 ;
        RECT 41.525 115.200 41.755 115.340 ;
        RECT 42.345 115.420 42.515 116.180 ;
        RECT 42.685 115.760 42.935 116.310 ;
        RECT 43.105 115.930 43.575 116.310 ;
        RECT 43.745 116.245 45.130 116.415 ;
        RECT 45.300 116.075 45.630 116.315 ;
        RECT 42.685 115.590 43.235 115.760 ;
        RECT 42.345 115.260 42.895 115.420 ;
        RECT 40.935 114.840 41.345 115.170 ;
        RECT 41.995 115.090 42.895 115.260 ;
        RECT 41.995 114.810 42.245 115.090 ;
        RECT 43.065 114.920 43.235 115.590 ;
        RECT 42.490 114.750 43.235 114.920 ;
        RECT 40.165 114.640 41.155 114.670 ;
        RECT 42.490 114.640 42.740 114.750 ;
        RECT 40.165 114.500 42.740 114.640 ;
        RECT 43.405 114.580 43.575 115.930 ;
        RECT 43.745 115.905 45.630 116.075 ;
        RECT 43.745 114.855 43.925 115.905 ;
        RECT 45.300 115.850 45.630 115.905 ;
        RECT 44.095 115.405 45.130 115.735 ;
        RECT 44.095 114.660 44.265 115.405 ;
        RECT 44.435 114.830 44.765 115.185 ;
        RECT 44.095 114.580 44.730 114.660 ;
        RECT 40.165 114.460 40.365 114.500 ;
        RECT 40.985 114.470 42.740 114.500 ;
        RECT 39.585 113.735 39.835 114.460 ;
        RECT 40.035 114.000 40.365 114.460 ;
        RECT 40.565 113.735 40.815 114.330 ;
        RECT 41.465 113.735 41.795 114.300 ;
        RECT 42.490 114.255 42.740 114.470 ;
        RECT 42.940 114.410 44.730 114.580 ;
        RECT 42.940 114.255 43.270 114.410 ;
        RECT 43.865 113.735 44.195 114.240 ;
        RECT 44.960 113.735 45.290 115.235 ;
        RECT 45.460 115.115 45.630 115.850 ;
        RECT 45.800 116.135 46.560 116.385 ;
        RECT 45.800 115.465 45.970 116.135 ;
        RECT 46.730 115.965 46.900 116.555 ;
        RECT 47.225 116.135 47.555 116.895 ;
        RECT 48.095 115.965 48.425 116.595 ;
        RECT 48.655 116.135 48.905 116.895 ;
        RECT 46.170 115.635 46.900 115.965 ;
        RECT 47.070 115.795 48.670 115.965 ;
        RECT 47.070 115.635 47.400 115.795 ;
        RECT 45.800 115.295 46.130 115.465 ;
        RECT 45.460 114.225 45.790 115.115 ;
        RECT 45.960 114.505 46.130 115.295 ;
        RECT 46.445 114.675 46.775 115.635 ;
        RECT 48.000 115.465 48.330 115.625 ;
        RECT 46.945 115.295 48.330 115.465 ;
        RECT 46.945 114.505 47.115 115.295 ;
        RECT 48.500 115.125 48.670 115.795 ;
        RECT 49.085 115.595 49.415 116.630 ;
        RECT 47.285 114.725 47.825 115.060 ;
        RECT 47.995 114.955 48.670 115.125 ;
        RECT 48.865 115.265 49.415 115.595 ;
        RECT 49.645 115.850 49.975 116.630 ;
        RECT 50.155 115.850 50.405 116.895 ;
        RECT 51.130 116.320 51.460 116.610 ;
        RECT 51.130 116.150 51.855 116.320 ;
        RECT 52.030 116.150 52.280 116.895 ;
        RECT 47.995 114.535 48.165 114.955 ;
        RECT 45.960 114.175 47.115 114.505 ;
        RECT 47.285 113.735 47.615 114.535 ;
        RECT 47.800 114.075 48.165 114.535 ;
        RECT 48.335 113.735 48.665 114.785 ;
        RECT 48.865 114.075 49.035 115.265 ;
        RECT 49.645 115.095 49.905 115.850 ;
        RECT 49.205 114.000 49.905 115.095 ;
        RECT 50.075 113.735 50.405 115.160 ;
        RECT 51.125 114.810 51.515 115.980 ;
        RECT 51.685 114.670 51.855 116.150 ;
        RECT 52.455 116.010 52.840 116.630 ;
        RECT 53.010 116.180 53.340 116.895 ;
        RECT 53.510 116.480 55.435 116.650 ;
        RECT 55.915 116.585 56.310 116.895 ;
        RECT 53.510 116.180 54.035 116.480 ;
        RECT 55.265 116.415 55.435 116.480 ;
        RECT 56.480 116.555 58.420 116.725 ;
        RECT 56.480 116.415 56.650 116.555 ;
        RECT 52.025 114.840 52.285 115.850 ;
        RECT 52.455 115.840 53.695 116.010 ;
        RECT 52.455 115.170 52.625 115.840 ;
        RECT 52.795 115.340 53.275 115.670 ;
        RECT 53.445 115.430 53.695 115.840 ;
        RECT 53.045 115.200 53.275 115.340 ;
        RECT 53.865 115.420 54.035 116.180 ;
        RECT 54.205 115.760 54.455 116.310 ;
        RECT 54.625 115.930 55.095 116.310 ;
        RECT 55.265 116.245 56.650 116.415 ;
        RECT 56.820 116.075 57.150 116.315 ;
        RECT 54.205 115.590 54.755 115.760 ;
        RECT 53.865 115.260 54.415 115.420 ;
        RECT 52.455 114.840 52.865 115.170 ;
        RECT 53.515 115.090 54.415 115.260 ;
        RECT 53.515 114.810 53.765 115.090 ;
        RECT 54.585 114.920 54.755 115.590 ;
        RECT 54.010 114.750 54.755 114.920 ;
        RECT 51.685 114.640 52.675 114.670 ;
        RECT 54.010 114.640 54.260 114.750 ;
        RECT 51.685 114.500 54.260 114.640 ;
        RECT 54.925 114.580 55.095 115.930 ;
        RECT 55.265 115.905 57.150 116.075 ;
        RECT 55.265 114.855 55.445 115.905 ;
        RECT 56.820 115.850 57.150 115.905 ;
        RECT 55.615 115.405 56.650 115.735 ;
        RECT 55.615 114.660 55.785 115.405 ;
        RECT 55.955 114.830 56.285 115.185 ;
        RECT 55.615 114.580 56.250 114.660 ;
        RECT 51.685 114.460 51.885 114.500 ;
        RECT 52.505 114.470 54.260 114.500 ;
        RECT 51.105 113.735 51.355 114.460 ;
        RECT 51.555 114.000 51.885 114.460 ;
        RECT 52.085 113.735 52.335 114.330 ;
        RECT 52.985 113.735 53.315 114.300 ;
        RECT 54.010 114.255 54.260 114.470 ;
        RECT 54.460 114.410 56.250 114.580 ;
        RECT 54.460 114.255 54.790 114.410 ;
        RECT 55.385 113.735 55.715 114.240 ;
        RECT 56.480 113.735 56.810 115.235 ;
        RECT 56.980 115.115 57.150 115.850 ;
        RECT 57.320 116.135 58.080 116.385 ;
        RECT 57.320 115.465 57.490 116.135 ;
        RECT 58.250 115.965 58.420 116.555 ;
        RECT 58.745 116.135 59.075 116.895 ;
        RECT 59.615 115.965 59.945 116.595 ;
        RECT 60.175 116.135 60.425 116.895 ;
        RECT 57.690 115.635 58.420 115.965 ;
        RECT 58.590 115.795 60.190 115.965 ;
        RECT 58.590 115.635 58.920 115.795 ;
        RECT 57.320 115.295 57.650 115.465 ;
        RECT 56.980 114.225 57.310 115.115 ;
        RECT 57.480 114.505 57.650 115.295 ;
        RECT 57.965 114.675 58.295 115.635 ;
        RECT 59.520 115.465 59.850 115.625 ;
        RECT 58.465 115.295 59.850 115.465 ;
        RECT 58.465 114.505 58.635 115.295 ;
        RECT 60.020 115.125 60.190 115.795 ;
        RECT 60.605 115.595 60.935 116.630 ;
        RECT 58.805 114.725 59.345 115.060 ;
        RECT 59.515 114.955 60.190 115.125 ;
        RECT 60.385 115.265 60.935 115.595 ;
        RECT 61.165 115.850 61.495 116.630 ;
        RECT 61.675 115.850 61.925 116.895 ;
        RECT 62.130 115.875 62.430 116.895 ;
        RECT 59.515 114.535 59.685 114.955 ;
        RECT 57.480 114.175 58.635 114.505 ;
        RECT 58.805 113.735 59.135 114.535 ;
        RECT 59.320 114.075 59.685 114.535 ;
        RECT 59.855 113.735 60.185 114.785 ;
        RECT 60.385 114.075 60.555 115.265 ;
        RECT 61.165 115.095 61.425 115.850 ;
        RECT 62.690 115.395 63.260 116.895 ;
        RECT 63.970 116.175 64.300 116.895 ;
        RECT 65.005 116.170 65.380 116.500 ;
        RECT 65.550 116.170 65.880 116.895 ;
        RECT 60.725 114.000 61.425 115.095 ;
        RECT 61.595 113.735 61.925 115.160 ;
        RECT 62.130 113.735 62.430 114.775 ;
        RECT 62.615 113.735 62.945 115.050 ;
        RECT 63.665 113.735 64.235 115.730 ;
        RECT 65.005 115.400 65.175 116.170 ;
        RECT 66.050 116.000 66.380 116.630 ;
        RECT 66.560 116.170 66.730 116.895 ;
        RECT 66.910 116.000 67.240 116.630 ;
        RECT 67.420 116.170 67.670 116.895 ;
        RECT 67.940 116.175 68.270 116.895 ;
        RECT 65.345 115.570 65.745 115.900 ;
        RECT 66.050 115.830 67.265 116.000 ;
        RECT 65.915 115.400 66.925 115.630 ;
        RECT 65.005 115.230 66.925 115.400 ;
        RECT 65.005 114.000 65.385 115.230 ;
        RECT 67.095 115.060 67.265 115.830 ;
        RECT 65.555 113.735 65.805 115.060 ;
        RECT 66.005 114.890 67.265 115.060 ;
        RECT 66.005 114.000 66.335 114.890 ;
        RECT 66.535 113.735 66.785 114.720 ;
        RECT 66.985 114.000 67.265 114.890 ;
        RECT 67.435 113.735 67.685 115.160 ;
        RECT 68.005 113.735 68.575 115.730 ;
        RECT 68.980 115.395 69.550 116.895 ;
        RECT 69.295 113.735 69.625 115.050 ;
        RECT 10.200 113.565 69.720 113.735 ;
        RECT 10.295 112.250 10.625 113.565 ;
        RECT 10.370 110.405 10.940 111.905 ;
        RECT 11.345 111.570 11.915 113.565 ;
        RECT 12.235 112.270 12.565 113.565 ;
        RECT 13.105 113.210 13.435 113.300 ;
        RECT 12.765 112.270 13.435 113.210 ;
        RECT 13.675 112.270 14.005 113.565 ;
        RECT 14.545 113.210 14.875 113.300 ;
        RECT 14.205 112.270 14.875 113.210 ;
        RECT 15.115 112.440 15.445 113.300 ;
        RECT 15.645 112.610 15.815 113.565 ;
        RECT 16.015 113.115 16.345 113.300 ;
        RECT 16.575 113.285 16.910 113.565 ;
        RECT 18.800 113.285 19.130 113.565 ;
        RECT 17.080 113.115 18.460 113.285 ;
        RECT 19.780 113.225 20.840 113.395 ;
        RECT 19.780 113.115 19.950 113.225 ;
        RECT 16.015 112.945 17.250 113.115 ;
        RECT 18.290 112.945 19.950 113.115 ;
        RECT 15.115 112.270 15.845 112.440 ;
        RECT 12.245 111.620 12.575 112.100 ;
        RECT 12.765 111.450 12.935 112.270 ;
        RECT 13.105 111.620 13.435 112.100 ;
        RECT 13.685 111.620 14.015 112.100 ;
        RECT 14.205 111.450 14.375 112.270 ;
        RECT 14.545 111.620 14.875 112.100 ;
        RECT 15.125 111.620 15.505 112.100 ;
        RECT 15.675 111.870 15.845 112.270 ;
        RECT 16.015 112.140 16.475 112.945 ;
        RECT 16.870 112.345 17.250 112.675 ;
        RECT 16.305 112.000 16.475 112.140 ;
        RECT 15.675 111.450 16.135 111.870 ;
        RECT 11.650 110.405 11.980 111.125 ;
        RECT 12.255 110.405 12.505 111.450 ;
        RECT 12.685 110.670 12.935 111.450 ;
        RECT 13.115 110.405 13.445 111.450 ;
        RECT 13.695 110.405 13.945 111.450 ;
        RECT 14.125 110.670 14.375 111.450 ;
        RECT 14.555 110.405 14.885 111.450 ;
        RECT 15.115 111.280 16.135 111.450 ;
        RECT 15.115 110.670 15.365 111.280 ;
        RECT 15.545 110.405 15.795 111.110 ;
        RECT 15.965 110.745 16.135 111.280 ;
        RECT 16.305 111.670 16.760 112.000 ;
        RECT 16.305 110.915 16.475 111.670 ;
        RECT 16.970 111.445 17.250 112.345 ;
        RECT 17.420 111.560 17.590 112.945 ;
        RECT 17.760 112.775 18.120 112.945 ;
        RECT 17.760 112.605 19.140 112.775 ;
        RECT 17.760 111.900 17.930 112.605 ;
        RECT 18.100 112.070 18.760 112.400 ;
        RECT 17.760 111.730 18.420 111.900 ;
        RECT 17.420 111.390 17.975 111.560 ;
        RECT 16.645 111.050 17.655 111.220 ;
        RECT 16.645 110.745 16.815 111.050 ;
        RECT 15.965 110.575 16.815 110.745 ;
        RECT 16.985 110.405 17.315 110.880 ;
        RECT 17.485 110.765 17.655 111.050 ;
        RECT 18.155 110.935 18.420 111.730 ;
        RECT 18.590 111.180 18.760 112.070 ;
        RECT 18.970 112.275 19.140 112.605 ;
        RECT 19.335 112.445 19.610 112.775 ;
        RECT 18.970 111.945 19.270 112.275 ;
        RECT 18.930 111.520 19.260 111.735 ;
        RECT 19.440 111.520 19.610 112.445 ;
        RECT 19.780 111.860 19.950 112.945 ;
        RECT 20.120 112.200 20.290 113.055 ;
        RECT 20.510 112.370 20.840 113.225 ;
        RECT 21.200 112.840 21.530 113.565 ;
        RECT 20.120 112.030 20.820 112.200 ;
        RECT 19.780 111.690 20.480 111.860 ;
        RECT 18.930 111.350 20.000 111.520 ;
        RECT 20.170 111.470 20.480 111.690 ;
        RECT 20.650 111.720 20.820 112.030 ;
        RECT 21.050 112.180 21.380 112.560 ;
        RECT 21.760 112.180 22.010 113.020 ;
        RECT 22.210 112.350 22.540 113.565 ;
        RECT 22.715 112.350 23.075 113.300 ;
        RECT 23.250 112.525 23.550 113.565 ;
        RECT 21.050 112.010 22.735 112.180 ;
        RECT 21.050 111.890 21.380 112.010 ;
        RECT 21.875 111.720 22.205 111.840 ;
        RECT 20.650 111.550 22.205 111.720 ;
        RECT 18.590 111.010 19.660 111.180 ;
        RECT 18.590 110.765 18.760 111.010 ;
        RECT 17.485 110.595 18.760 110.765 ;
        RECT 19.070 110.405 19.320 110.840 ;
        RECT 19.490 110.745 19.660 111.010 ;
        RECT 19.830 110.915 20.000 111.350 ;
        RECT 20.650 111.300 20.820 111.550 ;
        RECT 21.875 111.510 22.205 111.550 ;
        RECT 22.375 111.670 22.735 112.010 ;
        RECT 20.220 111.050 20.820 111.300 ;
        RECT 20.565 110.745 20.895 110.830 ;
        RECT 19.490 110.575 20.895 110.745 ;
        RECT 21.230 110.405 21.560 111.380 ;
        RECT 22.375 111.340 22.545 111.670 ;
        RECT 22.905 111.450 23.075 112.350 ;
        RECT 23.755 112.440 24.085 113.300 ;
        RECT 24.285 112.610 24.455 113.565 ;
        RECT 24.655 113.115 24.985 113.300 ;
        RECT 25.215 113.285 25.550 113.565 ;
        RECT 27.440 113.285 27.770 113.565 ;
        RECT 25.720 113.115 27.100 113.285 ;
        RECT 28.420 113.225 29.480 113.395 ;
        RECT 28.420 113.115 28.590 113.225 ;
        RECT 24.655 112.945 25.890 113.115 ;
        RECT 26.930 112.945 28.590 113.115 ;
        RECT 23.755 112.270 24.485 112.440 ;
        RECT 23.765 111.620 24.145 112.100 ;
        RECT 24.315 111.870 24.485 112.270 ;
        RECT 24.655 112.140 25.115 112.945 ;
        RECT 25.510 112.345 25.890 112.675 ;
        RECT 24.945 112.000 25.115 112.140 ;
        RECT 24.315 111.450 24.775 111.870 ;
        RECT 21.790 111.170 22.545 111.340 ;
        RECT 21.790 110.670 22.040 111.170 ;
        RECT 22.220 110.405 22.535 111.000 ;
        RECT 22.715 110.670 23.075 111.450 ;
        RECT 23.250 110.405 23.550 111.425 ;
        RECT 23.755 111.280 24.775 111.450 ;
        RECT 23.755 110.670 24.005 111.280 ;
        RECT 24.185 110.405 24.435 111.110 ;
        RECT 24.605 110.745 24.775 111.280 ;
        RECT 24.945 111.670 25.400 112.000 ;
        RECT 24.945 110.915 25.115 111.670 ;
        RECT 25.610 111.445 25.890 112.345 ;
        RECT 26.060 111.560 26.230 112.945 ;
        RECT 26.400 112.775 26.760 112.945 ;
        RECT 26.400 112.605 27.780 112.775 ;
        RECT 26.400 111.900 26.570 112.605 ;
        RECT 26.740 112.070 27.400 112.400 ;
        RECT 26.400 111.730 27.060 111.900 ;
        RECT 26.060 111.390 26.615 111.560 ;
        RECT 25.285 111.050 26.295 111.220 ;
        RECT 25.285 110.745 25.455 111.050 ;
        RECT 24.605 110.575 25.455 110.745 ;
        RECT 25.625 110.405 25.955 110.880 ;
        RECT 26.125 110.765 26.295 111.050 ;
        RECT 26.795 110.935 27.060 111.730 ;
        RECT 27.230 111.180 27.400 112.070 ;
        RECT 27.610 112.275 27.780 112.605 ;
        RECT 27.975 112.445 28.250 112.775 ;
        RECT 27.610 111.945 27.910 112.275 ;
        RECT 27.570 111.520 27.900 111.735 ;
        RECT 28.080 111.520 28.250 112.445 ;
        RECT 28.420 111.860 28.590 112.945 ;
        RECT 28.760 112.200 28.930 113.055 ;
        RECT 29.150 112.370 29.480 113.225 ;
        RECT 29.840 112.840 30.170 113.565 ;
        RECT 28.760 112.030 29.460 112.200 ;
        RECT 28.420 111.690 29.120 111.860 ;
        RECT 27.570 111.350 28.640 111.520 ;
        RECT 28.810 111.470 29.120 111.690 ;
        RECT 29.290 111.720 29.460 112.030 ;
        RECT 29.690 112.180 30.020 112.560 ;
        RECT 30.400 112.180 30.650 113.020 ;
        RECT 30.850 112.350 31.180 113.565 ;
        RECT 31.355 112.350 31.715 113.300 ;
        RECT 29.690 112.010 31.375 112.180 ;
        RECT 29.690 111.890 30.020 112.010 ;
        RECT 30.515 111.720 30.845 111.840 ;
        RECT 29.290 111.550 30.845 111.720 ;
        RECT 27.230 111.010 28.300 111.180 ;
        RECT 27.230 110.765 27.400 111.010 ;
        RECT 26.125 110.595 27.400 110.765 ;
        RECT 27.710 110.405 27.960 110.840 ;
        RECT 28.130 110.745 28.300 111.010 ;
        RECT 28.470 110.915 28.640 111.350 ;
        RECT 29.290 111.300 29.460 111.550 ;
        RECT 30.515 111.510 30.845 111.550 ;
        RECT 31.015 111.670 31.375 112.010 ;
        RECT 28.860 111.050 29.460 111.300 ;
        RECT 29.205 110.745 29.535 110.830 ;
        RECT 28.130 110.575 29.535 110.745 ;
        RECT 29.870 110.405 30.200 111.380 ;
        RECT 31.015 111.340 31.185 111.670 ;
        RECT 31.545 111.450 31.715 112.350 ;
        RECT 32.395 112.140 32.725 113.565 ;
        RECT 32.895 112.205 33.595 113.300 ;
        RECT 32.895 111.450 33.155 112.205 ;
        RECT 33.765 112.035 33.935 113.225 ;
        RECT 34.135 112.515 34.465 113.565 ;
        RECT 34.635 112.765 35.000 113.225 ;
        RECT 35.185 112.765 35.515 113.565 ;
        RECT 35.685 112.795 36.840 113.125 ;
        RECT 34.635 112.345 34.805 112.765 ;
        RECT 30.430 111.170 31.185 111.340 ;
        RECT 30.430 110.670 30.680 111.170 ;
        RECT 30.860 110.405 31.175 111.000 ;
        RECT 31.355 110.670 31.715 111.450 ;
        RECT 32.395 110.405 32.645 111.450 ;
        RECT 32.825 110.670 33.155 111.450 ;
        RECT 33.385 111.705 33.935 112.035 ;
        RECT 34.130 112.175 34.805 112.345 ;
        RECT 34.975 112.240 35.515 112.575 ;
        RECT 33.385 110.670 33.715 111.705 ;
        RECT 34.130 111.505 34.300 112.175 ;
        RECT 35.685 112.005 35.855 112.795 ;
        RECT 34.470 111.835 35.855 112.005 ;
        RECT 34.470 111.675 34.800 111.835 ;
        RECT 36.025 111.665 36.355 112.625 ;
        RECT 36.670 112.005 36.840 112.795 ;
        RECT 37.010 112.185 37.340 113.075 ;
        RECT 36.670 111.835 37.000 112.005 ;
        RECT 35.400 111.505 35.730 111.665 ;
        RECT 34.130 111.335 35.730 111.505 ;
        RECT 35.900 111.335 36.630 111.665 ;
        RECT 33.895 110.405 34.145 111.165 ;
        RECT 34.375 110.705 34.705 111.335 ;
        RECT 35.245 110.405 35.575 111.165 ;
        RECT 35.900 110.745 36.070 111.335 ;
        RECT 36.830 111.165 37.000 111.835 ;
        RECT 36.240 110.915 37.000 111.165 ;
        RECT 37.170 111.450 37.340 112.185 ;
        RECT 37.510 112.065 37.840 113.565 ;
        RECT 38.605 113.060 38.935 113.565 ;
        RECT 39.530 112.890 39.860 113.045 ;
        RECT 38.070 112.720 39.860 112.890 ;
        RECT 40.060 112.830 40.310 113.045 ;
        RECT 41.005 113.000 41.335 113.565 ;
        RECT 41.985 112.970 42.235 113.565 ;
        RECT 42.435 112.840 42.765 113.300 ;
        RECT 42.965 112.840 43.215 113.565 ;
        RECT 40.060 112.800 41.815 112.830 ;
        RECT 42.435 112.800 42.635 112.840 ;
        RECT 38.070 112.640 38.705 112.720 ;
        RECT 38.035 112.115 38.365 112.470 ;
        RECT 38.535 111.895 38.705 112.640 ;
        RECT 37.670 111.565 38.705 111.895 ;
        RECT 37.170 111.395 37.500 111.450 ;
        RECT 38.875 111.395 39.055 112.445 ;
        RECT 37.170 111.225 39.055 111.395 ;
        RECT 39.225 111.370 39.395 112.720 ;
        RECT 40.060 112.660 42.635 112.800 ;
        RECT 40.060 112.550 40.310 112.660 ;
        RECT 41.645 112.630 42.635 112.660 ;
        RECT 39.565 112.380 40.310 112.550 ;
        RECT 39.565 111.710 39.735 112.380 ;
        RECT 40.555 112.210 40.805 112.490 ;
        RECT 39.905 112.040 40.805 112.210 ;
        RECT 41.455 112.130 41.865 112.460 ;
        RECT 39.905 111.880 40.455 112.040 ;
        RECT 39.565 111.540 40.115 111.710 ;
        RECT 37.170 110.985 37.500 111.225 ;
        RECT 37.670 110.885 39.055 111.055 ;
        RECT 39.225 110.990 39.695 111.370 ;
        RECT 39.865 110.990 40.115 111.540 ;
        RECT 40.285 111.120 40.455 111.880 ;
        RECT 41.045 111.960 41.275 112.100 ;
        RECT 40.625 111.460 40.875 111.870 ;
        RECT 41.045 111.630 41.525 111.960 ;
        RECT 41.695 111.460 41.865 112.130 ;
        RECT 40.625 111.290 41.865 111.460 ;
        RECT 42.035 111.450 42.295 112.460 ;
        RECT 37.670 110.745 37.840 110.885 ;
        RECT 35.900 110.575 37.840 110.745 ;
        RECT 38.885 110.820 39.055 110.885 ;
        RECT 40.285 110.820 40.810 111.120 ;
        RECT 38.010 110.405 38.405 110.715 ;
        RECT 38.885 110.650 40.810 110.820 ;
        RECT 40.980 110.405 41.310 111.120 ;
        RECT 41.480 110.670 41.865 111.290 ;
        RECT 42.465 111.150 42.635 112.630 ;
        RECT 42.805 111.320 43.195 112.490 ;
        RECT 47.255 112.250 47.585 113.565 ;
        RECT 42.040 110.405 42.290 111.150 ;
        RECT 42.465 110.980 43.190 111.150 ;
        RECT 42.860 110.690 43.190 110.980 ;
        RECT 47.330 110.405 47.900 111.905 ;
        RECT 48.305 111.570 48.875 113.565 ;
        RECT 49.170 112.525 49.470 113.565 ;
        RECT 53.495 112.250 53.825 113.565 ;
        RECT 48.610 110.405 48.940 111.125 ;
        RECT 49.170 110.405 49.470 111.425 ;
        RECT 53.570 110.405 54.140 111.905 ;
        RECT 54.545 111.570 55.115 113.565 ;
        RECT 56.865 112.840 57.115 113.565 ;
        RECT 57.315 112.840 57.645 113.300 ;
        RECT 57.845 112.970 58.095 113.565 ;
        RECT 58.745 113.000 59.075 113.565 ;
        RECT 61.145 113.060 61.475 113.565 ;
        RECT 57.445 112.800 57.645 112.840 ;
        RECT 59.770 112.830 60.020 113.045 ;
        RECT 58.265 112.800 60.020 112.830 ;
        RECT 57.445 112.660 60.020 112.800 ;
        RECT 60.220 112.890 60.550 113.045 ;
        RECT 60.220 112.720 62.010 112.890 ;
        RECT 57.445 112.630 58.435 112.660 ;
        RECT 56.885 111.320 57.275 112.490 ;
        RECT 57.445 111.150 57.615 112.630 ;
        RECT 59.770 112.550 60.020 112.660 ;
        RECT 57.785 111.450 58.045 112.460 ;
        RECT 58.215 112.130 58.625 112.460 ;
        RECT 59.275 112.210 59.525 112.490 ;
        RECT 59.770 112.380 60.515 112.550 ;
        RECT 58.215 111.460 58.385 112.130 ;
        RECT 58.805 111.960 59.035 112.100 ;
        RECT 59.275 112.040 60.175 112.210 ;
        RECT 58.555 111.630 59.035 111.960 ;
        RECT 59.625 111.880 60.175 112.040 ;
        RECT 59.205 111.460 59.455 111.870 ;
        RECT 58.215 111.290 59.455 111.460 ;
        RECT 54.850 110.405 55.180 111.125 ;
        RECT 56.890 110.980 57.615 111.150 ;
        RECT 56.890 110.690 57.220 110.980 ;
        RECT 57.790 110.405 58.040 111.150 ;
        RECT 58.215 110.670 58.600 111.290 ;
        RECT 59.625 111.120 59.795 111.880 ;
        RECT 60.345 111.710 60.515 112.380 ;
        RECT 58.770 110.405 59.100 111.120 ;
        RECT 59.270 110.820 59.795 111.120 ;
        RECT 59.965 111.540 60.515 111.710 ;
        RECT 59.965 110.990 60.215 111.540 ;
        RECT 60.685 111.370 60.855 112.720 ;
        RECT 61.375 112.640 62.010 112.720 ;
        RECT 60.385 110.990 60.855 111.370 ;
        RECT 61.025 111.395 61.205 112.445 ;
        RECT 61.375 111.895 61.545 112.640 ;
        RECT 61.715 112.115 62.045 112.470 ;
        RECT 62.240 112.065 62.570 113.565 ;
        RECT 62.740 112.185 63.070 113.075 ;
        RECT 63.240 112.795 64.395 113.125 ;
        RECT 61.375 111.565 62.410 111.895 ;
        RECT 62.740 111.450 62.910 112.185 ;
        RECT 63.240 112.005 63.410 112.795 ;
        RECT 62.580 111.395 62.910 111.450 ;
        RECT 61.025 111.225 62.910 111.395 ;
        RECT 61.025 110.885 62.410 111.055 ;
        RECT 62.580 110.985 62.910 111.225 ;
        RECT 63.080 111.835 63.410 112.005 ;
        RECT 63.080 111.165 63.250 111.835 ;
        RECT 63.725 111.665 64.055 112.625 ;
        RECT 64.225 112.005 64.395 112.795 ;
        RECT 64.565 112.765 64.895 113.565 ;
        RECT 65.080 112.765 65.445 113.225 ;
        RECT 64.565 112.240 65.105 112.575 ;
        RECT 65.275 112.345 65.445 112.765 ;
        RECT 65.615 112.515 65.945 113.565 ;
        RECT 65.275 112.175 65.950 112.345 ;
        RECT 64.225 111.835 65.610 112.005 ;
        RECT 65.280 111.675 65.610 111.835 ;
        RECT 63.450 111.335 64.180 111.665 ;
        RECT 64.350 111.505 64.680 111.665 ;
        RECT 65.780 111.505 65.950 112.175 ;
        RECT 66.145 112.035 66.315 113.225 ;
        RECT 66.485 112.205 67.185 113.300 ;
        RECT 66.145 111.705 66.695 112.035 ;
        RECT 64.350 111.335 65.950 111.505 ;
        RECT 63.080 110.915 63.840 111.165 ;
        RECT 61.025 110.820 61.195 110.885 ;
        RECT 59.270 110.650 61.195 110.820 ;
        RECT 62.240 110.745 62.410 110.885 ;
        RECT 64.010 110.745 64.180 111.335 ;
        RECT 61.675 110.405 62.070 110.715 ;
        RECT 62.240 110.575 64.180 110.745 ;
        RECT 64.505 110.405 64.835 111.165 ;
        RECT 65.375 110.705 65.705 111.335 ;
        RECT 65.935 110.405 66.185 111.165 ;
        RECT 66.365 110.670 66.695 111.705 ;
        RECT 66.925 111.450 67.185 112.205 ;
        RECT 67.355 112.140 67.685 113.565 ;
        RECT 68.005 111.570 68.575 113.565 ;
        RECT 69.295 112.250 69.625 113.565 ;
        RECT 66.925 110.670 67.255 111.450 ;
        RECT 67.435 110.405 67.685 111.450 ;
        RECT 67.940 110.405 68.270 111.125 ;
        RECT 68.980 110.405 69.550 111.905 ;
        RECT 10.200 110.235 69.720 110.405 ;
        RECT 10.370 108.735 10.940 110.235 ;
        RECT 11.650 109.515 11.980 110.235 ;
        RECT 10.295 107.075 10.625 108.390 ;
        RECT 11.345 107.075 11.915 109.070 ;
        RECT 12.290 108.735 12.860 110.235 ;
        RECT 13.570 109.515 13.900 110.235 ;
        RECT 15.115 109.360 15.445 109.970 ;
        RECT 15.615 109.640 16.305 110.235 ;
        RECT 16.475 109.530 16.805 109.970 ;
        RECT 15.115 109.190 16.395 109.360 ;
        RECT 12.215 107.075 12.545 108.390 ;
        RECT 13.265 107.075 13.835 109.070 ;
        RECT 15.125 108.540 15.835 109.020 ;
        RECT 16.005 108.690 16.395 109.190 ;
        RECT 16.005 108.370 16.175 108.690 ;
        RECT 16.565 108.500 16.805 109.530 ;
        RECT 15.345 108.200 16.175 108.370 ;
        RECT 15.345 107.340 15.675 108.200 ;
        RECT 15.845 107.075 16.175 108.030 ;
        RECT 16.345 107.340 16.805 108.500 ;
        RECT 20.875 109.530 21.205 109.970 ;
        RECT 21.375 109.640 22.065 110.235 ;
        RECT 20.875 108.500 21.115 109.530 ;
        RECT 22.235 109.360 22.565 109.970 ;
        RECT 21.285 109.190 22.565 109.360 ;
        RECT 23.755 109.530 24.085 109.970 ;
        RECT 24.255 109.640 24.945 110.235 ;
        RECT 21.285 108.690 21.675 109.190 ;
        RECT 20.875 107.340 21.335 108.500 ;
        RECT 21.505 108.370 21.675 108.690 ;
        RECT 21.845 108.540 22.555 109.020 ;
        RECT 23.755 108.500 23.995 109.530 ;
        RECT 25.115 109.360 25.445 109.970 ;
        RECT 24.165 109.190 25.445 109.360 ;
        RECT 24.165 108.690 24.555 109.190 ;
        RECT 21.505 108.200 22.335 108.370 ;
        RECT 21.505 107.075 21.835 108.030 ;
        RECT 22.005 107.340 22.335 108.200 ;
        RECT 23.755 107.340 24.215 108.500 ;
        RECT 24.385 108.370 24.555 108.690 ;
        RECT 24.725 108.540 25.435 109.020 ;
        RECT 25.730 108.735 26.300 110.235 ;
        RECT 27.010 109.515 27.340 110.235 ;
        RECT 27.595 109.360 27.860 109.780 ;
        RECT 28.030 109.530 28.700 110.235 ;
        RECT 27.595 109.190 29.165 109.360 ;
        RECT 29.335 109.190 29.735 109.970 ;
        RECT 24.385 108.200 25.215 108.370 ;
        RECT 24.385 107.075 24.715 108.030 ;
        RECT 24.885 107.340 25.215 108.200 ;
        RECT 25.655 107.075 25.985 108.390 ;
        RECT 26.705 107.075 27.275 109.070 ;
        RECT 28.995 109.020 29.165 109.190 ;
        RECT 27.585 108.540 28.315 109.020 ;
        RECT 28.495 108.540 28.825 108.970 ;
        RECT 28.995 108.690 29.395 109.020 ;
        RECT 28.995 108.370 29.165 108.690 ;
        RECT 27.595 108.200 29.165 108.370 ;
        RECT 27.595 107.620 27.925 108.200 ;
        RECT 29.565 108.030 29.735 109.190 ;
        RECT 30.050 108.735 30.620 110.235 ;
        RECT 31.330 109.515 31.660 110.235 ;
        RECT 31.915 109.530 32.245 109.970 ;
        RECT 32.415 109.640 33.105 110.235 ;
        RECT 28.130 107.075 28.395 108.030 ;
        RECT 28.565 107.860 29.735 108.030 ;
        RECT 28.565 107.340 29.045 107.860 ;
        RECT 29.215 107.075 29.550 107.670 ;
        RECT 29.975 107.075 30.305 108.390 ;
        RECT 31.025 107.075 31.595 109.070 ;
        RECT 31.915 108.500 32.155 109.530 ;
        RECT 33.275 109.360 33.605 109.970 ;
        RECT 32.325 109.190 33.605 109.360 ;
        RECT 32.325 108.690 32.715 109.190 ;
        RECT 31.915 107.340 32.375 108.500 ;
        RECT 32.545 108.370 32.715 108.690 ;
        RECT 32.885 108.540 33.595 109.020 ;
        RECT 33.890 108.735 34.460 110.235 ;
        RECT 35.170 109.515 35.500 110.235 ;
        RECT 36.210 109.215 36.510 110.235 ;
        RECT 37.195 109.310 37.525 109.870 ;
        RECT 37.705 109.480 38.035 110.235 ;
        RECT 37.195 109.140 37.995 109.310 ;
        RECT 38.205 109.140 38.535 109.970 ;
        RECT 38.715 109.190 38.965 110.235 ;
        RECT 44.890 109.660 45.220 109.950 ;
        RECT 44.890 109.490 45.615 109.660 ;
        RECT 45.790 109.490 46.040 110.235 ;
        RECT 32.545 108.200 33.375 108.370 ;
        RECT 32.545 107.075 32.875 108.030 ;
        RECT 33.045 107.340 33.375 108.200 ;
        RECT 33.815 107.075 34.145 108.390 ;
        RECT 34.865 107.075 35.435 109.070 ;
        RECT 37.205 108.540 37.655 108.970 ;
        RECT 36.210 107.075 36.510 108.115 ;
        RECT 37.195 108.000 37.550 108.370 ;
        RECT 37.825 108.000 37.995 109.140 ;
        RECT 38.165 108.170 38.535 109.140 ;
        RECT 38.705 108.690 39.375 109.020 ;
        RECT 38.705 108.000 38.875 108.690 ;
        RECT 37.195 107.830 38.875 108.000 ;
        RECT 37.195 107.440 37.550 107.830 ;
        RECT 37.755 107.075 38.085 107.660 ;
        RECT 39.060 107.585 39.365 108.500 ;
        RECT 44.885 108.150 45.275 109.320 ;
        RECT 45.445 108.010 45.615 109.490 ;
        RECT 46.215 109.350 46.600 109.970 ;
        RECT 46.770 109.520 47.100 110.235 ;
        RECT 47.270 109.820 49.195 109.990 ;
        RECT 49.675 109.925 50.070 110.235 ;
        RECT 47.270 109.520 47.795 109.820 ;
        RECT 49.025 109.755 49.195 109.820 ;
        RECT 50.240 109.895 52.180 110.065 ;
        RECT 50.240 109.755 50.410 109.895 ;
        RECT 45.785 108.180 46.045 109.190 ;
        RECT 46.215 109.180 47.455 109.350 ;
        RECT 46.215 108.510 46.385 109.180 ;
        RECT 46.555 108.680 47.035 109.010 ;
        RECT 47.205 108.770 47.455 109.180 ;
        RECT 46.805 108.540 47.035 108.680 ;
        RECT 47.625 108.760 47.795 109.520 ;
        RECT 47.965 109.100 48.215 109.650 ;
        RECT 48.385 109.270 48.855 109.650 ;
        RECT 49.025 109.585 50.410 109.755 ;
        RECT 50.580 109.415 50.910 109.655 ;
        RECT 47.965 108.930 48.515 109.100 ;
        RECT 47.625 108.600 48.175 108.760 ;
        RECT 46.215 108.180 46.625 108.510 ;
        RECT 47.275 108.430 48.175 108.600 ;
        RECT 47.275 108.150 47.525 108.430 ;
        RECT 48.345 108.260 48.515 108.930 ;
        RECT 47.770 108.090 48.515 108.260 ;
        RECT 45.445 107.980 46.435 108.010 ;
        RECT 47.770 107.980 48.020 108.090 ;
        RECT 45.445 107.840 48.020 107.980 ;
        RECT 48.685 107.920 48.855 109.270 ;
        RECT 49.025 109.245 50.910 109.415 ;
        RECT 49.025 108.195 49.205 109.245 ;
        RECT 50.580 109.190 50.910 109.245 ;
        RECT 49.375 108.745 50.410 109.075 ;
        RECT 49.375 108.000 49.545 108.745 ;
        RECT 49.715 108.170 50.045 108.525 ;
        RECT 49.375 107.920 50.010 108.000 ;
        RECT 45.445 107.800 45.645 107.840 ;
        RECT 46.265 107.810 48.020 107.840 ;
        RECT 38.655 107.075 39.365 107.585 ;
        RECT 44.865 107.075 45.115 107.800 ;
        RECT 45.315 107.340 45.645 107.800 ;
        RECT 45.845 107.075 46.095 107.670 ;
        RECT 46.745 107.075 47.075 107.640 ;
        RECT 47.770 107.595 48.020 107.810 ;
        RECT 48.220 107.750 50.010 107.920 ;
        RECT 48.220 107.595 48.550 107.750 ;
        RECT 49.145 107.075 49.475 107.580 ;
        RECT 50.240 107.075 50.570 108.575 ;
        RECT 50.740 108.455 50.910 109.190 ;
        RECT 51.080 109.475 51.840 109.725 ;
        RECT 51.080 108.805 51.250 109.475 ;
        RECT 52.010 109.305 52.180 109.895 ;
        RECT 52.505 109.475 52.835 110.235 ;
        RECT 53.375 109.305 53.705 109.935 ;
        RECT 53.935 109.475 54.185 110.235 ;
        RECT 51.450 108.975 52.180 109.305 ;
        RECT 52.350 109.135 53.950 109.305 ;
        RECT 52.350 108.975 52.680 109.135 ;
        RECT 51.080 108.635 51.410 108.805 ;
        RECT 50.740 107.565 51.070 108.455 ;
        RECT 51.240 107.845 51.410 108.635 ;
        RECT 51.725 108.015 52.055 108.975 ;
        RECT 53.280 108.805 53.610 108.965 ;
        RECT 52.225 108.635 53.610 108.805 ;
        RECT 52.225 107.845 52.395 108.635 ;
        RECT 53.780 108.465 53.950 109.135 ;
        RECT 54.365 108.935 54.695 109.970 ;
        RECT 52.565 108.065 53.105 108.400 ;
        RECT 53.275 108.295 53.950 108.465 ;
        RECT 54.145 108.605 54.695 108.935 ;
        RECT 54.925 109.190 55.255 109.970 ;
        RECT 55.435 109.190 55.685 110.235 ;
        RECT 53.275 107.875 53.445 108.295 ;
        RECT 51.240 107.515 52.395 107.845 ;
        RECT 52.565 107.075 52.895 107.875 ;
        RECT 53.080 107.415 53.445 107.875 ;
        RECT 53.615 107.075 53.945 108.125 ;
        RECT 54.145 107.415 54.315 108.605 ;
        RECT 54.925 108.435 55.185 109.190 ;
        RECT 55.970 108.735 56.540 110.235 ;
        RECT 57.250 109.515 57.580 110.235 ;
        RECT 59.245 109.510 59.620 109.840 ;
        RECT 59.790 109.510 60.120 110.235 ;
        RECT 54.485 107.340 55.185 108.435 ;
        RECT 55.355 107.075 55.685 108.500 ;
        RECT 55.895 107.075 56.225 108.390 ;
        RECT 56.945 107.075 57.515 109.070 ;
        RECT 59.245 108.740 59.415 109.510 ;
        RECT 60.290 109.340 60.620 109.970 ;
        RECT 60.800 109.510 60.970 110.235 ;
        RECT 61.150 109.340 61.480 109.970 ;
        RECT 61.660 109.510 61.910 110.235 ;
        RECT 59.585 108.910 59.985 109.240 ;
        RECT 60.290 109.170 61.505 109.340 ;
        RECT 62.130 109.215 62.430 110.235 ;
        RECT 60.155 108.740 61.165 108.970 ;
        RECT 59.245 108.570 61.165 108.740 ;
        RECT 59.245 107.340 59.625 108.570 ;
        RECT 61.335 108.400 61.505 109.170 ;
        RECT 62.690 108.735 63.260 110.235 ;
        RECT 63.970 109.515 64.300 110.235 ;
        RECT 65.005 109.510 65.380 109.840 ;
        RECT 65.550 109.510 65.880 110.235 ;
        RECT 59.795 107.075 60.045 108.400 ;
        RECT 60.245 108.230 61.505 108.400 ;
        RECT 60.245 107.340 60.575 108.230 ;
        RECT 60.775 107.075 61.025 108.060 ;
        RECT 61.225 107.340 61.505 108.230 ;
        RECT 61.675 107.075 61.925 108.500 ;
        RECT 62.130 107.075 62.430 108.115 ;
        RECT 62.615 107.075 62.945 108.390 ;
        RECT 63.665 107.075 64.235 109.070 ;
        RECT 65.005 108.740 65.175 109.510 ;
        RECT 66.050 109.340 66.380 109.970 ;
        RECT 66.560 109.510 66.730 110.235 ;
        RECT 66.910 109.340 67.240 109.970 ;
        RECT 67.420 109.510 67.670 110.235 ;
        RECT 67.940 109.515 68.270 110.235 ;
        RECT 65.345 108.910 65.745 109.240 ;
        RECT 66.050 109.170 67.265 109.340 ;
        RECT 65.915 108.740 66.925 108.970 ;
        RECT 65.005 108.570 66.925 108.740 ;
        RECT 65.005 107.340 65.385 108.570 ;
        RECT 67.095 108.400 67.265 109.170 ;
        RECT 65.555 107.075 65.805 108.400 ;
        RECT 66.005 108.230 67.265 108.400 ;
        RECT 66.005 107.340 66.335 108.230 ;
        RECT 66.535 107.075 66.785 108.060 ;
        RECT 66.985 107.340 67.265 108.230 ;
        RECT 67.435 107.075 67.685 108.500 ;
        RECT 68.005 107.075 68.575 109.070 ;
        RECT 68.980 108.735 69.550 110.235 ;
        RECT 69.295 107.075 69.625 108.390 ;
        RECT 10.200 106.905 69.720 107.075 ;
        RECT 10.295 105.590 10.625 106.905 ;
        RECT 10.370 103.745 10.940 105.245 ;
        RECT 11.345 104.910 11.915 106.905 ;
        RECT 12.240 105.690 12.570 106.905 ;
        RECT 12.750 105.520 12.970 106.640 ;
        RECT 13.160 105.690 13.490 106.905 ;
        RECT 13.670 105.520 13.880 106.640 ;
        RECT 14.060 105.690 14.390 106.905 ;
        RECT 14.570 105.520 14.775 106.640 ;
        RECT 14.960 105.690 15.290 106.905 ;
        RECT 15.475 105.520 15.680 106.640 ;
        RECT 15.860 105.690 16.190 106.905 ;
        RECT 16.370 105.520 16.580 106.640 ;
        RECT 16.760 105.690 17.090 106.905 ;
        RECT 17.290 105.520 17.490 106.640 ;
        RECT 17.660 105.690 17.990 106.905 ;
        RECT 18.175 105.520 18.380 106.640 ;
        RECT 18.560 105.690 18.890 106.905 ;
        RECT 19.060 105.780 19.290 106.640 ;
        RECT 19.470 105.950 19.720 106.905 ;
        RECT 19.920 105.780 20.250 106.640 ;
        RECT 20.450 105.950 20.620 106.905 ;
        RECT 20.820 105.780 21.150 106.640 ;
        RECT 12.750 105.490 12.995 105.520 ;
        RECT 11.650 103.745 11.980 104.465 ;
        RECT 12.235 103.745 12.565 104.405 ;
        RECT 12.745 104.010 12.995 105.490 ;
        RECT 13.670 105.350 13.925 105.520 ;
        RECT 14.570 105.350 14.855 105.520 ;
        RECT 15.475 105.350 15.785 105.520 ;
        RECT 16.370 105.350 16.695 105.520 ;
        RECT 17.290 105.350 17.550 105.520 ;
        RECT 18.175 105.350 18.445 105.520 ;
        RECT 13.165 104.850 13.495 105.180 ;
        RECT 13.165 103.745 13.495 104.340 ;
        RECT 13.675 104.010 13.925 105.350 ;
        RECT 14.095 104.850 14.425 105.180 ;
        RECT 14.095 103.745 14.425 104.340 ;
        RECT 14.605 104.010 14.855 105.350 ;
        RECT 15.025 104.850 15.355 105.180 ;
        RECT 15.025 103.745 15.355 104.340 ;
        RECT 15.535 104.010 15.785 105.350 ;
        RECT 15.965 104.850 16.295 105.180 ;
        RECT 15.955 103.745 16.285 104.340 ;
        RECT 16.465 104.010 16.695 105.350 ;
        RECT 16.880 104.850 17.210 105.180 ;
        RECT 17.380 104.405 17.550 105.350 ;
        RECT 17.720 104.850 18.050 105.180 ;
        RECT 16.885 103.745 17.210 104.400 ;
        RECT 17.380 104.010 17.645 104.405 ;
        RECT 17.825 103.745 18.050 104.385 ;
        RECT 18.220 104.010 18.445 105.350 ;
        RECT 18.615 104.850 18.885 105.180 ;
        RECT 18.685 103.745 18.855 104.340 ;
        RECT 19.060 104.010 19.330 105.780 ;
        RECT 19.585 105.610 21.150 105.780 ;
        RECT 21.350 105.610 21.600 106.905 ;
        RECT 23.250 105.865 23.550 106.905 ;
        RECT 19.585 105.070 19.755 105.610 ;
        RECT 23.965 105.600 24.295 106.905 ;
        RECT 24.585 105.780 25.165 106.640 ;
        RECT 25.395 106.120 25.725 106.640 ;
        RECT 25.895 106.310 26.335 106.905 ;
        RECT 26.505 106.120 26.835 106.640 ;
        RECT 25.395 105.950 26.835 106.120 ;
        RECT 24.585 105.610 26.835 105.780 ;
        RECT 19.510 104.840 19.755 105.070 ;
        RECT 19.925 105.010 21.595 105.440 ;
        RECT 23.745 104.840 24.415 105.275 ;
        RECT 19.585 104.810 19.755 104.840 ;
        RECT 19.585 104.640 21.175 104.810 ;
        RECT 19.535 103.745 19.865 104.470 ;
        RECT 20.045 104.010 20.295 104.640 ;
        RECT 20.495 103.745 20.745 104.470 ;
        RECT 20.925 104.010 21.175 104.640 ;
        RECT 21.355 103.745 21.605 104.470 ;
        RECT 23.250 103.745 23.550 104.765 ;
        RECT 24.585 104.700 24.755 105.610 ;
        RECT 26.155 105.355 26.485 105.440 ;
        RECT 24.925 105.025 26.485 105.355 ;
        RECT 26.155 105.010 26.485 105.025 ;
        RECT 26.665 105.310 26.835 105.610 ;
        RECT 27.005 105.480 27.395 106.640 ;
        RECT 26.665 104.980 27.055 105.310 ;
        RECT 23.815 103.745 24.415 104.650 ;
        RECT 24.585 104.370 25.280 104.700 ;
        RECT 25.460 103.745 25.790 104.855 ;
        RECT 27.225 104.810 27.395 105.480 ;
        RECT 26.165 104.640 27.395 104.810 ;
        RECT 27.565 105.480 28.085 106.640 ;
        RECT 28.255 105.610 28.585 106.905 ;
        RECT 29.210 105.650 29.540 106.520 ;
        RECT 29.895 105.760 30.225 106.905 ;
        RECT 28.975 105.480 29.540 105.650 ;
        RECT 30.395 105.590 30.725 106.640 ;
        RECT 27.565 104.790 27.735 105.480 ;
        RECT 27.905 104.960 28.305 105.290 ;
        RECT 28.475 105.010 28.805 105.440 ;
        RECT 28.135 104.840 28.305 104.960 ;
        RECT 28.975 104.840 29.145 105.480 ;
        RECT 30.010 105.420 30.725 105.590 ;
        RECT 30.955 105.480 31.415 106.640 ;
        RECT 31.585 105.950 31.915 106.905 ;
        RECT 32.085 105.780 32.415 106.640 ;
        RECT 31.585 105.610 32.415 105.780 ;
        RECT 30.010 105.290 30.180 105.420 ;
        RECT 29.315 104.960 30.180 105.290 ;
        RECT 26.165 104.075 26.610 104.640 ;
        RECT 26.850 103.745 27.180 104.405 ;
        RECT 27.565 104.010 27.965 104.790 ;
        RECT 28.135 104.670 29.145 104.840 ;
        RECT 28.160 103.745 28.575 104.500 ;
        RECT 28.795 104.200 29.145 104.670 ;
        RECT 29.315 103.745 29.840 104.790 ;
        RECT 30.010 104.670 30.180 104.960 ;
        RECT 30.385 104.840 30.715 105.210 ;
        RECT 30.010 104.340 30.725 104.670 ;
        RECT 30.955 104.450 31.195 105.480 ;
        RECT 31.585 105.290 31.755 105.610 ;
        RECT 32.875 105.480 33.205 106.905 ;
        RECT 33.375 105.545 34.075 106.640 ;
        RECT 31.365 104.790 31.755 105.290 ;
        RECT 31.925 104.960 32.635 105.440 ;
        RECT 33.375 104.790 33.635 105.545 ;
        RECT 34.245 105.375 34.415 106.565 ;
        RECT 34.615 105.855 34.945 106.905 ;
        RECT 35.115 106.105 35.480 106.565 ;
        RECT 35.665 106.105 35.995 106.905 ;
        RECT 36.165 106.135 37.320 106.465 ;
        RECT 35.115 105.685 35.285 106.105 ;
        RECT 31.365 104.620 32.645 104.790 ;
        RECT 30.955 104.010 31.285 104.450 ;
        RECT 31.455 103.745 32.145 104.340 ;
        RECT 32.315 104.010 32.645 104.620 ;
        RECT 32.875 103.745 33.125 104.790 ;
        RECT 33.305 104.010 33.635 104.790 ;
        RECT 33.865 105.045 34.415 105.375 ;
        RECT 34.610 105.515 35.285 105.685 ;
        RECT 35.455 105.580 35.995 105.915 ;
        RECT 33.865 104.010 34.195 105.045 ;
        RECT 34.610 104.845 34.780 105.515 ;
        RECT 36.165 105.345 36.335 106.135 ;
        RECT 34.950 105.175 36.335 105.345 ;
        RECT 34.950 105.015 35.280 105.175 ;
        RECT 36.505 105.005 36.835 105.965 ;
        RECT 37.150 105.345 37.320 106.135 ;
        RECT 37.490 105.525 37.820 106.415 ;
        RECT 37.150 105.175 37.480 105.345 ;
        RECT 35.880 104.845 36.210 105.005 ;
        RECT 34.610 104.675 36.210 104.845 ;
        RECT 36.380 104.675 37.110 105.005 ;
        RECT 34.375 103.745 34.625 104.505 ;
        RECT 34.855 104.045 35.185 104.675 ;
        RECT 35.725 103.745 36.055 104.505 ;
        RECT 36.380 104.085 36.550 104.675 ;
        RECT 37.310 104.505 37.480 105.175 ;
        RECT 36.720 104.255 37.480 104.505 ;
        RECT 37.650 104.790 37.820 105.525 ;
        RECT 37.990 105.405 38.320 106.905 ;
        RECT 39.085 106.400 39.415 106.905 ;
        RECT 40.010 106.230 40.340 106.385 ;
        RECT 38.550 106.060 40.340 106.230 ;
        RECT 40.540 106.170 40.790 106.385 ;
        RECT 41.485 106.340 41.815 106.905 ;
        RECT 42.465 106.310 42.715 106.905 ;
        RECT 42.915 106.180 43.245 106.640 ;
        RECT 43.445 106.180 43.695 106.905 ;
        RECT 40.540 106.140 42.295 106.170 ;
        RECT 42.915 106.140 43.115 106.180 ;
        RECT 38.550 105.980 39.185 106.060 ;
        RECT 38.515 105.455 38.845 105.810 ;
        RECT 39.015 105.235 39.185 105.980 ;
        RECT 38.150 104.905 39.185 105.235 ;
        RECT 37.650 104.735 37.980 104.790 ;
        RECT 39.355 104.735 39.535 105.785 ;
        RECT 37.650 104.565 39.535 104.735 ;
        RECT 39.705 104.710 39.875 106.060 ;
        RECT 40.540 106.000 43.115 106.140 ;
        RECT 40.540 105.890 40.790 106.000 ;
        RECT 42.125 105.970 43.115 106.000 ;
        RECT 40.045 105.720 40.790 105.890 ;
        RECT 40.045 105.050 40.215 105.720 ;
        RECT 41.035 105.550 41.285 105.830 ;
        RECT 40.385 105.380 41.285 105.550 ;
        RECT 41.935 105.470 42.345 105.800 ;
        RECT 40.385 105.220 40.935 105.380 ;
        RECT 40.045 104.880 40.595 105.050 ;
        RECT 37.650 104.325 37.980 104.565 ;
        RECT 38.150 104.225 39.535 104.395 ;
        RECT 39.705 104.330 40.175 104.710 ;
        RECT 40.345 104.330 40.595 104.880 ;
        RECT 40.765 104.460 40.935 105.220 ;
        RECT 41.525 105.300 41.755 105.440 ;
        RECT 41.105 104.800 41.355 105.210 ;
        RECT 41.525 104.970 42.005 105.300 ;
        RECT 42.175 104.800 42.345 105.470 ;
        RECT 41.105 104.630 42.345 104.800 ;
        RECT 42.515 104.790 42.775 105.800 ;
        RECT 38.150 104.085 38.320 104.225 ;
        RECT 36.380 103.915 38.320 104.085 ;
        RECT 39.365 104.160 39.535 104.225 ;
        RECT 40.765 104.160 41.290 104.460 ;
        RECT 38.490 103.745 38.885 104.055 ;
        RECT 39.365 103.990 41.290 104.160 ;
        RECT 41.460 103.745 41.790 104.460 ;
        RECT 41.960 104.010 42.345 104.630 ;
        RECT 42.945 104.490 43.115 105.970 ;
        RECT 43.285 104.660 43.675 105.830 ;
        RECT 43.895 105.590 44.225 106.905 ;
        RECT 42.520 103.745 42.770 104.490 ;
        RECT 42.945 104.320 43.670 104.490 ;
        RECT 43.340 104.030 43.670 104.320 ;
        RECT 43.970 103.745 44.540 105.245 ;
        RECT 44.945 104.910 45.515 106.905 ;
        RECT 46.795 106.150 47.150 106.540 ;
        RECT 47.355 106.320 47.685 106.905 ;
        RECT 48.255 106.395 48.965 106.905 ;
        RECT 46.795 105.980 48.475 106.150 ;
        RECT 46.795 105.610 47.150 105.980 ;
        RECT 46.805 105.010 47.255 105.440 ;
        RECT 47.425 104.840 47.595 105.980 ;
        RECT 47.765 104.840 48.135 105.810 ;
        RECT 48.305 105.290 48.475 105.980 ;
        RECT 48.660 105.480 48.965 106.395 ;
        RECT 49.170 105.865 49.470 106.905 ;
        RECT 49.665 106.180 49.915 106.905 ;
        RECT 50.115 106.180 50.445 106.640 ;
        RECT 50.645 106.310 50.895 106.905 ;
        RECT 51.545 106.340 51.875 106.905 ;
        RECT 53.945 106.400 54.275 106.905 ;
        RECT 50.245 106.140 50.445 106.180 ;
        RECT 52.570 106.170 52.820 106.385 ;
        RECT 51.065 106.140 52.820 106.170 ;
        RECT 50.245 106.000 52.820 106.140 ;
        RECT 53.020 106.230 53.350 106.385 ;
        RECT 53.020 106.060 54.810 106.230 ;
        RECT 50.245 105.970 51.235 106.000 ;
        RECT 48.305 104.960 48.975 105.290 ;
        RECT 46.795 104.670 47.595 104.840 ;
        RECT 45.250 103.745 45.580 104.465 ;
        RECT 46.795 104.110 47.125 104.670 ;
        RECT 47.305 103.745 47.635 104.500 ;
        RECT 47.805 104.010 48.135 104.840 ;
        RECT 48.315 103.745 48.565 104.790 ;
        RECT 49.170 103.745 49.470 104.765 ;
        RECT 49.685 104.660 50.075 105.830 ;
        RECT 50.245 104.490 50.415 105.970 ;
        RECT 52.570 105.890 52.820 106.000 ;
        RECT 50.585 104.790 50.845 105.800 ;
        RECT 51.015 105.470 51.425 105.800 ;
        RECT 52.075 105.550 52.325 105.830 ;
        RECT 52.570 105.720 53.315 105.890 ;
        RECT 51.015 104.800 51.185 105.470 ;
        RECT 51.605 105.300 51.835 105.440 ;
        RECT 52.075 105.380 52.975 105.550 ;
        RECT 51.355 104.970 51.835 105.300 ;
        RECT 52.425 105.220 52.975 105.380 ;
        RECT 52.005 104.800 52.255 105.210 ;
        RECT 51.015 104.630 52.255 104.800 ;
        RECT 49.690 104.320 50.415 104.490 ;
        RECT 49.690 104.030 50.020 104.320 ;
        RECT 50.590 103.745 50.840 104.490 ;
        RECT 51.015 104.010 51.400 104.630 ;
        RECT 52.425 104.460 52.595 105.220 ;
        RECT 53.145 105.050 53.315 105.720 ;
        RECT 51.570 103.745 51.900 104.460 ;
        RECT 52.070 104.160 52.595 104.460 ;
        RECT 52.765 104.880 53.315 105.050 ;
        RECT 52.765 104.330 53.015 104.880 ;
        RECT 53.485 104.710 53.655 106.060 ;
        RECT 54.175 105.980 54.810 106.060 ;
        RECT 53.185 104.330 53.655 104.710 ;
        RECT 53.825 104.735 54.005 105.785 ;
        RECT 54.175 105.235 54.345 105.980 ;
        RECT 54.515 105.455 54.845 105.810 ;
        RECT 55.040 105.405 55.370 106.905 ;
        RECT 55.540 105.525 55.870 106.415 ;
        RECT 56.040 106.135 57.195 106.465 ;
        RECT 54.175 104.905 55.210 105.235 ;
        RECT 55.540 104.790 55.710 105.525 ;
        RECT 56.040 105.345 56.210 106.135 ;
        RECT 55.380 104.735 55.710 104.790 ;
        RECT 53.825 104.565 55.710 104.735 ;
        RECT 53.825 104.225 55.210 104.395 ;
        RECT 55.380 104.325 55.710 104.565 ;
        RECT 55.880 105.175 56.210 105.345 ;
        RECT 55.880 104.505 56.050 105.175 ;
        RECT 56.525 105.005 56.855 105.965 ;
        RECT 57.025 105.345 57.195 106.135 ;
        RECT 57.365 106.105 57.695 106.905 ;
        RECT 57.880 106.105 58.245 106.565 ;
        RECT 57.365 105.580 57.905 105.915 ;
        RECT 58.075 105.685 58.245 106.105 ;
        RECT 58.415 105.855 58.745 106.905 ;
        RECT 58.075 105.515 58.750 105.685 ;
        RECT 57.025 105.175 58.410 105.345 ;
        RECT 58.080 105.015 58.410 105.175 ;
        RECT 56.250 104.675 56.980 105.005 ;
        RECT 57.150 104.845 57.480 105.005 ;
        RECT 58.580 104.845 58.750 105.515 ;
        RECT 58.945 105.375 59.115 106.565 ;
        RECT 59.285 105.545 59.985 106.640 ;
        RECT 58.945 105.045 59.495 105.375 ;
        RECT 57.150 104.675 58.750 104.845 ;
        RECT 55.880 104.255 56.640 104.505 ;
        RECT 53.825 104.160 53.995 104.225 ;
        RECT 52.070 103.990 53.995 104.160 ;
        RECT 55.040 104.085 55.210 104.225 ;
        RECT 56.810 104.085 56.980 104.675 ;
        RECT 54.475 103.745 54.870 104.055 ;
        RECT 55.040 103.915 56.980 104.085 ;
        RECT 57.305 103.745 57.635 104.505 ;
        RECT 58.175 104.045 58.505 104.675 ;
        RECT 58.735 103.745 58.985 104.505 ;
        RECT 59.165 104.010 59.495 105.045 ;
        RECT 59.725 104.790 59.985 105.545 ;
        RECT 60.155 105.480 60.485 106.905 ;
        RECT 62.125 105.410 62.505 106.640 ;
        RECT 62.675 105.580 62.925 106.905 ;
        RECT 63.125 105.750 63.455 106.640 ;
        RECT 63.655 105.920 63.905 106.905 ;
        RECT 64.105 105.750 64.385 106.640 ;
        RECT 63.125 105.580 64.385 105.750 ;
        RECT 62.125 105.240 64.045 105.410 ;
        RECT 59.725 104.010 60.055 104.790 ;
        RECT 60.235 103.745 60.485 104.790 ;
        RECT 62.125 104.470 62.295 105.240 ;
        RECT 62.465 104.740 62.865 105.070 ;
        RECT 63.035 105.010 64.045 105.240 ;
        RECT 64.215 104.810 64.385 105.580 ;
        RECT 64.555 105.480 64.805 106.905 ;
        RECT 63.170 104.640 64.385 104.810 ;
        RECT 65.005 105.410 65.385 106.640 ;
        RECT 65.555 105.580 65.805 106.905 ;
        RECT 66.005 105.750 66.335 106.640 ;
        RECT 66.535 105.920 66.785 106.905 ;
        RECT 66.985 105.750 67.265 106.640 ;
        RECT 66.005 105.580 67.265 105.750 ;
        RECT 65.005 105.240 66.925 105.410 ;
        RECT 62.125 104.140 62.500 104.470 ;
        RECT 62.670 103.745 63.000 104.470 ;
        RECT 63.170 104.010 63.500 104.640 ;
        RECT 63.680 103.745 63.850 104.470 ;
        RECT 64.030 104.010 64.360 104.640 ;
        RECT 65.005 104.470 65.175 105.240 ;
        RECT 65.345 104.740 65.745 105.070 ;
        RECT 65.915 105.010 66.925 105.240 ;
        RECT 67.095 104.810 67.265 105.580 ;
        RECT 67.435 105.480 67.685 106.905 ;
        RECT 68.005 104.910 68.575 106.905 ;
        RECT 69.295 105.590 69.625 106.905 ;
        RECT 66.050 104.640 67.265 104.810 ;
        RECT 64.540 103.745 64.790 104.470 ;
        RECT 65.005 104.140 65.380 104.470 ;
        RECT 65.550 103.745 65.880 104.470 ;
        RECT 66.050 104.010 66.380 104.640 ;
        RECT 66.560 103.745 66.730 104.470 ;
        RECT 66.910 104.010 67.240 104.640 ;
        RECT 67.420 103.745 67.670 104.470 ;
        RECT 67.940 103.745 68.270 104.465 ;
        RECT 68.980 103.745 69.550 105.245 ;
        RECT 10.200 103.575 69.720 103.745 ;
        RECT 10.370 102.075 10.940 103.575 ;
        RECT 11.650 102.855 11.980 103.575 ;
        RECT 13.675 102.700 13.925 103.310 ;
        RECT 14.105 102.870 14.355 103.575 ;
        RECT 14.525 103.235 15.375 103.405 ;
        RECT 14.525 102.700 14.695 103.235 ;
        RECT 13.675 102.530 14.695 102.700 ;
        RECT 10.295 100.415 10.625 101.730 ;
        RECT 11.345 100.415 11.915 102.410 ;
        RECT 13.685 101.880 14.065 102.360 ;
        RECT 14.235 102.110 14.695 102.530 ;
        RECT 14.865 102.310 15.035 103.065 ;
        RECT 15.205 102.930 15.375 103.235 ;
        RECT 15.545 103.100 15.875 103.575 ;
        RECT 16.045 103.215 17.320 103.385 ;
        RECT 16.045 102.930 16.215 103.215 ;
        RECT 15.205 102.760 16.215 102.930 ;
        RECT 14.235 101.710 14.405 102.110 ;
        RECT 14.865 101.980 15.320 102.310 ;
        RECT 14.865 101.840 15.035 101.980 ;
        RECT 13.675 101.540 14.405 101.710 ;
        RECT 13.675 100.680 14.005 101.540 ;
        RECT 14.205 100.415 14.375 101.370 ;
        RECT 14.575 101.035 15.035 101.840 ;
        RECT 15.530 101.635 15.810 102.535 ;
        RECT 15.430 101.305 15.810 101.635 ;
        RECT 15.980 102.420 16.535 102.590 ;
        RECT 15.980 101.035 16.150 102.420 ;
        RECT 16.715 102.250 16.980 103.045 ;
        RECT 16.320 102.080 16.980 102.250 ;
        RECT 17.150 102.970 17.320 103.215 ;
        RECT 17.630 103.140 17.880 103.575 ;
        RECT 18.050 103.235 19.455 103.405 ;
        RECT 18.050 102.970 18.220 103.235 ;
        RECT 19.125 103.150 19.455 103.235 ;
        RECT 17.150 102.800 18.220 102.970 ;
        RECT 16.320 101.375 16.490 102.080 ;
        RECT 17.150 101.910 17.320 102.800 ;
        RECT 18.390 102.630 18.560 103.065 ;
        RECT 18.780 102.680 19.380 102.930 ;
        RECT 17.490 102.460 18.560 102.630 ;
        RECT 17.490 102.245 17.820 102.460 ;
        RECT 16.660 101.580 17.320 101.910 ;
        RECT 17.530 101.705 17.830 102.035 ;
        RECT 17.530 101.375 17.700 101.705 ;
        RECT 18.000 101.535 18.170 102.460 ;
        RECT 18.730 102.290 19.040 102.510 ;
        RECT 16.320 101.205 17.700 101.375 ;
        RECT 17.895 101.205 18.170 101.535 ;
        RECT 18.340 102.120 19.040 102.290 ;
        RECT 19.210 102.430 19.380 102.680 ;
        RECT 19.790 102.600 20.120 103.575 ;
        RECT 20.350 102.810 20.600 103.310 ;
        RECT 20.780 102.980 21.095 103.575 ;
        RECT 20.350 102.640 21.105 102.810 ;
        RECT 20.435 102.430 20.765 102.470 ;
        RECT 19.210 102.260 20.765 102.430 ;
        RECT 16.320 101.035 16.680 101.205 ;
        RECT 18.340 101.035 18.510 102.120 ;
        RECT 19.210 101.950 19.380 102.260 ;
        RECT 20.435 102.140 20.765 102.260 ;
        RECT 20.935 102.310 21.105 102.640 ;
        RECT 21.275 102.530 21.635 103.310 ;
        RECT 22.305 102.990 23.035 103.405 ;
        RECT 14.575 100.865 15.810 101.035 ;
        RECT 16.850 100.865 18.510 101.035 ;
        RECT 18.680 101.780 19.380 101.950 ;
        RECT 19.610 101.970 19.940 102.090 ;
        RECT 20.935 101.970 21.295 102.310 ;
        RECT 19.610 101.800 21.295 101.970 ;
        RECT 18.680 100.925 18.850 101.780 ;
        RECT 14.575 100.680 14.905 100.865 ;
        RECT 15.640 100.695 17.020 100.865 ;
        RECT 18.340 100.755 18.510 100.865 ;
        RECT 19.070 100.755 19.400 101.610 ;
        RECT 19.610 101.420 19.940 101.800 ;
        RECT 15.135 100.415 15.470 100.695 ;
        RECT 17.360 100.415 17.690 100.695 ;
        RECT 18.340 100.585 19.400 100.755 ;
        RECT 19.760 100.415 20.090 101.140 ;
        RECT 20.320 100.960 20.570 101.800 ;
        RECT 21.465 101.630 21.635 102.530 ;
        RECT 22.460 101.810 22.790 102.820 ;
        RECT 23.540 102.650 23.870 103.575 ;
        RECT 24.040 102.480 24.515 103.190 ;
        RECT 24.715 102.700 24.965 103.310 ;
        RECT 25.145 102.870 25.395 103.575 ;
        RECT 25.565 103.235 26.415 103.405 ;
        RECT 25.565 102.700 25.735 103.235 ;
        RECT 24.715 102.530 25.735 102.700 ;
        RECT 23.275 101.980 23.605 102.480 ;
        RECT 23.780 101.980 24.175 102.310 ;
        RECT 23.780 101.810 23.950 101.980 ;
        RECT 24.345 101.810 24.515 102.480 ;
        RECT 24.725 101.880 25.105 102.360 ;
        RECT 25.275 102.110 25.735 102.530 ;
        RECT 25.905 102.310 26.075 103.065 ;
        RECT 26.245 102.930 26.415 103.235 ;
        RECT 26.585 103.100 26.915 103.575 ;
        RECT 27.085 103.215 28.360 103.385 ;
        RECT 27.085 102.930 27.255 103.215 ;
        RECT 26.245 102.760 27.255 102.930 ;
        RECT 22.460 101.640 23.950 101.810 ;
        RECT 20.770 100.415 21.100 101.630 ;
        RECT 21.275 100.680 21.635 101.630 ;
        RECT 22.550 100.415 22.885 101.470 ;
        RECT 23.055 100.660 23.385 101.640 ;
        RECT 23.590 100.415 23.920 101.470 ;
        RECT 24.120 100.680 24.515 101.810 ;
        RECT 25.275 101.710 25.445 102.110 ;
        RECT 25.905 101.980 26.360 102.310 ;
        RECT 25.905 101.840 26.075 101.980 ;
        RECT 24.715 101.540 25.445 101.710 ;
        RECT 24.715 100.680 25.045 101.540 ;
        RECT 25.245 100.415 25.415 101.370 ;
        RECT 25.615 101.035 26.075 101.840 ;
        RECT 26.570 101.635 26.850 102.535 ;
        RECT 26.470 101.305 26.850 101.635 ;
        RECT 27.020 102.420 27.575 102.590 ;
        RECT 27.020 101.035 27.190 102.420 ;
        RECT 27.755 102.250 28.020 103.045 ;
        RECT 27.360 102.080 28.020 102.250 ;
        RECT 28.190 102.970 28.360 103.215 ;
        RECT 28.670 103.140 28.920 103.575 ;
        RECT 29.090 103.235 30.495 103.405 ;
        RECT 29.090 102.970 29.260 103.235 ;
        RECT 30.165 103.150 30.495 103.235 ;
        RECT 28.190 102.800 29.260 102.970 ;
        RECT 27.360 101.375 27.530 102.080 ;
        RECT 28.190 101.910 28.360 102.800 ;
        RECT 29.430 102.630 29.600 103.065 ;
        RECT 29.820 102.680 30.420 102.930 ;
        RECT 28.530 102.460 29.600 102.630 ;
        RECT 28.530 102.245 28.860 102.460 ;
        RECT 27.700 101.580 28.360 101.910 ;
        RECT 28.570 101.705 28.870 102.035 ;
        RECT 28.570 101.375 28.740 101.705 ;
        RECT 29.040 101.535 29.210 102.460 ;
        RECT 29.770 102.290 30.080 102.510 ;
        RECT 27.360 101.205 28.740 101.375 ;
        RECT 28.935 101.205 29.210 101.535 ;
        RECT 29.380 102.120 30.080 102.290 ;
        RECT 30.250 102.430 30.420 102.680 ;
        RECT 30.830 102.600 31.160 103.575 ;
        RECT 31.390 102.810 31.640 103.310 ;
        RECT 31.820 102.980 32.135 103.575 ;
        RECT 31.390 102.640 32.145 102.810 ;
        RECT 31.475 102.430 31.805 102.470 ;
        RECT 30.250 102.260 31.805 102.430 ;
        RECT 27.360 101.035 27.720 101.205 ;
        RECT 29.380 101.035 29.550 102.120 ;
        RECT 30.250 101.950 30.420 102.260 ;
        RECT 31.475 102.140 31.805 102.260 ;
        RECT 31.975 102.310 32.145 102.640 ;
        RECT 32.315 102.530 32.675 103.310 ;
        RECT 25.615 100.865 26.850 101.035 ;
        RECT 27.890 100.865 29.550 101.035 ;
        RECT 29.720 101.780 30.420 101.950 ;
        RECT 30.650 101.970 30.980 102.090 ;
        RECT 31.975 101.970 32.335 102.310 ;
        RECT 30.650 101.800 32.335 101.970 ;
        RECT 29.720 100.925 29.890 101.780 ;
        RECT 25.615 100.680 25.945 100.865 ;
        RECT 26.680 100.695 28.060 100.865 ;
        RECT 29.380 100.755 29.550 100.865 ;
        RECT 30.110 100.755 30.440 101.610 ;
        RECT 30.650 101.420 30.980 101.800 ;
        RECT 26.175 100.415 26.510 100.695 ;
        RECT 28.400 100.415 28.730 100.695 ;
        RECT 29.380 100.585 30.440 100.755 ;
        RECT 30.800 100.415 31.130 101.140 ;
        RECT 31.360 100.960 31.610 101.800 ;
        RECT 32.505 101.630 32.675 102.530 ;
        RECT 32.930 102.075 33.500 103.575 ;
        RECT 34.210 102.855 34.540 103.575 ;
        RECT 36.210 102.555 36.510 103.575 ;
        RECT 31.810 100.415 32.140 101.630 ;
        RECT 32.315 100.680 32.675 101.630 ;
        RECT 32.855 100.415 33.185 101.730 ;
        RECT 33.905 100.415 34.475 102.410 ;
        RECT 40.610 102.075 41.180 103.575 ;
        RECT 41.890 102.855 42.220 103.575 ;
        RECT 43.450 103.000 43.780 103.290 ;
        RECT 43.450 102.830 44.175 103.000 ;
        RECT 44.350 102.830 44.600 103.575 ;
        RECT 36.210 100.415 36.510 101.455 ;
        RECT 40.535 100.415 40.865 101.730 ;
        RECT 41.585 100.415 42.155 102.410 ;
        RECT 43.445 101.490 43.835 102.660 ;
        RECT 44.005 101.350 44.175 102.830 ;
        RECT 44.775 102.690 45.160 103.310 ;
        RECT 45.330 102.860 45.660 103.575 ;
        RECT 45.830 103.160 47.755 103.330 ;
        RECT 48.235 103.265 48.630 103.575 ;
        RECT 45.830 102.860 46.355 103.160 ;
        RECT 47.585 103.095 47.755 103.160 ;
        RECT 48.800 103.235 50.740 103.405 ;
        RECT 48.800 103.095 48.970 103.235 ;
        RECT 44.345 101.520 44.605 102.530 ;
        RECT 44.775 102.520 46.015 102.690 ;
        RECT 44.775 101.850 44.945 102.520 ;
        RECT 45.115 102.020 45.595 102.350 ;
        RECT 45.765 102.110 46.015 102.520 ;
        RECT 45.365 101.880 45.595 102.020 ;
        RECT 46.185 102.100 46.355 102.860 ;
        RECT 46.525 102.440 46.775 102.990 ;
        RECT 46.945 102.610 47.415 102.990 ;
        RECT 47.585 102.925 48.970 103.095 ;
        RECT 49.140 102.755 49.470 102.995 ;
        RECT 46.525 102.270 47.075 102.440 ;
        RECT 46.185 101.940 46.735 102.100 ;
        RECT 44.775 101.520 45.185 101.850 ;
        RECT 45.835 101.770 46.735 101.940 ;
        RECT 45.835 101.490 46.085 101.770 ;
        RECT 46.905 101.600 47.075 102.270 ;
        RECT 46.330 101.430 47.075 101.600 ;
        RECT 44.005 101.320 44.995 101.350 ;
        RECT 46.330 101.320 46.580 101.430 ;
        RECT 44.005 101.180 46.580 101.320 ;
        RECT 47.245 101.260 47.415 102.610 ;
        RECT 47.585 102.585 49.470 102.755 ;
        RECT 47.585 101.535 47.765 102.585 ;
        RECT 49.140 102.530 49.470 102.585 ;
        RECT 47.935 102.085 48.970 102.415 ;
        RECT 47.935 101.340 48.105 102.085 ;
        RECT 48.275 101.510 48.605 101.865 ;
        RECT 47.935 101.260 48.570 101.340 ;
        RECT 44.005 101.140 44.205 101.180 ;
        RECT 44.825 101.150 46.580 101.180 ;
        RECT 43.425 100.415 43.675 101.140 ;
        RECT 43.875 100.680 44.205 101.140 ;
        RECT 44.405 100.415 44.655 101.010 ;
        RECT 45.305 100.415 45.635 100.980 ;
        RECT 46.330 100.935 46.580 101.150 ;
        RECT 46.780 101.090 48.570 101.260 ;
        RECT 46.780 100.935 47.110 101.090 ;
        RECT 47.705 100.415 48.035 100.920 ;
        RECT 48.800 100.415 49.130 101.915 ;
        RECT 49.300 101.795 49.470 102.530 ;
        RECT 49.640 102.815 50.400 103.065 ;
        RECT 49.640 102.145 49.810 102.815 ;
        RECT 50.570 102.645 50.740 103.235 ;
        RECT 51.065 102.815 51.395 103.575 ;
        RECT 51.935 102.645 52.265 103.275 ;
        RECT 52.495 102.815 52.745 103.575 ;
        RECT 50.010 102.315 50.740 102.645 ;
        RECT 50.910 102.475 52.510 102.645 ;
        RECT 50.910 102.315 51.240 102.475 ;
        RECT 49.640 101.975 49.970 102.145 ;
        RECT 49.300 100.905 49.630 101.795 ;
        RECT 49.800 101.185 49.970 101.975 ;
        RECT 50.285 101.355 50.615 102.315 ;
        RECT 51.840 102.145 52.170 102.305 ;
        RECT 50.785 101.975 52.170 102.145 ;
        RECT 50.785 101.185 50.955 101.975 ;
        RECT 52.340 101.805 52.510 102.475 ;
        RECT 52.925 102.275 53.255 103.310 ;
        RECT 51.125 101.405 51.665 101.740 ;
        RECT 51.835 101.635 52.510 101.805 ;
        RECT 52.705 101.945 53.255 102.275 ;
        RECT 53.485 102.530 53.815 103.310 ;
        RECT 53.995 102.530 54.245 103.575 ;
        RECT 59.245 102.850 59.620 103.180 ;
        RECT 59.790 102.850 60.120 103.575 ;
        RECT 51.835 101.215 52.005 101.635 ;
        RECT 49.800 100.855 50.955 101.185 ;
        RECT 51.125 100.415 51.455 101.215 ;
        RECT 51.640 100.755 52.005 101.215 ;
        RECT 52.175 100.415 52.505 101.465 ;
        RECT 52.705 100.755 52.875 101.945 ;
        RECT 53.485 101.775 53.745 102.530 ;
        RECT 59.245 102.080 59.415 102.850 ;
        RECT 60.290 102.680 60.620 103.310 ;
        RECT 60.800 102.850 60.970 103.575 ;
        RECT 61.150 102.680 61.480 103.310 ;
        RECT 61.660 102.850 61.910 103.575 ;
        RECT 59.585 102.250 59.985 102.580 ;
        RECT 60.290 102.510 61.505 102.680 ;
        RECT 62.130 102.555 62.430 103.575 ;
        RECT 60.155 102.080 61.165 102.310 ;
        RECT 59.245 101.910 61.165 102.080 ;
        RECT 53.045 100.680 53.745 101.775 ;
        RECT 53.915 100.415 54.245 101.840 ;
        RECT 59.245 100.680 59.625 101.910 ;
        RECT 61.335 101.740 61.505 102.510 ;
        RECT 63.090 102.530 63.445 103.310 ;
        RECT 63.615 102.720 63.945 103.575 ;
        RECT 64.125 102.550 64.805 102.860 ;
        RECT 63.090 101.840 63.260 102.530 ;
        RECT 63.620 102.380 64.805 102.550 ;
        RECT 65.005 102.850 65.380 103.180 ;
        RECT 65.550 102.850 65.880 103.575 ;
        RECT 63.620 102.360 63.790 102.380 ;
        RECT 63.430 102.030 63.790 102.360 ;
        RECT 59.795 100.415 60.045 101.740 ;
        RECT 60.245 101.570 61.505 101.740 ;
        RECT 60.245 100.680 60.575 101.570 ;
        RECT 60.775 100.415 61.025 101.400 ;
        RECT 61.225 100.680 61.505 101.570 ;
        RECT 61.675 100.415 61.925 101.840 ;
        RECT 62.130 100.415 62.430 101.455 ;
        RECT 63.090 100.680 63.450 101.840 ;
        RECT 63.620 101.710 63.790 102.030 ;
        RECT 64.010 101.880 64.795 102.210 ;
        RECT 65.005 102.080 65.175 102.850 ;
        RECT 66.050 102.680 66.380 103.310 ;
        RECT 66.560 102.850 66.730 103.575 ;
        RECT 66.910 102.680 67.240 103.310 ;
        RECT 67.420 102.850 67.670 103.575 ;
        RECT 67.940 102.855 68.270 103.575 ;
        RECT 65.345 102.250 65.745 102.580 ;
        RECT 66.050 102.510 67.265 102.680 ;
        RECT 65.915 102.080 66.925 102.310 ;
        RECT 65.005 101.910 66.925 102.080 ;
        RECT 63.620 101.540 64.450 101.710 ;
        RECT 63.620 100.415 63.950 101.370 ;
        RECT 64.120 100.680 64.450 101.540 ;
        RECT 65.005 100.680 65.385 101.910 ;
        RECT 67.095 101.740 67.265 102.510 ;
        RECT 65.555 100.415 65.805 101.740 ;
        RECT 66.005 101.570 67.265 101.740 ;
        RECT 66.005 100.680 66.335 101.570 ;
        RECT 66.535 100.415 66.785 101.400 ;
        RECT 66.985 100.680 67.265 101.570 ;
        RECT 67.435 100.415 67.685 101.840 ;
        RECT 68.005 100.415 68.575 102.410 ;
        RECT 68.980 102.075 69.550 103.575 ;
        RECT 233.850 103.400 234.350 103.900 ;
        RECT 69.295 100.415 69.625 101.730 ;
        RECT 10.200 100.245 69.720 100.415 ;
        RECT 10.295 98.930 10.625 100.245 ;
        RECT 10.370 97.085 10.940 98.585 ;
        RECT 11.345 98.250 11.915 100.245 ;
        RECT 12.215 98.930 12.545 100.245 ;
        RECT 11.650 97.085 11.980 97.805 ;
        RECT 12.290 97.085 12.860 98.585 ;
        RECT 13.265 98.250 13.835 100.245 ;
        RECT 15.595 98.820 16.055 99.980 ;
        RECT 16.225 99.290 16.555 100.245 ;
        RECT 16.725 99.120 17.055 99.980 ;
        RECT 16.225 98.950 17.055 99.120 ;
        RECT 18.955 99.230 19.285 99.700 ;
        RECT 19.490 99.400 19.820 100.245 ;
        RECT 19.990 99.905 21.965 100.075 ;
        RECT 19.990 99.230 20.160 99.905 ;
        RECT 18.955 99.060 20.160 99.230 ;
        RECT 18.955 98.950 19.285 99.060 ;
        RECT 13.570 97.085 13.900 97.805 ;
        RECT 15.595 97.790 15.835 98.820 ;
        RECT 16.225 98.630 16.395 98.950 ;
        RECT 16.005 98.130 16.395 98.630 ;
        RECT 16.565 98.300 17.275 98.780 ;
        RECT 18.955 98.130 19.125 98.950 ;
        RECT 20.905 98.890 21.235 99.735 ;
        RECT 19.345 98.350 19.675 98.780 ;
        RECT 19.845 98.720 21.235 98.890 ;
        RECT 16.005 97.960 17.285 98.130 ;
        RECT 15.595 97.350 15.925 97.790 ;
        RECT 16.095 97.085 16.785 97.680 ;
        RECT 16.955 97.350 17.285 97.960 ;
        RECT 18.955 97.540 19.285 98.130 ;
        RECT 19.465 97.680 19.675 98.130 ;
        RECT 19.845 98.020 20.015 98.720 ;
        RECT 21.795 98.650 21.965 99.905 ;
        RECT 22.135 98.820 22.465 100.245 ;
        RECT 22.635 98.820 23.075 99.980 ;
        RECT 23.250 99.205 23.550 100.245 ;
        RECT 23.735 98.930 24.065 100.245 ;
        RECT 20.185 98.220 20.525 98.550 ;
        RECT 19.845 97.850 20.185 98.020 ;
        RECT 19.465 97.085 19.845 97.680 ;
        RECT 20.015 97.640 20.185 97.850 ;
        RECT 20.355 97.980 20.525 98.220 ;
        RECT 20.725 98.180 21.115 98.550 ;
        RECT 21.295 97.980 21.625 98.550 ;
        RECT 21.795 98.320 22.195 98.650 ;
        RECT 22.365 98.300 22.735 98.630 ;
        RECT 22.365 98.150 22.535 98.300 ;
        RECT 20.355 97.810 21.625 97.980 ;
        RECT 21.795 97.980 22.535 98.150 ;
        RECT 22.905 98.130 23.075 98.820 ;
        RECT 21.795 97.640 21.965 97.980 ;
        RECT 20.015 97.390 21.965 97.640 ;
        RECT 22.135 97.085 22.465 97.810 ;
        RECT 22.705 97.350 23.075 98.130 ;
        RECT 23.250 97.085 23.550 98.105 ;
        RECT 23.810 97.085 24.380 98.585 ;
        RECT 24.785 98.250 25.355 100.245 ;
        RECT 25.675 98.820 26.135 99.980 ;
        RECT 26.305 99.290 26.635 100.245 ;
        RECT 26.805 99.120 27.135 99.980 ;
        RECT 26.305 98.950 27.135 99.120 ;
        RECT 25.090 97.085 25.420 97.805 ;
        RECT 25.675 97.790 25.915 98.820 ;
        RECT 26.305 98.630 26.475 98.950 ;
        RECT 27.565 98.820 27.955 99.980 ;
        RECT 28.125 99.460 28.455 99.980 ;
        RECT 28.625 99.650 29.065 100.245 ;
        RECT 29.235 99.460 29.565 99.980 ;
        RECT 28.125 99.290 29.565 99.460 ;
        RECT 29.795 99.120 30.375 99.980 ;
        RECT 28.125 98.950 30.375 99.120 ;
        RECT 26.085 98.130 26.475 98.630 ;
        RECT 26.645 98.300 27.355 98.780 ;
        RECT 27.565 98.150 27.735 98.820 ;
        RECT 28.125 98.650 28.295 98.950 ;
        RECT 27.905 98.320 28.295 98.650 ;
        RECT 28.475 98.695 28.805 98.780 ;
        RECT 28.475 98.365 30.035 98.695 ;
        RECT 28.475 98.350 28.805 98.365 ;
        RECT 26.085 97.960 27.365 98.130 ;
        RECT 27.565 97.980 28.795 98.150 ;
        RECT 25.675 97.350 26.005 97.790 ;
        RECT 26.175 97.085 26.865 97.680 ;
        RECT 27.035 97.350 27.365 97.960 ;
        RECT 27.780 97.085 28.110 97.745 ;
        RECT 28.350 97.415 28.795 97.980 ;
        RECT 29.170 97.085 29.500 98.195 ;
        RECT 30.205 98.040 30.375 98.950 ;
        RECT 30.665 98.940 30.995 100.245 ;
        RECT 31.915 98.820 32.245 100.245 ;
        RECT 32.415 98.885 33.115 99.980 ;
        RECT 30.545 98.180 31.215 98.615 ;
        RECT 32.415 98.130 32.675 98.885 ;
        RECT 33.285 98.715 33.455 99.905 ;
        RECT 33.655 99.195 33.985 100.245 ;
        RECT 34.155 99.445 34.520 99.905 ;
        RECT 34.705 99.445 35.035 100.245 ;
        RECT 35.205 99.475 36.360 99.805 ;
        RECT 34.155 99.025 34.325 99.445 ;
        RECT 29.680 97.710 30.375 98.040 ;
        RECT 30.545 97.085 31.145 97.990 ;
        RECT 31.915 97.085 32.165 98.130 ;
        RECT 32.345 97.350 32.675 98.130 ;
        RECT 32.905 98.385 33.455 98.715 ;
        RECT 33.650 98.855 34.325 99.025 ;
        RECT 34.495 98.920 35.035 99.255 ;
        RECT 32.905 97.350 33.235 98.385 ;
        RECT 33.650 98.185 33.820 98.855 ;
        RECT 35.205 98.685 35.375 99.475 ;
        RECT 33.990 98.515 35.375 98.685 ;
        RECT 33.990 98.355 34.320 98.515 ;
        RECT 35.545 98.345 35.875 99.305 ;
        RECT 36.190 98.685 36.360 99.475 ;
        RECT 36.530 98.865 36.860 99.755 ;
        RECT 36.190 98.515 36.520 98.685 ;
        RECT 34.920 98.185 35.250 98.345 ;
        RECT 33.650 98.015 35.250 98.185 ;
        RECT 35.420 98.015 36.150 98.345 ;
        RECT 33.415 97.085 33.665 97.845 ;
        RECT 33.895 97.385 34.225 98.015 ;
        RECT 34.765 97.085 35.095 97.845 ;
        RECT 35.420 97.425 35.590 98.015 ;
        RECT 36.350 97.845 36.520 98.515 ;
        RECT 35.760 97.595 36.520 97.845 ;
        RECT 36.690 98.130 36.860 98.865 ;
        RECT 37.030 98.745 37.360 100.245 ;
        RECT 38.125 99.740 38.455 100.245 ;
        RECT 39.050 99.570 39.380 99.725 ;
        RECT 37.590 99.400 39.380 99.570 ;
        RECT 39.580 99.510 39.830 99.725 ;
        RECT 40.525 99.680 40.855 100.245 ;
        RECT 41.505 99.650 41.755 100.245 ;
        RECT 41.955 99.520 42.285 99.980 ;
        RECT 42.485 99.520 42.735 100.245 ;
        RECT 39.580 99.480 41.335 99.510 ;
        RECT 41.955 99.480 42.155 99.520 ;
        RECT 37.590 99.320 38.225 99.400 ;
        RECT 37.555 98.795 37.885 99.150 ;
        RECT 38.055 98.575 38.225 99.320 ;
        RECT 37.190 98.245 38.225 98.575 ;
        RECT 36.690 98.075 37.020 98.130 ;
        RECT 38.395 98.075 38.575 99.125 ;
        RECT 36.690 97.905 38.575 98.075 ;
        RECT 38.745 98.050 38.915 99.400 ;
        RECT 39.580 99.340 42.155 99.480 ;
        RECT 39.580 99.230 39.830 99.340 ;
        RECT 41.165 99.310 42.155 99.340 ;
        RECT 39.085 99.060 39.830 99.230 ;
        RECT 39.085 98.390 39.255 99.060 ;
        RECT 40.075 98.890 40.325 99.170 ;
        RECT 39.425 98.720 40.325 98.890 ;
        RECT 40.975 98.810 41.385 99.140 ;
        RECT 39.425 98.560 39.975 98.720 ;
        RECT 39.085 98.220 39.635 98.390 ;
        RECT 36.690 97.665 37.020 97.905 ;
        RECT 37.190 97.565 38.575 97.735 ;
        RECT 38.745 97.670 39.215 98.050 ;
        RECT 39.385 97.670 39.635 98.220 ;
        RECT 39.805 97.800 39.975 98.560 ;
        RECT 40.565 98.640 40.795 98.780 ;
        RECT 40.145 98.140 40.395 98.550 ;
        RECT 40.565 98.310 41.045 98.640 ;
        RECT 41.215 98.140 41.385 98.810 ;
        RECT 40.145 97.970 41.385 98.140 ;
        RECT 41.555 98.130 41.815 99.140 ;
        RECT 37.190 97.425 37.360 97.565 ;
        RECT 35.420 97.255 37.360 97.425 ;
        RECT 38.405 97.500 38.575 97.565 ;
        RECT 39.805 97.500 40.330 97.800 ;
        RECT 37.530 97.085 37.925 97.395 ;
        RECT 38.405 97.330 40.330 97.500 ;
        RECT 40.500 97.085 40.830 97.800 ;
        RECT 41.000 97.350 41.385 97.970 ;
        RECT 41.985 97.830 42.155 99.310 ;
        RECT 42.325 98.000 42.715 99.170 ;
        RECT 46.775 98.930 47.105 100.245 ;
        RECT 41.560 97.085 41.810 97.830 ;
        RECT 41.985 97.660 42.710 97.830 ;
        RECT 42.380 97.370 42.710 97.660 ;
        RECT 46.850 97.085 47.420 98.585 ;
        RECT 47.825 98.250 48.395 100.245 ;
        RECT 49.170 99.205 49.470 100.245 ;
        RECT 50.125 98.750 50.505 99.980 ;
        RECT 50.675 98.920 50.925 100.245 ;
        RECT 51.125 99.090 51.455 99.980 ;
        RECT 51.655 99.260 51.905 100.245 ;
        RECT 52.105 99.090 52.385 99.980 ;
        RECT 51.125 98.920 52.385 99.090 ;
        RECT 50.125 98.580 52.045 98.750 ;
        RECT 48.130 97.085 48.460 97.805 ;
        RECT 49.170 97.085 49.470 98.105 ;
        RECT 50.125 97.810 50.295 98.580 ;
        RECT 50.465 98.080 50.865 98.410 ;
        RECT 51.035 98.350 52.045 98.580 ;
        RECT 52.215 98.150 52.385 98.920 ;
        RECT 52.555 98.820 52.805 100.245 ;
        RECT 51.170 97.980 52.385 98.150 ;
        RECT 53.965 98.750 54.345 99.980 ;
        RECT 54.515 98.920 54.765 100.245 ;
        RECT 54.965 99.090 55.295 99.980 ;
        RECT 55.495 99.260 55.745 100.245 ;
        RECT 55.945 99.090 56.225 99.980 ;
        RECT 54.965 98.920 56.225 99.090 ;
        RECT 53.965 98.580 55.885 98.750 ;
        RECT 50.125 97.480 50.500 97.810 ;
        RECT 50.670 97.085 51.000 97.810 ;
        RECT 51.170 97.350 51.500 97.980 ;
        RECT 51.680 97.085 51.850 97.810 ;
        RECT 52.030 97.350 52.360 97.980 ;
        RECT 53.965 97.810 54.135 98.580 ;
        RECT 54.305 98.080 54.705 98.410 ;
        RECT 54.875 98.350 55.885 98.580 ;
        RECT 56.055 98.150 56.225 98.920 ;
        RECT 56.395 98.820 56.645 100.245 ;
        RECT 56.865 99.520 57.115 100.245 ;
        RECT 57.315 99.520 57.645 99.980 ;
        RECT 57.845 99.650 58.095 100.245 ;
        RECT 58.745 99.680 59.075 100.245 ;
        RECT 61.145 99.740 61.475 100.245 ;
        RECT 57.445 99.480 57.645 99.520 ;
        RECT 59.770 99.510 60.020 99.725 ;
        RECT 58.265 99.480 60.020 99.510 ;
        RECT 57.445 99.340 60.020 99.480 ;
        RECT 60.220 99.570 60.550 99.725 ;
        RECT 60.220 99.400 62.010 99.570 ;
        RECT 57.445 99.310 58.435 99.340 ;
        RECT 55.010 97.980 56.225 98.150 ;
        RECT 56.885 98.000 57.275 99.170 ;
        RECT 52.540 97.085 52.790 97.810 ;
        RECT 53.965 97.480 54.340 97.810 ;
        RECT 54.510 97.085 54.840 97.810 ;
        RECT 55.010 97.350 55.340 97.980 ;
        RECT 55.520 97.085 55.690 97.810 ;
        RECT 55.870 97.350 56.200 97.980 ;
        RECT 57.445 97.830 57.615 99.310 ;
        RECT 59.770 99.230 60.020 99.340 ;
        RECT 57.785 98.130 58.045 99.140 ;
        RECT 58.215 98.810 58.625 99.140 ;
        RECT 59.275 98.890 59.525 99.170 ;
        RECT 59.770 99.060 60.515 99.230 ;
        RECT 58.215 98.140 58.385 98.810 ;
        RECT 58.805 98.640 59.035 98.780 ;
        RECT 59.275 98.720 60.175 98.890 ;
        RECT 58.555 98.310 59.035 98.640 ;
        RECT 59.625 98.560 60.175 98.720 ;
        RECT 59.205 98.140 59.455 98.550 ;
        RECT 58.215 97.970 59.455 98.140 ;
        RECT 56.380 97.085 56.630 97.810 ;
        RECT 56.890 97.660 57.615 97.830 ;
        RECT 56.890 97.370 57.220 97.660 ;
        RECT 57.790 97.085 58.040 97.830 ;
        RECT 58.215 97.350 58.600 97.970 ;
        RECT 59.625 97.800 59.795 98.560 ;
        RECT 60.345 98.390 60.515 99.060 ;
        RECT 58.770 97.085 59.100 97.800 ;
        RECT 59.270 97.500 59.795 97.800 ;
        RECT 59.965 98.220 60.515 98.390 ;
        RECT 59.965 97.670 60.215 98.220 ;
        RECT 60.685 98.050 60.855 99.400 ;
        RECT 61.375 99.320 62.010 99.400 ;
        RECT 60.385 97.670 60.855 98.050 ;
        RECT 61.025 98.075 61.205 99.125 ;
        RECT 61.375 98.575 61.545 99.320 ;
        RECT 61.715 98.795 62.045 99.150 ;
        RECT 62.240 98.745 62.570 100.245 ;
        RECT 62.740 98.865 63.070 99.755 ;
        RECT 63.240 99.475 64.395 99.805 ;
        RECT 61.375 98.245 62.410 98.575 ;
        RECT 62.740 98.130 62.910 98.865 ;
        RECT 63.240 98.685 63.410 99.475 ;
        RECT 62.580 98.075 62.910 98.130 ;
        RECT 61.025 97.905 62.910 98.075 ;
        RECT 61.025 97.565 62.410 97.735 ;
        RECT 62.580 97.665 62.910 97.905 ;
        RECT 63.080 98.515 63.410 98.685 ;
        RECT 63.080 97.845 63.250 98.515 ;
        RECT 63.725 98.345 64.055 99.305 ;
        RECT 64.225 98.685 64.395 99.475 ;
        RECT 64.565 99.445 64.895 100.245 ;
        RECT 65.080 99.445 65.445 99.905 ;
        RECT 64.565 98.920 65.105 99.255 ;
        RECT 65.275 99.025 65.445 99.445 ;
        RECT 65.615 99.195 65.945 100.245 ;
        RECT 65.275 98.855 65.950 99.025 ;
        RECT 64.225 98.515 65.610 98.685 ;
        RECT 65.280 98.355 65.610 98.515 ;
        RECT 63.450 98.015 64.180 98.345 ;
        RECT 64.350 98.185 64.680 98.345 ;
        RECT 65.780 98.185 65.950 98.855 ;
        RECT 66.145 98.715 66.315 99.905 ;
        RECT 66.485 98.885 67.185 99.980 ;
        RECT 66.145 98.385 66.695 98.715 ;
        RECT 64.350 98.015 65.950 98.185 ;
        RECT 63.080 97.595 63.840 97.845 ;
        RECT 61.025 97.500 61.195 97.565 ;
        RECT 59.270 97.330 61.195 97.500 ;
        RECT 62.240 97.425 62.410 97.565 ;
        RECT 64.010 97.425 64.180 98.015 ;
        RECT 61.675 97.085 62.070 97.395 ;
        RECT 62.240 97.255 64.180 97.425 ;
        RECT 64.505 97.085 64.835 97.845 ;
        RECT 65.375 97.385 65.705 98.015 ;
        RECT 65.935 97.085 66.185 97.845 ;
        RECT 66.365 97.350 66.695 98.385 ;
        RECT 66.925 98.130 67.185 98.885 ;
        RECT 67.355 98.820 67.685 100.245 ;
        RECT 68.005 98.250 68.575 100.245 ;
        RECT 69.295 98.930 69.625 100.245 ;
        RECT 66.925 97.350 67.255 98.130 ;
        RECT 67.435 97.085 67.685 98.130 ;
        RECT 67.940 97.085 68.270 97.805 ;
        RECT 68.980 97.085 69.550 98.585 ;
        RECT 10.200 96.915 69.720 97.085 ;
        RECT 10.370 95.415 10.940 96.915 ;
        RECT 11.650 96.195 11.980 96.915 ;
        RECT 10.295 93.755 10.625 95.070 ;
        RECT 11.345 93.755 11.915 95.750 ;
        RECT 23.810 95.415 24.380 96.915 ;
        RECT 25.090 96.195 25.420 96.915 ;
        RECT 27.115 96.210 27.365 96.915 ;
        RECT 27.545 96.210 27.885 96.650 ;
        RECT 23.735 93.755 24.065 95.070 ;
        RECT 24.785 93.755 25.355 95.750 ;
        RECT 27.215 95.370 27.545 96.040 ;
        RECT 27.215 94.680 27.385 95.370 ;
        RECT 27.715 95.180 27.885 96.210 ;
        RECT 28.055 96.190 28.305 96.915 ;
        RECT 28.475 96.190 28.835 96.650 ;
        RECT 27.555 94.850 27.885 95.180 ;
        RECT 28.085 94.850 28.495 95.990 ;
        RECT 28.665 94.680 28.835 96.190 ;
        RECT 29.035 95.890 29.715 96.200 ;
        RECT 29.895 96.060 30.225 96.915 ;
        RECT 29.035 95.720 30.220 95.890 ;
        RECT 30.395 95.870 30.750 96.650 ;
        RECT 30.050 95.700 30.220 95.720 ;
        RECT 29.045 95.220 29.830 95.550 ;
        RECT 30.050 95.370 30.410 95.700 ;
        RECT 30.050 95.050 30.220 95.370 ;
        RECT 30.580 95.180 30.750 95.870 ;
        RECT 27.215 94.510 28.835 94.680 ;
        RECT 27.105 93.755 27.435 94.340 ;
        RECT 28.005 93.755 28.335 94.340 ;
        RECT 28.535 94.020 28.835 94.510 ;
        RECT 29.390 94.880 30.220 95.050 ;
        RECT 29.390 94.020 29.720 94.880 ;
        RECT 29.890 93.755 30.220 94.710 ;
        RECT 30.390 94.020 30.750 95.180 ;
        RECT 30.955 96.210 31.285 96.650 ;
        RECT 31.455 96.320 32.145 96.915 ;
        RECT 30.955 95.180 31.195 96.210 ;
        RECT 32.315 96.040 32.645 96.650 ;
        RECT 31.365 95.870 32.645 96.040 ;
        RECT 32.875 95.990 33.205 96.550 ;
        RECT 33.385 96.160 33.715 96.915 ;
        RECT 31.365 95.370 31.755 95.870 ;
        RECT 32.875 95.820 33.675 95.990 ;
        RECT 33.885 95.820 34.215 96.650 ;
        RECT 34.395 95.870 34.645 96.915 ;
        RECT 36.210 95.895 36.510 96.915 ;
        RECT 38.170 96.340 38.500 96.630 ;
        RECT 38.170 96.170 38.895 96.340 ;
        RECT 39.070 96.170 39.320 96.915 ;
        RECT 30.955 94.020 31.415 95.180 ;
        RECT 31.585 95.050 31.755 95.370 ;
        RECT 31.925 95.220 32.635 95.700 ;
        RECT 32.885 95.220 33.335 95.650 ;
        RECT 31.585 94.880 32.415 95.050 ;
        RECT 31.585 93.755 31.915 94.710 ;
        RECT 32.085 94.020 32.415 94.880 ;
        RECT 32.875 94.680 33.230 95.050 ;
        RECT 33.505 94.680 33.675 95.820 ;
        RECT 33.845 94.850 34.215 95.820 ;
        RECT 34.385 95.370 35.055 95.700 ;
        RECT 34.385 94.680 34.555 95.370 ;
        RECT 32.875 94.510 34.555 94.680 ;
        RECT 32.875 94.120 33.230 94.510 ;
        RECT 33.435 93.755 33.765 94.340 ;
        RECT 34.740 94.265 35.045 95.180 ;
        RECT 38.165 94.830 38.555 96.000 ;
        RECT 34.335 93.755 35.045 94.265 ;
        RECT 36.210 93.755 36.510 94.795 ;
        RECT 38.725 94.690 38.895 96.170 ;
        RECT 39.495 96.030 39.880 96.650 ;
        RECT 40.050 96.200 40.380 96.915 ;
        RECT 40.550 96.500 42.475 96.670 ;
        RECT 42.955 96.605 43.350 96.915 ;
        RECT 40.550 96.200 41.075 96.500 ;
        RECT 42.305 96.435 42.475 96.500 ;
        RECT 43.520 96.575 45.460 96.745 ;
        RECT 43.520 96.435 43.690 96.575 ;
        RECT 39.065 94.860 39.325 95.870 ;
        RECT 39.495 95.860 40.735 96.030 ;
        RECT 39.495 95.190 39.665 95.860 ;
        RECT 39.835 95.360 40.315 95.690 ;
        RECT 40.485 95.450 40.735 95.860 ;
        RECT 40.085 95.220 40.315 95.360 ;
        RECT 40.905 95.440 41.075 96.200 ;
        RECT 41.245 95.780 41.495 96.330 ;
        RECT 41.665 95.950 42.135 96.330 ;
        RECT 42.305 96.265 43.690 96.435 ;
        RECT 43.860 96.095 44.190 96.335 ;
        RECT 41.245 95.610 41.795 95.780 ;
        RECT 40.905 95.280 41.455 95.440 ;
        RECT 39.495 94.860 39.905 95.190 ;
        RECT 40.555 95.110 41.455 95.280 ;
        RECT 40.555 94.830 40.805 95.110 ;
        RECT 41.625 94.940 41.795 95.610 ;
        RECT 41.050 94.770 41.795 94.940 ;
        RECT 38.725 94.660 39.715 94.690 ;
        RECT 41.050 94.660 41.300 94.770 ;
        RECT 38.725 94.520 41.300 94.660 ;
        RECT 41.965 94.600 42.135 95.950 ;
        RECT 42.305 95.925 44.190 96.095 ;
        RECT 42.305 94.875 42.485 95.925 ;
        RECT 43.860 95.870 44.190 95.925 ;
        RECT 42.655 95.425 43.690 95.755 ;
        RECT 42.655 94.680 42.825 95.425 ;
        RECT 42.995 94.850 43.325 95.205 ;
        RECT 42.655 94.600 43.290 94.680 ;
        RECT 38.725 94.480 38.925 94.520 ;
        RECT 39.545 94.490 41.300 94.520 ;
        RECT 38.145 93.755 38.395 94.480 ;
        RECT 38.595 94.020 38.925 94.480 ;
        RECT 39.125 93.755 39.375 94.350 ;
        RECT 40.025 93.755 40.355 94.320 ;
        RECT 41.050 94.275 41.300 94.490 ;
        RECT 41.500 94.430 43.290 94.600 ;
        RECT 41.500 94.275 41.830 94.430 ;
        RECT 42.425 93.755 42.755 94.260 ;
        RECT 43.520 93.755 43.850 95.255 ;
        RECT 44.020 95.135 44.190 95.870 ;
        RECT 44.360 96.155 45.120 96.405 ;
        RECT 44.360 95.485 44.530 96.155 ;
        RECT 45.290 95.985 45.460 96.575 ;
        RECT 45.785 96.155 46.115 96.915 ;
        RECT 46.655 95.985 46.985 96.615 ;
        RECT 47.215 96.155 47.465 96.915 ;
        RECT 44.730 95.655 45.460 95.985 ;
        RECT 45.630 95.815 47.230 95.985 ;
        RECT 45.630 95.655 45.960 95.815 ;
        RECT 44.360 95.315 44.690 95.485 ;
        RECT 44.020 94.245 44.350 95.135 ;
        RECT 44.520 94.525 44.690 95.315 ;
        RECT 45.005 94.695 45.335 95.655 ;
        RECT 46.560 95.485 46.890 95.645 ;
        RECT 45.505 95.315 46.890 95.485 ;
        RECT 45.505 94.525 45.675 95.315 ;
        RECT 47.060 95.145 47.230 95.815 ;
        RECT 47.645 95.615 47.975 96.650 ;
        RECT 45.845 94.745 46.385 95.080 ;
        RECT 46.555 94.975 47.230 95.145 ;
        RECT 47.425 95.285 47.975 95.615 ;
        RECT 48.205 95.870 48.535 96.650 ;
        RECT 48.715 95.870 48.965 96.915 ;
        RECT 49.195 95.870 49.445 96.915 ;
        RECT 49.625 95.870 49.955 96.650 ;
        RECT 46.555 94.555 46.725 94.975 ;
        RECT 44.520 94.195 45.675 94.525 ;
        RECT 45.845 93.755 46.175 94.555 ;
        RECT 46.360 94.095 46.725 94.555 ;
        RECT 46.895 93.755 47.225 94.805 ;
        RECT 47.425 94.095 47.595 95.285 ;
        RECT 48.205 95.115 48.465 95.870 ;
        RECT 47.765 94.020 48.465 95.115 ;
        RECT 48.635 93.755 48.965 95.180 ;
        RECT 49.195 93.755 49.525 95.180 ;
        RECT 49.695 95.115 49.955 95.870 ;
        RECT 50.185 95.615 50.515 96.650 ;
        RECT 50.695 96.155 50.945 96.915 ;
        RECT 51.175 95.985 51.505 96.615 ;
        RECT 52.045 96.155 52.375 96.915 ;
        RECT 52.700 96.575 54.640 96.745 ;
        RECT 54.810 96.605 55.205 96.915 ;
        RECT 52.700 95.985 52.870 96.575 ;
        RECT 54.470 96.435 54.640 96.575 ;
        RECT 55.685 96.500 57.610 96.670 ;
        RECT 55.685 96.435 55.855 96.500 ;
        RECT 53.040 96.155 53.800 96.405 ;
        RECT 50.930 95.815 52.530 95.985 ;
        RECT 50.185 95.285 50.735 95.615 ;
        RECT 49.695 94.020 50.395 95.115 ;
        RECT 50.565 94.095 50.735 95.285 ;
        RECT 50.930 95.145 51.100 95.815 ;
        RECT 52.200 95.655 52.530 95.815 ;
        RECT 52.700 95.655 53.430 95.985 ;
        RECT 51.270 95.485 51.600 95.645 ;
        RECT 51.270 95.315 52.655 95.485 ;
        RECT 50.930 94.975 51.605 95.145 ;
        RECT 50.935 93.755 51.265 94.805 ;
        RECT 51.435 94.555 51.605 94.975 ;
        RECT 51.775 94.745 52.315 95.080 ;
        RECT 51.435 94.095 51.800 94.555 ;
        RECT 51.985 93.755 52.315 94.555 ;
        RECT 52.485 94.525 52.655 95.315 ;
        RECT 52.825 94.695 53.155 95.655 ;
        RECT 53.630 95.485 53.800 96.155 ;
        RECT 53.470 95.315 53.800 95.485 ;
        RECT 53.970 96.095 54.300 96.335 ;
        RECT 54.470 96.265 55.855 96.435 ;
        RECT 53.970 95.925 55.855 96.095 ;
        RECT 53.970 95.870 54.300 95.925 ;
        RECT 53.470 94.525 53.640 95.315 ;
        RECT 53.970 95.135 54.140 95.870 ;
        RECT 54.470 95.425 55.505 95.755 ;
        RECT 52.485 94.195 53.640 94.525 ;
        RECT 53.810 94.245 54.140 95.135 ;
        RECT 54.310 93.755 54.640 95.255 ;
        RECT 54.835 94.850 55.165 95.205 ;
        RECT 55.335 94.680 55.505 95.425 ;
        RECT 55.675 94.875 55.855 95.925 ;
        RECT 56.025 95.950 56.495 96.330 ;
        RECT 54.870 94.600 55.505 94.680 ;
        RECT 56.025 94.600 56.195 95.950 ;
        RECT 56.665 95.780 56.915 96.330 ;
        RECT 56.365 95.610 56.915 95.780 ;
        RECT 57.085 96.200 57.610 96.500 ;
        RECT 57.780 96.200 58.110 96.915 ;
        RECT 56.365 94.940 56.535 95.610 ;
        RECT 57.085 95.440 57.255 96.200 ;
        RECT 58.280 96.030 58.665 96.650 ;
        RECT 58.840 96.170 59.090 96.915 ;
        RECT 59.660 96.340 59.990 96.630 ;
        RECT 59.265 96.170 59.990 96.340 ;
        RECT 57.425 95.860 58.665 96.030 ;
        RECT 57.425 95.450 57.675 95.860 ;
        RECT 56.705 95.280 57.255 95.440 ;
        RECT 57.845 95.360 58.325 95.690 ;
        RECT 56.705 95.110 57.605 95.280 ;
        RECT 57.845 95.220 58.075 95.360 ;
        RECT 58.495 95.190 58.665 95.860 ;
        RECT 56.365 94.770 57.110 94.940 ;
        RECT 57.355 94.830 57.605 95.110 ;
        RECT 58.255 94.860 58.665 95.190 ;
        RECT 58.835 94.860 59.095 95.870 ;
        RECT 56.860 94.660 57.110 94.770 ;
        RECT 59.265 94.690 59.435 96.170 ;
        RECT 59.605 94.830 59.995 96.000 ;
        RECT 60.290 95.415 60.860 96.915 ;
        RECT 61.570 96.195 61.900 96.915 ;
        RECT 62.130 95.895 62.430 96.915 ;
        RECT 58.445 94.660 59.435 94.690 ;
        RECT 54.870 94.430 56.660 94.600 ;
        RECT 56.330 94.275 56.660 94.430 ;
        RECT 56.860 94.520 59.435 94.660 ;
        RECT 56.860 94.490 58.615 94.520 ;
        RECT 56.860 94.275 57.110 94.490 ;
        RECT 59.235 94.480 59.435 94.520 ;
        RECT 55.405 93.755 55.735 94.260 ;
        RECT 57.805 93.755 58.135 94.320 ;
        RECT 58.785 93.755 59.035 94.350 ;
        RECT 59.235 94.020 59.565 94.480 ;
        RECT 59.765 93.755 60.015 94.480 ;
        RECT 60.215 93.755 60.545 95.070 ;
        RECT 61.265 93.755 61.835 95.750 ;
        RECT 62.690 95.415 63.260 96.915 ;
        RECT 63.970 96.195 64.300 96.915 ;
        RECT 65.005 96.190 65.380 96.520 ;
        RECT 65.550 96.190 65.880 96.915 ;
        RECT 62.130 93.755 62.430 94.795 ;
        RECT 62.615 93.755 62.945 95.070 ;
        RECT 63.665 93.755 64.235 95.750 ;
        RECT 65.005 95.420 65.175 96.190 ;
        RECT 66.050 96.020 66.380 96.650 ;
        RECT 66.560 96.190 66.730 96.915 ;
        RECT 66.910 96.020 67.240 96.650 ;
        RECT 67.420 96.190 67.670 96.915 ;
        RECT 67.940 96.195 68.270 96.915 ;
        RECT 65.345 95.590 65.745 95.920 ;
        RECT 66.050 95.850 67.265 96.020 ;
        RECT 65.915 95.420 66.925 95.650 ;
        RECT 65.005 95.250 66.925 95.420 ;
        RECT 65.005 94.020 65.385 95.250 ;
        RECT 67.095 95.080 67.265 95.850 ;
        RECT 65.555 93.755 65.805 95.080 ;
        RECT 66.005 94.910 67.265 95.080 ;
        RECT 66.005 94.020 66.335 94.910 ;
        RECT 66.535 93.755 66.785 94.740 ;
        RECT 66.985 94.020 67.265 94.910 ;
        RECT 67.435 93.755 67.685 95.180 ;
        RECT 68.005 93.755 68.575 95.750 ;
        RECT 68.980 95.415 69.550 96.915 ;
        RECT 69.295 93.755 69.625 95.070 ;
        RECT 10.200 93.585 69.720 93.755 ;
        RECT 10.295 92.270 10.625 93.585 ;
        RECT 10.370 90.425 10.940 91.925 ;
        RECT 11.345 91.590 11.915 93.585 ;
        RECT 19.895 92.270 20.225 93.585 ;
        RECT 11.650 90.425 11.980 91.145 ;
        RECT 19.970 90.425 20.540 91.925 ;
        RECT 20.945 91.590 21.515 93.585 ;
        RECT 23.250 92.545 23.550 93.585 ;
        RECT 23.745 93.000 24.075 93.585 ;
        RECT 24.645 93.000 24.975 93.585 ;
        RECT 25.175 92.830 25.475 93.320 ;
        RECT 23.855 92.660 25.475 92.830 ;
        RECT 23.855 91.970 24.025 92.660 ;
        RECT 24.195 92.160 24.525 92.490 ;
        RECT 21.250 90.425 21.580 91.145 ;
        RECT 23.250 90.425 23.550 91.445 ;
        RECT 23.855 91.300 24.185 91.970 ;
        RECT 24.355 91.130 24.525 92.160 ;
        RECT 24.725 91.350 25.135 92.490 ;
        RECT 25.305 91.150 25.475 92.660 ;
        RECT 25.675 92.160 26.005 93.585 ;
        RECT 26.175 92.225 26.875 93.320 ;
        RECT 26.175 91.470 26.435 92.225 ;
        RECT 27.045 92.055 27.215 93.245 ;
        RECT 27.415 92.535 27.745 93.585 ;
        RECT 27.915 92.785 28.280 93.245 ;
        RECT 28.465 92.785 28.795 93.585 ;
        RECT 28.965 92.815 30.120 93.145 ;
        RECT 27.915 92.365 28.085 92.785 ;
        RECT 23.755 90.425 24.005 91.130 ;
        RECT 24.185 90.690 24.525 91.130 ;
        RECT 24.695 90.425 24.945 91.150 ;
        RECT 25.115 90.690 25.475 91.150 ;
        RECT 25.675 90.425 25.925 91.470 ;
        RECT 26.105 90.690 26.435 91.470 ;
        RECT 26.665 91.725 27.215 92.055 ;
        RECT 27.410 92.195 28.085 92.365 ;
        RECT 28.255 92.260 28.795 92.595 ;
        RECT 26.665 90.690 26.995 91.725 ;
        RECT 27.410 91.525 27.580 92.195 ;
        RECT 28.965 92.025 29.135 92.815 ;
        RECT 27.750 91.855 29.135 92.025 ;
        RECT 27.750 91.695 28.080 91.855 ;
        RECT 29.305 91.685 29.635 92.645 ;
        RECT 29.950 92.025 30.120 92.815 ;
        RECT 30.290 92.205 30.620 93.095 ;
        RECT 29.950 91.855 30.280 92.025 ;
        RECT 28.680 91.525 29.010 91.685 ;
        RECT 27.410 91.355 29.010 91.525 ;
        RECT 29.180 91.355 29.910 91.685 ;
        RECT 27.175 90.425 27.425 91.185 ;
        RECT 27.655 90.725 27.985 91.355 ;
        RECT 28.525 90.425 28.855 91.185 ;
        RECT 29.180 90.765 29.350 91.355 ;
        RECT 30.110 91.185 30.280 91.855 ;
        RECT 29.520 90.935 30.280 91.185 ;
        RECT 30.450 91.470 30.620 92.205 ;
        RECT 30.790 92.085 31.120 93.585 ;
        RECT 31.885 93.080 32.215 93.585 ;
        RECT 32.810 92.910 33.140 93.065 ;
        RECT 31.350 92.740 33.140 92.910 ;
        RECT 33.340 92.850 33.590 93.065 ;
        RECT 34.285 93.020 34.615 93.585 ;
        RECT 35.265 92.990 35.515 93.585 ;
        RECT 35.715 92.860 36.045 93.320 ;
        RECT 36.245 92.860 36.495 93.585 ;
        RECT 33.340 92.820 35.095 92.850 ;
        RECT 35.715 92.820 35.915 92.860 ;
        RECT 31.350 92.660 31.985 92.740 ;
        RECT 31.315 92.135 31.645 92.490 ;
        RECT 31.815 91.915 31.985 92.660 ;
        RECT 30.950 91.585 31.985 91.915 ;
        RECT 30.450 91.415 30.780 91.470 ;
        RECT 32.155 91.415 32.335 92.465 ;
        RECT 30.450 91.245 32.335 91.415 ;
        RECT 32.505 91.390 32.675 92.740 ;
        RECT 33.340 92.680 35.915 92.820 ;
        RECT 33.340 92.570 33.590 92.680 ;
        RECT 34.925 92.650 35.915 92.680 ;
        RECT 32.845 92.400 33.590 92.570 ;
        RECT 32.845 91.730 33.015 92.400 ;
        RECT 33.835 92.230 34.085 92.510 ;
        RECT 33.185 92.060 34.085 92.230 ;
        RECT 34.735 92.150 35.145 92.480 ;
        RECT 33.185 91.900 33.735 92.060 ;
        RECT 32.845 91.560 33.395 91.730 ;
        RECT 30.450 91.005 30.780 91.245 ;
        RECT 30.950 90.905 32.335 91.075 ;
        RECT 32.505 91.010 32.975 91.390 ;
        RECT 33.145 91.010 33.395 91.560 ;
        RECT 33.565 91.140 33.735 91.900 ;
        RECT 34.325 91.980 34.555 92.120 ;
        RECT 33.905 91.480 34.155 91.890 ;
        RECT 34.325 91.650 34.805 91.980 ;
        RECT 34.975 91.480 35.145 92.150 ;
        RECT 33.905 91.310 35.145 91.480 ;
        RECT 35.315 91.470 35.575 92.480 ;
        RECT 30.950 90.765 31.120 90.905 ;
        RECT 29.180 90.595 31.120 90.765 ;
        RECT 32.165 90.840 32.335 90.905 ;
        RECT 33.565 90.840 34.090 91.140 ;
        RECT 31.290 90.425 31.685 90.735 ;
        RECT 32.165 90.670 34.090 90.840 ;
        RECT 34.260 90.425 34.590 91.140 ;
        RECT 34.760 90.690 35.145 91.310 ;
        RECT 35.745 91.170 35.915 92.650 ;
        RECT 36.085 91.340 36.475 92.510 ;
        RECT 36.715 92.160 37.045 93.585 ;
        RECT 37.215 92.225 37.915 93.320 ;
        RECT 37.215 91.470 37.475 92.225 ;
        RECT 38.085 92.055 38.255 93.245 ;
        RECT 38.455 92.535 38.785 93.585 ;
        RECT 38.955 92.785 39.320 93.245 ;
        RECT 39.505 92.785 39.835 93.585 ;
        RECT 40.005 92.815 41.160 93.145 ;
        RECT 38.955 92.365 39.125 92.785 ;
        RECT 35.320 90.425 35.570 91.170 ;
        RECT 35.745 91.000 36.470 91.170 ;
        RECT 36.140 90.710 36.470 91.000 ;
        RECT 36.715 90.425 36.965 91.470 ;
        RECT 37.145 90.690 37.475 91.470 ;
        RECT 37.705 91.725 38.255 92.055 ;
        RECT 38.450 92.195 39.125 92.365 ;
        RECT 39.295 92.260 39.835 92.595 ;
        RECT 37.705 90.690 38.035 91.725 ;
        RECT 38.450 91.525 38.620 92.195 ;
        RECT 40.005 92.025 40.175 92.815 ;
        RECT 38.790 91.855 40.175 92.025 ;
        RECT 38.790 91.695 39.120 91.855 ;
        RECT 40.345 91.685 40.675 92.645 ;
        RECT 40.990 92.025 41.160 92.815 ;
        RECT 41.330 92.205 41.660 93.095 ;
        RECT 40.990 91.855 41.320 92.025 ;
        RECT 39.720 91.525 40.050 91.685 ;
        RECT 38.450 91.355 40.050 91.525 ;
        RECT 40.220 91.355 40.950 91.685 ;
        RECT 38.215 90.425 38.465 91.185 ;
        RECT 38.695 90.725 39.025 91.355 ;
        RECT 39.565 90.425 39.895 91.185 ;
        RECT 40.220 90.765 40.390 91.355 ;
        RECT 41.150 91.185 41.320 91.855 ;
        RECT 40.560 90.935 41.320 91.185 ;
        RECT 41.490 91.470 41.660 92.205 ;
        RECT 41.830 92.085 42.160 93.585 ;
        RECT 42.925 93.080 43.255 93.585 ;
        RECT 43.850 92.910 44.180 93.065 ;
        RECT 42.390 92.740 44.180 92.910 ;
        RECT 44.380 92.850 44.630 93.065 ;
        RECT 45.325 93.020 45.655 93.585 ;
        RECT 46.305 92.990 46.555 93.585 ;
        RECT 46.755 92.860 47.085 93.320 ;
        RECT 47.285 92.860 47.535 93.585 ;
        RECT 44.380 92.820 46.135 92.850 ;
        RECT 46.755 92.820 46.955 92.860 ;
        RECT 42.390 92.660 43.025 92.740 ;
        RECT 42.355 92.135 42.685 92.490 ;
        RECT 42.855 91.915 43.025 92.660 ;
        RECT 41.990 91.585 43.025 91.915 ;
        RECT 41.490 91.415 41.820 91.470 ;
        RECT 43.195 91.415 43.375 92.465 ;
        RECT 41.490 91.245 43.375 91.415 ;
        RECT 43.545 91.390 43.715 92.740 ;
        RECT 44.380 92.680 46.955 92.820 ;
        RECT 44.380 92.570 44.630 92.680 ;
        RECT 45.965 92.650 46.955 92.680 ;
        RECT 43.885 92.400 44.630 92.570 ;
        RECT 43.885 91.730 44.055 92.400 ;
        RECT 44.875 92.230 45.125 92.510 ;
        RECT 44.225 92.060 45.125 92.230 ;
        RECT 45.775 92.150 46.185 92.480 ;
        RECT 44.225 91.900 44.775 92.060 ;
        RECT 43.885 91.560 44.435 91.730 ;
        RECT 41.490 91.005 41.820 91.245 ;
        RECT 41.990 90.905 43.375 91.075 ;
        RECT 43.545 91.010 44.015 91.390 ;
        RECT 44.185 91.010 44.435 91.560 ;
        RECT 44.605 91.140 44.775 91.900 ;
        RECT 45.365 91.980 45.595 92.120 ;
        RECT 44.945 91.480 45.195 91.890 ;
        RECT 45.365 91.650 45.845 91.980 ;
        RECT 46.015 91.480 46.185 92.150 ;
        RECT 44.945 91.310 46.185 91.480 ;
        RECT 46.355 91.470 46.615 92.480 ;
        RECT 41.990 90.765 42.160 90.905 ;
        RECT 40.220 90.595 42.160 90.765 ;
        RECT 43.205 90.840 43.375 90.905 ;
        RECT 44.605 90.840 45.130 91.140 ;
        RECT 42.330 90.425 42.725 90.735 ;
        RECT 43.205 90.670 45.130 90.840 ;
        RECT 45.300 90.425 45.630 91.140 ;
        RECT 45.800 90.690 46.185 91.310 ;
        RECT 46.785 91.170 46.955 92.650 ;
        RECT 49.170 92.545 49.470 93.585 ;
        RECT 47.125 91.340 47.515 92.510 ;
        RECT 51.085 92.090 51.465 93.320 ;
        RECT 51.635 92.260 51.885 93.585 ;
        RECT 52.085 92.430 52.415 93.320 ;
        RECT 52.615 92.600 52.865 93.585 ;
        RECT 53.065 92.430 53.345 93.320 ;
        RECT 52.085 92.260 53.345 92.430 ;
        RECT 51.085 91.920 53.005 92.090 ;
        RECT 46.360 90.425 46.610 91.170 ;
        RECT 46.785 91.000 47.510 91.170 ;
        RECT 47.180 90.710 47.510 91.000 ;
        RECT 49.170 90.425 49.470 91.445 ;
        RECT 51.085 91.150 51.255 91.920 ;
        RECT 51.425 91.420 51.825 91.750 ;
        RECT 51.995 91.690 53.005 91.920 ;
        RECT 53.175 91.490 53.345 92.260 ;
        RECT 53.515 92.160 53.765 93.585 ;
        RECT 52.130 91.320 53.345 91.490 ;
        RECT 53.965 92.090 54.345 93.320 ;
        RECT 54.515 92.260 54.765 93.585 ;
        RECT 54.965 92.430 55.295 93.320 ;
        RECT 55.495 92.600 55.745 93.585 ;
        RECT 55.945 92.430 56.225 93.320 ;
        RECT 54.965 92.260 56.225 92.430 ;
        RECT 53.965 91.920 55.885 92.090 ;
        RECT 51.085 90.820 51.460 91.150 ;
        RECT 51.630 90.425 51.960 91.150 ;
        RECT 52.130 90.690 52.460 91.320 ;
        RECT 52.640 90.425 52.810 91.150 ;
        RECT 52.990 90.690 53.320 91.320 ;
        RECT 53.965 91.150 54.135 91.920 ;
        RECT 54.305 91.420 54.705 91.750 ;
        RECT 54.875 91.690 55.885 91.920 ;
        RECT 56.055 91.490 56.225 92.260 ;
        RECT 56.395 92.160 56.645 93.585 ;
        RECT 56.865 92.860 57.115 93.585 ;
        RECT 57.315 92.860 57.645 93.320 ;
        RECT 57.845 92.990 58.095 93.585 ;
        RECT 58.745 93.020 59.075 93.585 ;
        RECT 61.145 93.080 61.475 93.585 ;
        RECT 57.445 92.820 57.645 92.860 ;
        RECT 59.770 92.850 60.020 93.065 ;
        RECT 58.265 92.820 60.020 92.850 ;
        RECT 57.445 92.680 60.020 92.820 ;
        RECT 60.220 92.910 60.550 93.065 ;
        RECT 60.220 92.740 62.010 92.910 ;
        RECT 57.445 92.650 58.435 92.680 ;
        RECT 55.010 91.320 56.225 91.490 ;
        RECT 56.885 91.340 57.275 92.510 ;
        RECT 53.500 90.425 53.750 91.150 ;
        RECT 53.965 90.820 54.340 91.150 ;
        RECT 54.510 90.425 54.840 91.150 ;
        RECT 55.010 90.690 55.340 91.320 ;
        RECT 55.520 90.425 55.690 91.150 ;
        RECT 55.870 90.690 56.200 91.320 ;
        RECT 57.445 91.170 57.615 92.650 ;
        RECT 59.770 92.570 60.020 92.680 ;
        RECT 57.785 91.470 58.045 92.480 ;
        RECT 58.215 92.150 58.625 92.480 ;
        RECT 59.275 92.230 59.525 92.510 ;
        RECT 59.770 92.400 60.515 92.570 ;
        RECT 58.215 91.480 58.385 92.150 ;
        RECT 58.805 91.980 59.035 92.120 ;
        RECT 59.275 92.060 60.175 92.230 ;
        RECT 58.555 91.650 59.035 91.980 ;
        RECT 59.625 91.900 60.175 92.060 ;
        RECT 59.205 91.480 59.455 91.890 ;
        RECT 58.215 91.310 59.455 91.480 ;
        RECT 56.380 90.425 56.630 91.150 ;
        RECT 56.890 91.000 57.615 91.170 ;
        RECT 56.890 90.710 57.220 91.000 ;
        RECT 57.790 90.425 58.040 91.170 ;
        RECT 58.215 90.690 58.600 91.310 ;
        RECT 59.625 91.140 59.795 91.900 ;
        RECT 60.345 91.730 60.515 92.400 ;
        RECT 58.770 90.425 59.100 91.140 ;
        RECT 59.270 90.840 59.795 91.140 ;
        RECT 59.965 91.560 60.515 91.730 ;
        RECT 59.965 91.010 60.215 91.560 ;
        RECT 60.685 91.390 60.855 92.740 ;
        RECT 61.375 92.660 62.010 92.740 ;
        RECT 60.385 91.010 60.855 91.390 ;
        RECT 61.025 91.415 61.205 92.465 ;
        RECT 61.375 91.915 61.545 92.660 ;
        RECT 61.715 92.135 62.045 92.490 ;
        RECT 62.240 92.085 62.570 93.585 ;
        RECT 62.740 92.205 63.070 93.095 ;
        RECT 63.240 92.815 64.395 93.145 ;
        RECT 61.375 91.585 62.410 91.915 ;
        RECT 62.740 91.470 62.910 92.205 ;
        RECT 63.240 92.025 63.410 92.815 ;
        RECT 62.580 91.415 62.910 91.470 ;
        RECT 61.025 91.245 62.910 91.415 ;
        RECT 61.025 90.905 62.410 91.075 ;
        RECT 62.580 91.005 62.910 91.245 ;
        RECT 63.080 91.855 63.410 92.025 ;
        RECT 63.080 91.185 63.250 91.855 ;
        RECT 63.725 91.685 64.055 92.645 ;
        RECT 64.225 92.025 64.395 92.815 ;
        RECT 64.565 92.785 64.895 93.585 ;
        RECT 65.080 92.785 65.445 93.245 ;
        RECT 64.565 92.260 65.105 92.595 ;
        RECT 65.275 92.365 65.445 92.785 ;
        RECT 65.615 92.535 65.945 93.585 ;
        RECT 65.275 92.195 65.950 92.365 ;
        RECT 64.225 91.855 65.610 92.025 ;
        RECT 65.280 91.695 65.610 91.855 ;
        RECT 63.450 91.355 64.180 91.685 ;
        RECT 64.350 91.525 64.680 91.685 ;
        RECT 65.780 91.525 65.950 92.195 ;
        RECT 66.145 92.055 66.315 93.245 ;
        RECT 66.485 92.225 67.185 93.320 ;
        RECT 66.145 91.725 66.695 92.055 ;
        RECT 64.350 91.355 65.950 91.525 ;
        RECT 63.080 90.935 63.840 91.185 ;
        RECT 61.025 90.840 61.195 90.905 ;
        RECT 59.270 90.670 61.195 90.840 ;
        RECT 62.240 90.765 62.410 90.905 ;
        RECT 64.010 90.765 64.180 91.355 ;
        RECT 61.675 90.425 62.070 90.735 ;
        RECT 62.240 90.595 64.180 90.765 ;
        RECT 64.505 90.425 64.835 91.185 ;
        RECT 65.375 90.725 65.705 91.355 ;
        RECT 65.935 90.425 66.185 91.185 ;
        RECT 66.365 90.690 66.695 91.725 ;
        RECT 66.925 91.470 67.185 92.225 ;
        RECT 67.355 92.160 67.685 93.585 ;
        RECT 68.005 91.590 68.575 93.585 ;
        RECT 69.295 92.270 69.625 93.585 ;
        RECT 112.980 93.045 115.080 93.215 ;
        RECT 66.925 90.690 67.255 91.470 ;
        RECT 67.435 90.425 67.685 91.470 ;
        RECT 67.940 90.425 68.270 91.145 ;
        RECT 68.980 90.425 69.550 91.925 ;
        RECT 10.200 90.255 69.720 90.425 ;
        RECT 10.370 88.755 10.940 90.255 ;
        RECT 11.650 89.535 11.980 90.255 ;
        RECT 25.210 89.680 25.540 89.970 ;
        RECT 25.210 89.510 25.935 89.680 ;
        RECT 26.110 89.510 26.360 90.255 ;
        RECT 10.295 87.095 10.625 88.410 ;
        RECT 11.345 87.095 11.915 89.090 ;
        RECT 25.205 88.170 25.595 89.340 ;
        RECT 25.765 88.030 25.935 89.510 ;
        RECT 26.535 89.370 26.920 89.990 ;
        RECT 27.090 89.540 27.420 90.255 ;
        RECT 27.590 89.840 29.515 90.010 ;
        RECT 29.995 89.945 30.390 90.255 ;
        RECT 27.590 89.540 28.115 89.840 ;
        RECT 29.345 89.775 29.515 89.840 ;
        RECT 30.560 89.915 32.500 90.085 ;
        RECT 30.560 89.775 30.730 89.915 ;
        RECT 26.105 88.200 26.365 89.210 ;
        RECT 26.535 89.200 27.775 89.370 ;
        RECT 26.535 88.530 26.705 89.200 ;
        RECT 26.875 88.700 27.355 89.030 ;
        RECT 27.525 88.790 27.775 89.200 ;
        RECT 27.125 88.560 27.355 88.700 ;
        RECT 27.945 88.780 28.115 89.540 ;
        RECT 28.285 89.120 28.535 89.670 ;
        RECT 28.705 89.290 29.175 89.670 ;
        RECT 29.345 89.605 30.730 89.775 ;
        RECT 30.900 89.435 31.230 89.675 ;
        RECT 28.285 88.950 28.835 89.120 ;
        RECT 27.945 88.620 28.495 88.780 ;
        RECT 26.535 88.200 26.945 88.530 ;
        RECT 27.595 88.450 28.495 88.620 ;
        RECT 27.595 88.170 27.845 88.450 ;
        RECT 28.665 88.280 28.835 88.950 ;
        RECT 28.090 88.110 28.835 88.280 ;
        RECT 25.765 88.000 26.755 88.030 ;
        RECT 28.090 88.000 28.340 88.110 ;
        RECT 25.765 87.860 28.340 88.000 ;
        RECT 29.005 87.940 29.175 89.290 ;
        RECT 29.345 89.265 31.230 89.435 ;
        RECT 29.345 88.215 29.525 89.265 ;
        RECT 30.900 89.210 31.230 89.265 ;
        RECT 29.695 88.765 30.730 89.095 ;
        RECT 29.695 88.020 29.865 88.765 ;
        RECT 30.035 88.190 30.365 88.545 ;
        RECT 29.695 87.940 30.330 88.020 ;
        RECT 25.765 87.820 25.965 87.860 ;
        RECT 26.585 87.830 28.340 87.860 ;
        RECT 25.185 87.095 25.435 87.820 ;
        RECT 25.635 87.360 25.965 87.820 ;
        RECT 26.165 87.095 26.415 87.690 ;
        RECT 27.065 87.095 27.395 87.660 ;
        RECT 28.090 87.615 28.340 87.830 ;
        RECT 28.540 87.770 30.330 87.940 ;
        RECT 28.540 87.615 28.870 87.770 ;
        RECT 29.465 87.095 29.795 87.600 ;
        RECT 30.560 87.095 30.890 88.595 ;
        RECT 31.060 88.475 31.230 89.210 ;
        RECT 31.400 89.495 32.160 89.745 ;
        RECT 31.400 88.825 31.570 89.495 ;
        RECT 32.330 89.325 32.500 89.915 ;
        RECT 32.825 89.495 33.155 90.255 ;
        RECT 33.695 89.325 34.025 89.955 ;
        RECT 34.255 89.495 34.505 90.255 ;
        RECT 31.770 88.995 32.500 89.325 ;
        RECT 32.670 89.155 34.270 89.325 ;
        RECT 32.670 88.995 33.000 89.155 ;
        RECT 31.400 88.655 31.730 88.825 ;
        RECT 31.060 87.585 31.390 88.475 ;
        RECT 31.560 87.865 31.730 88.655 ;
        RECT 32.045 88.035 32.375 88.995 ;
        RECT 33.600 88.825 33.930 88.985 ;
        RECT 32.545 88.655 33.930 88.825 ;
        RECT 32.545 87.865 32.715 88.655 ;
        RECT 34.100 88.485 34.270 89.155 ;
        RECT 34.685 88.955 35.015 89.990 ;
        RECT 32.885 88.085 33.425 88.420 ;
        RECT 33.595 88.315 34.270 88.485 ;
        RECT 34.465 88.625 35.015 88.955 ;
        RECT 35.245 89.210 35.575 89.990 ;
        RECT 35.755 89.210 36.005 90.255 ;
        RECT 36.210 89.235 36.510 90.255 ;
        RECT 36.690 89.210 37.045 89.990 ;
        RECT 37.215 89.400 37.545 90.255 ;
        RECT 37.725 89.230 38.405 89.540 ;
        RECT 33.595 87.895 33.765 88.315 ;
        RECT 31.560 87.535 32.715 87.865 ;
        RECT 32.885 87.095 33.215 87.895 ;
        RECT 33.400 87.435 33.765 87.895 ;
        RECT 33.935 87.095 34.265 88.145 ;
        RECT 34.465 87.435 34.635 88.625 ;
        RECT 35.245 88.455 35.505 89.210 ;
        RECT 36.690 88.520 36.860 89.210 ;
        RECT 37.220 89.060 38.405 89.230 ;
        RECT 40.045 89.530 40.420 89.860 ;
        RECT 40.590 89.530 40.920 90.255 ;
        RECT 37.220 89.040 37.390 89.060 ;
        RECT 37.030 88.710 37.390 89.040 ;
        RECT 34.805 87.360 35.505 88.455 ;
        RECT 35.675 87.095 36.005 88.520 ;
        RECT 36.210 87.095 36.510 88.135 ;
        RECT 36.690 87.360 37.050 88.520 ;
        RECT 37.220 88.390 37.390 88.710 ;
        RECT 37.610 88.560 38.395 88.890 ;
        RECT 40.045 88.760 40.215 89.530 ;
        RECT 41.090 89.360 41.420 89.990 ;
        RECT 41.600 89.530 41.770 90.255 ;
        RECT 41.950 89.360 42.280 89.990 ;
        RECT 42.460 89.530 42.710 90.255 ;
        RECT 42.925 89.530 43.300 89.860 ;
        RECT 43.470 89.530 43.800 90.255 ;
        RECT 40.385 88.930 40.785 89.260 ;
        RECT 41.090 89.190 42.305 89.360 ;
        RECT 40.955 88.760 41.965 88.990 ;
        RECT 40.045 88.590 41.965 88.760 ;
        RECT 37.220 88.220 38.050 88.390 ;
        RECT 37.220 87.095 37.550 88.050 ;
        RECT 37.720 87.360 38.050 88.220 ;
        RECT 40.045 87.360 40.425 88.590 ;
        RECT 42.135 88.420 42.305 89.190 ;
        RECT 42.925 88.760 43.095 89.530 ;
        RECT 43.970 89.360 44.300 89.990 ;
        RECT 44.480 89.530 44.650 90.255 ;
        RECT 44.830 89.360 45.160 89.990 ;
        RECT 45.340 89.530 45.590 90.255 ;
        RECT 45.850 89.680 46.180 89.970 ;
        RECT 45.850 89.510 46.575 89.680 ;
        RECT 46.750 89.510 47.000 90.255 ;
        RECT 43.265 88.930 43.665 89.260 ;
        RECT 43.970 89.190 45.185 89.360 ;
        RECT 43.835 88.760 44.845 88.990 ;
        RECT 42.925 88.590 44.845 88.760 ;
        RECT 40.595 87.095 40.845 88.420 ;
        RECT 41.045 88.250 42.305 88.420 ;
        RECT 41.045 87.360 41.375 88.250 ;
        RECT 41.575 87.095 41.825 88.080 ;
        RECT 42.025 87.360 42.305 88.250 ;
        RECT 42.475 87.095 42.725 88.520 ;
        RECT 42.925 87.360 43.305 88.590 ;
        RECT 45.015 88.420 45.185 89.190 ;
        RECT 43.475 87.095 43.725 88.420 ;
        RECT 43.925 88.250 45.185 88.420 ;
        RECT 43.925 87.360 44.255 88.250 ;
        RECT 44.455 87.095 44.705 88.080 ;
        RECT 44.905 87.360 45.185 88.250 ;
        RECT 45.355 87.095 45.605 88.520 ;
        RECT 45.845 88.170 46.235 89.340 ;
        RECT 46.405 88.030 46.575 89.510 ;
        RECT 47.175 89.370 47.560 89.990 ;
        RECT 47.730 89.540 48.060 90.255 ;
        RECT 48.230 89.840 50.155 90.010 ;
        RECT 50.635 89.945 51.030 90.255 ;
        RECT 48.230 89.540 48.755 89.840 ;
        RECT 49.985 89.775 50.155 89.840 ;
        RECT 51.200 89.915 53.140 90.085 ;
        RECT 51.200 89.775 51.370 89.915 ;
        RECT 46.745 88.200 47.005 89.210 ;
        RECT 47.175 89.200 48.415 89.370 ;
        RECT 47.175 88.530 47.345 89.200 ;
        RECT 47.515 88.700 47.995 89.030 ;
        RECT 48.165 88.790 48.415 89.200 ;
        RECT 47.765 88.560 47.995 88.700 ;
        RECT 48.585 88.780 48.755 89.540 ;
        RECT 48.925 89.120 49.175 89.670 ;
        RECT 49.345 89.290 49.815 89.670 ;
        RECT 49.985 89.605 51.370 89.775 ;
        RECT 51.540 89.435 51.870 89.675 ;
        RECT 48.925 88.950 49.475 89.120 ;
        RECT 48.585 88.620 49.135 88.780 ;
        RECT 47.175 88.200 47.585 88.530 ;
        RECT 48.235 88.450 49.135 88.620 ;
        RECT 48.235 88.170 48.485 88.450 ;
        RECT 49.305 88.280 49.475 88.950 ;
        RECT 48.730 88.110 49.475 88.280 ;
        RECT 46.405 88.000 47.395 88.030 ;
        RECT 48.730 88.000 48.980 88.110 ;
        RECT 46.405 87.860 48.980 88.000 ;
        RECT 49.645 87.940 49.815 89.290 ;
        RECT 49.985 89.265 51.870 89.435 ;
        RECT 49.985 88.215 50.165 89.265 ;
        RECT 51.540 89.210 51.870 89.265 ;
        RECT 50.335 88.765 51.370 89.095 ;
        RECT 50.335 88.020 50.505 88.765 ;
        RECT 50.675 88.190 51.005 88.545 ;
        RECT 50.335 87.940 50.970 88.020 ;
        RECT 46.405 87.820 46.605 87.860 ;
        RECT 47.225 87.830 48.980 87.860 ;
        RECT 45.825 87.095 46.075 87.820 ;
        RECT 46.275 87.360 46.605 87.820 ;
        RECT 46.805 87.095 47.055 87.690 ;
        RECT 47.705 87.095 48.035 87.660 ;
        RECT 48.730 87.615 48.980 87.830 ;
        RECT 49.180 87.770 50.970 87.940 ;
        RECT 49.180 87.615 49.510 87.770 ;
        RECT 50.105 87.095 50.435 87.600 ;
        RECT 51.200 87.095 51.530 88.595 ;
        RECT 51.700 88.475 51.870 89.210 ;
        RECT 52.040 89.495 52.800 89.745 ;
        RECT 52.040 88.825 52.210 89.495 ;
        RECT 52.970 89.325 53.140 89.915 ;
        RECT 53.465 89.495 53.795 90.255 ;
        RECT 54.335 89.325 54.665 89.955 ;
        RECT 54.895 89.495 55.145 90.255 ;
        RECT 52.410 88.995 53.140 89.325 ;
        RECT 53.310 89.155 54.910 89.325 ;
        RECT 53.310 88.995 53.640 89.155 ;
        RECT 52.040 88.655 52.370 88.825 ;
        RECT 51.700 87.585 52.030 88.475 ;
        RECT 52.200 87.865 52.370 88.655 ;
        RECT 52.685 88.035 53.015 88.995 ;
        RECT 54.240 88.825 54.570 88.985 ;
        RECT 53.185 88.655 54.570 88.825 ;
        RECT 53.185 87.865 53.355 88.655 ;
        RECT 54.740 88.485 54.910 89.155 ;
        RECT 55.325 88.955 55.655 89.990 ;
        RECT 53.525 88.085 54.065 88.420 ;
        RECT 54.235 88.315 54.910 88.485 ;
        RECT 55.105 88.625 55.655 88.955 ;
        RECT 55.885 89.210 56.215 89.990 ;
        RECT 56.395 89.210 56.645 90.255 ;
        RECT 56.875 89.550 57.205 89.990 ;
        RECT 57.375 89.660 58.065 90.255 ;
        RECT 54.235 87.895 54.405 88.315 ;
        RECT 52.200 87.535 53.355 87.865 ;
        RECT 53.525 87.095 53.855 87.895 ;
        RECT 54.040 87.435 54.405 87.895 ;
        RECT 54.575 87.095 54.905 88.145 ;
        RECT 55.105 87.435 55.275 88.625 ;
        RECT 55.885 88.455 56.145 89.210 ;
        RECT 56.875 88.520 57.115 89.550 ;
        RECT 58.235 89.380 58.565 89.990 ;
        RECT 57.285 89.210 58.565 89.380 ;
        RECT 59.245 89.530 59.620 89.860 ;
        RECT 59.790 89.530 60.120 90.255 ;
        RECT 57.285 88.710 57.675 89.210 ;
        RECT 55.445 87.360 56.145 88.455 ;
        RECT 56.315 87.095 56.645 88.520 ;
        RECT 56.875 87.360 57.335 88.520 ;
        RECT 57.505 88.390 57.675 88.710 ;
        RECT 57.845 88.560 58.555 89.040 ;
        RECT 59.245 88.760 59.415 89.530 ;
        RECT 60.290 89.360 60.620 89.990 ;
        RECT 60.800 89.530 60.970 90.255 ;
        RECT 61.150 89.360 61.480 89.990 ;
        RECT 61.660 89.530 61.910 90.255 ;
        RECT 59.585 88.930 59.985 89.260 ;
        RECT 60.290 89.190 61.505 89.360 ;
        RECT 62.130 89.235 62.430 90.255 ;
        RECT 60.155 88.760 61.165 88.990 ;
        RECT 59.245 88.590 61.165 88.760 ;
        RECT 57.505 88.220 58.335 88.390 ;
        RECT 57.505 87.095 57.835 88.050 ;
        RECT 58.005 87.360 58.335 88.220 ;
        RECT 59.245 87.360 59.625 88.590 ;
        RECT 61.335 88.420 61.505 89.190 ;
        RECT 62.690 88.755 63.260 90.255 ;
        RECT 63.970 89.535 64.300 90.255 ;
        RECT 65.005 89.530 65.380 89.860 ;
        RECT 65.550 89.530 65.880 90.255 ;
        RECT 59.795 87.095 60.045 88.420 ;
        RECT 60.245 88.250 61.505 88.420 ;
        RECT 60.245 87.360 60.575 88.250 ;
        RECT 60.775 87.095 61.025 88.080 ;
        RECT 61.225 87.360 61.505 88.250 ;
        RECT 61.675 87.095 61.925 88.520 ;
        RECT 62.130 87.095 62.430 88.135 ;
        RECT 62.615 87.095 62.945 88.410 ;
        RECT 63.665 87.095 64.235 89.090 ;
        RECT 65.005 88.760 65.175 89.530 ;
        RECT 66.050 89.360 66.380 89.990 ;
        RECT 66.560 89.530 66.730 90.255 ;
        RECT 66.910 89.360 67.240 89.990 ;
        RECT 67.420 89.530 67.670 90.255 ;
        RECT 67.940 89.535 68.270 90.255 ;
        RECT 65.345 88.930 65.745 89.260 ;
        RECT 66.050 89.190 67.265 89.360 ;
        RECT 65.915 88.760 66.925 88.990 ;
        RECT 65.005 88.590 66.925 88.760 ;
        RECT 65.005 87.360 65.385 88.590 ;
        RECT 67.095 88.420 67.265 89.190 ;
        RECT 65.555 87.095 65.805 88.420 ;
        RECT 66.005 88.250 67.265 88.420 ;
        RECT 66.005 87.360 66.335 88.250 ;
        RECT 66.535 87.095 66.785 88.080 ;
        RECT 66.985 87.360 67.265 88.250 ;
        RECT 67.435 87.095 67.685 88.520 ;
        RECT 68.005 87.095 68.575 89.090 ;
        RECT 68.980 88.755 69.550 90.255 ;
        RECT 69.295 87.095 69.625 88.410 ;
        RECT 112.980 87.995 113.150 93.045 ;
        RECT 113.780 92.535 114.280 92.705 ;
        RECT 113.550 91.825 113.720 92.365 ;
        RECT 114.340 91.825 114.510 92.365 ;
        RECT 113.780 91.485 114.280 91.655 ;
        RECT 113.550 90.775 113.720 91.315 ;
        RECT 114.340 90.775 114.510 91.315 ;
        RECT 113.780 90.435 114.280 90.605 ;
        RECT 113.550 89.725 113.720 90.265 ;
        RECT 114.340 89.725 114.510 90.265 ;
        RECT 113.780 89.385 114.280 89.555 ;
        RECT 113.550 88.675 113.720 89.215 ;
        RECT 114.340 88.675 114.510 89.215 ;
        RECT 113.780 88.335 114.280 88.505 ;
        RECT 114.910 87.995 115.080 93.045 ;
        RECT 112.980 87.825 115.080 87.995 ;
        RECT 115.440 93.045 117.540 93.215 ;
        RECT 112.980 87.295 115.080 87.465 ;
        RECT 10.200 86.925 69.720 87.095 ;
        RECT 10.295 85.610 10.625 86.925 ;
        RECT 10.370 83.765 10.940 85.265 ;
        RECT 11.345 84.930 11.915 86.925 ;
        RECT 12.715 85.500 12.965 86.925 ;
        RECT 13.135 85.770 13.415 86.660 ;
        RECT 13.615 85.940 13.865 86.925 ;
        RECT 14.065 85.770 14.395 86.660 ;
        RECT 13.135 85.600 14.395 85.770 ;
        RECT 14.595 85.600 14.845 86.925 ;
        RECT 13.135 84.830 13.305 85.600 ;
        RECT 15.015 85.430 15.395 86.660 ;
        RECT 23.250 85.885 23.550 86.925 ;
        RECT 23.735 85.610 24.065 86.925 ;
        RECT 13.475 85.260 15.395 85.430 ;
        RECT 13.475 85.030 14.485 85.260 ;
        RECT 13.135 84.660 14.350 84.830 ;
        RECT 14.655 84.760 15.055 85.090 ;
        RECT 11.650 83.765 11.980 84.485 ;
        RECT 12.730 83.765 12.980 84.490 ;
        RECT 13.160 84.030 13.490 84.660 ;
        RECT 13.670 83.765 13.840 84.490 ;
        RECT 14.020 84.030 14.350 84.660 ;
        RECT 15.225 84.490 15.395 85.260 ;
        RECT 14.520 83.765 14.850 84.490 ;
        RECT 15.020 84.160 15.395 84.490 ;
        RECT 23.250 83.765 23.550 84.785 ;
        RECT 23.810 83.765 24.380 85.265 ;
        RECT 24.785 84.930 25.355 86.925 ;
        RECT 26.865 85.800 27.195 86.660 ;
        RECT 27.365 85.970 27.695 86.925 ;
        RECT 26.865 85.630 27.695 85.800 ;
        RECT 26.645 84.980 27.355 85.460 ;
        RECT 27.525 85.310 27.695 85.630 ;
        RECT 27.865 85.500 28.325 86.660 ;
        RECT 32.375 85.610 32.705 86.925 ;
        RECT 27.525 84.810 27.915 85.310 ;
        RECT 26.635 84.640 27.915 84.810 ;
        RECT 25.090 83.765 25.420 84.485 ;
        RECT 26.635 84.030 26.965 84.640 ;
        RECT 28.085 84.470 28.325 85.500 ;
        RECT 27.135 83.765 27.825 84.360 ;
        RECT 27.995 84.030 28.325 84.470 ;
        RECT 32.450 83.765 33.020 85.265 ;
        RECT 33.425 84.930 33.995 86.925 ;
        RECT 34.545 85.800 34.875 86.660 ;
        RECT 35.045 85.970 35.375 86.925 ;
        RECT 34.545 85.630 35.375 85.800 ;
        RECT 34.325 84.980 35.035 85.460 ;
        RECT 35.205 85.310 35.375 85.630 ;
        RECT 35.545 85.500 36.005 86.660 ;
        RECT 36.210 85.885 36.510 86.925 ;
        RECT 36.715 85.500 37.045 86.925 ;
        RECT 37.215 85.565 37.915 86.660 ;
        RECT 35.205 84.810 35.595 85.310 ;
        RECT 34.315 84.640 35.595 84.810 ;
        RECT 33.730 83.765 34.060 84.485 ;
        RECT 34.315 84.030 34.645 84.640 ;
        RECT 35.765 84.470 36.005 85.500 ;
        RECT 37.215 84.810 37.475 85.565 ;
        RECT 38.085 85.395 38.255 86.585 ;
        RECT 38.455 85.875 38.785 86.925 ;
        RECT 38.955 86.125 39.320 86.585 ;
        RECT 39.505 86.125 39.835 86.925 ;
        RECT 40.005 86.155 41.160 86.485 ;
        RECT 38.955 85.705 39.125 86.125 ;
        RECT 34.815 83.765 35.505 84.360 ;
        RECT 35.675 84.030 36.005 84.470 ;
        RECT 36.210 83.765 36.510 84.785 ;
        RECT 36.715 83.765 36.965 84.810 ;
        RECT 37.145 84.030 37.475 84.810 ;
        RECT 37.705 85.065 38.255 85.395 ;
        RECT 38.450 85.535 39.125 85.705 ;
        RECT 39.295 85.600 39.835 85.935 ;
        RECT 37.705 84.030 38.035 85.065 ;
        RECT 38.450 84.865 38.620 85.535 ;
        RECT 40.005 85.365 40.175 86.155 ;
        RECT 38.790 85.195 40.175 85.365 ;
        RECT 38.790 85.035 39.120 85.195 ;
        RECT 40.345 85.025 40.675 85.985 ;
        RECT 40.990 85.365 41.160 86.155 ;
        RECT 41.330 85.545 41.660 86.435 ;
        RECT 40.990 85.195 41.320 85.365 ;
        RECT 39.720 84.865 40.050 85.025 ;
        RECT 38.450 84.695 40.050 84.865 ;
        RECT 40.220 84.695 40.950 85.025 ;
        RECT 38.215 83.765 38.465 84.525 ;
        RECT 38.695 84.065 39.025 84.695 ;
        RECT 39.565 83.765 39.895 84.525 ;
        RECT 40.220 84.105 40.390 84.695 ;
        RECT 41.150 84.525 41.320 85.195 ;
        RECT 40.560 84.275 41.320 84.525 ;
        RECT 41.490 84.810 41.660 85.545 ;
        RECT 41.830 85.425 42.160 86.925 ;
        RECT 42.925 86.420 43.255 86.925 ;
        RECT 43.850 86.250 44.180 86.405 ;
        RECT 42.390 86.080 44.180 86.250 ;
        RECT 44.380 86.190 44.630 86.405 ;
        RECT 45.325 86.360 45.655 86.925 ;
        RECT 46.305 86.330 46.555 86.925 ;
        RECT 46.755 86.200 47.085 86.660 ;
        RECT 47.285 86.200 47.535 86.925 ;
        RECT 44.380 86.160 46.135 86.190 ;
        RECT 46.755 86.160 46.955 86.200 ;
        RECT 42.390 86.000 43.025 86.080 ;
        RECT 42.355 85.475 42.685 85.830 ;
        RECT 42.855 85.255 43.025 86.000 ;
        RECT 41.990 84.925 43.025 85.255 ;
        RECT 41.490 84.755 41.820 84.810 ;
        RECT 43.195 84.755 43.375 85.805 ;
        RECT 41.490 84.585 43.375 84.755 ;
        RECT 43.545 84.730 43.715 86.080 ;
        RECT 44.380 86.020 46.955 86.160 ;
        RECT 44.380 85.910 44.630 86.020 ;
        RECT 45.965 85.990 46.955 86.020 ;
        RECT 43.885 85.740 44.630 85.910 ;
        RECT 43.885 85.070 44.055 85.740 ;
        RECT 44.875 85.570 45.125 85.850 ;
        RECT 44.225 85.400 45.125 85.570 ;
        RECT 45.775 85.490 46.185 85.820 ;
        RECT 44.225 85.240 44.775 85.400 ;
        RECT 43.885 84.900 44.435 85.070 ;
        RECT 41.490 84.345 41.820 84.585 ;
        RECT 41.990 84.245 43.375 84.415 ;
        RECT 43.545 84.350 44.015 84.730 ;
        RECT 44.185 84.350 44.435 84.900 ;
        RECT 44.605 84.480 44.775 85.240 ;
        RECT 45.365 85.320 45.595 85.460 ;
        RECT 44.945 84.820 45.195 85.230 ;
        RECT 45.365 84.990 45.845 85.320 ;
        RECT 46.015 84.820 46.185 85.490 ;
        RECT 44.945 84.650 46.185 84.820 ;
        RECT 46.355 84.810 46.615 85.820 ;
        RECT 41.990 84.105 42.160 84.245 ;
        RECT 40.220 83.935 42.160 84.105 ;
        RECT 43.205 84.180 43.375 84.245 ;
        RECT 44.605 84.180 45.130 84.480 ;
        RECT 42.330 83.765 42.725 84.075 ;
        RECT 43.205 84.010 45.130 84.180 ;
        RECT 45.300 83.765 45.630 84.480 ;
        RECT 45.800 84.030 46.185 84.650 ;
        RECT 46.785 84.510 46.955 85.990 ;
        RECT 49.170 85.885 49.470 86.925 ;
        RECT 47.125 84.680 47.515 85.850 ;
        RECT 49.675 85.500 50.005 86.925 ;
        RECT 50.175 85.565 50.875 86.660 ;
        RECT 50.175 84.810 50.435 85.565 ;
        RECT 51.045 85.395 51.215 86.585 ;
        RECT 51.415 85.875 51.745 86.925 ;
        RECT 51.915 86.125 52.280 86.585 ;
        RECT 52.465 86.125 52.795 86.925 ;
        RECT 52.965 86.155 54.120 86.485 ;
        RECT 51.915 85.705 52.085 86.125 ;
        RECT 46.360 83.765 46.610 84.510 ;
        RECT 46.785 84.340 47.510 84.510 ;
        RECT 47.180 84.050 47.510 84.340 ;
        RECT 49.170 83.765 49.470 84.785 ;
        RECT 49.675 83.765 49.925 84.810 ;
        RECT 50.105 84.030 50.435 84.810 ;
        RECT 50.665 85.065 51.215 85.395 ;
        RECT 51.410 85.535 52.085 85.705 ;
        RECT 52.255 85.600 52.795 85.935 ;
        RECT 50.665 84.030 50.995 85.065 ;
        RECT 51.410 84.865 51.580 85.535 ;
        RECT 52.965 85.365 53.135 86.155 ;
        RECT 51.750 85.195 53.135 85.365 ;
        RECT 51.750 85.035 52.080 85.195 ;
        RECT 53.305 85.025 53.635 85.985 ;
        RECT 53.950 85.365 54.120 86.155 ;
        RECT 54.290 85.545 54.620 86.435 ;
        RECT 53.950 85.195 54.280 85.365 ;
        RECT 52.680 84.865 53.010 85.025 ;
        RECT 51.410 84.695 53.010 84.865 ;
        RECT 53.180 84.695 53.910 85.025 ;
        RECT 51.175 83.765 51.425 84.525 ;
        RECT 51.655 84.065 51.985 84.695 ;
        RECT 52.525 83.765 52.855 84.525 ;
        RECT 53.180 84.105 53.350 84.695 ;
        RECT 54.110 84.525 54.280 85.195 ;
        RECT 53.520 84.275 54.280 84.525 ;
        RECT 54.450 84.810 54.620 85.545 ;
        RECT 54.790 85.425 55.120 86.925 ;
        RECT 55.885 86.420 56.215 86.925 ;
        RECT 56.810 86.250 57.140 86.405 ;
        RECT 55.350 86.080 57.140 86.250 ;
        RECT 57.340 86.190 57.590 86.405 ;
        RECT 58.285 86.360 58.615 86.925 ;
        RECT 59.265 86.330 59.515 86.925 ;
        RECT 59.715 86.200 60.045 86.660 ;
        RECT 60.245 86.200 60.495 86.925 ;
        RECT 57.340 86.160 59.095 86.190 ;
        RECT 59.715 86.160 59.915 86.200 ;
        RECT 55.350 86.000 55.985 86.080 ;
        RECT 55.315 85.475 55.645 85.830 ;
        RECT 55.815 85.255 55.985 86.000 ;
        RECT 54.950 84.925 55.985 85.255 ;
        RECT 54.450 84.755 54.780 84.810 ;
        RECT 56.155 84.755 56.335 85.805 ;
        RECT 54.450 84.585 56.335 84.755 ;
        RECT 56.505 84.730 56.675 86.080 ;
        RECT 57.340 86.020 59.915 86.160 ;
        RECT 57.340 85.910 57.590 86.020 ;
        RECT 58.925 85.990 59.915 86.020 ;
        RECT 56.845 85.740 57.590 85.910 ;
        RECT 56.845 85.070 57.015 85.740 ;
        RECT 57.835 85.570 58.085 85.850 ;
        RECT 57.185 85.400 58.085 85.570 ;
        RECT 58.735 85.490 59.145 85.820 ;
        RECT 57.185 85.240 57.735 85.400 ;
        RECT 56.845 84.900 57.395 85.070 ;
        RECT 54.450 84.345 54.780 84.585 ;
        RECT 54.950 84.245 56.335 84.415 ;
        RECT 56.505 84.350 56.975 84.730 ;
        RECT 57.145 84.350 57.395 84.900 ;
        RECT 57.565 84.480 57.735 85.240 ;
        RECT 58.325 85.320 58.555 85.460 ;
        RECT 57.905 84.820 58.155 85.230 ;
        RECT 58.325 84.990 58.805 85.320 ;
        RECT 58.975 84.820 59.145 85.490 ;
        RECT 57.905 84.650 59.145 84.820 ;
        RECT 59.315 84.810 59.575 85.820 ;
        RECT 54.950 84.105 55.120 84.245 ;
        RECT 53.180 83.935 55.120 84.105 ;
        RECT 56.165 84.180 56.335 84.245 ;
        RECT 57.565 84.180 58.090 84.480 ;
        RECT 55.290 83.765 55.685 84.075 ;
        RECT 56.165 84.010 58.090 84.180 ;
        RECT 58.260 83.765 58.590 84.480 ;
        RECT 58.760 84.030 59.145 84.650 ;
        RECT 59.745 84.510 59.915 85.990 ;
        RECT 62.130 85.885 62.430 86.925 ;
        RECT 60.085 84.680 60.475 85.850 ;
        RECT 62.635 85.500 63.095 86.660 ;
        RECT 63.265 85.970 63.595 86.925 ;
        RECT 63.765 85.800 64.095 86.660 ;
        RECT 63.265 85.630 64.095 85.800 ;
        RECT 59.320 83.765 59.570 84.510 ;
        RECT 59.745 84.340 60.470 84.510 ;
        RECT 60.140 84.050 60.470 84.340 ;
        RECT 62.130 83.765 62.430 84.785 ;
        RECT 62.635 84.470 62.875 85.500 ;
        RECT 63.265 85.310 63.435 85.630 ;
        RECT 63.045 84.810 63.435 85.310 ;
        RECT 63.605 84.980 64.315 85.460 ;
        RECT 65.005 85.430 65.385 86.660 ;
        RECT 65.555 85.600 65.805 86.925 ;
        RECT 66.005 85.770 66.335 86.660 ;
        RECT 66.535 85.940 66.785 86.925 ;
        RECT 66.985 85.770 67.265 86.660 ;
        RECT 66.005 85.600 67.265 85.770 ;
        RECT 65.005 85.260 66.925 85.430 ;
        RECT 63.045 84.640 64.325 84.810 ;
        RECT 62.635 84.030 62.965 84.470 ;
        RECT 63.135 83.765 63.825 84.360 ;
        RECT 63.995 84.030 64.325 84.640 ;
        RECT 65.005 84.490 65.175 85.260 ;
        RECT 65.345 84.760 65.745 85.090 ;
        RECT 65.915 85.030 66.925 85.260 ;
        RECT 67.095 84.830 67.265 85.600 ;
        RECT 67.435 85.500 67.685 86.925 ;
        RECT 68.005 84.930 68.575 86.925 ;
        RECT 69.295 85.610 69.625 86.925 ;
        RECT 66.050 84.660 67.265 84.830 ;
        RECT 65.005 84.160 65.380 84.490 ;
        RECT 65.550 83.765 65.880 84.490 ;
        RECT 66.050 84.030 66.380 84.660 ;
        RECT 66.560 83.765 66.730 84.490 ;
        RECT 66.910 84.030 67.240 84.660 ;
        RECT 67.420 83.765 67.670 84.490 ;
        RECT 67.940 83.765 68.270 84.485 ;
        RECT 68.980 83.765 69.550 85.265 ;
        RECT 10.200 83.595 69.720 83.765 ;
        RECT 112.980 77.885 113.150 87.295 ;
        RECT 113.780 86.785 114.280 86.955 ;
        RECT 113.550 85.030 113.720 86.570 ;
        RECT 114.340 85.030 114.510 86.570 ;
        RECT 113.780 84.645 114.280 84.815 ;
        RECT 113.550 82.890 113.720 84.430 ;
        RECT 114.340 82.890 114.510 84.430 ;
        RECT 113.780 82.505 114.280 82.675 ;
        RECT 113.550 80.750 113.720 82.290 ;
        RECT 114.340 80.750 114.510 82.290 ;
        RECT 113.780 80.365 114.280 80.535 ;
        RECT 113.550 78.610 113.720 80.150 ;
        RECT 114.340 78.610 114.510 80.150 ;
        RECT 113.780 78.225 114.280 78.395 ;
        RECT 114.910 77.885 115.080 87.295 ;
        RECT 115.440 83.635 115.610 93.045 ;
        RECT 116.240 92.535 116.740 92.705 ;
        RECT 116.010 90.780 116.180 92.320 ;
        RECT 116.800 90.780 116.970 92.320 ;
        RECT 116.240 90.395 116.740 90.565 ;
        RECT 116.010 88.640 116.180 90.180 ;
        RECT 116.800 88.640 116.970 90.180 ;
        RECT 116.240 88.255 116.740 88.425 ;
        RECT 116.010 86.500 116.180 88.040 ;
        RECT 116.800 86.500 116.970 88.040 ;
        RECT 116.240 86.115 116.740 86.285 ;
        RECT 116.010 84.360 116.180 85.900 ;
        RECT 116.800 84.360 116.970 85.900 ;
        RECT 116.240 83.975 116.740 84.145 ;
        RECT 117.370 83.635 117.540 93.045 ;
        RECT 117.900 93.050 120.000 93.220 ;
        RECT 117.900 88.000 118.070 93.050 ;
        RECT 118.700 92.540 119.200 92.710 ;
        RECT 118.470 91.830 118.640 92.370 ;
        RECT 119.260 91.830 119.430 92.370 ;
        RECT 118.700 91.490 119.200 91.660 ;
        RECT 118.470 90.780 118.640 91.320 ;
        RECT 119.260 90.780 119.430 91.320 ;
        RECT 118.700 90.440 119.200 90.610 ;
        RECT 118.470 89.730 118.640 90.270 ;
        RECT 119.260 89.730 119.430 90.270 ;
        RECT 118.700 89.390 119.200 89.560 ;
        RECT 118.470 88.680 118.640 89.220 ;
        RECT 119.260 88.680 119.430 89.220 ;
        RECT 118.700 88.340 119.200 88.510 ;
        RECT 119.830 88.000 120.000 93.050 ;
        RECT 117.900 87.830 120.000 88.000 ;
        RECT 120.360 93.050 124.390 93.220 ;
        RECT 115.440 83.465 117.540 83.635 ;
        RECT 117.900 87.300 120.000 87.470 ;
        RECT 112.980 77.715 115.080 77.885 ;
        RECT 115.440 82.935 117.540 83.105 ;
        RECT 115.440 77.885 115.610 82.935 ;
        RECT 116.240 82.425 116.740 82.595 ;
        RECT 116.010 81.715 116.180 82.255 ;
        RECT 116.800 81.715 116.970 82.255 ;
        RECT 116.240 81.375 116.740 81.545 ;
        RECT 116.010 80.665 116.180 81.205 ;
        RECT 116.800 80.665 116.970 81.205 ;
        RECT 116.240 80.325 116.740 80.495 ;
        RECT 116.010 79.615 116.180 80.155 ;
        RECT 116.800 79.615 116.970 80.155 ;
        RECT 116.240 79.275 116.740 79.445 ;
        RECT 116.010 78.565 116.180 79.105 ;
        RECT 116.800 78.565 116.970 79.105 ;
        RECT 116.240 78.225 116.740 78.395 ;
        RECT 117.370 77.885 117.540 82.935 ;
        RECT 115.440 77.715 117.540 77.885 ;
        RECT 117.900 77.890 118.070 87.300 ;
        RECT 118.700 86.790 119.200 86.960 ;
        RECT 118.470 85.035 118.640 86.575 ;
        RECT 119.260 85.035 119.430 86.575 ;
        RECT 118.700 84.650 119.200 84.820 ;
        RECT 118.470 82.895 118.640 84.435 ;
        RECT 119.260 82.895 119.430 84.435 ;
        RECT 118.700 82.510 119.200 82.680 ;
        RECT 118.470 80.755 118.640 82.295 ;
        RECT 119.260 80.755 119.430 82.295 ;
        RECT 118.700 80.370 119.200 80.540 ;
        RECT 118.470 78.615 118.640 80.155 ;
        RECT 119.260 78.615 119.430 80.155 ;
        RECT 118.700 78.230 119.200 78.400 ;
        RECT 119.830 77.890 120.000 87.300 ;
        RECT 120.360 83.640 120.530 93.050 ;
        RECT 121.160 92.540 121.660 92.710 ;
        RECT 120.930 90.785 121.100 92.325 ;
        RECT 121.720 90.785 121.890 92.325 ;
        RECT 121.160 90.400 121.660 90.570 ;
        RECT 120.930 88.645 121.100 90.185 ;
        RECT 121.720 88.645 121.890 90.185 ;
        RECT 121.160 88.260 121.660 88.430 ;
        RECT 120.930 86.505 121.100 88.045 ;
        RECT 121.720 86.505 121.890 88.045 ;
        RECT 121.160 86.120 121.660 86.290 ;
        RECT 120.930 84.365 121.100 85.905 ;
        RECT 121.720 84.365 121.890 85.905 ;
        RECT 121.160 83.980 121.660 84.150 ;
        RECT 122.290 83.640 122.460 93.050 ;
        RECT 123.090 92.540 123.590 92.710 ;
        RECT 122.860 90.785 123.030 92.325 ;
        RECT 123.650 90.785 123.820 92.325 ;
        RECT 123.090 90.400 123.590 90.570 ;
        RECT 122.860 88.645 123.030 90.185 ;
        RECT 123.650 88.645 123.820 90.185 ;
        RECT 123.090 88.260 123.590 88.430 ;
        RECT 122.860 86.505 123.030 88.045 ;
        RECT 123.650 86.505 123.820 88.045 ;
        RECT 123.090 86.120 123.590 86.290 ;
        RECT 122.860 84.365 123.030 85.905 ;
        RECT 123.650 84.365 123.820 85.905 ;
        RECT 123.090 83.980 123.590 84.150 ;
        RECT 124.220 83.640 124.390 93.050 ;
        RECT 124.750 93.050 128.780 93.220 ;
        RECT 124.750 88.000 124.920 93.050 ;
        RECT 125.550 92.540 126.050 92.710 ;
        RECT 125.320 91.830 125.490 92.370 ;
        RECT 126.110 91.830 126.280 92.370 ;
        RECT 125.550 91.490 126.050 91.660 ;
        RECT 125.320 90.780 125.490 91.320 ;
        RECT 126.110 90.780 126.280 91.320 ;
        RECT 125.550 90.440 126.050 90.610 ;
        RECT 125.320 89.730 125.490 90.270 ;
        RECT 126.110 89.730 126.280 90.270 ;
        RECT 125.550 89.390 126.050 89.560 ;
        RECT 125.320 88.680 125.490 89.220 ;
        RECT 126.110 88.680 126.280 89.220 ;
        RECT 125.550 88.340 126.050 88.510 ;
        RECT 126.680 88.000 126.850 93.050 ;
        RECT 127.480 92.540 127.980 92.710 ;
        RECT 127.250 91.830 127.420 92.370 ;
        RECT 128.040 91.830 128.210 92.370 ;
        RECT 127.480 91.490 127.980 91.660 ;
        RECT 127.250 90.780 127.420 91.320 ;
        RECT 128.040 90.780 128.210 91.320 ;
        RECT 127.480 90.440 127.980 90.610 ;
        RECT 127.250 89.730 127.420 90.270 ;
        RECT 128.040 89.730 128.210 90.270 ;
        RECT 127.480 89.390 127.980 89.560 ;
        RECT 127.250 88.680 127.420 89.220 ;
        RECT 128.040 88.680 128.210 89.220 ;
        RECT 127.480 88.340 127.980 88.510 ;
        RECT 128.610 88.000 128.780 93.050 ;
        RECT 124.750 87.830 128.780 88.000 ;
        RECT 129.120 93.000 129.290 93.210 ;
        RECT 132.450 93.085 132.620 93.210 ;
        RECT 129.120 92.670 130.175 93.000 ;
        RECT 129.120 92.070 129.290 92.670 ;
        RECT 130.345 92.585 130.825 93.085 ;
        RECT 131.025 92.755 134.045 93.085 ;
        RECT 130.345 92.500 132.185 92.585 ;
        RECT 129.555 92.255 132.185 92.500 ;
        RECT 129.555 92.240 130.825 92.255 ;
        RECT 129.120 91.740 130.175 92.070 ;
        RECT 129.120 91.070 129.290 91.740 ;
        RECT 130.345 91.570 130.825 92.240 ;
        RECT 132.450 92.085 132.620 92.755 ;
        RECT 134.245 92.585 134.725 93.085 ;
        RECT 135.780 93.000 135.950 93.210 ;
        RECT 134.895 92.670 135.950 93.000 ;
        RECT 132.885 92.500 134.725 92.585 ;
        RECT 132.885 92.255 135.515 92.500 ;
        RECT 134.245 92.240 135.515 92.255 ;
        RECT 131.025 91.755 134.045 92.085 ;
        RECT 129.555 91.555 130.825 91.570 ;
        RECT 129.555 91.385 132.185 91.555 ;
        RECT 129.555 91.310 130.515 91.385 ;
        RECT 129.555 91.240 130.385 91.310 ;
        RECT 129.120 90.740 130.045 91.070 ;
        RECT 129.120 90.210 129.290 90.740 ;
        RECT 130.215 90.560 130.385 91.240 ;
        RECT 129.555 90.390 130.385 90.560 ;
        RECT 129.120 89.880 130.045 90.210 ;
        RECT 129.120 89.270 129.290 89.880 ;
        RECT 130.215 89.700 130.385 90.390 ;
        RECT 129.555 89.450 130.385 89.700 ;
        RECT 130.555 89.450 130.985 91.140 ;
        RECT 131.155 90.735 131.325 91.385 ;
        RECT 132.450 91.185 132.620 91.755 ;
        RECT 134.245 91.570 134.725 92.240 ;
        RECT 135.780 92.070 135.950 92.670 ;
        RECT 134.895 91.740 135.950 92.070 ;
        RECT 134.245 91.555 135.515 91.570 ;
        RECT 132.885 91.385 135.515 91.555 ;
        RECT 131.495 90.935 133.575 91.185 ;
        RECT 131.155 90.405 132.185 90.735 ;
        RECT 131.155 89.705 131.325 90.405 ;
        RECT 132.450 90.235 132.620 90.935 ;
        RECT 133.745 90.735 133.915 91.385 ;
        RECT 134.555 91.310 135.515 91.385 ;
        RECT 134.685 91.240 135.515 91.310 ;
        RECT 132.885 90.405 133.915 90.735 ;
        RECT 131.495 89.905 133.575 90.235 ;
        RECT 131.155 89.455 132.185 89.705 ;
        RECT 129.120 89.020 130.335 89.270 ;
        RECT 129.120 88.680 129.290 89.020 ;
        RECT 130.620 88.765 130.820 89.450 ;
        RECT 132.450 89.255 132.620 89.905 ;
        RECT 133.745 89.705 133.915 90.405 ;
        RECT 132.885 89.455 133.915 89.705 ;
        RECT 134.085 89.450 134.515 91.140 ;
        RECT 134.685 90.560 134.855 91.240 ;
        RECT 135.780 91.070 135.950 91.740 ;
        RECT 135.025 90.740 135.950 91.070 ;
        RECT 134.685 90.390 135.515 90.560 ;
        RECT 134.685 89.700 134.855 90.390 ;
        RECT 135.780 90.210 135.950 90.740 ;
        RECT 135.025 89.880 135.950 90.210 ;
        RECT 134.685 89.450 135.515 89.700 ;
        RECT 131.025 89.005 134.045 89.255 ;
        RECT 132.450 88.765 132.620 89.005 ;
        RECT 134.250 88.765 134.450 89.450 ;
        RECT 135.780 89.270 135.950 89.880 ;
        RECT 134.735 89.020 135.950 89.270 ;
        RECT 129.120 88.350 130.175 88.680 ;
        RECT 120.360 83.470 124.390 83.640 ;
        RECT 129.120 87.750 129.290 88.350 ;
        RECT 130.345 88.265 130.825 88.765 ;
        RECT 131.025 88.435 134.045 88.765 ;
        RECT 130.345 88.180 132.185 88.265 ;
        RECT 129.555 87.935 132.185 88.180 ;
        RECT 129.555 87.920 130.825 87.935 ;
        RECT 129.120 87.420 130.175 87.750 ;
        RECT 129.120 86.750 129.290 87.420 ;
        RECT 130.345 87.250 130.825 87.920 ;
        RECT 132.450 87.765 132.620 88.435 ;
        RECT 134.245 88.265 134.725 88.765 ;
        RECT 135.780 88.680 135.950 89.020 ;
        RECT 134.895 88.350 135.950 88.680 ;
        RECT 132.885 88.180 134.725 88.265 ;
        RECT 132.885 87.935 135.515 88.180 ;
        RECT 134.245 87.920 135.515 87.935 ;
        RECT 131.025 87.435 134.045 87.765 ;
        RECT 129.555 87.235 130.825 87.250 ;
        RECT 129.555 87.065 132.185 87.235 ;
        RECT 129.555 86.990 130.515 87.065 ;
        RECT 129.555 86.920 130.385 86.990 ;
        RECT 129.120 86.420 130.045 86.750 ;
        RECT 129.120 85.890 129.290 86.420 ;
        RECT 130.215 86.240 130.385 86.920 ;
        RECT 129.555 86.070 130.385 86.240 ;
        RECT 129.120 85.560 130.045 85.890 ;
        RECT 129.120 84.950 129.290 85.560 ;
        RECT 130.215 85.380 130.385 86.070 ;
        RECT 129.555 85.130 130.385 85.380 ;
        RECT 130.555 85.130 130.985 86.820 ;
        RECT 131.155 86.415 131.325 87.065 ;
        RECT 132.450 86.865 132.620 87.435 ;
        RECT 134.245 87.250 134.725 87.920 ;
        RECT 135.780 87.750 135.950 88.350 ;
        RECT 136.990 93.045 139.090 93.215 ;
        RECT 136.990 87.995 137.160 93.045 ;
        RECT 137.790 92.535 138.290 92.705 ;
        RECT 137.560 91.825 137.730 92.365 ;
        RECT 138.350 91.825 138.520 92.365 ;
        RECT 137.790 91.485 138.290 91.655 ;
        RECT 137.560 90.775 137.730 91.315 ;
        RECT 138.350 90.775 138.520 91.315 ;
        RECT 137.790 90.435 138.290 90.605 ;
        RECT 137.560 89.725 137.730 90.265 ;
        RECT 138.350 89.725 138.520 90.265 ;
        RECT 137.790 89.385 138.290 89.555 ;
        RECT 137.560 88.675 137.730 89.215 ;
        RECT 138.350 88.675 138.520 89.215 ;
        RECT 137.790 88.335 138.290 88.505 ;
        RECT 138.920 87.995 139.090 93.045 ;
        RECT 136.990 87.825 139.090 87.995 ;
        RECT 139.450 93.045 141.550 93.215 ;
        RECT 134.895 87.420 135.950 87.750 ;
        RECT 134.245 87.235 135.515 87.250 ;
        RECT 132.885 87.065 135.515 87.235 ;
        RECT 131.495 86.615 133.575 86.865 ;
        RECT 131.155 86.085 132.185 86.415 ;
        RECT 131.155 85.385 131.325 86.085 ;
        RECT 132.450 85.915 132.620 86.615 ;
        RECT 133.745 86.415 133.915 87.065 ;
        RECT 134.555 86.990 135.515 87.065 ;
        RECT 134.685 86.920 135.515 86.990 ;
        RECT 132.885 86.085 133.915 86.415 ;
        RECT 131.495 85.585 133.575 85.915 ;
        RECT 131.155 85.135 132.185 85.385 ;
        RECT 129.120 84.700 130.335 84.950 ;
        RECT 129.120 84.480 129.290 84.700 ;
        RECT 129.120 84.180 130.310 84.480 ;
        RECT 129.120 83.975 129.290 84.180 ;
        RECT 129.120 83.645 130.045 83.975 ;
        RECT 130.620 83.965 130.820 85.130 ;
        RECT 132.450 84.935 132.620 85.585 ;
        RECT 133.745 85.385 133.915 86.085 ;
        RECT 132.885 85.135 133.915 85.385 ;
        RECT 134.085 85.130 134.515 86.820 ;
        RECT 134.685 86.240 134.855 86.920 ;
        RECT 135.780 86.750 135.950 87.420 ;
        RECT 135.025 86.420 135.950 86.750 ;
        RECT 134.685 86.070 135.515 86.240 ;
        RECT 134.685 85.380 134.855 86.070 ;
        RECT 135.780 85.890 135.950 86.420 ;
        RECT 135.025 85.560 135.950 85.890 ;
        RECT 134.685 85.130 135.515 85.380 ;
        RECT 131.025 84.685 134.045 84.935 ;
        RECT 132.450 84.480 132.620 84.685 ;
        RECT 131.410 84.180 133.660 84.480 ;
        RECT 132.450 83.970 132.620 84.180 ;
        RECT 130.215 83.735 131.325 83.965 ;
        RECT 117.900 77.720 120.000 77.890 ;
        RECT 129.120 83.065 129.290 83.645 ;
        RECT 130.215 83.465 130.385 83.735 ;
        RECT 131.155 83.520 131.325 83.735 ;
        RECT 131.495 83.720 133.575 83.970 ;
        RECT 134.255 83.965 134.455 85.130 ;
        RECT 135.780 84.950 135.950 85.560 ;
        RECT 134.735 84.700 135.950 84.950 ;
        RECT 135.780 84.480 135.950 84.700 ;
        RECT 134.760 84.180 135.950 84.480 ;
        RECT 135.780 83.975 135.950 84.180 ;
        RECT 133.745 83.735 134.855 83.965 ;
        RECT 129.555 83.295 130.385 83.465 ;
        RECT 129.120 82.735 130.045 83.065 ;
        RECT 129.120 82.135 129.290 82.735 ;
        RECT 130.215 82.555 130.385 83.295 ;
        RECT 129.555 82.305 130.385 82.555 ;
        RECT 129.120 81.805 130.335 82.135 ;
        RECT 130.555 81.815 130.985 83.490 ;
        RECT 131.155 83.190 132.185 83.520 ;
        RECT 131.155 82.620 131.325 83.190 ;
        RECT 132.450 82.990 132.620 83.720 ;
        RECT 133.745 83.520 133.915 83.735 ;
        RECT 132.885 83.190 133.915 83.520 ;
        RECT 131.495 82.820 133.575 82.990 ;
        RECT 131.155 82.290 132.185 82.620 ;
        RECT 132.450 82.090 132.620 82.820 ;
        RECT 133.745 82.620 133.915 83.190 ;
        RECT 132.885 82.290 133.915 82.620 ;
        RECT 131.155 81.840 133.915 82.090 ;
        RECT 129.120 81.065 129.290 81.805 ;
        RECT 130.620 81.565 130.820 81.815 ;
        RECT 129.555 81.235 132.185 81.565 ;
        RECT 132.450 81.065 132.620 81.840 ;
        RECT 134.085 81.815 134.515 83.490 ;
        RECT 134.685 83.465 134.855 83.735 ;
        RECT 135.025 83.645 135.950 83.975 ;
        RECT 134.685 83.295 135.515 83.465 ;
        RECT 134.685 82.555 134.855 83.295 ;
        RECT 135.780 83.065 135.950 83.645 ;
        RECT 135.025 82.735 135.950 83.065 ;
        RECT 134.685 82.305 135.515 82.555 ;
        RECT 135.780 82.135 135.950 82.735 ;
        RECT 134.250 81.565 134.450 81.815 ;
        RECT 134.735 81.805 135.950 82.135 ;
        RECT 132.885 81.235 135.515 81.565 ;
        RECT 135.780 81.065 135.950 81.805 ;
        RECT 129.120 80.735 130.335 81.065 ;
        RECT 129.120 80.160 129.290 80.735 ;
        RECT 130.505 80.375 130.985 81.065 ;
        RECT 131.155 80.735 133.915 81.065 ;
        RECT 129.120 79.860 130.310 80.160 ;
        RECT 129.120 79.145 129.290 79.860 ;
        RECT 130.570 79.645 130.770 80.375 ;
        RECT 132.450 80.160 132.620 80.735 ;
        RECT 134.085 80.375 134.565 81.065 ;
        RECT 134.735 80.735 135.950 81.065 ;
        RECT 131.410 79.860 133.660 80.160 ;
        RECT 129.555 79.315 132.185 79.645 ;
        RECT 132.450 79.145 132.620 79.860 ;
        RECT 134.300 79.645 134.500 80.375 ;
        RECT 135.780 80.160 135.950 80.735 ;
        RECT 134.760 79.860 135.950 80.160 ;
        RECT 132.885 79.315 135.515 79.645 ;
        RECT 135.780 79.145 135.950 79.860 ;
        RECT 129.120 78.815 130.335 79.145 ;
        RECT 129.120 77.350 129.290 78.815 ;
        RECT 130.505 78.455 130.985 79.145 ;
        RECT 131.155 78.815 133.915 79.145 ;
        RECT 132.450 78.225 132.620 78.815 ;
        RECT 134.085 78.455 134.565 79.145 ;
        RECT 134.735 78.815 135.950 79.145 ;
        RECT 129.555 77.840 130.215 78.170 ;
        RECT 130.385 77.895 130.755 78.225 ;
        RECT 131.025 77.895 134.045 78.225 ;
        RECT 134.315 77.895 134.685 78.225 ;
        RECT 135.780 78.200 135.950 78.815 ;
        RECT 130.045 77.725 130.215 77.840 ;
        RECT 130.045 77.555 132.185 77.725 ;
        RECT 130.385 77.495 132.185 77.555 ;
        RECT 129.120 77.020 130.215 77.350 ;
        RECT 132.450 77.325 132.620 77.895 ;
        RECT 134.855 77.870 135.950 78.200 ;
        RECT 132.885 77.665 134.685 77.725 ;
        RECT 132.885 77.495 135.025 77.665 ;
        RECT 134.855 77.380 135.025 77.495 ;
        RECT 129.120 76.265 129.290 77.020 ;
        RECT 130.385 76.995 130.755 77.325 ;
        RECT 131.025 76.995 134.045 77.325 ;
        RECT 134.315 76.995 134.685 77.325 ;
        RECT 134.855 77.050 135.515 77.380 ;
        RECT 130.490 76.765 130.690 76.995 ;
        RECT 129.555 76.435 132.185 76.765 ;
        RECT 132.450 76.265 132.620 76.995 ;
        RECT 135.780 76.890 135.950 77.870 ;
        RECT 136.990 87.295 139.090 87.465 ;
        RECT 136.990 77.885 137.160 87.295 ;
        RECT 137.790 86.785 138.290 86.955 ;
        RECT 137.560 85.030 137.730 86.570 ;
        RECT 138.350 85.030 138.520 86.570 ;
        RECT 137.790 84.645 138.290 84.815 ;
        RECT 137.560 82.890 137.730 84.430 ;
        RECT 138.350 82.890 138.520 84.430 ;
        RECT 137.790 82.505 138.290 82.675 ;
        RECT 137.560 80.750 137.730 82.290 ;
        RECT 138.350 80.750 138.520 82.290 ;
        RECT 137.790 80.365 138.290 80.535 ;
        RECT 137.560 78.610 137.730 80.150 ;
        RECT 138.350 78.610 138.520 80.150 ;
        RECT 137.790 78.225 138.290 78.395 ;
        RECT 138.920 77.885 139.090 87.295 ;
        RECT 139.450 83.635 139.620 93.045 ;
        RECT 140.250 92.535 140.750 92.705 ;
        RECT 140.020 90.780 140.190 92.320 ;
        RECT 140.810 90.780 140.980 92.320 ;
        RECT 140.250 90.395 140.750 90.565 ;
        RECT 140.020 88.640 140.190 90.180 ;
        RECT 140.810 88.640 140.980 90.180 ;
        RECT 140.250 88.255 140.750 88.425 ;
        RECT 140.020 86.500 140.190 88.040 ;
        RECT 140.810 86.500 140.980 88.040 ;
        RECT 140.250 86.115 140.750 86.285 ;
        RECT 140.020 84.360 140.190 85.900 ;
        RECT 140.810 84.360 140.980 85.900 ;
        RECT 140.250 83.975 140.750 84.145 ;
        RECT 141.380 83.635 141.550 93.045 ;
        RECT 141.910 93.050 144.010 93.220 ;
        RECT 141.910 88.000 142.080 93.050 ;
        RECT 142.710 92.540 143.210 92.710 ;
        RECT 142.480 91.830 142.650 92.370 ;
        RECT 143.270 91.830 143.440 92.370 ;
        RECT 142.710 91.490 143.210 91.660 ;
        RECT 142.480 90.780 142.650 91.320 ;
        RECT 143.270 90.780 143.440 91.320 ;
        RECT 142.710 90.440 143.210 90.610 ;
        RECT 142.480 89.730 142.650 90.270 ;
        RECT 143.270 89.730 143.440 90.270 ;
        RECT 142.710 89.390 143.210 89.560 ;
        RECT 142.480 88.680 142.650 89.220 ;
        RECT 143.270 88.680 143.440 89.220 ;
        RECT 142.710 88.340 143.210 88.510 ;
        RECT 143.840 88.000 144.010 93.050 ;
        RECT 141.910 87.830 144.010 88.000 ;
        RECT 144.370 93.050 148.400 93.220 ;
        RECT 139.450 83.465 141.550 83.635 ;
        RECT 141.910 87.300 144.010 87.470 ;
        RECT 136.990 77.715 139.090 77.885 ;
        RECT 139.450 82.935 141.550 83.105 ;
        RECT 139.450 77.885 139.620 82.935 ;
        RECT 140.250 82.425 140.750 82.595 ;
        RECT 140.020 81.715 140.190 82.255 ;
        RECT 140.810 81.715 140.980 82.255 ;
        RECT 140.250 81.375 140.750 81.545 ;
        RECT 140.020 80.665 140.190 81.205 ;
        RECT 140.810 80.665 140.980 81.205 ;
        RECT 140.250 80.325 140.750 80.495 ;
        RECT 140.020 79.615 140.190 80.155 ;
        RECT 140.810 79.615 140.980 80.155 ;
        RECT 140.250 79.275 140.750 79.445 ;
        RECT 140.020 78.565 140.190 79.105 ;
        RECT 140.810 78.565 140.980 79.105 ;
        RECT 140.250 78.225 140.750 78.395 ;
        RECT 141.380 77.885 141.550 82.935 ;
        RECT 139.450 77.715 141.550 77.885 ;
        RECT 141.910 77.890 142.080 87.300 ;
        RECT 142.710 86.790 143.210 86.960 ;
        RECT 142.480 85.035 142.650 86.575 ;
        RECT 143.270 85.035 143.440 86.575 ;
        RECT 142.710 84.650 143.210 84.820 ;
        RECT 142.480 82.895 142.650 84.435 ;
        RECT 143.270 82.895 143.440 84.435 ;
        RECT 142.710 82.510 143.210 82.680 ;
        RECT 142.480 80.755 142.650 82.295 ;
        RECT 143.270 80.755 143.440 82.295 ;
        RECT 142.710 80.370 143.210 80.540 ;
        RECT 142.480 78.615 142.650 80.155 ;
        RECT 143.270 78.615 143.440 80.155 ;
        RECT 142.710 78.230 143.210 78.400 ;
        RECT 143.840 77.890 144.010 87.300 ;
        RECT 144.370 83.640 144.540 93.050 ;
        RECT 145.170 92.540 145.670 92.710 ;
        RECT 144.940 90.785 145.110 92.325 ;
        RECT 145.730 90.785 145.900 92.325 ;
        RECT 145.170 90.400 145.670 90.570 ;
        RECT 144.940 88.645 145.110 90.185 ;
        RECT 145.730 88.645 145.900 90.185 ;
        RECT 145.170 88.260 145.670 88.430 ;
        RECT 144.940 86.505 145.110 88.045 ;
        RECT 145.730 86.505 145.900 88.045 ;
        RECT 145.170 86.120 145.670 86.290 ;
        RECT 144.940 84.365 145.110 85.905 ;
        RECT 145.730 84.365 145.900 85.905 ;
        RECT 145.170 83.980 145.670 84.150 ;
        RECT 146.300 83.640 146.470 93.050 ;
        RECT 147.100 92.540 147.600 92.710 ;
        RECT 146.870 90.785 147.040 92.325 ;
        RECT 147.660 90.785 147.830 92.325 ;
        RECT 147.100 90.400 147.600 90.570 ;
        RECT 146.870 88.645 147.040 90.185 ;
        RECT 147.660 88.645 147.830 90.185 ;
        RECT 147.100 88.260 147.600 88.430 ;
        RECT 146.870 86.505 147.040 88.045 ;
        RECT 147.660 86.505 147.830 88.045 ;
        RECT 147.100 86.120 147.600 86.290 ;
        RECT 146.870 84.365 147.040 85.905 ;
        RECT 147.660 84.365 147.830 85.905 ;
        RECT 147.100 83.980 147.600 84.150 ;
        RECT 148.230 83.640 148.400 93.050 ;
        RECT 148.760 93.050 152.790 93.220 ;
        RECT 148.760 88.000 148.930 93.050 ;
        RECT 149.560 92.540 150.060 92.710 ;
        RECT 149.330 91.830 149.500 92.370 ;
        RECT 150.120 91.830 150.290 92.370 ;
        RECT 149.560 91.490 150.060 91.660 ;
        RECT 149.330 90.780 149.500 91.320 ;
        RECT 150.120 90.780 150.290 91.320 ;
        RECT 149.560 90.440 150.060 90.610 ;
        RECT 149.330 89.730 149.500 90.270 ;
        RECT 150.120 89.730 150.290 90.270 ;
        RECT 149.560 89.390 150.060 89.560 ;
        RECT 149.330 88.680 149.500 89.220 ;
        RECT 150.120 88.680 150.290 89.220 ;
        RECT 149.560 88.340 150.060 88.510 ;
        RECT 150.690 88.000 150.860 93.050 ;
        RECT 151.490 92.540 151.990 92.710 ;
        RECT 151.260 91.830 151.430 92.370 ;
        RECT 152.050 91.830 152.220 92.370 ;
        RECT 151.490 91.490 151.990 91.660 ;
        RECT 151.260 90.780 151.430 91.320 ;
        RECT 152.050 90.780 152.220 91.320 ;
        RECT 151.490 90.440 151.990 90.610 ;
        RECT 151.260 89.730 151.430 90.270 ;
        RECT 152.050 89.730 152.220 90.270 ;
        RECT 151.490 89.390 151.990 89.560 ;
        RECT 151.260 88.680 151.430 89.220 ;
        RECT 152.050 88.680 152.220 89.220 ;
        RECT 151.490 88.340 151.990 88.510 ;
        RECT 152.620 88.000 152.790 93.050 ;
        RECT 148.760 87.830 152.790 88.000 ;
        RECT 153.130 93.000 153.300 93.210 ;
        RECT 156.460 93.085 156.630 93.210 ;
        RECT 153.130 92.670 154.185 93.000 ;
        RECT 153.130 92.070 153.300 92.670 ;
        RECT 154.355 92.585 154.835 93.085 ;
        RECT 155.035 92.755 158.055 93.085 ;
        RECT 154.355 92.500 156.195 92.585 ;
        RECT 153.565 92.255 156.195 92.500 ;
        RECT 153.565 92.240 154.835 92.255 ;
        RECT 153.130 91.740 154.185 92.070 ;
        RECT 153.130 91.070 153.300 91.740 ;
        RECT 154.355 91.570 154.835 92.240 ;
        RECT 156.460 92.085 156.630 92.755 ;
        RECT 158.255 92.585 158.735 93.085 ;
        RECT 159.790 93.000 159.960 93.210 ;
        RECT 158.905 92.670 159.960 93.000 ;
        RECT 156.895 92.500 158.735 92.585 ;
        RECT 156.895 92.255 159.525 92.500 ;
        RECT 158.255 92.240 159.525 92.255 ;
        RECT 155.035 91.755 158.055 92.085 ;
        RECT 153.565 91.555 154.835 91.570 ;
        RECT 153.565 91.385 156.195 91.555 ;
        RECT 153.565 91.310 154.525 91.385 ;
        RECT 153.565 91.240 154.395 91.310 ;
        RECT 153.130 90.740 154.055 91.070 ;
        RECT 153.130 90.210 153.300 90.740 ;
        RECT 154.225 90.560 154.395 91.240 ;
        RECT 153.565 90.390 154.395 90.560 ;
        RECT 153.130 89.880 154.055 90.210 ;
        RECT 153.130 89.270 153.300 89.880 ;
        RECT 154.225 89.700 154.395 90.390 ;
        RECT 153.565 89.450 154.395 89.700 ;
        RECT 154.565 89.450 154.995 91.140 ;
        RECT 155.165 90.735 155.335 91.385 ;
        RECT 156.460 91.185 156.630 91.755 ;
        RECT 158.255 91.570 158.735 92.240 ;
        RECT 159.790 92.070 159.960 92.670 ;
        RECT 158.905 91.740 159.960 92.070 ;
        RECT 158.255 91.555 159.525 91.570 ;
        RECT 156.895 91.385 159.525 91.555 ;
        RECT 155.505 90.935 157.585 91.185 ;
        RECT 155.165 90.405 156.195 90.735 ;
        RECT 155.165 89.705 155.335 90.405 ;
        RECT 156.460 90.235 156.630 90.935 ;
        RECT 157.755 90.735 157.925 91.385 ;
        RECT 158.565 91.310 159.525 91.385 ;
        RECT 158.695 91.240 159.525 91.310 ;
        RECT 156.895 90.405 157.925 90.735 ;
        RECT 155.505 89.905 157.585 90.235 ;
        RECT 155.165 89.455 156.195 89.705 ;
        RECT 153.130 89.020 154.345 89.270 ;
        RECT 153.130 88.680 153.300 89.020 ;
        RECT 154.630 88.765 154.830 89.450 ;
        RECT 156.460 89.255 156.630 89.905 ;
        RECT 157.755 89.705 157.925 90.405 ;
        RECT 156.895 89.455 157.925 89.705 ;
        RECT 158.095 89.450 158.525 91.140 ;
        RECT 158.695 90.560 158.865 91.240 ;
        RECT 159.790 91.070 159.960 91.740 ;
        RECT 159.035 90.740 159.960 91.070 ;
        RECT 158.695 90.390 159.525 90.560 ;
        RECT 158.695 89.700 158.865 90.390 ;
        RECT 159.790 90.210 159.960 90.740 ;
        RECT 159.035 89.880 159.960 90.210 ;
        RECT 158.695 89.450 159.525 89.700 ;
        RECT 155.035 89.005 158.055 89.255 ;
        RECT 156.460 88.765 156.630 89.005 ;
        RECT 158.260 88.765 158.460 89.450 ;
        RECT 159.790 89.270 159.960 89.880 ;
        RECT 158.745 89.020 159.960 89.270 ;
        RECT 153.130 88.350 154.185 88.680 ;
        RECT 144.370 83.470 148.400 83.640 ;
        RECT 153.130 87.750 153.300 88.350 ;
        RECT 154.355 88.265 154.835 88.765 ;
        RECT 155.035 88.435 158.055 88.765 ;
        RECT 154.355 88.180 156.195 88.265 ;
        RECT 153.565 87.935 156.195 88.180 ;
        RECT 153.565 87.920 154.835 87.935 ;
        RECT 153.130 87.420 154.185 87.750 ;
        RECT 153.130 86.750 153.300 87.420 ;
        RECT 154.355 87.250 154.835 87.920 ;
        RECT 156.460 87.765 156.630 88.435 ;
        RECT 158.255 88.265 158.735 88.765 ;
        RECT 159.790 88.680 159.960 89.020 ;
        RECT 158.905 88.350 159.960 88.680 ;
        RECT 156.895 88.180 158.735 88.265 ;
        RECT 156.895 87.935 159.525 88.180 ;
        RECT 158.255 87.920 159.525 87.935 ;
        RECT 155.035 87.435 158.055 87.765 ;
        RECT 153.565 87.235 154.835 87.250 ;
        RECT 153.565 87.065 156.195 87.235 ;
        RECT 153.565 86.990 154.525 87.065 ;
        RECT 153.565 86.920 154.395 86.990 ;
        RECT 153.130 86.420 154.055 86.750 ;
        RECT 153.130 85.890 153.300 86.420 ;
        RECT 154.225 86.240 154.395 86.920 ;
        RECT 153.565 86.070 154.395 86.240 ;
        RECT 153.130 85.560 154.055 85.890 ;
        RECT 153.130 84.950 153.300 85.560 ;
        RECT 154.225 85.380 154.395 86.070 ;
        RECT 153.565 85.130 154.395 85.380 ;
        RECT 154.565 85.130 154.995 86.820 ;
        RECT 155.165 86.415 155.335 87.065 ;
        RECT 156.460 86.865 156.630 87.435 ;
        RECT 158.255 87.250 158.735 87.920 ;
        RECT 159.790 87.750 159.960 88.350 ;
        RECT 161.000 93.045 163.100 93.215 ;
        RECT 161.000 87.995 161.170 93.045 ;
        RECT 161.800 92.535 162.300 92.705 ;
        RECT 161.570 91.825 161.740 92.365 ;
        RECT 162.360 91.825 162.530 92.365 ;
        RECT 161.800 91.485 162.300 91.655 ;
        RECT 161.570 90.775 161.740 91.315 ;
        RECT 162.360 90.775 162.530 91.315 ;
        RECT 161.800 90.435 162.300 90.605 ;
        RECT 161.570 89.725 161.740 90.265 ;
        RECT 162.360 89.725 162.530 90.265 ;
        RECT 161.800 89.385 162.300 89.555 ;
        RECT 161.570 88.675 161.740 89.215 ;
        RECT 162.360 88.675 162.530 89.215 ;
        RECT 161.800 88.335 162.300 88.505 ;
        RECT 162.930 87.995 163.100 93.045 ;
        RECT 161.000 87.825 163.100 87.995 ;
        RECT 163.460 93.045 165.560 93.215 ;
        RECT 158.905 87.420 159.960 87.750 ;
        RECT 158.255 87.235 159.525 87.250 ;
        RECT 156.895 87.065 159.525 87.235 ;
        RECT 155.505 86.615 157.585 86.865 ;
        RECT 155.165 86.085 156.195 86.415 ;
        RECT 155.165 85.385 155.335 86.085 ;
        RECT 156.460 85.915 156.630 86.615 ;
        RECT 157.755 86.415 157.925 87.065 ;
        RECT 158.565 86.990 159.525 87.065 ;
        RECT 158.695 86.920 159.525 86.990 ;
        RECT 156.895 86.085 157.925 86.415 ;
        RECT 155.505 85.585 157.585 85.915 ;
        RECT 155.165 85.135 156.195 85.385 ;
        RECT 153.130 84.700 154.345 84.950 ;
        RECT 153.130 84.480 153.300 84.700 ;
        RECT 153.130 84.180 154.320 84.480 ;
        RECT 153.130 83.975 153.300 84.180 ;
        RECT 153.130 83.645 154.055 83.975 ;
        RECT 154.630 83.965 154.830 85.130 ;
        RECT 156.460 84.935 156.630 85.585 ;
        RECT 157.755 85.385 157.925 86.085 ;
        RECT 156.895 85.135 157.925 85.385 ;
        RECT 158.095 85.130 158.525 86.820 ;
        RECT 158.695 86.240 158.865 86.920 ;
        RECT 159.790 86.750 159.960 87.420 ;
        RECT 159.035 86.420 159.960 86.750 ;
        RECT 158.695 86.070 159.525 86.240 ;
        RECT 158.695 85.380 158.865 86.070 ;
        RECT 159.790 85.890 159.960 86.420 ;
        RECT 159.035 85.560 159.960 85.890 ;
        RECT 158.695 85.130 159.525 85.380 ;
        RECT 155.035 84.685 158.055 84.935 ;
        RECT 156.460 84.480 156.630 84.685 ;
        RECT 155.420 84.180 157.670 84.480 ;
        RECT 156.460 83.970 156.630 84.180 ;
        RECT 154.225 83.735 155.335 83.965 ;
        RECT 141.910 77.720 144.010 77.890 ;
        RECT 153.130 83.065 153.300 83.645 ;
        RECT 154.225 83.465 154.395 83.735 ;
        RECT 155.165 83.520 155.335 83.735 ;
        RECT 155.505 83.720 157.585 83.970 ;
        RECT 158.265 83.965 158.465 85.130 ;
        RECT 159.790 84.950 159.960 85.560 ;
        RECT 158.745 84.700 159.960 84.950 ;
        RECT 159.790 84.480 159.960 84.700 ;
        RECT 158.770 84.180 159.960 84.480 ;
        RECT 159.790 83.975 159.960 84.180 ;
        RECT 157.755 83.735 158.865 83.965 ;
        RECT 153.565 83.295 154.395 83.465 ;
        RECT 153.130 82.735 154.055 83.065 ;
        RECT 153.130 82.135 153.300 82.735 ;
        RECT 154.225 82.555 154.395 83.295 ;
        RECT 153.565 82.305 154.395 82.555 ;
        RECT 153.130 81.805 154.345 82.135 ;
        RECT 154.565 81.815 154.995 83.490 ;
        RECT 155.165 83.190 156.195 83.520 ;
        RECT 155.165 82.620 155.335 83.190 ;
        RECT 156.460 82.990 156.630 83.720 ;
        RECT 157.755 83.520 157.925 83.735 ;
        RECT 156.895 83.190 157.925 83.520 ;
        RECT 155.505 82.820 157.585 82.990 ;
        RECT 155.165 82.290 156.195 82.620 ;
        RECT 156.460 82.090 156.630 82.820 ;
        RECT 157.755 82.620 157.925 83.190 ;
        RECT 156.895 82.290 157.925 82.620 ;
        RECT 155.165 81.840 157.925 82.090 ;
        RECT 153.130 81.065 153.300 81.805 ;
        RECT 154.630 81.565 154.830 81.815 ;
        RECT 153.565 81.235 156.195 81.565 ;
        RECT 156.460 81.065 156.630 81.840 ;
        RECT 158.095 81.815 158.525 83.490 ;
        RECT 158.695 83.465 158.865 83.735 ;
        RECT 159.035 83.645 159.960 83.975 ;
        RECT 158.695 83.295 159.525 83.465 ;
        RECT 158.695 82.555 158.865 83.295 ;
        RECT 159.790 83.065 159.960 83.645 ;
        RECT 159.035 82.735 159.960 83.065 ;
        RECT 158.695 82.305 159.525 82.555 ;
        RECT 159.790 82.135 159.960 82.735 ;
        RECT 158.260 81.565 158.460 81.815 ;
        RECT 158.745 81.805 159.960 82.135 ;
        RECT 156.895 81.235 159.525 81.565 ;
        RECT 159.790 81.065 159.960 81.805 ;
        RECT 153.130 80.735 154.345 81.065 ;
        RECT 153.130 80.160 153.300 80.735 ;
        RECT 154.515 80.375 154.995 81.065 ;
        RECT 155.165 80.735 157.925 81.065 ;
        RECT 153.130 79.860 154.320 80.160 ;
        RECT 153.130 79.145 153.300 79.860 ;
        RECT 154.580 79.645 154.780 80.375 ;
        RECT 156.460 80.160 156.630 80.735 ;
        RECT 158.095 80.375 158.575 81.065 ;
        RECT 158.745 80.735 159.960 81.065 ;
        RECT 155.420 79.860 157.670 80.160 ;
        RECT 153.565 79.315 156.195 79.645 ;
        RECT 156.460 79.145 156.630 79.860 ;
        RECT 158.310 79.645 158.510 80.375 ;
        RECT 159.790 80.160 159.960 80.735 ;
        RECT 158.770 79.860 159.960 80.160 ;
        RECT 156.895 79.315 159.525 79.645 ;
        RECT 159.790 79.145 159.960 79.860 ;
        RECT 153.130 78.815 154.345 79.145 ;
        RECT 153.130 77.350 153.300 78.815 ;
        RECT 154.515 78.455 154.995 79.145 ;
        RECT 155.165 78.815 157.925 79.145 ;
        RECT 156.460 78.225 156.630 78.815 ;
        RECT 158.095 78.455 158.575 79.145 ;
        RECT 158.745 78.815 159.960 79.145 ;
        RECT 153.565 77.840 154.225 78.170 ;
        RECT 154.395 77.895 154.765 78.225 ;
        RECT 155.035 77.895 158.055 78.225 ;
        RECT 158.325 77.895 158.695 78.225 ;
        RECT 159.790 78.200 159.960 78.815 ;
        RECT 154.055 77.725 154.225 77.840 ;
        RECT 154.055 77.555 156.195 77.725 ;
        RECT 154.395 77.495 156.195 77.555 ;
        RECT 153.130 77.020 154.225 77.350 ;
        RECT 156.460 77.325 156.630 77.895 ;
        RECT 158.865 77.870 159.960 78.200 ;
        RECT 156.895 77.665 158.695 77.725 ;
        RECT 156.895 77.495 159.035 77.665 ;
        RECT 158.865 77.380 159.035 77.495 ;
        RECT 129.120 75.935 130.335 76.265 ;
        RECT 129.120 75.450 129.290 75.935 ;
        RECT 130.505 75.575 130.985 76.265 ;
        RECT 131.155 75.935 132.620 76.265 ;
        RECT 132.450 75.450 132.620 75.935 ;
        RECT 153.130 76.265 153.300 77.020 ;
        RECT 154.395 76.995 154.765 77.325 ;
        RECT 155.035 76.995 158.055 77.325 ;
        RECT 158.325 76.995 158.695 77.325 ;
        RECT 158.865 77.050 159.525 77.380 ;
        RECT 154.500 76.765 154.700 76.995 ;
        RECT 153.565 76.435 156.195 76.765 ;
        RECT 156.460 76.265 156.630 76.995 ;
        RECT 159.790 76.890 159.960 77.870 ;
        RECT 161.000 87.295 163.100 87.465 ;
        RECT 161.000 77.885 161.170 87.295 ;
        RECT 161.800 86.785 162.300 86.955 ;
        RECT 161.570 85.030 161.740 86.570 ;
        RECT 162.360 85.030 162.530 86.570 ;
        RECT 161.800 84.645 162.300 84.815 ;
        RECT 161.570 82.890 161.740 84.430 ;
        RECT 162.360 82.890 162.530 84.430 ;
        RECT 161.800 82.505 162.300 82.675 ;
        RECT 161.570 80.750 161.740 82.290 ;
        RECT 162.360 80.750 162.530 82.290 ;
        RECT 161.800 80.365 162.300 80.535 ;
        RECT 161.570 78.610 161.740 80.150 ;
        RECT 162.360 78.610 162.530 80.150 ;
        RECT 161.800 78.225 162.300 78.395 ;
        RECT 162.930 77.885 163.100 87.295 ;
        RECT 163.460 83.635 163.630 93.045 ;
        RECT 164.260 92.535 164.760 92.705 ;
        RECT 164.030 90.780 164.200 92.320 ;
        RECT 164.820 90.780 164.990 92.320 ;
        RECT 164.260 90.395 164.760 90.565 ;
        RECT 164.030 88.640 164.200 90.180 ;
        RECT 164.820 88.640 164.990 90.180 ;
        RECT 164.260 88.255 164.760 88.425 ;
        RECT 164.030 86.500 164.200 88.040 ;
        RECT 164.820 86.500 164.990 88.040 ;
        RECT 164.260 86.115 164.760 86.285 ;
        RECT 164.030 84.360 164.200 85.900 ;
        RECT 164.820 84.360 164.990 85.900 ;
        RECT 164.260 83.975 164.760 84.145 ;
        RECT 165.390 83.635 165.560 93.045 ;
        RECT 165.920 93.050 168.020 93.220 ;
        RECT 165.920 88.000 166.090 93.050 ;
        RECT 166.720 92.540 167.220 92.710 ;
        RECT 166.490 91.830 166.660 92.370 ;
        RECT 167.280 91.830 167.450 92.370 ;
        RECT 166.720 91.490 167.220 91.660 ;
        RECT 166.490 90.780 166.660 91.320 ;
        RECT 167.280 90.780 167.450 91.320 ;
        RECT 166.720 90.440 167.220 90.610 ;
        RECT 166.490 89.730 166.660 90.270 ;
        RECT 167.280 89.730 167.450 90.270 ;
        RECT 166.720 89.390 167.220 89.560 ;
        RECT 166.490 88.680 166.660 89.220 ;
        RECT 167.280 88.680 167.450 89.220 ;
        RECT 166.720 88.340 167.220 88.510 ;
        RECT 167.850 88.000 168.020 93.050 ;
        RECT 165.920 87.830 168.020 88.000 ;
        RECT 168.380 93.050 172.410 93.220 ;
        RECT 163.460 83.465 165.560 83.635 ;
        RECT 165.920 87.300 168.020 87.470 ;
        RECT 161.000 77.715 163.100 77.885 ;
        RECT 163.460 82.935 165.560 83.105 ;
        RECT 163.460 77.885 163.630 82.935 ;
        RECT 164.260 82.425 164.760 82.595 ;
        RECT 164.030 81.715 164.200 82.255 ;
        RECT 164.820 81.715 164.990 82.255 ;
        RECT 164.260 81.375 164.760 81.545 ;
        RECT 164.030 80.665 164.200 81.205 ;
        RECT 164.820 80.665 164.990 81.205 ;
        RECT 164.260 80.325 164.760 80.495 ;
        RECT 164.030 79.615 164.200 80.155 ;
        RECT 164.820 79.615 164.990 80.155 ;
        RECT 164.260 79.275 164.760 79.445 ;
        RECT 164.030 78.565 164.200 79.105 ;
        RECT 164.820 78.565 164.990 79.105 ;
        RECT 164.260 78.225 164.760 78.395 ;
        RECT 165.390 77.885 165.560 82.935 ;
        RECT 163.460 77.715 165.560 77.885 ;
        RECT 165.920 77.890 166.090 87.300 ;
        RECT 166.720 86.790 167.220 86.960 ;
        RECT 166.490 85.035 166.660 86.575 ;
        RECT 167.280 85.035 167.450 86.575 ;
        RECT 166.720 84.650 167.220 84.820 ;
        RECT 166.490 82.895 166.660 84.435 ;
        RECT 167.280 82.895 167.450 84.435 ;
        RECT 166.720 82.510 167.220 82.680 ;
        RECT 166.490 80.755 166.660 82.295 ;
        RECT 167.280 80.755 167.450 82.295 ;
        RECT 166.720 80.370 167.220 80.540 ;
        RECT 166.490 78.615 166.660 80.155 ;
        RECT 167.280 78.615 167.450 80.155 ;
        RECT 166.720 78.230 167.220 78.400 ;
        RECT 167.850 77.890 168.020 87.300 ;
        RECT 168.380 83.640 168.550 93.050 ;
        RECT 169.180 92.540 169.680 92.710 ;
        RECT 168.950 90.785 169.120 92.325 ;
        RECT 169.740 90.785 169.910 92.325 ;
        RECT 169.180 90.400 169.680 90.570 ;
        RECT 168.950 88.645 169.120 90.185 ;
        RECT 169.740 88.645 169.910 90.185 ;
        RECT 169.180 88.260 169.680 88.430 ;
        RECT 168.950 86.505 169.120 88.045 ;
        RECT 169.740 86.505 169.910 88.045 ;
        RECT 169.180 86.120 169.680 86.290 ;
        RECT 168.950 84.365 169.120 85.905 ;
        RECT 169.740 84.365 169.910 85.905 ;
        RECT 169.180 83.980 169.680 84.150 ;
        RECT 170.310 83.640 170.480 93.050 ;
        RECT 171.110 92.540 171.610 92.710 ;
        RECT 170.880 90.785 171.050 92.325 ;
        RECT 171.670 90.785 171.840 92.325 ;
        RECT 171.110 90.400 171.610 90.570 ;
        RECT 170.880 88.645 171.050 90.185 ;
        RECT 171.670 88.645 171.840 90.185 ;
        RECT 171.110 88.260 171.610 88.430 ;
        RECT 170.880 86.505 171.050 88.045 ;
        RECT 171.670 86.505 171.840 88.045 ;
        RECT 171.110 86.120 171.610 86.290 ;
        RECT 170.880 84.365 171.050 85.905 ;
        RECT 171.670 84.365 171.840 85.905 ;
        RECT 171.110 83.980 171.610 84.150 ;
        RECT 172.240 83.640 172.410 93.050 ;
        RECT 172.770 93.050 176.800 93.220 ;
        RECT 172.770 88.000 172.940 93.050 ;
        RECT 173.570 92.540 174.070 92.710 ;
        RECT 173.340 91.830 173.510 92.370 ;
        RECT 174.130 91.830 174.300 92.370 ;
        RECT 173.570 91.490 174.070 91.660 ;
        RECT 173.340 90.780 173.510 91.320 ;
        RECT 174.130 90.780 174.300 91.320 ;
        RECT 173.570 90.440 174.070 90.610 ;
        RECT 173.340 89.730 173.510 90.270 ;
        RECT 174.130 89.730 174.300 90.270 ;
        RECT 173.570 89.390 174.070 89.560 ;
        RECT 173.340 88.680 173.510 89.220 ;
        RECT 174.130 88.680 174.300 89.220 ;
        RECT 173.570 88.340 174.070 88.510 ;
        RECT 174.700 88.000 174.870 93.050 ;
        RECT 175.500 92.540 176.000 92.710 ;
        RECT 175.270 91.830 175.440 92.370 ;
        RECT 176.060 91.830 176.230 92.370 ;
        RECT 175.500 91.490 176.000 91.660 ;
        RECT 175.270 90.780 175.440 91.320 ;
        RECT 176.060 90.780 176.230 91.320 ;
        RECT 175.500 90.440 176.000 90.610 ;
        RECT 175.270 89.730 175.440 90.270 ;
        RECT 176.060 89.730 176.230 90.270 ;
        RECT 175.500 89.390 176.000 89.560 ;
        RECT 175.270 88.680 175.440 89.220 ;
        RECT 176.060 88.680 176.230 89.220 ;
        RECT 175.500 88.340 176.000 88.510 ;
        RECT 176.630 88.000 176.800 93.050 ;
        RECT 172.770 87.830 176.800 88.000 ;
        RECT 177.140 93.000 177.310 93.210 ;
        RECT 180.470 93.085 180.640 93.210 ;
        RECT 177.140 92.670 178.195 93.000 ;
        RECT 177.140 92.070 177.310 92.670 ;
        RECT 178.365 92.585 178.845 93.085 ;
        RECT 179.045 92.755 182.065 93.085 ;
        RECT 178.365 92.500 180.205 92.585 ;
        RECT 177.575 92.255 180.205 92.500 ;
        RECT 177.575 92.240 178.845 92.255 ;
        RECT 177.140 91.740 178.195 92.070 ;
        RECT 177.140 91.070 177.310 91.740 ;
        RECT 178.365 91.570 178.845 92.240 ;
        RECT 180.470 92.085 180.640 92.755 ;
        RECT 182.265 92.585 182.745 93.085 ;
        RECT 183.800 93.000 183.970 93.210 ;
        RECT 182.915 92.670 183.970 93.000 ;
        RECT 180.905 92.500 182.745 92.585 ;
        RECT 180.905 92.255 183.535 92.500 ;
        RECT 182.265 92.240 183.535 92.255 ;
        RECT 179.045 91.755 182.065 92.085 ;
        RECT 177.575 91.555 178.845 91.570 ;
        RECT 177.575 91.385 180.205 91.555 ;
        RECT 177.575 91.310 178.535 91.385 ;
        RECT 177.575 91.240 178.405 91.310 ;
        RECT 177.140 90.740 178.065 91.070 ;
        RECT 177.140 90.210 177.310 90.740 ;
        RECT 178.235 90.560 178.405 91.240 ;
        RECT 177.575 90.390 178.405 90.560 ;
        RECT 177.140 89.880 178.065 90.210 ;
        RECT 177.140 89.270 177.310 89.880 ;
        RECT 178.235 89.700 178.405 90.390 ;
        RECT 177.575 89.450 178.405 89.700 ;
        RECT 178.575 89.450 179.005 91.140 ;
        RECT 179.175 90.735 179.345 91.385 ;
        RECT 180.470 91.185 180.640 91.755 ;
        RECT 182.265 91.570 182.745 92.240 ;
        RECT 183.800 92.070 183.970 92.670 ;
        RECT 182.915 91.740 183.970 92.070 ;
        RECT 182.265 91.555 183.535 91.570 ;
        RECT 180.905 91.385 183.535 91.555 ;
        RECT 179.515 90.935 181.595 91.185 ;
        RECT 179.175 90.405 180.205 90.735 ;
        RECT 179.175 89.705 179.345 90.405 ;
        RECT 180.470 90.235 180.640 90.935 ;
        RECT 181.765 90.735 181.935 91.385 ;
        RECT 182.575 91.310 183.535 91.385 ;
        RECT 182.705 91.240 183.535 91.310 ;
        RECT 180.905 90.405 181.935 90.735 ;
        RECT 179.515 89.905 181.595 90.235 ;
        RECT 179.175 89.455 180.205 89.705 ;
        RECT 177.140 89.020 178.355 89.270 ;
        RECT 177.140 88.680 177.310 89.020 ;
        RECT 178.640 88.765 178.840 89.450 ;
        RECT 180.470 89.255 180.640 89.905 ;
        RECT 181.765 89.705 181.935 90.405 ;
        RECT 180.905 89.455 181.935 89.705 ;
        RECT 182.105 89.450 182.535 91.140 ;
        RECT 182.705 90.560 182.875 91.240 ;
        RECT 183.800 91.070 183.970 91.740 ;
        RECT 183.045 90.740 183.970 91.070 ;
        RECT 182.705 90.390 183.535 90.560 ;
        RECT 182.705 89.700 182.875 90.390 ;
        RECT 183.800 90.210 183.970 90.740 ;
        RECT 183.045 89.880 183.970 90.210 ;
        RECT 182.705 89.450 183.535 89.700 ;
        RECT 179.045 89.005 182.065 89.255 ;
        RECT 180.470 88.765 180.640 89.005 ;
        RECT 182.270 88.765 182.470 89.450 ;
        RECT 183.800 89.270 183.970 89.880 ;
        RECT 182.755 89.020 183.970 89.270 ;
        RECT 177.140 88.350 178.195 88.680 ;
        RECT 168.380 83.470 172.410 83.640 ;
        RECT 177.140 87.750 177.310 88.350 ;
        RECT 178.365 88.265 178.845 88.765 ;
        RECT 179.045 88.435 182.065 88.765 ;
        RECT 178.365 88.180 180.205 88.265 ;
        RECT 177.575 87.935 180.205 88.180 ;
        RECT 177.575 87.920 178.845 87.935 ;
        RECT 177.140 87.420 178.195 87.750 ;
        RECT 177.140 86.750 177.310 87.420 ;
        RECT 178.365 87.250 178.845 87.920 ;
        RECT 180.470 87.765 180.640 88.435 ;
        RECT 182.265 88.265 182.745 88.765 ;
        RECT 183.800 88.680 183.970 89.020 ;
        RECT 182.915 88.350 183.970 88.680 ;
        RECT 180.905 88.180 182.745 88.265 ;
        RECT 180.905 87.935 183.535 88.180 ;
        RECT 182.265 87.920 183.535 87.935 ;
        RECT 179.045 87.435 182.065 87.765 ;
        RECT 177.575 87.235 178.845 87.250 ;
        RECT 177.575 87.065 180.205 87.235 ;
        RECT 177.575 86.990 178.535 87.065 ;
        RECT 177.575 86.920 178.405 86.990 ;
        RECT 177.140 86.420 178.065 86.750 ;
        RECT 177.140 85.890 177.310 86.420 ;
        RECT 178.235 86.240 178.405 86.920 ;
        RECT 177.575 86.070 178.405 86.240 ;
        RECT 177.140 85.560 178.065 85.890 ;
        RECT 177.140 84.950 177.310 85.560 ;
        RECT 178.235 85.380 178.405 86.070 ;
        RECT 177.575 85.130 178.405 85.380 ;
        RECT 178.575 85.130 179.005 86.820 ;
        RECT 179.175 86.415 179.345 87.065 ;
        RECT 180.470 86.865 180.640 87.435 ;
        RECT 182.265 87.250 182.745 87.920 ;
        RECT 183.800 87.750 183.970 88.350 ;
        RECT 185.010 93.045 187.110 93.215 ;
        RECT 185.010 87.995 185.180 93.045 ;
        RECT 185.810 92.535 186.310 92.705 ;
        RECT 185.580 91.825 185.750 92.365 ;
        RECT 186.370 91.825 186.540 92.365 ;
        RECT 185.810 91.485 186.310 91.655 ;
        RECT 185.580 90.775 185.750 91.315 ;
        RECT 186.370 90.775 186.540 91.315 ;
        RECT 185.810 90.435 186.310 90.605 ;
        RECT 185.580 89.725 185.750 90.265 ;
        RECT 186.370 89.725 186.540 90.265 ;
        RECT 185.810 89.385 186.310 89.555 ;
        RECT 185.580 88.675 185.750 89.215 ;
        RECT 186.370 88.675 186.540 89.215 ;
        RECT 185.810 88.335 186.310 88.505 ;
        RECT 186.940 87.995 187.110 93.045 ;
        RECT 185.010 87.825 187.110 87.995 ;
        RECT 187.470 93.045 189.570 93.215 ;
        RECT 182.915 87.420 183.970 87.750 ;
        RECT 182.265 87.235 183.535 87.250 ;
        RECT 180.905 87.065 183.535 87.235 ;
        RECT 179.515 86.615 181.595 86.865 ;
        RECT 179.175 86.085 180.205 86.415 ;
        RECT 179.175 85.385 179.345 86.085 ;
        RECT 180.470 85.915 180.640 86.615 ;
        RECT 181.765 86.415 181.935 87.065 ;
        RECT 182.575 86.990 183.535 87.065 ;
        RECT 182.705 86.920 183.535 86.990 ;
        RECT 180.905 86.085 181.935 86.415 ;
        RECT 179.515 85.585 181.595 85.915 ;
        RECT 179.175 85.135 180.205 85.385 ;
        RECT 177.140 84.700 178.355 84.950 ;
        RECT 177.140 84.480 177.310 84.700 ;
        RECT 177.140 84.180 178.330 84.480 ;
        RECT 177.140 83.975 177.310 84.180 ;
        RECT 177.140 83.645 178.065 83.975 ;
        RECT 178.640 83.965 178.840 85.130 ;
        RECT 180.470 84.935 180.640 85.585 ;
        RECT 181.765 85.385 181.935 86.085 ;
        RECT 180.905 85.135 181.935 85.385 ;
        RECT 182.105 85.130 182.535 86.820 ;
        RECT 182.705 86.240 182.875 86.920 ;
        RECT 183.800 86.750 183.970 87.420 ;
        RECT 183.045 86.420 183.970 86.750 ;
        RECT 182.705 86.070 183.535 86.240 ;
        RECT 182.705 85.380 182.875 86.070 ;
        RECT 183.800 85.890 183.970 86.420 ;
        RECT 183.045 85.560 183.970 85.890 ;
        RECT 182.705 85.130 183.535 85.380 ;
        RECT 179.045 84.685 182.065 84.935 ;
        RECT 180.470 84.480 180.640 84.685 ;
        RECT 179.430 84.180 181.680 84.480 ;
        RECT 180.470 83.970 180.640 84.180 ;
        RECT 178.235 83.735 179.345 83.965 ;
        RECT 165.920 77.720 168.020 77.890 ;
        RECT 177.140 83.065 177.310 83.645 ;
        RECT 178.235 83.465 178.405 83.735 ;
        RECT 179.175 83.520 179.345 83.735 ;
        RECT 179.515 83.720 181.595 83.970 ;
        RECT 182.275 83.965 182.475 85.130 ;
        RECT 183.800 84.950 183.970 85.560 ;
        RECT 182.755 84.700 183.970 84.950 ;
        RECT 183.800 84.480 183.970 84.700 ;
        RECT 182.780 84.180 183.970 84.480 ;
        RECT 183.800 83.975 183.970 84.180 ;
        RECT 181.765 83.735 182.875 83.965 ;
        RECT 177.575 83.295 178.405 83.465 ;
        RECT 177.140 82.735 178.065 83.065 ;
        RECT 177.140 82.135 177.310 82.735 ;
        RECT 178.235 82.555 178.405 83.295 ;
        RECT 177.575 82.305 178.405 82.555 ;
        RECT 177.140 81.805 178.355 82.135 ;
        RECT 178.575 81.815 179.005 83.490 ;
        RECT 179.175 83.190 180.205 83.520 ;
        RECT 179.175 82.620 179.345 83.190 ;
        RECT 180.470 82.990 180.640 83.720 ;
        RECT 181.765 83.520 181.935 83.735 ;
        RECT 180.905 83.190 181.935 83.520 ;
        RECT 179.515 82.820 181.595 82.990 ;
        RECT 179.175 82.290 180.205 82.620 ;
        RECT 180.470 82.090 180.640 82.820 ;
        RECT 181.765 82.620 181.935 83.190 ;
        RECT 180.905 82.290 181.935 82.620 ;
        RECT 179.175 81.840 181.935 82.090 ;
        RECT 177.140 81.065 177.310 81.805 ;
        RECT 178.640 81.565 178.840 81.815 ;
        RECT 177.575 81.235 180.205 81.565 ;
        RECT 180.470 81.065 180.640 81.840 ;
        RECT 182.105 81.815 182.535 83.490 ;
        RECT 182.705 83.465 182.875 83.735 ;
        RECT 183.045 83.645 183.970 83.975 ;
        RECT 182.705 83.295 183.535 83.465 ;
        RECT 182.705 82.555 182.875 83.295 ;
        RECT 183.800 83.065 183.970 83.645 ;
        RECT 183.045 82.735 183.970 83.065 ;
        RECT 182.705 82.305 183.535 82.555 ;
        RECT 183.800 82.135 183.970 82.735 ;
        RECT 182.270 81.565 182.470 81.815 ;
        RECT 182.755 81.805 183.970 82.135 ;
        RECT 180.905 81.235 183.535 81.565 ;
        RECT 183.800 81.065 183.970 81.805 ;
        RECT 177.140 80.735 178.355 81.065 ;
        RECT 177.140 80.160 177.310 80.735 ;
        RECT 178.525 80.375 179.005 81.065 ;
        RECT 179.175 80.735 181.935 81.065 ;
        RECT 177.140 79.860 178.330 80.160 ;
        RECT 177.140 79.145 177.310 79.860 ;
        RECT 178.590 79.645 178.790 80.375 ;
        RECT 180.470 80.160 180.640 80.735 ;
        RECT 182.105 80.375 182.585 81.065 ;
        RECT 182.755 80.735 183.970 81.065 ;
        RECT 179.430 79.860 181.680 80.160 ;
        RECT 177.575 79.315 180.205 79.645 ;
        RECT 180.470 79.145 180.640 79.860 ;
        RECT 182.320 79.645 182.520 80.375 ;
        RECT 183.800 80.160 183.970 80.735 ;
        RECT 182.780 79.860 183.970 80.160 ;
        RECT 180.905 79.315 183.535 79.645 ;
        RECT 183.800 79.145 183.970 79.860 ;
        RECT 177.140 78.815 178.355 79.145 ;
        RECT 177.140 77.350 177.310 78.815 ;
        RECT 178.525 78.455 179.005 79.145 ;
        RECT 179.175 78.815 181.935 79.145 ;
        RECT 180.470 78.225 180.640 78.815 ;
        RECT 182.105 78.455 182.585 79.145 ;
        RECT 182.755 78.815 183.970 79.145 ;
        RECT 177.575 77.840 178.235 78.170 ;
        RECT 178.405 77.895 178.775 78.225 ;
        RECT 179.045 77.895 182.065 78.225 ;
        RECT 182.335 77.895 182.705 78.225 ;
        RECT 183.800 78.200 183.970 78.815 ;
        RECT 178.065 77.725 178.235 77.840 ;
        RECT 178.065 77.555 180.205 77.725 ;
        RECT 178.405 77.495 180.205 77.555 ;
        RECT 177.140 77.020 178.235 77.350 ;
        RECT 180.470 77.325 180.640 77.895 ;
        RECT 182.875 77.870 183.970 78.200 ;
        RECT 180.905 77.665 182.705 77.725 ;
        RECT 180.905 77.495 183.045 77.665 ;
        RECT 182.875 77.380 183.045 77.495 ;
        RECT 153.130 75.935 154.345 76.265 ;
        RECT 153.130 75.450 153.300 75.935 ;
        RECT 154.515 75.575 154.995 76.265 ;
        RECT 155.165 75.935 156.630 76.265 ;
        RECT 156.460 75.450 156.630 75.935 ;
        RECT 177.140 76.265 177.310 77.020 ;
        RECT 178.405 76.995 178.775 77.325 ;
        RECT 179.045 76.995 182.065 77.325 ;
        RECT 182.335 76.995 182.705 77.325 ;
        RECT 182.875 77.050 183.535 77.380 ;
        RECT 178.510 76.765 178.710 76.995 ;
        RECT 177.575 76.435 180.205 76.765 ;
        RECT 180.470 76.265 180.640 76.995 ;
        RECT 183.800 76.890 183.970 77.870 ;
        RECT 185.010 87.295 187.110 87.465 ;
        RECT 185.010 77.885 185.180 87.295 ;
        RECT 185.810 86.785 186.310 86.955 ;
        RECT 185.580 85.030 185.750 86.570 ;
        RECT 186.370 85.030 186.540 86.570 ;
        RECT 185.810 84.645 186.310 84.815 ;
        RECT 185.580 82.890 185.750 84.430 ;
        RECT 186.370 82.890 186.540 84.430 ;
        RECT 185.810 82.505 186.310 82.675 ;
        RECT 185.580 80.750 185.750 82.290 ;
        RECT 186.370 80.750 186.540 82.290 ;
        RECT 185.810 80.365 186.310 80.535 ;
        RECT 185.580 78.610 185.750 80.150 ;
        RECT 186.370 78.610 186.540 80.150 ;
        RECT 185.810 78.225 186.310 78.395 ;
        RECT 186.940 77.885 187.110 87.295 ;
        RECT 187.470 83.635 187.640 93.045 ;
        RECT 188.270 92.535 188.770 92.705 ;
        RECT 188.040 90.780 188.210 92.320 ;
        RECT 188.830 90.780 189.000 92.320 ;
        RECT 188.270 90.395 188.770 90.565 ;
        RECT 188.040 88.640 188.210 90.180 ;
        RECT 188.830 88.640 189.000 90.180 ;
        RECT 188.270 88.255 188.770 88.425 ;
        RECT 188.040 86.500 188.210 88.040 ;
        RECT 188.830 86.500 189.000 88.040 ;
        RECT 188.270 86.115 188.770 86.285 ;
        RECT 188.040 84.360 188.210 85.900 ;
        RECT 188.830 84.360 189.000 85.900 ;
        RECT 188.270 83.975 188.770 84.145 ;
        RECT 189.400 83.635 189.570 93.045 ;
        RECT 189.930 93.050 192.030 93.220 ;
        RECT 189.930 88.000 190.100 93.050 ;
        RECT 190.730 92.540 191.230 92.710 ;
        RECT 190.500 91.830 190.670 92.370 ;
        RECT 191.290 91.830 191.460 92.370 ;
        RECT 190.730 91.490 191.230 91.660 ;
        RECT 190.500 90.780 190.670 91.320 ;
        RECT 191.290 90.780 191.460 91.320 ;
        RECT 190.730 90.440 191.230 90.610 ;
        RECT 190.500 89.730 190.670 90.270 ;
        RECT 191.290 89.730 191.460 90.270 ;
        RECT 190.730 89.390 191.230 89.560 ;
        RECT 190.500 88.680 190.670 89.220 ;
        RECT 191.290 88.680 191.460 89.220 ;
        RECT 190.730 88.340 191.230 88.510 ;
        RECT 191.860 88.000 192.030 93.050 ;
        RECT 189.930 87.830 192.030 88.000 ;
        RECT 192.390 93.050 196.420 93.220 ;
        RECT 187.470 83.465 189.570 83.635 ;
        RECT 189.930 87.300 192.030 87.470 ;
        RECT 185.010 77.715 187.110 77.885 ;
        RECT 187.470 82.935 189.570 83.105 ;
        RECT 187.470 77.885 187.640 82.935 ;
        RECT 188.270 82.425 188.770 82.595 ;
        RECT 188.040 81.715 188.210 82.255 ;
        RECT 188.830 81.715 189.000 82.255 ;
        RECT 188.270 81.375 188.770 81.545 ;
        RECT 188.040 80.665 188.210 81.205 ;
        RECT 188.830 80.665 189.000 81.205 ;
        RECT 188.270 80.325 188.770 80.495 ;
        RECT 188.040 79.615 188.210 80.155 ;
        RECT 188.830 79.615 189.000 80.155 ;
        RECT 188.270 79.275 188.770 79.445 ;
        RECT 188.040 78.565 188.210 79.105 ;
        RECT 188.830 78.565 189.000 79.105 ;
        RECT 188.270 78.225 188.770 78.395 ;
        RECT 189.400 77.885 189.570 82.935 ;
        RECT 187.470 77.715 189.570 77.885 ;
        RECT 189.930 77.890 190.100 87.300 ;
        RECT 190.730 86.790 191.230 86.960 ;
        RECT 190.500 85.035 190.670 86.575 ;
        RECT 191.290 85.035 191.460 86.575 ;
        RECT 190.730 84.650 191.230 84.820 ;
        RECT 190.500 82.895 190.670 84.435 ;
        RECT 191.290 82.895 191.460 84.435 ;
        RECT 190.730 82.510 191.230 82.680 ;
        RECT 190.500 80.755 190.670 82.295 ;
        RECT 191.290 80.755 191.460 82.295 ;
        RECT 190.730 80.370 191.230 80.540 ;
        RECT 190.500 78.615 190.670 80.155 ;
        RECT 191.290 78.615 191.460 80.155 ;
        RECT 190.730 78.230 191.230 78.400 ;
        RECT 191.860 77.890 192.030 87.300 ;
        RECT 192.390 83.640 192.560 93.050 ;
        RECT 193.190 92.540 193.690 92.710 ;
        RECT 192.960 90.785 193.130 92.325 ;
        RECT 193.750 90.785 193.920 92.325 ;
        RECT 193.190 90.400 193.690 90.570 ;
        RECT 192.960 88.645 193.130 90.185 ;
        RECT 193.750 88.645 193.920 90.185 ;
        RECT 193.190 88.260 193.690 88.430 ;
        RECT 192.960 86.505 193.130 88.045 ;
        RECT 193.750 86.505 193.920 88.045 ;
        RECT 193.190 86.120 193.690 86.290 ;
        RECT 192.960 84.365 193.130 85.905 ;
        RECT 193.750 84.365 193.920 85.905 ;
        RECT 193.190 83.980 193.690 84.150 ;
        RECT 194.320 83.640 194.490 93.050 ;
        RECT 195.120 92.540 195.620 92.710 ;
        RECT 194.890 90.785 195.060 92.325 ;
        RECT 195.680 90.785 195.850 92.325 ;
        RECT 195.120 90.400 195.620 90.570 ;
        RECT 194.890 88.645 195.060 90.185 ;
        RECT 195.680 88.645 195.850 90.185 ;
        RECT 195.120 88.260 195.620 88.430 ;
        RECT 194.890 86.505 195.060 88.045 ;
        RECT 195.680 86.505 195.850 88.045 ;
        RECT 195.120 86.120 195.620 86.290 ;
        RECT 194.890 84.365 195.060 85.905 ;
        RECT 195.680 84.365 195.850 85.905 ;
        RECT 195.120 83.980 195.620 84.150 ;
        RECT 196.250 83.640 196.420 93.050 ;
        RECT 196.780 93.050 200.810 93.220 ;
        RECT 196.780 88.000 196.950 93.050 ;
        RECT 197.580 92.540 198.080 92.710 ;
        RECT 197.350 91.830 197.520 92.370 ;
        RECT 198.140 91.830 198.310 92.370 ;
        RECT 197.580 91.490 198.080 91.660 ;
        RECT 197.350 90.780 197.520 91.320 ;
        RECT 198.140 90.780 198.310 91.320 ;
        RECT 197.580 90.440 198.080 90.610 ;
        RECT 197.350 89.730 197.520 90.270 ;
        RECT 198.140 89.730 198.310 90.270 ;
        RECT 197.580 89.390 198.080 89.560 ;
        RECT 197.350 88.680 197.520 89.220 ;
        RECT 198.140 88.680 198.310 89.220 ;
        RECT 197.580 88.340 198.080 88.510 ;
        RECT 198.710 88.000 198.880 93.050 ;
        RECT 199.510 92.540 200.010 92.710 ;
        RECT 199.280 91.830 199.450 92.370 ;
        RECT 200.070 91.830 200.240 92.370 ;
        RECT 199.510 91.490 200.010 91.660 ;
        RECT 199.280 90.780 199.450 91.320 ;
        RECT 200.070 90.780 200.240 91.320 ;
        RECT 199.510 90.440 200.010 90.610 ;
        RECT 199.280 89.730 199.450 90.270 ;
        RECT 200.070 89.730 200.240 90.270 ;
        RECT 199.510 89.390 200.010 89.560 ;
        RECT 199.280 88.680 199.450 89.220 ;
        RECT 200.070 88.680 200.240 89.220 ;
        RECT 199.510 88.340 200.010 88.510 ;
        RECT 200.640 88.000 200.810 93.050 ;
        RECT 196.780 87.830 200.810 88.000 ;
        RECT 201.150 93.000 201.320 93.210 ;
        RECT 204.480 93.085 204.650 93.210 ;
        RECT 201.150 92.670 202.205 93.000 ;
        RECT 201.150 92.070 201.320 92.670 ;
        RECT 202.375 92.585 202.855 93.085 ;
        RECT 203.055 92.755 206.075 93.085 ;
        RECT 202.375 92.500 204.215 92.585 ;
        RECT 201.585 92.255 204.215 92.500 ;
        RECT 201.585 92.240 202.855 92.255 ;
        RECT 201.150 91.740 202.205 92.070 ;
        RECT 201.150 91.070 201.320 91.740 ;
        RECT 202.375 91.570 202.855 92.240 ;
        RECT 204.480 92.085 204.650 92.755 ;
        RECT 206.275 92.585 206.755 93.085 ;
        RECT 207.810 93.000 207.980 93.210 ;
        RECT 206.925 92.670 207.980 93.000 ;
        RECT 204.915 92.500 206.755 92.585 ;
        RECT 204.915 92.255 207.545 92.500 ;
        RECT 206.275 92.240 207.545 92.255 ;
        RECT 203.055 91.755 206.075 92.085 ;
        RECT 201.585 91.555 202.855 91.570 ;
        RECT 201.585 91.385 204.215 91.555 ;
        RECT 201.585 91.310 202.545 91.385 ;
        RECT 201.585 91.240 202.415 91.310 ;
        RECT 201.150 90.740 202.075 91.070 ;
        RECT 201.150 90.210 201.320 90.740 ;
        RECT 202.245 90.560 202.415 91.240 ;
        RECT 201.585 90.390 202.415 90.560 ;
        RECT 201.150 89.880 202.075 90.210 ;
        RECT 201.150 89.270 201.320 89.880 ;
        RECT 202.245 89.700 202.415 90.390 ;
        RECT 201.585 89.450 202.415 89.700 ;
        RECT 202.585 89.450 203.015 91.140 ;
        RECT 203.185 90.735 203.355 91.385 ;
        RECT 204.480 91.185 204.650 91.755 ;
        RECT 206.275 91.570 206.755 92.240 ;
        RECT 207.810 92.070 207.980 92.670 ;
        RECT 206.925 91.740 207.980 92.070 ;
        RECT 206.275 91.555 207.545 91.570 ;
        RECT 204.915 91.385 207.545 91.555 ;
        RECT 203.525 90.935 205.605 91.185 ;
        RECT 203.185 90.405 204.215 90.735 ;
        RECT 203.185 89.705 203.355 90.405 ;
        RECT 204.480 90.235 204.650 90.935 ;
        RECT 205.775 90.735 205.945 91.385 ;
        RECT 206.585 91.310 207.545 91.385 ;
        RECT 206.715 91.240 207.545 91.310 ;
        RECT 204.915 90.405 205.945 90.735 ;
        RECT 203.525 89.905 205.605 90.235 ;
        RECT 203.185 89.455 204.215 89.705 ;
        RECT 201.150 89.020 202.365 89.270 ;
        RECT 201.150 88.680 201.320 89.020 ;
        RECT 202.650 88.765 202.850 89.450 ;
        RECT 204.480 89.255 204.650 89.905 ;
        RECT 205.775 89.705 205.945 90.405 ;
        RECT 204.915 89.455 205.945 89.705 ;
        RECT 206.115 89.450 206.545 91.140 ;
        RECT 206.715 90.560 206.885 91.240 ;
        RECT 207.810 91.070 207.980 91.740 ;
        RECT 207.055 90.740 207.980 91.070 ;
        RECT 206.715 90.390 207.545 90.560 ;
        RECT 206.715 89.700 206.885 90.390 ;
        RECT 207.810 90.210 207.980 90.740 ;
        RECT 207.055 89.880 207.980 90.210 ;
        RECT 206.715 89.450 207.545 89.700 ;
        RECT 203.055 89.005 206.075 89.255 ;
        RECT 204.480 88.765 204.650 89.005 ;
        RECT 206.280 88.765 206.480 89.450 ;
        RECT 207.810 89.270 207.980 89.880 ;
        RECT 206.765 89.020 207.980 89.270 ;
        RECT 201.150 88.350 202.205 88.680 ;
        RECT 192.390 83.470 196.420 83.640 ;
        RECT 201.150 87.750 201.320 88.350 ;
        RECT 202.375 88.265 202.855 88.765 ;
        RECT 203.055 88.435 206.075 88.765 ;
        RECT 202.375 88.180 204.215 88.265 ;
        RECT 201.585 87.935 204.215 88.180 ;
        RECT 201.585 87.920 202.855 87.935 ;
        RECT 201.150 87.420 202.205 87.750 ;
        RECT 201.150 86.750 201.320 87.420 ;
        RECT 202.375 87.250 202.855 87.920 ;
        RECT 204.480 87.765 204.650 88.435 ;
        RECT 206.275 88.265 206.755 88.765 ;
        RECT 207.810 88.680 207.980 89.020 ;
        RECT 206.925 88.350 207.980 88.680 ;
        RECT 204.915 88.180 206.755 88.265 ;
        RECT 204.915 87.935 207.545 88.180 ;
        RECT 206.275 87.920 207.545 87.935 ;
        RECT 203.055 87.435 206.075 87.765 ;
        RECT 201.585 87.235 202.855 87.250 ;
        RECT 201.585 87.065 204.215 87.235 ;
        RECT 201.585 86.990 202.545 87.065 ;
        RECT 201.585 86.920 202.415 86.990 ;
        RECT 201.150 86.420 202.075 86.750 ;
        RECT 201.150 85.890 201.320 86.420 ;
        RECT 202.245 86.240 202.415 86.920 ;
        RECT 201.585 86.070 202.415 86.240 ;
        RECT 201.150 85.560 202.075 85.890 ;
        RECT 201.150 84.950 201.320 85.560 ;
        RECT 202.245 85.380 202.415 86.070 ;
        RECT 201.585 85.130 202.415 85.380 ;
        RECT 202.585 85.130 203.015 86.820 ;
        RECT 203.185 86.415 203.355 87.065 ;
        RECT 204.480 86.865 204.650 87.435 ;
        RECT 206.275 87.250 206.755 87.920 ;
        RECT 207.810 87.750 207.980 88.350 ;
        RECT 209.020 93.045 211.120 93.215 ;
        RECT 209.020 87.995 209.190 93.045 ;
        RECT 209.820 92.535 210.320 92.705 ;
        RECT 209.590 91.825 209.760 92.365 ;
        RECT 210.380 91.825 210.550 92.365 ;
        RECT 209.820 91.485 210.320 91.655 ;
        RECT 209.590 90.775 209.760 91.315 ;
        RECT 210.380 90.775 210.550 91.315 ;
        RECT 209.820 90.435 210.320 90.605 ;
        RECT 209.590 89.725 209.760 90.265 ;
        RECT 210.380 89.725 210.550 90.265 ;
        RECT 209.820 89.385 210.320 89.555 ;
        RECT 209.590 88.675 209.760 89.215 ;
        RECT 210.380 88.675 210.550 89.215 ;
        RECT 209.820 88.335 210.320 88.505 ;
        RECT 210.950 87.995 211.120 93.045 ;
        RECT 209.020 87.825 211.120 87.995 ;
        RECT 211.480 93.045 213.580 93.215 ;
        RECT 206.925 87.420 207.980 87.750 ;
        RECT 206.275 87.235 207.545 87.250 ;
        RECT 204.915 87.065 207.545 87.235 ;
        RECT 203.525 86.615 205.605 86.865 ;
        RECT 203.185 86.085 204.215 86.415 ;
        RECT 203.185 85.385 203.355 86.085 ;
        RECT 204.480 85.915 204.650 86.615 ;
        RECT 205.775 86.415 205.945 87.065 ;
        RECT 206.585 86.990 207.545 87.065 ;
        RECT 206.715 86.920 207.545 86.990 ;
        RECT 204.915 86.085 205.945 86.415 ;
        RECT 203.525 85.585 205.605 85.915 ;
        RECT 203.185 85.135 204.215 85.385 ;
        RECT 201.150 84.700 202.365 84.950 ;
        RECT 201.150 84.480 201.320 84.700 ;
        RECT 201.150 84.180 202.340 84.480 ;
        RECT 201.150 83.975 201.320 84.180 ;
        RECT 201.150 83.645 202.075 83.975 ;
        RECT 202.650 83.965 202.850 85.130 ;
        RECT 204.480 84.935 204.650 85.585 ;
        RECT 205.775 85.385 205.945 86.085 ;
        RECT 204.915 85.135 205.945 85.385 ;
        RECT 206.115 85.130 206.545 86.820 ;
        RECT 206.715 86.240 206.885 86.920 ;
        RECT 207.810 86.750 207.980 87.420 ;
        RECT 207.055 86.420 207.980 86.750 ;
        RECT 206.715 86.070 207.545 86.240 ;
        RECT 206.715 85.380 206.885 86.070 ;
        RECT 207.810 85.890 207.980 86.420 ;
        RECT 207.055 85.560 207.980 85.890 ;
        RECT 206.715 85.130 207.545 85.380 ;
        RECT 203.055 84.685 206.075 84.935 ;
        RECT 204.480 84.480 204.650 84.685 ;
        RECT 203.440 84.180 205.690 84.480 ;
        RECT 204.480 83.970 204.650 84.180 ;
        RECT 202.245 83.735 203.355 83.965 ;
        RECT 189.930 77.720 192.030 77.890 ;
        RECT 201.150 83.065 201.320 83.645 ;
        RECT 202.245 83.465 202.415 83.735 ;
        RECT 203.185 83.520 203.355 83.735 ;
        RECT 203.525 83.720 205.605 83.970 ;
        RECT 206.285 83.965 206.485 85.130 ;
        RECT 207.810 84.950 207.980 85.560 ;
        RECT 206.765 84.700 207.980 84.950 ;
        RECT 207.810 84.480 207.980 84.700 ;
        RECT 206.790 84.180 207.980 84.480 ;
        RECT 207.810 83.975 207.980 84.180 ;
        RECT 205.775 83.735 206.885 83.965 ;
        RECT 201.585 83.295 202.415 83.465 ;
        RECT 201.150 82.735 202.075 83.065 ;
        RECT 201.150 82.135 201.320 82.735 ;
        RECT 202.245 82.555 202.415 83.295 ;
        RECT 201.585 82.305 202.415 82.555 ;
        RECT 201.150 81.805 202.365 82.135 ;
        RECT 202.585 81.815 203.015 83.490 ;
        RECT 203.185 83.190 204.215 83.520 ;
        RECT 203.185 82.620 203.355 83.190 ;
        RECT 204.480 82.990 204.650 83.720 ;
        RECT 205.775 83.520 205.945 83.735 ;
        RECT 204.915 83.190 205.945 83.520 ;
        RECT 203.525 82.820 205.605 82.990 ;
        RECT 203.185 82.290 204.215 82.620 ;
        RECT 204.480 82.090 204.650 82.820 ;
        RECT 205.775 82.620 205.945 83.190 ;
        RECT 204.915 82.290 205.945 82.620 ;
        RECT 203.185 81.840 205.945 82.090 ;
        RECT 201.150 81.065 201.320 81.805 ;
        RECT 202.650 81.565 202.850 81.815 ;
        RECT 201.585 81.235 204.215 81.565 ;
        RECT 204.480 81.065 204.650 81.840 ;
        RECT 206.115 81.815 206.545 83.490 ;
        RECT 206.715 83.465 206.885 83.735 ;
        RECT 207.055 83.645 207.980 83.975 ;
        RECT 206.715 83.295 207.545 83.465 ;
        RECT 206.715 82.555 206.885 83.295 ;
        RECT 207.810 83.065 207.980 83.645 ;
        RECT 207.055 82.735 207.980 83.065 ;
        RECT 206.715 82.305 207.545 82.555 ;
        RECT 207.810 82.135 207.980 82.735 ;
        RECT 206.280 81.565 206.480 81.815 ;
        RECT 206.765 81.805 207.980 82.135 ;
        RECT 204.915 81.235 207.545 81.565 ;
        RECT 207.810 81.065 207.980 81.805 ;
        RECT 201.150 80.735 202.365 81.065 ;
        RECT 201.150 80.160 201.320 80.735 ;
        RECT 202.535 80.375 203.015 81.065 ;
        RECT 203.185 80.735 205.945 81.065 ;
        RECT 201.150 79.860 202.340 80.160 ;
        RECT 201.150 79.145 201.320 79.860 ;
        RECT 202.600 79.645 202.800 80.375 ;
        RECT 204.480 80.160 204.650 80.735 ;
        RECT 206.115 80.375 206.595 81.065 ;
        RECT 206.765 80.735 207.980 81.065 ;
        RECT 203.440 79.860 205.690 80.160 ;
        RECT 201.585 79.315 204.215 79.645 ;
        RECT 204.480 79.145 204.650 79.860 ;
        RECT 206.330 79.645 206.530 80.375 ;
        RECT 207.810 80.160 207.980 80.735 ;
        RECT 206.790 79.860 207.980 80.160 ;
        RECT 204.915 79.315 207.545 79.645 ;
        RECT 207.810 79.145 207.980 79.860 ;
        RECT 201.150 78.815 202.365 79.145 ;
        RECT 201.150 77.350 201.320 78.815 ;
        RECT 202.535 78.455 203.015 79.145 ;
        RECT 203.185 78.815 205.945 79.145 ;
        RECT 204.480 78.225 204.650 78.815 ;
        RECT 206.115 78.455 206.595 79.145 ;
        RECT 206.765 78.815 207.980 79.145 ;
        RECT 201.585 77.840 202.245 78.170 ;
        RECT 202.415 77.895 202.785 78.225 ;
        RECT 203.055 77.895 206.075 78.225 ;
        RECT 206.345 77.895 206.715 78.225 ;
        RECT 207.810 78.200 207.980 78.815 ;
        RECT 202.075 77.725 202.245 77.840 ;
        RECT 202.075 77.555 204.215 77.725 ;
        RECT 202.415 77.495 204.215 77.555 ;
        RECT 201.150 77.020 202.245 77.350 ;
        RECT 204.480 77.325 204.650 77.895 ;
        RECT 206.885 77.870 207.980 78.200 ;
        RECT 204.915 77.665 206.715 77.725 ;
        RECT 204.915 77.495 207.055 77.665 ;
        RECT 206.885 77.380 207.055 77.495 ;
        RECT 177.140 75.935 178.355 76.265 ;
        RECT 177.140 75.450 177.310 75.935 ;
        RECT 178.525 75.575 179.005 76.265 ;
        RECT 179.175 75.935 180.640 76.265 ;
        RECT 180.470 75.450 180.640 75.935 ;
        RECT 201.150 76.265 201.320 77.020 ;
        RECT 202.415 76.995 202.785 77.325 ;
        RECT 203.055 76.995 206.075 77.325 ;
        RECT 206.345 76.995 206.715 77.325 ;
        RECT 206.885 77.050 207.545 77.380 ;
        RECT 202.520 76.765 202.720 76.995 ;
        RECT 201.585 76.435 204.215 76.765 ;
        RECT 204.480 76.265 204.650 76.995 ;
        RECT 207.810 76.890 207.980 77.870 ;
        RECT 209.020 87.295 211.120 87.465 ;
        RECT 209.020 77.885 209.190 87.295 ;
        RECT 209.820 86.785 210.320 86.955 ;
        RECT 209.590 85.030 209.760 86.570 ;
        RECT 210.380 85.030 210.550 86.570 ;
        RECT 209.820 84.645 210.320 84.815 ;
        RECT 209.590 82.890 209.760 84.430 ;
        RECT 210.380 82.890 210.550 84.430 ;
        RECT 209.820 82.505 210.320 82.675 ;
        RECT 209.590 80.750 209.760 82.290 ;
        RECT 210.380 80.750 210.550 82.290 ;
        RECT 209.820 80.365 210.320 80.535 ;
        RECT 209.590 78.610 209.760 80.150 ;
        RECT 210.380 78.610 210.550 80.150 ;
        RECT 209.820 78.225 210.320 78.395 ;
        RECT 210.950 77.885 211.120 87.295 ;
        RECT 211.480 83.635 211.650 93.045 ;
        RECT 212.280 92.535 212.780 92.705 ;
        RECT 212.050 90.780 212.220 92.320 ;
        RECT 212.840 90.780 213.010 92.320 ;
        RECT 212.280 90.395 212.780 90.565 ;
        RECT 212.050 88.640 212.220 90.180 ;
        RECT 212.840 88.640 213.010 90.180 ;
        RECT 212.280 88.255 212.780 88.425 ;
        RECT 212.050 86.500 212.220 88.040 ;
        RECT 212.840 86.500 213.010 88.040 ;
        RECT 212.280 86.115 212.780 86.285 ;
        RECT 212.050 84.360 212.220 85.900 ;
        RECT 212.840 84.360 213.010 85.900 ;
        RECT 212.280 83.975 212.780 84.145 ;
        RECT 213.410 83.635 213.580 93.045 ;
        RECT 213.940 93.050 216.040 93.220 ;
        RECT 213.940 88.000 214.110 93.050 ;
        RECT 214.740 92.540 215.240 92.710 ;
        RECT 214.510 91.830 214.680 92.370 ;
        RECT 215.300 91.830 215.470 92.370 ;
        RECT 214.740 91.490 215.240 91.660 ;
        RECT 214.510 90.780 214.680 91.320 ;
        RECT 215.300 90.780 215.470 91.320 ;
        RECT 214.740 90.440 215.240 90.610 ;
        RECT 214.510 89.730 214.680 90.270 ;
        RECT 215.300 89.730 215.470 90.270 ;
        RECT 214.740 89.390 215.240 89.560 ;
        RECT 214.510 88.680 214.680 89.220 ;
        RECT 215.300 88.680 215.470 89.220 ;
        RECT 214.740 88.340 215.240 88.510 ;
        RECT 215.870 88.000 216.040 93.050 ;
        RECT 213.940 87.830 216.040 88.000 ;
        RECT 216.400 93.050 220.430 93.220 ;
        RECT 211.480 83.465 213.580 83.635 ;
        RECT 213.940 87.300 216.040 87.470 ;
        RECT 209.020 77.715 211.120 77.885 ;
        RECT 211.480 82.935 213.580 83.105 ;
        RECT 211.480 77.885 211.650 82.935 ;
        RECT 212.280 82.425 212.780 82.595 ;
        RECT 212.050 81.715 212.220 82.255 ;
        RECT 212.840 81.715 213.010 82.255 ;
        RECT 212.280 81.375 212.780 81.545 ;
        RECT 212.050 80.665 212.220 81.205 ;
        RECT 212.840 80.665 213.010 81.205 ;
        RECT 212.280 80.325 212.780 80.495 ;
        RECT 212.050 79.615 212.220 80.155 ;
        RECT 212.840 79.615 213.010 80.155 ;
        RECT 212.280 79.275 212.780 79.445 ;
        RECT 212.050 78.565 212.220 79.105 ;
        RECT 212.840 78.565 213.010 79.105 ;
        RECT 212.280 78.225 212.780 78.395 ;
        RECT 213.410 77.885 213.580 82.935 ;
        RECT 211.480 77.715 213.580 77.885 ;
        RECT 213.940 77.890 214.110 87.300 ;
        RECT 214.740 86.790 215.240 86.960 ;
        RECT 214.510 85.035 214.680 86.575 ;
        RECT 215.300 85.035 215.470 86.575 ;
        RECT 214.740 84.650 215.240 84.820 ;
        RECT 214.510 82.895 214.680 84.435 ;
        RECT 215.300 82.895 215.470 84.435 ;
        RECT 214.740 82.510 215.240 82.680 ;
        RECT 214.510 80.755 214.680 82.295 ;
        RECT 215.300 80.755 215.470 82.295 ;
        RECT 214.740 80.370 215.240 80.540 ;
        RECT 214.510 78.615 214.680 80.155 ;
        RECT 215.300 78.615 215.470 80.155 ;
        RECT 214.740 78.230 215.240 78.400 ;
        RECT 215.870 77.890 216.040 87.300 ;
        RECT 216.400 83.640 216.570 93.050 ;
        RECT 217.200 92.540 217.700 92.710 ;
        RECT 216.970 90.785 217.140 92.325 ;
        RECT 217.760 90.785 217.930 92.325 ;
        RECT 217.200 90.400 217.700 90.570 ;
        RECT 216.970 88.645 217.140 90.185 ;
        RECT 217.760 88.645 217.930 90.185 ;
        RECT 217.200 88.260 217.700 88.430 ;
        RECT 216.970 86.505 217.140 88.045 ;
        RECT 217.760 86.505 217.930 88.045 ;
        RECT 217.200 86.120 217.700 86.290 ;
        RECT 216.970 84.365 217.140 85.905 ;
        RECT 217.760 84.365 217.930 85.905 ;
        RECT 217.200 83.980 217.700 84.150 ;
        RECT 218.330 83.640 218.500 93.050 ;
        RECT 219.130 92.540 219.630 92.710 ;
        RECT 218.900 90.785 219.070 92.325 ;
        RECT 219.690 90.785 219.860 92.325 ;
        RECT 219.130 90.400 219.630 90.570 ;
        RECT 218.900 88.645 219.070 90.185 ;
        RECT 219.690 88.645 219.860 90.185 ;
        RECT 219.130 88.260 219.630 88.430 ;
        RECT 218.900 86.505 219.070 88.045 ;
        RECT 219.690 86.505 219.860 88.045 ;
        RECT 219.130 86.120 219.630 86.290 ;
        RECT 218.900 84.365 219.070 85.905 ;
        RECT 219.690 84.365 219.860 85.905 ;
        RECT 219.130 83.980 219.630 84.150 ;
        RECT 220.260 83.640 220.430 93.050 ;
        RECT 220.790 93.050 224.820 93.220 ;
        RECT 220.790 88.000 220.960 93.050 ;
        RECT 221.590 92.540 222.090 92.710 ;
        RECT 221.360 91.830 221.530 92.370 ;
        RECT 222.150 91.830 222.320 92.370 ;
        RECT 221.590 91.490 222.090 91.660 ;
        RECT 221.360 90.780 221.530 91.320 ;
        RECT 222.150 90.780 222.320 91.320 ;
        RECT 221.590 90.440 222.090 90.610 ;
        RECT 221.360 89.730 221.530 90.270 ;
        RECT 222.150 89.730 222.320 90.270 ;
        RECT 221.590 89.390 222.090 89.560 ;
        RECT 221.360 88.680 221.530 89.220 ;
        RECT 222.150 88.680 222.320 89.220 ;
        RECT 221.590 88.340 222.090 88.510 ;
        RECT 222.720 88.000 222.890 93.050 ;
        RECT 223.520 92.540 224.020 92.710 ;
        RECT 223.290 91.830 223.460 92.370 ;
        RECT 224.080 91.830 224.250 92.370 ;
        RECT 223.520 91.490 224.020 91.660 ;
        RECT 223.290 90.780 223.460 91.320 ;
        RECT 224.080 90.780 224.250 91.320 ;
        RECT 223.520 90.440 224.020 90.610 ;
        RECT 223.290 89.730 223.460 90.270 ;
        RECT 224.080 89.730 224.250 90.270 ;
        RECT 223.520 89.390 224.020 89.560 ;
        RECT 223.290 88.680 223.460 89.220 ;
        RECT 224.080 88.680 224.250 89.220 ;
        RECT 223.520 88.340 224.020 88.510 ;
        RECT 224.650 88.000 224.820 93.050 ;
        RECT 220.790 87.830 224.820 88.000 ;
        RECT 225.160 93.000 225.330 93.210 ;
        RECT 228.490 93.085 228.660 93.210 ;
        RECT 225.160 92.670 226.215 93.000 ;
        RECT 225.160 92.070 225.330 92.670 ;
        RECT 226.385 92.585 226.865 93.085 ;
        RECT 227.065 92.755 230.085 93.085 ;
        RECT 226.385 92.500 228.225 92.585 ;
        RECT 225.595 92.255 228.225 92.500 ;
        RECT 225.595 92.240 226.865 92.255 ;
        RECT 225.160 91.740 226.215 92.070 ;
        RECT 225.160 91.070 225.330 91.740 ;
        RECT 226.385 91.570 226.865 92.240 ;
        RECT 228.490 92.085 228.660 92.755 ;
        RECT 230.285 92.585 230.765 93.085 ;
        RECT 231.820 93.000 231.990 93.210 ;
        RECT 230.935 92.670 231.990 93.000 ;
        RECT 228.925 92.500 230.765 92.585 ;
        RECT 228.925 92.255 231.555 92.500 ;
        RECT 230.285 92.240 231.555 92.255 ;
        RECT 227.065 91.755 230.085 92.085 ;
        RECT 225.595 91.555 226.865 91.570 ;
        RECT 225.595 91.385 228.225 91.555 ;
        RECT 225.595 91.310 226.555 91.385 ;
        RECT 225.595 91.240 226.425 91.310 ;
        RECT 225.160 90.740 226.085 91.070 ;
        RECT 225.160 90.210 225.330 90.740 ;
        RECT 226.255 90.560 226.425 91.240 ;
        RECT 225.595 90.390 226.425 90.560 ;
        RECT 225.160 89.880 226.085 90.210 ;
        RECT 225.160 89.270 225.330 89.880 ;
        RECT 226.255 89.700 226.425 90.390 ;
        RECT 225.595 89.450 226.425 89.700 ;
        RECT 226.595 89.450 227.025 91.140 ;
        RECT 227.195 90.735 227.365 91.385 ;
        RECT 228.490 91.185 228.660 91.755 ;
        RECT 230.285 91.570 230.765 92.240 ;
        RECT 231.820 92.070 231.990 92.670 ;
        RECT 230.935 91.740 231.990 92.070 ;
        RECT 230.285 91.555 231.555 91.570 ;
        RECT 228.925 91.385 231.555 91.555 ;
        RECT 227.535 90.935 229.615 91.185 ;
        RECT 227.195 90.405 228.225 90.735 ;
        RECT 227.195 89.705 227.365 90.405 ;
        RECT 228.490 90.235 228.660 90.935 ;
        RECT 229.785 90.735 229.955 91.385 ;
        RECT 230.595 91.310 231.555 91.385 ;
        RECT 230.725 91.240 231.555 91.310 ;
        RECT 228.925 90.405 229.955 90.735 ;
        RECT 227.535 89.905 229.615 90.235 ;
        RECT 227.195 89.455 228.225 89.705 ;
        RECT 225.160 89.020 226.375 89.270 ;
        RECT 225.160 88.680 225.330 89.020 ;
        RECT 226.660 88.765 226.860 89.450 ;
        RECT 228.490 89.255 228.660 89.905 ;
        RECT 229.785 89.705 229.955 90.405 ;
        RECT 228.925 89.455 229.955 89.705 ;
        RECT 230.125 89.450 230.555 91.140 ;
        RECT 230.725 90.560 230.895 91.240 ;
        RECT 231.820 91.070 231.990 91.740 ;
        RECT 231.065 90.740 231.990 91.070 ;
        RECT 230.725 90.390 231.555 90.560 ;
        RECT 230.725 89.700 230.895 90.390 ;
        RECT 231.820 90.210 231.990 90.740 ;
        RECT 231.065 89.880 231.990 90.210 ;
        RECT 230.725 89.450 231.555 89.700 ;
        RECT 227.065 89.005 230.085 89.255 ;
        RECT 228.490 88.765 228.660 89.005 ;
        RECT 230.290 88.765 230.490 89.450 ;
        RECT 231.820 89.270 231.990 89.880 ;
        RECT 230.775 89.020 231.990 89.270 ;
        RECT 225.160 88.350 226.215 88.680 ;
        RECT 216.400 83.470 220.430 83.640 ;
        RECT 225.160 87.750 225.330 88.350 ;
        RECT 226.385 88.265 226.865 88.765 ;
        RECT 227.065 88.435 230.085 88.765 ;
        RECT 226.385 88.180 228.225 88.265 ;
        RECT 225.595 87.935 228.225 88.180 ;
        RECT 225.595 87.920 226.865 87.935 ;
        RECT 225.160 87.420 226.215 87.750 ;
        RECT 225.160 86.750 225.330 87.420 ;
        RECT 226.385 87.250 226.865 87.920 ;
        RECT 228.490 87.765 228.660 88.435 ;
        RECT 230.285 88.265 230.765 88.765 ;
        RECT 231.820 88.680 231.990 89.020 ;
        RECT 230.935 88.350 231.990 88.680 ;
        RECT 228.925 88.180 230.765 88.265 ;
        RECT 228.925 87.935 231.555 88.180 ;
        RECT 230.285 87.920 231.555 87.935 ;
        RECT 227.065 87.435 230.085 87.765 ;
        RECT 225.595 87.235 226.865 87.250 ;
        RECT 225.595 87.065 228.225 87.235 ;
        RECT 225.595 86.990 226.555 87.065 ;
        RECT 225.595 86.920 226.425 86.990 ;
        RECT 225.160 86.420 226.085 86.750 ;
        RECT 225.160 85.890 225.330 86.420 ;
        RECT 226.255 86.240 226.425 86.920 ;
        RECT 225.595 86.070 226.425 86.240 ;
        RECT 225.160 85.560 226.085 85.890 ;
        RECT 225.160 84.950 225.330 85.560 ;
        RECT 226.255 85.380 226.425 86.070 ;
        RECT 225.595 85.130 226.425 85.380 ;
        RECT 226.595 85.130 227.025 86.820 ;
        RECT 227.195 86.415 227.365 87.065 ;
        RECT 228.490 86.865 228.660 87.435 ;
        RECT 230.285 87.250 230.765 87.920 ;
        RECT 231.820 87.750 231.990 88.350 ;
        RECT 233.035 93.045 235.135 93.215 ;
        RECT 233.035 87.995 233.205 93.045 ;
        RECT 233.835 92.535 234.335 92.705 ;
        RECT 233.605 91.825 233.775 92.365 ;
        RECT 234.395 91.825 234.565 92.365 ;
        RECT 233.835 91.485 234.335 91.655 ;
        RECT 233.605 90.775 233.775 91.315 ;
        RECT 234.395 90.775 234.565 91.315 ;
        RECT 233.835 90.435 234.335 90.605 ;
        RECT 233.605 89.725 233.775 90.265 ;
        RECT 234.395 89.725 234.565 90.265 ;
        RECT 233.835 89.385 234.335 89.555 ;
        RECT 233.605 88.675 233.775 89.215 ;
        RECT 234.395 88.675 234.565 89.215 ;
        RECT 233.835 88.335 234.335 88.505 ;
        RECT 234.965 87.995 235.135 93.045 ;
        RECT 233.035 87.825 235.135 87.995 ;
        RECT 235.495 93.045 237.595 93.215 ;
        RECT 230.935 87.420 231.990 87.750 ;
        RECT 230.285 87.235 231.555 87.250 ;
        RECT 228.925 87.065 231.555 87.235 ;
        RECT 227.535 86.615 229.615 86.865 ;
        RECT 227.195 86.085 228.225 86.415 ;
        RECT 227.195 85.385 227.365 86.085 ;
        RECT 228.490 85.915 228.660 86.615 ;
        RECT 229.785 86.415 229.955 87.065 ;
        RECT 230.595 86.990 231.555 87.065 ;
        RECT 230.725 86.920 231.555 86.990 ;
        RECT 228.925 86.085 229.955 86.415 ;
        RECT 227.535 85.585 229.615 85.915 ;
        RECT 227.195 85.135 228.225 85.385 ;
        RECT 225.160 84.700 226.375 84.950 ;
        RECT 225.160 84.480 225.330 84.700 ;
        RECT 225.160 84.180 226.350 84.480 ;
        RECT 225.160 83.975 225.330 84.180 ;
        RECT 225.160 83.645 226.085 83.975 ;
        RECT 226.660 83.965 226.860 85.130 ;
        RECT 228.490 84.935 228.660 85.585 ;
        RECT 229.785 85.385 229.955 86.085 ;
        RECT 228.925 85.135 229.955 85.385 ;
        RECT 230.125 85.130 230.555 86.820 ;
        RECT 230.725 86.240 230.895 86.920 ;
        RECT 231.820 86.750 231.990 87.420 ;
        RECT 231.065 86.420 231.990 86.750 ;
        RECT 230.725 86.070 231.555 86.240 ;
        RECT 230.725 85.380 230.895 86.070 ;
        RECT 231.820 85.890 231.990 86.420 ;
        RECT 231.065 85.560 231.990 85.890 ;
        RECT 230.725 85.130 231.555 85.380 ;
        RECT 227.065 84.685 230.085 84.935 ;
        RECT 228.490 84.480 228.660 84.685 ;
        RECT 227.450 84.180 229.700 84.480 ;
        RECT 228.490 83.970 228.660 84.180 ;
        RECT 226.255 83.735 227.365 83.965 ;
        RECT 213.940 77.720 216.040 77.890 ;
        RECT 225.160 83.065 225.330 83.645 ;
        RECT 226.255 83.465 226.425 83.735 ;
        RECT 227.195 83.520 227.365 83.735 ;
        RECT 227.535 83.720 229.615 83.970 ;
        RECT 230.295 83.965 230.495 85.130 ;
        RECT 231.820 84.950 231.990 85.560 ;
        RECT 230.775 84.700 231.990 84.950 ;
        RECT 231.820 84.480 231.990 84.700 ;
        RECT 230.800 84.180 231.990 84.480 ;
        RECT 231.820 83.975 231.990 84.180 ;
        RECT 229.785 83.735 230.895 83.965 ;
        RECT 225.595 83.295 226.425 83.465 ;
        RECT 225.160 82.735 226.085 83.065 ;
        RECT 225.160 82.135 225.330 82.735 ;
        RECT 226.255 82.555 226.425 83.295 ;
        RECT 225.595 82.305 226.425 82.555 ;
        RECT 225.160 81.805 226.375 82.135 ;
        RECT 226.595 81.815 227.025 83.490 ;
        RECT 227.195 83.190 228.225 83.520 ;
        RECT 227.195 82.620 227.365 83.190 ;
        RECT 228.490 82.990 228.660 83.720 ;
        RECT 229.785 83.520 229.955 83.735 ;
        RECT 228.925 83.190 229.955 83.520 ;
        RECT 227.535 82.820 229.615 82.990 ;
        RECT 227.195 82.290 228.225 82.620 ;
        RECT 228.490 82.090 228.660 82.820 ;
        RECT 229.785 82.620 229.955 83.190 ;
        RECT 228.925 82.290 229.955 82.620 ;
        RECT 227.195 81.840 229.955 82.090 ;
        RECT 225.160 81.065 225.330 81.805 ;
        RECT 226.660 81.565 226.860 81.815 ;
        RECT 225.595 81.235 228.225 81.565 ;
        RECT 228.490 81.065 228.660 81.840 ;
        RECT 230.125 81.815 230.555 83.490 ;
        RECT 230.725 83.465 230.895 83.735 ;
        RECT 231.065 83.645 231.990 83.975 ;
        RECT 230.725 83.295 231.555 83.465 ;
        RECT 230.725 82.555 230.895 83.295 ;
        RECT 231.820 83.065 231.990 83.645 ;
        RECT 231.065 82.735 231.990 83.065 ;
        RECT 230.725 82.305 231.555 82.555 ;
        RECT 231.820 82.135 231.990 82.735 ;
        RECT 230.290 81.565 230.490 81.815 ;
        RECT 230.775 81.805 231.990 82.135 ;
        RECT 228.925 81.235 231.555 81.565 ;
        RECT 231.820 81.065 231.990 81.805 ;
        RECT 225.160 80.735 226.375 81.065 ;
        RECT 225.160 80.160 225.330 80.735 ;
        RECT 226.545 80.375 227.025 81.065 ;
        RECT 227.195 80.735 229.955 81.065 ;
        RECT 225.160 79.860 226.350 80.160 ;
        RECT 225.160 79.145 225.330 79.860 ;
        RECT 226.610 79.645 226.810 80.375 ;
        RECT 228.490 80.160 228.660 80.735 ;
        RECT 230.125 80.375 230.605 81.065 ;
        RECT 230.775 80.735 231.990 81.065 ;
        RECT 227.450 79.860 229.700 80.160 ;
        RECT 225.595 79.315 228.225 79.645 ;
        RECT 228.490 79.145 228.660 79.860 ;
        RECT 230.340 79.645 230.540 80.375 ;
        RECT 231.820 80.160 231.990 80.735 ;
        RECT 230.800 79.860 231.990 80.160 ;
        RECT 228.925 79.315 231.555 79.645 ;
        RECT 231.820 79.145 231.990 79.860 ;
        RECT 225.160 78.815 226.375 79.145 ;
        RECT 225.160 77.350 225.330 78.815 ;
        RECT 226.545 78.455 227.025 79.145 ;
        RECT 227.195 78.815 229.955 79.145 ;
        RECT 228.490 78.225 228.660 78.815 ;
        RECT 230.125 78.455 230.605 79.145 ;
        RECT 230.775 78.815 231.990 79.145 ;
        RECT 225.595 77.840 226.255 78.170 ;
        RECT 226.425 77.895 226.795 78.225 ;
        RECT 227.065 77.895 230.085 78.225 ;
        RECT 230.355 77.895 230.725 78.225 ;
        RECT 231.820 78.200 231.990 78.815 ;
        RECT 226.085 77.725 226.255 77.840 ;
        RECT 226.085 77.555 228.225 77.725 ;
        RECT 226.425 77.495 228.225 77.555 ;
        RECT 225.160 77.020 226.255 77.350 ;
        RECT 228.490 77.325 228.660 77.895 ;
        RECT 230.895 77.870 231.990 78.200 ;
        RECT 228.925 77.665 230.725 77.725 ;
        RECT 228.925 77.495 231.065 77.665 ;
        RECT 230.895 77.380 231.065 77.495 ;
        RECT 201.150 75.935 202.365 76.265 ;
        RECT 201.150 75.450 201.320 75.935 ;
        RECT 202.535 75.575 203.015 76.265 ;
        RECT 203.185 75.935 204.650 76.265 ;
        RECT 204.480 75.450 204.650 75.935 ;
        RECT 225.160 76.265 225.330 77.020 ;
        RECT 226.425 76.995 226.795 77.325 ;
        RECT 227.065 76.995 230.085 77.325 ;
        RECT 230.355 76.995 230.725 77.325 ;
        RECT 230.895 77.050 231.555 77.380 ;
        RECT 226.530 76.765 226.730 76.995 ;
        RECT 225.595 76.435 228.225 76.765 ;
        RECT 228.490 76.265 228.660 76.995 ;
        RECT 231.820 76.890 231.990 77.870 ;
        RECT 233.035 87.295 235.135 87.465 ;
        RECT 233.035 77.885 233.205 87.295 ;
        RECT 233.835 86.785 234.335 86.955 ;
        RECT 233.605 85.030 233.775 86.570 ;
        RECT 234.395 85.030 234.565 86.570 ;
        RECT 233.835 84.645 234.335 84.815 ;
        RECT 233.605 82.890 233.775 84.430 ;
        RECT 234.395 82.890 234.565 84.430 ;
        RECT 233.835 82.505 234.335 82.675 ;
        RECT 233.605 80.750 233.775 82.290 ;
        RECT 234.395 80.750 234.565 82.290 ;
        RECT 233.835 80.365 234.335 80.535 ;
        RECT 233.605 78.610 233.775 80.150 ;
        RECT 234.395 78.610 234.565 80.150 ;
        RECT 233.835 78.225 234.335 78.395 ;
        RECT 234.965 77.885 235.135 87.295 ;
        RECT 235.495 83.635 235.665 93.045 ;
        RECT 236.295 92.535 236.795 92.705 ;
        RECT 236.065 90.780 236.235 92.320 ;
        RECT 236.855 90.780 237.025 92.320 ;
        RECT 236.295 90.395 236.795 90.565 ;
        RECT 236.065 88.640 236.235 90.180 ;
        RECT 236.855 88.640 237.025 90.180 ;
        RECT 236.295 88.255 236.795 88.425 ;
        RECT 236.065 86.500 236.235 88.040 ;
        RECT 236.855 86.500 237.025 88.040 ;
        RECT 236.295 86.115 236.795 86.285 ;
        RECT 236.065 84.360 236.235 85.900 ;
        RECT 236.855 84.360 237.025 85.900 ;
        RECT 236.295 83.975 236.795 84.145 ;
        RECT 237.425 83.635 237.595 93.045 ;
        RECT 237.955 93.050 240.055 93.220 ;
        RECT 237.955 88.000 238.125 93.050 ;
        RECT 238.755 92.540 239.255 92.710 ;
        RECT 238.525 91.830 238.695 92.370 ;
        RECT 239.315 91.830 239.485 92.370 ;
        RECT 238.755 91.490 239.255 91.660 ;
        RECT 238.525 90.780 238.695 91.320 ;
        RECT 239.315 90.780 239.485 91.320 ;
        RECT 238.755 90.440 239.255 90.610 ;
        RECT 238.525 89.730 238.695 90.270 ;
        RECT 239.315 89.730 239.485 90.270 ;
        RECT 238.755 89.390 239.255 89.560 ;
        RECT 238.525 88.680 238.695 89.220 ;
        RECT 239.315 88.680 239.485 89.220 ;
        RECT 238.755 88.340 239.255 88.510 ;
        RECT 239.885 88.000 240.055 93.050 ;
        RECT 237.955 87.830 240.055 88.000 ;
        RECT 240.415 93.050 244.445 93.220 ;
        RECT 235.495 83.465 237.595 83.635 ;
        RECT 237.955 87.300 240.055 87.470 ;
        RECT 233.035 77.715 235.135 77.885 ;
        RECT 235.495 82.935 237.595 83.105 ;
        RECT 235.495 77.885 235.665 82.935 ;
        RECT 236.295 82.425 236.795 82.595 ;
        RECT 236.065 81.715 236.235 82.255 ;
        RECT 236.855 81.715 237.025 82.255 ;
        RECT 236.295 81.375 236.795 81.545 ;
        RECT 236.065 80.665 236.235 81.205 ;
        RECT 236.855 80.665 237.025 81.205 ;
        RECT 236.295 80.325 236.795 80.495 ;
        RECT 236.065 79.615 236.235 80.155 ;
        RECT 236.855 79.615 237.025 80.155 ;
        RECT 236.295 79.275 236.795 79.445 ;
        RECT 236.065 78.565 236.235 79.105 ;
        RECT 236.855 78.565 237.025 79.105 ;
        RECT 236.295 78.225 236.795 78.395 ;
        RECT 237.425 77.885 237.595 82.935 ;
        RECT 235.495 77.715 237.595 77.885 ;
        RECT 237.955 77.890 238.125 87.300 ;
        RECT 238.755 86.790 239.255 86.960 ;
        RECT 238.525 85.035 238.695 86.575 ;
        RECT 239.315 85.035 239.485 86.575 ;
        RECT 238.755 84.650 239.255 84.820 ;
        RECT 238.525 82.895 238.695 84.435 ;
        RECT 239.315 82.895 239.485 84.435 ;
        RECT 238.755 82.510 239.255 82.680 ;
        RECT 238.525 80.755 238.695 82.295 ;
        RECT 239.315 80.755 239.485 82.295 ;
        RECT 238.755 80.370 239.255 80.540 ;
        RECT 238.525 78.615 238.695 80.155 ;
        RECT 239.315 78.615 239.485 80.155 ;
        RECT 238.755 78.230 239.255 78.400 ;
        RECT 239.885 77.890 240.055 87.300 ;
        RECT 240.415 83.640 240.585 93.050 ;
        RECT 241.215 92.540 241.715 92.710 ;
        RECT 240.985 90.785 241.155 92.325 ;
        RECT 241.775 90.785 241.945 92.325 ;
        RECT 241.215 90.400 241.715 90.570 ;
        RECT 240.985 88.645 241.155 90.185 ;
        RECT 241.775 88.645 241.945 90.185 ;
        RECT 241.215 88.260 241.715 88.430 ;
        RECT 240.985 86.505 241.155 88.045 ;
        RECT 241.775 86.505 241.945 88.045 ;
        RECT 241.215 86.120 241.715 86.290 ;
        RECT 240.985 84.365 241.155 85.905 ;
        RECT 241.775 84.365 241.945 85.905 ;
        RECT 241.215 83.980 241.715 84.150 ;
        RECT 242.345 83.640 242.515 93.050 ;
        RECT 243.145 92.540 243.645 92.710 ;
        RECT 242.915 90.785 243.085 92.325 ;
        RECT 243.705 90.785 243.875 92.325 ;
        RECT 243.145 90.400 243.645 90.570 ;
        RECT 242.915 88.645 243.085 90.185 ;
        RECT 243.705 88.645 243.875 90.185 ;
        RECT 243.145 88.260 243.645 88.430 ;
        RECT 242.915 86.505 243.085 88.045 ;
        RECT 243.705 86.505 243.875 88.045 ;
        RECT 243.145 86.120 243.645 86.290 ;
        RECT 242.915 84.365 243.085 85.905 ;
        RECT 243.705 84.365 243.875 85.905 ;
        RECT 243.145 83.980 243.645 84.150 ;
        RECT 244.275 83.640 244.445 93.050 ;
        RECT 244.805 93.050 248.835 93.220 ;
        RECT 244.805 88.000 244.975 93.050 ;
        RECT 245.605 92.540 246.105 92.710 ;
        RECT 245.375 91.830 245.545 92.370 ;
        RECT 246.165 91.830 246.335 92.370 ;
        RECT 245.605 91.490 246.105 91.660 ;
        RECT 245.375 90.780 245.545 91.320 ;
        RECT 246.165 90.780 246.335 91.320 ;
        RECT 245.605 90.440 246.105 90.610 ;
        RECT 245.375 89.730 245.545 90.270 ;
        RECT 246.165 89.730 246.335 90.270 ;
        RECT 245.605 89.390 246.105 89.560 ;
        RECT 245.375 88.680 245.545 89.220 ;
        RECT 246.165 88.680 246.335 89.220 ;
        RECT 245.605 88.340 246.105 88.510 ;
        RECT 246.735 88.000 246.905 93.050 ;
        RECT 247.535 92.540 248.035 92.710 ;
        RECT 247.305 91.830 247.475 92.370 ;
        RECT 248.095 91.830 248.265 92.370 ;
        RECT 247.535 91.490 248.035 91.660 ;
        RECT 247.305 90.780 247.475 91.320 ;
        RECT 248.095 90.780 248.265 91.320 ;
        RECT 247.535 90.440 248.035 90.610 ;
        RECT 247.305 89.730 247.475 90.270 ;
        RECT 248.095 89.730 248.265 90.270 ;
        RECT 247.535 89.390 248.035 89.560 ;
        RECT 247.305 88.680 247.475 89.220 ;
        RECT 248.095 88.680 248.265 89.220 ;
        RECT 247.535 88.340 248.035 88.510 ;
        RECT 248.665 88.000 248.835 93.050 ;
        RECT 244.805 87.830 248.835 88.000 ;
        RECT 249.175 93.000 249.345 93.210 ;
        RECT 252.505 93.085 252.675 93.210 ;
        RECT 249.175 92.670 250.230 93.000 ;
        RECT 249.175 92.070 249.345 92.670 ;
        RECT 250.400 92.585 250.880 93.085 ;
        RECT 251.080 92.755 254.100 93.085 ;
        RECT 250.400 92.500 252.240 92.585 ;
        RECT 249.610 92.255 252.240 92.500 ;
        RECT 249.610 92.240 250.880 92.255 ;
        RECT 249.175 91.740 250.230 92.070 ;
        RECT 249.175 91.070 249.345 91.740 ;
        RECT 250.400 91.570 250.880 92.240 ;
        RECT 252.505 92.085 252.675 92.755 ;
        RECT 254.300 92.585 254.780 93.085 ;
        RECT 255.835 93.000 256.005 93.210 ;
        RECT 254.950 92.670 256.005 93.000 ;
        RECT 252.940 92.500 254.780 92.585 ;
        RECT 252.940 92.255 255.570 92.500 ;
        RECT 254.300 92.240 255.570 92.255 ;
        RECT 251.080 91.755 254.100 92.085 ;
        RECT 249.610 91.555 250.880 91.570 ;
        RECT 249.610 91.385 252.240 91.555 ;
        RECT 249.610 91.310 250.570 91.385 ;
        RECT 249.610 91.240 250.440 91.310 ;
        RECT 249.175 90.740 250.100 91.070 ;
        RECT 249.175 90.210 249.345 90.740 ;
        RECT 250.270 90.560 250.440 91.240 ;
        RECT 249.610 90.390 250.440 90.560 ;
        RECT 249.175 89.880 250.100 90.210 ;
        RECT 249.175 89.270 249.345 89.880 ;
        RECT 250.270 89.700 250.440 90.390 ;
        RECT 249.610 89.450 250.440 89.700 ;
        RECT 250.610 89.450 251.040 91.140 ;
        RECT 251.210 90.735 251.380 91.385 ;
        RECT 252.505 91.185 252.675 91.755 ;
        RECT 254.300 91.570 254.780 92.240 ;
        RECT 255.835 92.070 256.005 92.670 ;
        RECT 254.950 91.740 256.005 92.070 ;
        RECT 254.300 91.555 255.570 91.570 ;
        RECT 252.940 91.385 255.570 91.555 ;
        RECT 251.550 90.935 253.630 91.185 ;
        RECT 251.210 90.405 252.240 90.735 ;
        RECT 251.210 89.705 251.380 90.405 ;
        RECT 252.505 90.235 252.675 90.935 ;
        RECT 253.800 90.735 253.970 91.385 ;
        RECT 254.610 91.310 255.570 91.385 ;
        RECT 254.740 91.240 255.570 91.310 ;
        RECT 252.940 90.405 253.970 90.735 ;
        RECT 251.550 89.905 253.630 90.235 ;
        RECT 251.210 89.455 252.240 89.705 ;
        RECT 249.175 89.020 250.390 89.270 ;
        RECT 249.175 88.680 249.345 89.020 ;
        RECT 250.675 88.765 250.875 89.450 ;
        RECT 252.505 89.255 252.675 89.905 ;
        RECT 253.800 89.705 253.970 90.405 ;
        RECT 252.940 89.455 253.970 89.705 ;
        RECT 254.140 89.450 254.570 91.140 ;
        RECT 254.740 90.560 254.910 91.240 ;
        RECT 255.835 91.070 256.005 91.740 ;
        RECT 255.080 90.740 256.005 91.070 ;
        RECT 254.740 90.390 255.570 90.560 ;
        RECT 254.740 89.700 254.910 90.390 ;
        RECT 255.835 90.210 256.005 90.740 ;
        RECT 255.080 89.880 256.005 90.210 ;
        RECT 254.740 89.450 255.570 89.700 ;
        RECT 251.080 89.005 254.100 89.255 ;
        RECT 252.505 88.765 252.675 89.005 ;
        RECT 254.305 88.765 254.505 89.450 ;
        RECT 255.835 89.270 256.005 89.880 ;
        RECT 254.790 89.020 256.005 89.270 ;
        RECT 249.175 88.350 250.230 88.680 ;
        RECT 240.415 83.470 244.445 83.640 ;
        RECT 249.175 87.750 249.345 88.350 ;
        RECT 250.400 88.265 250.880 88.765 ;
        RECT 251.080 88.435 254.100 88.765 ;
        RECT 250.400 88.180 252.240 88.265 ;
        RECT 249.610 87.935 252.240 88.180 ;
        RECT 249.610 87.920 250.880 87.935 ;
        RECT 249.175 87.420 250.230 87.750 ;
        RECT 249.175 86.750 249.345 87.420 ;
        RECT 250.400 87.250 250.880 87.920 ;
        RECT 252.505 87.765 252.675 88.435 ;
        RECT 254.300 88.265 254.780 88.765 ;
        RECT 255.835 88.680 256.005 89.020 ;
        RECT 254.950 88.350 256.005 88.680 ;
        RECT 252.940 88.180 254.780 88.265 ;
        RECT 252.940 87.935 255.570 88.180 ;
        RECT 254.300 87.920 255.570 87.935 ;
        RECT 251.080 87.435 254.100 87.765 ;
        RECT 249.610 87.235 250.880 87.250 ;
        RECT 249.610 87.065 252.240 87.235 ;
        RECT 249.610 86.990 250.570 87.065 ;
        RECT 249.610 86.920 250.440 86.990 ;
        RECT 249.175 86.420 250.100 86.750 ;
        RECT 249.175 85.890 249.345 86.420 ;
        RECT 250.270 86.240 250.440 86.920 ;
        RECT 249.610 86.070 250.440 86.240 ;
        RECT 249.175 85.560 250.100 85.890 ;
        RECT 249.175 84.950 249.345 85.560 ;
        RECT 250.270 85.380 250.440 86.070 ;
        RECT 249.610 85.130 250.440 85.380 ;
        RECT 250.610 85.130 251.040 86.820 ;
        RECT 251.210 86.415 251.380 87.065 ;
        RECT 252.505 86.865 252.675 87.435 ;
        RECT 254.300 87.250 254.780 87.920 ;
        RECT 255.835 87.750 256.005 88.350 ;
        RECT 257.090 93.045 259.190 93.215 ;
        RECT 257.090 87.995 257.260 93.045 ;
        RECT 257.890 92.535 258.390 92.705 ;
        RECT 257.660 91.825 257.830 92.365 ;
        RECT 258.450 91.825 258.620 92.365 ;
        RECT 257.890 91.485 258.390 91.655 ;
        RECT 257.660 90.775 257.830 91.315 ;
        RECT 258.450 90.775 258.620 91.315 ;
        RECT 257.890 90.435 258.390 90.605 ;
        RECT 257.660 89.725 257.830 90.265 ;
        RECT 258.450 89.725 258.620 90.265 ;
        RECT 257.890 89.385 258.390 89.555 ;
        RECT 257.660 88.675 257.830 89.215 ;
        RECT 258.450 88.675 258.620 89.215 ;
        RECT 257.890 88.335 258.390 88.505 ;
        RECT 259.020 87.995 259.190 93.045 ;
        RECT 257.090 87.825 259.190 87.995 ;
        RECT 259.550 93.045 261.650 93.215 ;
        RECT 254.950 87.420 256.005 87.750 ;
        RECT 254.300 87.235 255.570 87.250 ;
        RECT 252.940 87.065 255.570 87.235 ;
        RECT 251.550 86.615 253.630 86.865 ;
        RECT 251.210 86.085 252.240 86.415 ;
        RECT 251.210 85.385 251.380 86.085 ;
        RECT 252.505 85.915 252.675 86.615 ;
        RECT 253.800 86.415 253.970 87.065 ;
        RECT 254.610 86.990 255.570 87.065 ;
        RECT 254.740 86.920 255.570 86.990 ;
        RECT 252.940 86.085 253.970 86.415 ;
        RECT 251.550 85.585 253.630 85.915 ;
        RECT 251.210 85.135 252.240 85.385 ;
        RECT 249.175 84.700 250.390 84.950 ;
        RECT 249.175 84.480 249.345 84.700 ;
        RECT 249.175 84.180 250.365 84.480 ;
        RECT 249.175 83.975 249.345 84.180 ;
        RECT 249.175 83.645 250.100 83.975 ;
        RECT 250.675 83.965 250.875 85.130 ;
        RECT 252.505 84.935 252.675 85.585 ;
        RECT 253.800 85.385 253.970 86.085 ;
        RECT 252.940 85.135 253.970 85.385 ;
        RECT 254.140 85.130 254.570 86.820 ;
        RECT 254.740 86.240 254.910 86.920 ;
        RECT 255.835 86.750 256.005 87.420 ;
        RECT 255.080 86.420 256.005 86.750 ;
        RECT 254.740 86.070 255.570 86.240 ;
        RECT 254.740 85.380 254.910 86.070 ;
        RECT 255.835 85.890 256.005 86.420 ;
        RECT 255.080 85.560 256.005 85.890 ;
        RECT 254.740 85.130 255.570 85.380 ;
        RECT 251.080 84.685 254.100 84.935 ;
        RECT 252.505 84.480 252.675 84.685 ;
        RECT 251.465 84.180 253.715 84.480 ;
        RECT 252.505 83.970 252.675 84.180 ;
        RECT 250.270 83.735 251.380 83.965 ;
        RECT 237.955 77.720 240.055 77.890 ;
        RECT 249.175 83.065 249.345 83.645 ;
        RECT 250.270 83.465 250.440 83.735 ;
        RECT 251.210 83.520 251.380 83.735 ;
        RECT 251.550 83.720 253.630 83.970 ;
        RECT 254.310 83.965 254.510 85.130 ;
        RECT 255.835 84.950 256.005 85.560 ;
        RECT 254.790 84.700 256.005 84.950 ;
        RECT 255.835 84.480 256.005 84.700 ;
        RECT 254.815 84.180 256.005 84.480 ;
        RECT 255.835 83.975 256.005 84.180 ;
        RECT 253.800 83.735 254.910 83.965 ;
        RECT 249.610 83.295 250.440 83.465 ;
        RECT 249.175 82.735 250.100 83.065 ;
        RECT 249.175 82.135 249.345 82.735 ;
        RECT 250.270 82.555 250.440 83.295 ;
        RECT 249.610 82.305 250.440 82.555 ;
        RECT 249.175 81.805 250.390 82.135 ;
        RECT 250.610 81.815 251.040 83.490 ;
        RECT 251.210 83.190 252.240 83.520 ;
        RECT 251.210 82.620 251.380 83.190 ;
        RECT 252.505 82.990 252.675 83.720 ;
        RECT 253.800 83.520 253.970 83.735 ;
        RECT 252.940 83.190 253.970 83.520 ;
        RECT 251.550 82.820 253.630 82.990 ;
        RECT 251.210 82.290 252.240 82.620 ;
        RECT 252.505 82.090 252.675 82.820 ;
        RECT 253.800 82.620 253.970 83.190 ;
        RECT 252.940 82.290 253.970 82.620 ;
        RECT 251.210 81.840 253.970 82.090 ;
        RECT 249.175 81.065 249.345 81.805 ;
        RECT 250.675 81.565 250.875 81.815 ;
        RECT 249.610 81.235 252.240 81.565 ;
        RECT 252.505 81.065 252.675 81.840 ;
        RECT 254.140 81.815 254.570 83.490 ;
        RECT 254.740 83.465 254.910 83.735 ;
        RECT 255.080 83.645 256.005 83.975 ;
        RECT 254.740 83.295 255.570 83.465 ;
        RECT 254.740 82.555 254.910 83.295 ;
        RECT 255.835 83.065 256.005 83.645 ;
        RECT 255.080 82.735 256.005 83.065 ;
        RECT 254.740 82.305 255.570 82.555 ;
        RECT 255.835 82.135 256.005 82.735 ;
        RECT 254.305 81.565 254.505 81.815 ;
        RECT 254.790 81.805 256.005 82.135 ;
        RECT 252.940 81.235 255.570 81.565 ;
        RECT 255.835 81.065 256.005 81.805 ;
        RECT 249.175 80.735 250.390 81.065 ;
        RECT 249.175 80.160 249.345 80.735 ;
        RECT 250.560 80.375 251.040 81.065 ;
        RECT 251.210 80.735 253.970 81.065 ;
        RECT 249.175 79.860 250.365 80.160 ;
        RECT 249.175 79.145 249.345 79.860 ;
        RECT 250.625 79.645 250.825 80.375 ;
        RECT 252.505 80.160 252.675 80.735 ;
        RECT 254.140 80.375 254.620 81.065 ;
        RECT 254.790 80.735 256.005 81.065 ;
        RECT 251.465 79.860 253.715 80.160 ;
        RECT 249.610 79.315 252.240 79.645 ;
        RECT 252.505 79.145 252.675 79.860 ;
        RECT 254.355 79.645 254.555 80.375 ;
        RECT 255.835 80.160 256.005 80.735 ;
        RECT 254.815 79.860 256.005 80.160 ;
        RECT 252.940 79.315 255.570 79.645 ;
        RECT 255.835 79.145 256.005 79.860 ;
        RECT 249.175 78.815 250.390 79.145 ;
        RECT 249.175 77.350 249.345 78.815 ;
        RECT 250.560 78.455 251.040 79.145 ;
        RECT 251.210 78.815 253.970 79.145 ;
        RECT 252.505 78.225 252.675 78.815 ;
        RECT 254.140 78.455 254.620 79.145 ;
        RECT 254.790 78.815 256.005 79.145 ;
        RECT 249.610 77.840 250.270 78.170 ;
        RECT 250.440 77.895 250.810 78.225 ;
        RECT 251.080 77.895 254.100 78.225 ;
        RECT 254.370 77.895 254.740 78.225 ;
        RECT 255.835 78.200 256.005 78.815 ;
        RECT 250.100 77.725 250.270 77.840 ;
        RECT 250.100 77.555 252.240 77.725 ;
        RECT 250.440 77.495 252.240 77.555 ;
        RECT 249.175 77.020 250.270 77.350 ;
        RECT 252.505 77.325 252.675 77.895 ;
        RECT 254.910 77.870 256.005 78.200 ;
        RECT 252.940 77.665 254.740 77.725 ;
        RECT 252.940 77.495 255.080 77.665 ;
        RECT 254.910 77.380 255.080 77.495 ;
        RECT 225.160 75.935 226.375 76.265 ;
        RECT 225.160 75.450 225.330 75.935 ;
        RECT 226.545 75.575 227.025 76.265 ;
        RECT 227.195 75.935 228.660 76.265 ;
        RECT 228.490 75.450 228.660 75.935 ;
        RECT 249.175 76.265 249.345 77.020 ;
        RECT 250.440 76.995 250.810 77.325 ;
        RECT 251.080 76.995 254.100 77.325 ;
        RECT 254.370 76.995 254.740 77.325 ;
        RECT 254.910 77.050 255.570 77.380 ;
        RECT 250.545 76.765 250.745 76.995 ;
        RECT 249.610 76.435 252.240 76.765 ;
        RECT 252.505 76.265 252.675 76.995 ;
        RECT 255.835 76.890 256.005 77.870 ;
        RECT 257.090 87.295 259.190 87.465 ;
        RECT 257.090 77.885 257.260 87.295 ;
        RECT 257.890 86.785 258.390 86.955 ;
        RECT 257.660 85.030 257.830 86.570 ;
        RECT 258.450 85.030 258.620 86.570 ;
        RECT 257.890 84.645 258.390 84.815 ;
        RECT 257.660 82.890 257.830 84.430 ;
        RECT 258.450 82.890 258.620 84.430 ;
        RECT 257.890 82.505 258.390 82.675 ;
        RECT 257.660 80.750 257.830 82.290 ;
        RECT 258.450 80.750 258.620 82.290 ;
        RECT 257.890 80.365 258.390 80.535 ;
        RECT 257.660 78.610 257.830 80.150 ;
        RECT 258.450 78.610 258.620 80.150 ;
        RECT 257.890 78.225 258.390 78.395 ;
        RECT 259.020 77.885 259.190 87.295 ;
        RECT 259.550 83.635 259.720 93.045 ;
        RECT 260.350 92.535 260.850 92.705 ;
        RECT 260.120 90.780 260.290 92.320 ;
        RECT 260.910 90.780 261.080 92.320 ;
        RECT 260.350 90.395 260.850 90.565 ;
        RECT 260.120 88.640 260.290 90.180 ;
        RECT 260.910 88.640 261.080 90.180 ;
        RECT 260.350 88.255 260.850 88.425 ;
        RECT 260.120 86.500 260.290 88.040 ;
        RECT 260.910 86.500 261.080 88.040 ;
        RECT 260.350 86.115 260.850 86.285 ;
        RECT 260.120 84.360 260.290 85.900 ;
        RECT 260.910 84.360 261.080 85.900 ;
        RECT 260.350 83.975 260.850 84.145 ;
        RECT 261.480 83.635 261.650 93.045 ;
        RECT 262.010 93.050 264.110 93.220 ;
        RECT 262.010 88.000 262.180 93.050 ;
        RECT 262.810 92.540 263.310 92.710 ;
        RECT 262.580 91.830 262.750 92.370 ;
        RECT 263.370 91.830 263.540 92.370 ;
        RECT 262.810 91.490 263.310 91.660 ;
        RECT 262.580 90.780 262.750 91.320 ;
        RECT 263.370 90.780 263.540 91.320 ;
        RECT 262.810 90.440 263.310 90.610 ;
        RECT 262.580 89.730 262.750 90.270 ;
        RECT 263.370 89.730 263.540 90.270 ;
        RECT 262.810 89.390 263.310 89.560 ;
        RECT 262.580 88.680 262.750 89.220 ;
        RECT 263.370 88.680 263.540 89.220 ;
        RECT 262.810 88.340 263.310 88.510 ;
        RECT 263.940 88.000 264.110 93.050 ;
        RECT 262.010 87.830 264.110 88.000 ;
        RECT 264.470 93.050 268.500 93.220 ;
        RECT 259.550 83.465 261.650 83.635 ;
        RECT 262.010 87.300 264.110 87.470 ;
        RECT 257.090 77.715 259.190 77.885 ;
        RECT 259.550 82.935 261.650 83.105 ;
        RECT 259.550 77.885 259.720 82.935 ;
        RECT 260.350 82.425 260.850 82.595 ;
        RECT 260.120 81.715 260.290 82.255 ;
        RECT 260.910 81.715 261.080 82.255 ;
        RECT 260.350 81.375 260.850 81.545 ;
        RECT 260.120 80.665 260.290 81.205 ;
        RECT 260.910 80.665 261.080 81.205 ;
        RECT 260.350 80.325 260.850 80.495 ;
        RECT 260.120 79.615 260.290 80.155 ;
        RECT 260.910 79.615 261.080 80.155 ;
        RECT 260.350 79.275 260.850 79.445 ;
        RECT 260.120 78.565 260.290 79.105 ;
        RECT 260.910 78.565 261.080 79.105 ;
        RECT 260.350 78.225 260.850 78.395 ;
        RECT 261.480 77.885 261.650 82.935 ;
        RECT 259.550 77.715 261.650 77.885 ;
        RECT 262.010 77.890 262.180 87.300 ;
        RECT 262.810 86.790 263.310 86.960 ;
        RECT 262.580 85.035 262.750 86.575 ;
        RECT 263.370 85.035 263.540 86.575 ;
        RECT 262.810 84.650 263.310 84.820 ;
        RECT 262.580 82.895 262.750 84.435 ;
        RECT 263.370 82.895 263.540 84.435 ;
        RECT 262.810 82.510 263.310 82.680 ;
        RECT 262.580 80.755 262.750 82.295 ;
        RECT 263.370 80.755 263.540 82.295 ;
        RECT 262.810 80.370 263.310 80.540 ;
        RECT 262.580 78.615 262.750 80.155 ;
        RECT 263.370 78.615 263.540 80.155 ;
        RECT 262.810 78.230 263.310 78.400 ;
        RECT 263.940 77.890 264.110 87.300 ;
        RECT 264.470 83.640 264.640 93.050 ;
        RECT 265.270 92.540 265.770 92.710 ;
        RECT 265.040 90.785 265.210 92.325 ;
        RECT 265.830 90.785 266.000 92.325 ;
        RECT 265.270 90.400 265.770 90.570 ;
        RECT 265.040 88.645 265.210 90.185 ;
        RECT 265.830 88.645 266.000 90.185 ;
        RECT 265.270 88.260 265.770 88.430 ;
        RECT 265.040 86.505 265.210 88.045 ;
        RECT 265.830 86.505 266.000 88.045 ;
        RECT 265.270 86.120 265.770 86.290 ;
        RECT 265.040 84.365 265.210 85.905 ;
        RECT 265.830 84.365 266.000 85.905 ;
        RECT 265.270 83.980 265.770 84.150 ;
        RECT 266.400 83.640 266.570 93.050 ;
        RECT 267.200 92.540 267.700 92.710 ;
        RECT 266.970 90.785 267.140 92.325 ;
        RECT 267.760 90.785 267.930 92.325 ;
        RECT 267.200 90.400 267.700 90.570 ;
        RECT 266.970 88.645 267.140 90.185 ;
        RECT 267.760 88.645 267.930 90.185 ;
        RECT 267.200 88.260 267.700 88.430 ;
        RECT 266.970 86.505 267.140 88.045 ;
        RECT 267.760 86.505 267.930 88.045 ;
        RECT 267.200 86.120 267.700 86.290 ;
        RECT 266.970 84.365 267.140 85.905 ;
        RECT 267.760 84.365 267.930 85.905 ;
        RECT 267.200 83.980 267.700 84.150 ;
        RECT 268.330 83.640 268.500 93.050 ;
        RECT 268.860 93.050 272.890 93.220 ;
        RECT 268.860 88.000 269.030 93.050 ;
        RECT 269.660 92.540 270.160 92.710 ;
        RECT 269.430 91.830 269.600 92.370 ;
        RECT 270.220 91.830 270.390 92.370 ;
        RECT 269.660 91.490 270.160 91.660 ;
        RECT 269.430 90.780 269.600 91.320 ;
        RECT 270.220 90.780 270.390 91.320 ;
        RECT 269.660 90.440 270.160 90.610 ;
        RECT 269.430 89.730 269.600 90.270 ;
        RECT 270.220 89.730 270.390 90.270 ;
        RECT 269.660 89.390 270.160 89.560 ;
        RECT 269.430 88.680 269.600 89.220 ;
        RECT 270.220 88.680 270.390 89.220 ;
        RECT 269.660 88.340 270.160 88.510 ;
        RECT 270.790 88.000 270.960 93.050 ;
        RECT 271.590 92.540 272.090 92.710 ;
        RECT 271.360 91.830 271.530 92.370 ;
        RECT 272.150 91.830 272.320 92.370 ;
        RECT 271.590 91.490 272.090 91.660 ;
        RECT 271.360 90.780 271.530 91.320 ;
        RECT 272.150 90.780 272.320 91.320 ;
        RECT 271.590 90.440 272.090 90.610 ;
        RECT 271.360 89.730 271.530 90.270 ;
        RECT 272.150 89.730 272.320 90.270 ;
        RECT 271.590 89.390 272.090 89.560 ;
        RECT 271.360 88.680 271.530 89.220 ;
        RECT 272.150 88.680 272.320 89.220 ;
        RECT 271.590 88.340 272.090 88.510 ;
        RECT 272.720 88.000 272.890 93.050 ;
        RECT 268.860 87.830 272.890 88.000 ;
        RECT 273.230 93.000 273.400 93.210 ;
        RECT 276.560 93.085 276.730 93.210 ;
        RECT 273.230 92.670 274.285 93.000 ;
        RECT 273.230 92.070 273.400 92.670 ;
        RECT 274.455 92.585 274.935 93.085 ;
        RECT 275.135 92.755 278.155 93.085 ;
        RECT 274.455 92.500 276.295 92.585 ;
        RECT 273.665 92.255 276.295 92.500 ;
        RECT 273.665 92.240 274.935 92.255 ;
        RECT 273.230 91.740 274.285 92.070 ;
        RECT 273.230 91.070 273.400 91.740 ;
        RECT 274.455 91.570 274.935 92.240 ;
        RECT 276.560 92.085 276.730 92.755 ;
        RECT 278.355 92.585 278.835 93.085 ;
        RECT 279.890 93.000 280.060 93.210 ;
        RECT 279.005 92.670 280.060 93.000 ;
        RECT 276.995 92.500 278.835 92.585 ;
        RECT 276.995 92.255 279.625 92.500 ;
        RECT 278.355 92.240 279.625 92.255 ;
        RECT 275.135 91.755 278.155 92.085 ;
        RECT 273.665 91.555 274.935 91.570 ;
        RECT 273.665 91.385 276.295 91.555 ;
        RECT 273.665 91.310 274.625 91.385 ;
        RECT 273.665 91.240 274.495 91.310 ;
        RECT 273.230 90.740 274.155 91.070 ;
        RECT 273.230 90.210 273.400 90.740 ;
        RECT 274.325 90.560 274.495 91.240 ;
        RECT 273.665 90.390 274.495 90.560 ;
        RECT 273.230 89.880 274.155 90.210 ;
        RECT 273.230 89.270 273.400 89.880 ;
        RECT 274.325 89.700 274.495 90.390 ;
        RECT 273.665 89.450 274.495 89.700 ;
        RECT 274.665 89.450 275.095 91.140 ;
        RECT 275.265 90.735 275.435 91.385 ;
        RECT 276.560 91.185 276.730 91.755 ;
        RECT 278.355 91.570 278.835 92.240 ;
        RECT 279.890 92.070 280.060 92.670 ;
        RECT 279.005 91.740 280.060 92.070 ;
        RECT 278.355 91.555 279.625 91.570 ;
        RECT 276.995 91.385 279.625 91.555 ;
        RECT 275.605 90.935 277.685 91.185 ;
        RECT 275.265 90.405 276.295 90.735 ;
        RECT 275.265 89.705 275.435 90.405 ;
        RECT 276.560 90.235 276.730 90.935 ;
        RECT 277.855 90.735 278.025 91.385 ;
        RECT 278.665 91.310 279.625 91.385 ;
        RECT 278.795 91.240 279.625 91.310 ;
        RECT 276.995 90.405 278.025 90.735 ;
        RECT 275.605 89.905 277.685 90.235 ;
        RECT 275.265 89.455 276.295 89.705 ;
        RECT 273.230 89.020 274.445 89.270 ;
        RECT 273.230 88.680 273.400 89.020 ;
        RECT 274.730 88.765 274.930 89.450 ;
        RECT 276.560 89.255 276.730 89.905 ;
        RECT 277.855 89.705 278.025 90.405 ;
        RECT 276.995 89.455 278.025 89.705 ;
        RECT 278.195 89.450 278.625 91.140 ;
        RECT 278.795 90.560 278.965 91.240 ;
        RECT 279.890 91.070 280.060 91.740 ;
        RECT 279.135 90.740 280.060 91.070 ;
        RECT 278.795 90.390 279.625 90.560 ;
        RECT 278.795 89.700 278.965 90.390 ;
        RECT 279.890 90.210 280.060 90.740 ;
        RECT 279.135 89.880 280.060 90.210 ;
        RECT 278.795 89.450 279.625 89.700 ;
        RECT 275.135 89.005 278.155 89.255 ;
        RECT 276.560 88.765 276.730 89.005 ;
        RECT 278.360 88.765 278.560 89.450 ;
        RECT 279.890 89.270 280.060 89.880 ;
        RECT 278.845 89.020 280.060 89.270 ;
        RECT 273.230 88.350 274.285 88.680 ;
        RECT 264.470 83.470 268.500 83.640 ;
        RECT 273.230 87.750 273.400 88.350 ;
        RECT 274.455 88.265 274.935 88.765 ;
        RECT 275.135 88.435 278.155 88.765 ;
        RECT 274.455 88.180 276.295 88.265 ;
        RECT 273.665 87.935 276.295 88.180 ;
        RECT 273.665 87.920 274.935 87.935 ;
        RECT 273.230 87.420 274.285 87.750 ;
        RECT 273.230 86.750 273.400 87.420 ;
        RECT 274.455 87.250 274.935 87.920 ;
        RECT 276.560 87.765 276.730 88.435 ;
        RECT 278.355 88.265 278.835 88.765 ;
        RECT 279.890 88.680 280.060 89.020 ;
        RECT 279.005 88.350 280.060 88.680 ;
        RECT 276.995 88.180 278.835 88.265 ;
        RECT 276.995 87.935 279.625 88.180 ;
        RECT 278.355 87.920 279.625 87.935 ;
        RECT 275.135 87.435 278.155 87.765 ;
        RECT 273.665 87.235 274.935 87.250 ;
        RECT 273.665 87.065 276.295 87.235 ;
        RECT 273.665 86.990 274.625 87.065 ;
        RECT 273.665 86.920 274.495 86.990 ;
        RECT 273.230 86.420 274.155 86.750 ;
        RECT 273.230 85.890 273.400 86.420 ;
        RECT 274.325 86.240 274.495 86.920 ;
        RECT 273.665 86.070 274.495 86.240 ;
        RECT 273.230 85.560 274.155 85.890 ;
        RECT 273.230 84.950 273.400 85.560 ;
        RECT 274.325 85.380 274.495 86.070 ;
        RECT 273.665 85.130 274.495 85.380 ;
        RECT 274.665 85.130 275.095 86.820 ;
        RECT 275.265 86.415 275.435 87.065 ;
        RECT 276.560 86.865 276.730 87.435 ;
        RECT 278.355 87.250 278.835 87.920 ;
        RECT 279.890 87.750 280.060 88.350 ;
        RECT 281.050 93.045 283.150 93.215 ;
        RECT 281.050 87.995 281.220 93.045 ;
        RECT 281.850 92.535 282.350 92.705 ;
        RECT 281.620 91.825 281.790 92.365 ;
        RECT 282.410 91.825 282.580 92.365 ;
        RECT 281.850 91.485 282.350 91.655 ;
        RECT 281.620 90.775 281.790 91.315 ;
        RECT 282.410 90.775 282.580 91.315 ;
        RECT 281.850 90.435 282.350 90.605 ;
        RECT 281.620 89.725 281.790 90.265 ;
        RECT 282.410 89.725 282.580 90.265 ;
        RECT 281.850 89.385 282.350 89.555 ;
        RECT 281.620 88.675 281.790 89.215 ;
        RECT 282.410 88.675 282.580 89.215 ;
        RECT 281.850 88.335 282.350 88.505 ;
        RECT 282.980 87.995 283.150 93.045 ;
        RECT 281.050 87.825 283.150 87.995 ;
        RECT 283.510 93.045 285.610 93.215 ;
        RECT 279.005 87.420 280.060 87.750 ;
        RECT 278.355 87.235 279.625 87.250 ;
        RECT 276.995 87.065 279.625 87.235 ;
        RECT 275.605 86.615 277.685 86.865 ;
        RECT 275.265 86.085 276.295 86.415 ;
        RECT 275.265 85.385 275.435 86.085 ;
        RECT 276.560 85.915 276.730 86.615 ;
        RECT 277.855 86.415 278.025 87.065 ;
        RECT 278.665 86.990 279.625 87.065 ;
        RECT 278.795 86.920 279.625 86.990 ;
        RECT 276.995 86.085 278.025 86.415 ;
        RECT 275.605 85.585 277.685 85.915 ;
        RECT 275.265 85.135 276.295 85.385 ;
        RECT 273.230 84.700 274.445 84.950 ;
        RECT 273.230 84.480 273.400 84.700 ;
        RECT 273.230 84.180 274.420 84.480 ;
        RECT 273.230 83.975 273.400 84.180 ;
        RECT 273.230 83.645 274.155 83.975 ;
        RECT 274.730 83.965 274.930 85.130 ;
        RECT 276.560 84.935 276.730 85.585 ;
        RECT 277.855 85.385 278.025 86.085 ;
        RECT 276.995 85.135 278.025 85.385 ;
        RECT 278.195 85.130 278.625 86.820 ;
        RECT 278.795 86.240 278.965 86.920 ;
        RECT 279.890 86.750 280.060 87.420 ;
        RECT 279.135 86.420 280.060 86.750 ;
        RECT 278.795 86.070 279.625 86.240 ;
        RECT 278.795 85.380 278.965 86.070 ;
        RECT 279.890 85.890 280.060 86.420 ;
        RECT 279.135 85.560 280.060 85.890 ;
        RECT 278.795 85.130 279.625 85.380 ;
        RECT 275.135 84.685 278.155 84.935 ;
        RECT 276.560 84.480 276.730 84.685 ;
        RECT 275.520 84.180 277.770 84.480 ;
        RECT 276.560 83.970 276.730 84.180 ;
        RECT 274.325 83.735 275.435 83.965 ;
        RECT 262.010 77.720 264.110 77.890 ;
        RECT 273.230 83.065 273.400 83.645 ;
        RECT 274.325 83.465 274.495 83.735 ;
        RECT 275.265 83.520 275.435 83.735 ;
        RECT 275.605 83.720 277.685 83.970 ;
        RECT 278.365 83.965 278.565 85.130 ;
        RECT 279.890 84.950 280.060 85.560 ;
        RECT 278.845 84.700 280.060 84.950 ;
        RECT 279.890 84.480 280.060 84.700 ;
        RECT 278.870 84.180 280.060 84.480 ;
        RECT 279.890 83.975 280.060 84.180 ;
        RECT 277.855 83.735 278.965 83.965 ;
        RECT 273.665 83.295 274.495 83.465 ;
        RECT 273.230 82.735 274.155 83.065 ;
        RECT 273.230 82.135 273.400 82.735 ;
        RECT 274.325 82.555 274.495 83.295 ;
        RECT 273.665 82.305 274.495 82.555 ;
        RECT 273.230 81.805 274.445 82.135 ;
        RECT 274.665 81.815 275.095 83.490 ;
        RECT 275.265 83.190 276.295 83.520 ;
        RECT 275.265 82.620 275.435 83.190 ;
        RECT 276.560 82.990 276.730 83.720 ;
        RECT 277.855 83.520 278.025 83.735 ;
        RECT 276.995 83.190 278.025 83.520 ;
        RECT 275.605 82.820 277.685 82.990 ;
        RECT 275.265 82.290 276.295 82.620 ;
        RECT 276.560 82.090 276.730 82.820 ;
        RECT 277.855 82.620 278.025 83.190 ;
        RECT 276.995 82.290 278.025 82.620 ;
        RECT 275.265 81.840 278.025 82.090 ;
        RECT 273.230 81.065 273.400 81.805 ;
        RECT 274.730 81.565 274.930 81.815 ;
        RECT 273.665 81.235 276.295 81.565 ;
        RECT 276.560 81.065 276.730 81.840 ;
        RECT 278.195 81.815 278.625 83.490 ;
        RECT 278.795 83.465 278.965 83.735 ;
        RECT 279.135 83.645 280.060 83.975 ;
        RECT 278.795 83.295 279.625 83.465 ;
        RECT 278.795 82.555 278.965 83.295 ;
        RECT 279.890 83.065 280.060 83.645 ;
        RECT 279.135 82.735 280.060 83.065 ;
        RECT 278.795 82.305 279.625 82.555 ;
        RECT 279.890 82.135 280.060 82.735 ;
        RECT 278.360 81.565 278.560 81.815 ;
        RECT 278.845 81.805 280.060 82.135 ;
        RECT 276.995 81.235 279.625 81.565 ;
        RECT 279.890 81.065 280.060 81.805 ;
        RECT 273.230 80.735 274.445 81.065 ;
        RECT 273.230 80.160 273.400 80.735 ;
        RECT 274.615 80.375 275.095 81.065 ;
        RECT 275.265 80.735 278.025 81.065 ;
        RECT 273.230 79.860 274.420 80.160 ;
        RECT 273.230 79.145 273.400 79.860 ;
        RECT 274.680 79.645 274.880 80.375 ;
        RECT 276.560 80.160 276.730 80.735 ;
        RECT 278.195 80.375 278.675 81.065 ;
        RECT 278.845 80.735 280.060 81.065 ;
        RECT 275.520 79.860 277.770 80.160 ;
        RECT 273.665 79.315 276.295 79.645 ;
        RECT 276.560 79.145 276.730 79.860 ;
        RECT 278.410 79.645 278.610 80.375 ;
        RECT 279.890 80.160 280.060 80.735 ;
        RECT 278.870 79.860 280.060 80.160 ;
        RECT 276.995 79.315 279.625 79.645 ;
        RECT 279.890 79.145 280.060 79.860 ;
        RECT 273.230 78.815 274.445 79.145 ;
        RECT 273.230 77.350 273.400 78.815 ;
        RECT 274.615 78.455 275.095 79.145 ;
        RECT 275.265 78.815 278.025 79.145 ;
        RECT 276.560 78.225 276.730 78.815 ;
        RECT 278.195 78.455 278.675 79.145 ;
        RECT 278.845 78.815 280.060 79.145 ;
        RECT 273.665 77.840 274.325 78.170 ;
        RECT 274.495 77.895 274.865 78.225 ;
        RECT 275.135 77.895 278.155 78.225 ;
        RECT 278.425 77.895 278.795 78.225 ;
        RECT 279.890 78.200 280.060 78.815 ;
        RECT 274.155 77.725 274.325 77.840 ;
        RECT 274.155 77.555 276.295 77.725 ;
        RECT 274.495 77.495 276.295 77.555 ;
        RECT 273.230 77.020 274.325 77.350 ;
        RECT 276.560 77.325 276.730 77.895 ;
        RECT 278.965 77.870 280.060 78.200 ;
        RECT 276.995 77.665 278.795 77.725 ;
        RECT 276.995 77.495 279.135 77.665 ;
        RECT 278.965 77.380 279.135 77.495 ;
        RECT 249.175 75.935 250.390 76.265 ;
        RECT 249.175 75.450 249.345 75.935 ;
        RECT 250.560 75.575 251.040 76.265 ;
        RECT 251.210 75.935 252.675 76.265 ;
        RECT 252.505 75.450 252.675 75.935 ;
        RECT 273.230 76.265 273.400 77.020 ;
        RECT 274.495 76.995 274.865 77.325 ;
        RECT 275.135 76.995 278.155 77.325 ;
        RECT 278.425 76.995 278.795 77.325 ;
        RECT 278.965 77.050 279.625 77.380 ;
        RECT 274.600 76.765 274.800 76.995 ;
        RECT 273.665 76.435 276.295 76.765 ;
        RECT 276.560 76.265 276.730 76.995 ;
        RECT 279.890 76.890 280.060 77.870 ;
        RECT 281.050 87.295 283.150 87.465 ;
        RECT 281.050 77.885 281.220 87.295 ;
        RECT 281.850 86.785 282.350 86.955 ;
        RECT 281.620 85.030 281.790 86.570 ;
        RECT 282.410 85.030 282.580 86.570 ;
        RECT 281.850 84.645 282.350 84.815 ;
        RECT 281.620 82.890 281.790 84.430 ;
        RECT 282.410 82.890 282.580 84.430 ;
        RECT 281.850 82.505 282.350 82.675 ;
        RECT 281.620 80.750 281.790 82.290 ;
        RECT 282.410 80.750 282.580 82.290 ;
        RECT 281.850 80.365 282.350 80.535 ;
        RECT 281.620 78.610 281.790 80.150 ;
        RECT 282.410 78.610 282.580 80.150 ;
        RECT 281.850 78.225 282.350 78.395 ;
        RECT 282.980 77.885 283.150 87.295 ;
        RECT 283.510 83.635 283.680 93.045 ;
        RECT 284.310 92.535 284.810 92.705 ;
        RECT 284.080 90.780 284.250 92.320 ;
        RECT 284.870 90.780 285.040 92.320 ;
        RECT 284.310 90.395 284.810 90.565 ;
        RECT 284.080 88.640 284.250 90.180 ;
        RECT 284.870 88.640 285.040 90.180 ;
        RECT 284.310 88.255 284.810 88.425 ;
        RECT 284.080 86.500 284.250 88.040 ;
        RECT 284.870 86.500 285.040 88.040 ;
        RECT 284.310 86.115 284.810 86.285 ;
        RECT 284.080 84.360 284.250 85.900 ;
        RECT 284.870 84.360 285.040 85.900 ;
        RECT 284.310 83.975 284.810 84.145 ;
        RECT 285.440 83.635 285.610 93.045 ;
        RECT 285.970 93.050 288.070 93.220 ;
        RECT 285.970 88.000 286.140 93.050 ;
        RECT 286.770 92.540 287.270 92.710 ;
        RECT 286.540 91.830 286.710 92.370 ;
        RECT 287.330 91.830 287.500 92.370 ;
        RECT 286.770 91.490 287.270 91.660 ;
        RECT 286.540 90.780 286.710 91.320 ;
        RECT 287.330 90.780 287.500 91.320 ;
        RECT 286.770 90.440 287.270 90.610 ;
        RECT 286.540 89.730 286.710 90.270 ;
        RECT 287.330 89.730 287.500 90.270 ;
        RECT 286.770 89.390 287.270 89.560 ;
        RECT 286.540 88.680 286.710 89.220 ;
        RECT 287.330 88.680 287.500 89.220 ;
        RECT 286.770 88.340 287.270 88.510 ;
        RECT 287.900 88.000 288.070 93.050 ;
        RECT 285.970 87.830 288.070 88.000 ;
        RECT 288.430 93.050 292.460 93.220 ;
        RECT 283.510 83.465 285.610 83.635 ;
        RECT 285.970 87.300 288.070 87.470 ;
        RECT 281.050 77.715 283.150 77.885 ;
        RECT 283.510 82.935 285.610 83.105 ;
        RECT 283.510 77.885 283.680 82.935 ;
        RECT 284.310 82.425 284.810 82.595 ;
        RECT 284.080 81.715 284.250 82.255 ;
        RECT 284.870 81.715 285.040 82.255 ;
        RECT 284.310 81.375 284.810 81.545 ;
        RECT 284.080 80.665 284.250 81.205 ;
        RECT 284.870 80.665 285.040 81.205 ;
        RECT 284.310 80.325 284.810 80.495 ;
        RECT 284.080 79.615 284.250 80.155 ;
        RECT 284.870 79.615 285.040 80.155 ;
        RECT 284.310 79.275 284.810 79.445 ;
        RECT 284.080 78.565 284.250 79.105 ;
        RECT 284.870 78.565 285.040 79.105 ;
        RECT 284.310 78.225 284.810 78.395 ;
        RECT 285.440 77.885 285.610 82.935 ;
        RECT 283.510 77.715 285.610 77.885 ;
        RECT 285.970 77.890 286.140 87.300 ;
        RECT 286.770 86.790 287.270 86.960 ;
        RECT 286.540 85.035 286.710 86.575 ;
        RECT 287.330 85.035 287.500 86.575 ;
        RECT 286.770 84.650 287.270 84.820 ;
        RECT 286.540 82.895 286.710 84.435 ;
        RECT 287.330 82.895 287.500 84.435 ;
        RECT 286.770 82.510 287.270 82.680 ;
        RECT 286.540 80.755 286.710 82.295 ;
        RECT 287.330 80.755 287.500 82.295 ;
        RECT 286.770 80.370 287.270 80.540 ;
        RECT 286.540 78.615 286.710 80.155 ;
        RECT 287.330 78.615 287.500 80.155 ;
        RECT 286.770 78.230 287.270 78.400 ;
        RECT 287.900 77.890 288.070 87.300 ;
        RECT 288.430 83.640 288.600 93.050 ;
        RECT 289.230 92.540 289.730 92.710 ;
        RECT 289.000 90.785 289.170 92.325 ;
        RECT 289.790 90.785 289.960 92.325 ;
        RECT 289.230 90.400 289.730 90.570 ;
        RECT 289.000 88.645 289.170 90.185 ;
        RECT 289.790 88.645 289.960 90.185 ;
        RECT 289.230 88.260 289.730 88.430 ;
        RECT 289.000 86.505 289.170 88.045 ;
        RECT 289.790 86.505 289.960 88.045 ;
        RECT 289.230 86.120 289.730 86.290 ;
        RECT 289.000 84.365 289.170 85.905 ;
        RECT 289.790 84.365 289.960 85.905 ;
        RECT 289.230 83.980 289.730 84.150 ;
        RECT 290.360 83.640 290.530 93.050 ;
        RECT 291.160 92.540 291.660 92.710 ;
        RECT 290.930 90.785 291.100 92.325 ;
        RECT 291.720 90.785 291.890 92.325 ;
        RECT 291.160 90.400 291.660 90.570 ;
        RECT 290.930 88.645 291.100 90.185 ;
        RECT 291.720 88.645 291.890 90.185 ;
        RECT 291.160 88.260 291.660 88.430 ;
        RECT 290.930 86.505 291.100 88.045 ;
        RECT 291.720 86.505 291.890 88.045 ;
        RECT 291.160 86.120 291.660 86.290 ;
        RECT 290.930 84.365 291.100 85.905 ;
        RECT 291.720 84.365 291.890 85.905 ;
        RECT 291.160 83.980 291.660 84.150 ;
        RECT 292.290 83.640 292.460 93.050 ;
        RECT 292.820 93.050 296.850 93.220 ;
        RECT 292.820 88.000 292.990 93.050 ;
        RECT 293.620 92.540 294.120 92.710 ;
        RECT 293.390 91.830 293.560 92.370 ;
        RECT 294.180 91.830 294.350 92.370 ;
        RECT 293.620 91.490 294.120 91.660 ;
        RECT 293.390 90.780 293.560 91.320 ;
        RECT 294.180 90.780 294.350 91.320 ;
        RECT 293.620 90.440 294.120 90.610 ;
        RECT 293.390 89.730 293.560 90.270 ;
        RECT 294.180 89.730 294.350 90.270 ;
        RECT 293.620 89.390 294.120 89.560 ;
        RECT 293.390 88.680 293.560 89.220 ;
        RECT 294.180 88.680 294.350 89.220 ;
        RECT 293.620 88.340 294.120 88.510 ;
        RECT 294.750 88.000 294.920 93.050 ;
        RECT 295.550 92.540 296.050 92.710 ;
        RECT 295.320 91.830 295.490 92.370 ;
        RECT 296.110 91.830 296.280 92.370 ;
        RECT 295.550 91.490 296.050 91.660 ;
        RECT 295.320 90.780 295.490 91.320 ;
        RECT 296.110 90.780 296.280 91.320 ;
        RECT 295.550 90.440 296.050 90.610 ;
        RECT 295.320 89.730 295.490 90.270 ;
        RECT 296.110 89.730 296.280 90.270 ;
        RECT 295.550 89.390 296.050 89.560 ;
        RECT 295.320 88.680 295.490 89.220 ;
        RECT 296.110 88.680 296.280 89.220 ;
        RECT 295.550 88.340 296.050 88.510 ;
        RECT 296.680 88.000 296.850 93.050 ;
        RECT 292.820 87.830 296.850 88.000 ;
        RECT 297.190 93.000 297.360 93.210 ;
        RECT 300.520 93.085 300.690 93.210 ;
        RECT 297.190 92.670 298.245 93.000 ;
        RECT 297.190 92.070 297.360 92.670 ;
        RECT 298.415 92.585 298.895 93.085 ;
        RECT 299.095 92.755 302.115 93.085 ;
        RECT 298.415 92.500 300.255 92.585 ;
        RECT 297.625 92.255 300.255 92.500 ;
        RECT 297.625 92.240 298.895 92.255 ;
        RECT 297.190 91.740 298.245 92.070 ;
        RECT 297.190 91.070 297.360 91.740 ;
        RECT 298.415 91.570 298.895 92.240 ;
        RECT 300.520 92.085 300.690 92.755 ;
        RECT 302.315 92.585 302.795 93.085 ;
        RECT 303.850 93.000 304.020 93.210 ;
        RECT 302.965 92.670 304.020 93.000 ;
        RECT 300.955 92.500 302.795 92.585 ;
        RECT 300.955 92.255 303.585 92.500 ;
        RECT 302.315 92.240 303.585 92.255 ;
        RECT 299.095 91.755 302.115 92.085 ;
        RECT 297.625 91.555 298.895 91.570 ;
        RECT 297.625 91.385 300.255 91.555 ;
        RECT 297.625 91.310 298.585 91.385 ;
        RECT 297.625 91.240 298.455 91.310 ;
        RECT 297.190 90.740 298.115 91.070 ;
        RECT 297.190 90.210 297.360 90.740 ;
        RECT 298.285 90.560 298.455 91.240 ;
        RECT 297.625 90.390 298.455 90.560 ;
        RECT 297.190 89.880 298.115 90.210 ;
        RECT 297.190 89.270 297.360 89.880 ;
        RECT 298.285 89.700 298.455 90.390 ;
        RECT 297.625 89.450 298.455 89.700 ;
        RECT 298.625 89.450 299.055 91.140 ;
        RECT 299.225 90.735 299.395 91.385 ;
        RECT 300.520 91.185 300.690 91.755 ;
        RECT 302.315 91.570 302.795 92.240 ;
        RECT 303.850 92.070 304.020 92.670 ;
        RECT 302.965 91.740 304.020 92.070 ;
        RECT 302.315 91.555 303.585 91.570 ;
        RECT 300.955 91.385 303.585 91.555 ;
        RECT 299.565 90.935 301.645 91.185 ;
        RECT 299.225 90.405 300.255 90.735 ;
        RECT 299.225 89.705 299.395 90.405 ;
        RECT 300.520 90.235 300.690 90.935 ;
        RECT 301.815 90.735 301.985 91.385 ;
        RECT 302.625 91.310 303.585 91.385 ;
        RECT 302.755 91.240 303.585 91.310 ;
        RECT 300.955 90.405 301.985 90.735 ;
        RECT 299.565 89.905 301.645 90.235 ;
        RECT 299.225 89.455 300.255 89.705 ;
        RECT 297.190 89.020 298.405 89.270 ;
        RECT 297.190 88.680 297.360 89.020 ;
        RECT 298.690 88.765 298.890 89.450 ;
        RECT 300.520 89.255 300.690 89.905 ;
        RECT 301.815 89.705 301.985 90.405 ;
        RECT 300.955 89.455 301.985 89.705 ;
        RECT 302.155 89.450 302.585 91.140 ;
        RECT 302.755 90.560 302.925 91.240 ;
        RECT 303.850 91.070 304.020 91.740 ;
        RECT 303.095 90.740 304.020 91.070 ;
        RECT 302.755 90.390 303.585 90.560 ;
        RECT 302.755 89.700 302.925 90.390 ;
        RECT 303.850 90.210 304.020 90.740 ;
        RECT 303.095 89.880 304.020 90.210 ;
        RECT 302.755 89.450 303.585 89.700 ;
        RECT 299.095 89.005 302.115 89.255 ;
        RECT 300.520 88.765 300.690 89.005 ;
        RECT 302.320 88.765 302.520 89.450 ;
        RECT 303.850 89.270 304.020 89.880 ;
        RECT 302.805 89.020 304.020 89.270 ;
        RECT 297.190 88.350 298.245 88.680 ;
        RECT 288.430 83.470 292.460 83.640 ;
        RECT 297.190 87.750 297.360 88.350 ;
        RECT 298.415 88.265 298.895 88.765 ;
        RECT 299.095 88.435 302.115 88.765 ;
        RECT 298.415 88.180 300.255 88.265 ;
        RECT 297.625 87.935 300.255 88.180 ;
        RECT 297.625 87.920 298.895 87.935 ;
        RECT 297.190 87.420 298.245 87.750 ;
        RECT 297.190 86.750 297.360 87.420 ;
        RECT 298.415 87.250 298.895 87.920 ;
        RECT 300.520 87.765 300.690 88.435 ;
        RECT 302.315 88.265 302.795 88.765 ;
        RECT 303.850 88.680 304.020 89.020 ;
        RECT 302.965 88.350 304.020 88.680 ;
        RECT 300.955 88.180 302.795 88.265 ;
        RECT 300.955 87.935 303.585 88.180 ;
        RECT 302.315 87.920 303.585 87.935 ;
        RECT 299.095 87.435 302.115 87.765 ;
        RECT 297.625 87.235 298.895 87.250 ;
        RECT 297.625 87.065 300.255 87.235 ;
        RECT 297.625 86.990 298.585 87.065 ;
        RECT 297.625 86.920 298.455 86.990 ;
        RECT 297.190 86.420 298.115 86.750 ;
        RECT 297.190 85.890 297.360 86.420 ;
        RECT 298.285 86.240 298.455 86.920 ;
        RECT 297.625 86.070 298.455 86.240 ;
        RECT 297.190 85.560 298.115 85.890 ;
        RECT 297.190 84.950 297.360 85.560 ;
        RECT 298.285 85.380 298.455 86.070 ;
        RECT 297.625 85.130 298.455 85.380 ;
        RECT 298.625 85.130 299.055 86.820 ;
        RECT 299.225 86.415 299.395 87.065 ;
        RECT 300.520 86.865 300.690 87.435 ;
        RECT 302.315 87.250 302.795 87.920 ;
        RECT 303.850 87.750 304.020 88.350 ;
        RECT 305.060 93.045 307.160 93.215 ;
        RECT 305.060 87.995 305.230 93.045 ;
        RECT 305.860 92.535 306.360 92.705 ;
        RECT 305.630 91.825 305.800 92.365 ;
        RECT 306.420 91.825 306.590 92.365 ;
        RECT 305.860 91.485 306.360 91.655 ;
        RECT 305.630 90.775 305.800 91.315 ;
        RECT 306.420 90.775 306.590 91.315 ;
        RECT 305.860 90.435 306.360 90.605 ;
        RECT 305.630 89.725 305.800 90.265 ;
        RECT 306.420 89.725 306.590 90.265 ;
        RECT 305.860 89.385 306.360 89.555 ;
        RECT 305.630 88.675 305.800 89.215 ;
        RECT 306.420 88.675 306.590 89.215 ;
        RECT 305.860 88.335 306.360 88.505 ;
        RECT 306.990 87.995 307.160 93.045 ;
        RECT 305.060 87.825 307.160 87.995 ;
        RECT 307.520 93.045 309.620 93.215 ;
        RECT 302.965 87.420 304.020 87.750 ;
        RECT 302.315 87.235 303.585 87.250 ;
        RECT 300.955 87.065 303.585 87.235 ;
        RECT 299.565 86.615 301.645 86.865 ;
        RECT 299.225 86.085 300.255 86.415 ;
        RECT 299.225 85.385 299.395 86.085 ;
        RECT 300.520 85.915 300.690 86.615 ;
        RECT 301.815 86.415 301.985 87.065 ;
        RECT 302.625 86.990 303.585 87.065 ;
        RECT 302.755 86.920 303.585 86.990 ;
        RECT 300.955 86.085 301.985 86.415 ;
        RECT 299.565 85.585 301.645 85.915 ;
        RECT 299.225 85.135 300.255 85.385 ;
        RECT 297.190 84.700 298.405 84.950 ;
        RECT 297.190 84.480 297.360 84.700 ;
        RECT 297.190 84.180 298.380 84.480 ;
        RECT 297.190 83.975 297.360 84.180 ;
        RECT 297.190 83.645 298.115 83.975 ;
        RECT 298.690 83.965 298.890 85.130 ;
        RECT 300.520 84.935 300.690 85.585 ;
        RECT 301.815 85.385 301.985 86.085 ;
        RECT 300.955 85.135 301.985 85.385 ;
        RECT 302.155 85.130 302.585 86.820 ;
        RECT 302.755 86.240 302.925 86.920 ;
        RECT 303.850 86.750 304.020 87.420 ;
        RECT 303.095 86.420 304.020 86.750 ;
        RECT 302.755 86.070 303.585 86.240 ;
        RECT 302.755 85.380 302.925 86.070 ;
        RECT 303.850 85.890 304.020 86.420 ;
        RECT 303.095 85.560 304.020 85.890 ;
        RECT 302.755 85.130 303.585 85.380 ;
        RECT 299.095 84.685 302.115 84.935 ;
        RECT 300.520 84.480 300.690 84.685 ;
        RECT 299.480 84.180 301.730 84.480 ;
        RECT 300.520 83.970 300.690 84.180 ;
        RECT 298.285 83.735 299.395 83.965 ;
        RECT 285.970 77.720 288.070 77.890 ;
        RECT 297.190 83.065 297.360 83.645 ;
        RECT 298.285 83.465 298.455 83.735 ;
        RECT 299.225 83.520 299.395 83.735 ;
        RECT 299.565 83.720 301.645 83.970 ;
        RECT 302.325 83.965 302.525 85.130 ;
        RECT 303.850 84.950 304.020 85.560 ;
        RECT 302.805 84.700 304.020 84.950 ;
        RECT 303.850 84.480 304.020 84.700 ;
        RECT 302.830 84.180 304.020 84.480 ;
        RECT 303.850 83.975 304.020 84.180 ;
        RECT 301.815 83.735 302.925 83.965 ;
        RECT 297.625 83.295 298.455 83.465 ;
        RECT 297.190 82.735 298.115 83.065 ;
        RECT 297.190 82.135 297.360 82.735 ;
        RECT 298.285 82.555 298.455 83.295 ;
        RECT 297.625 82.305 298.455 82.555 ;
        RECT 297.190 81.805 298.405 82.135 ;
        RECT 298.625 81.815 299.055 83.490 ;
        RECT 299.225 83.190 300.255 83.520 ;
        RECT 299.225 82.620 299.395 83.190 ;
        RECT 300.520 82.990 300.690 83.720 ;
        RECT 301.815 83.520 301.985 83.735 ;
        RECT 300.955 83.190 301.985 83.520 ;
        RECT 299.565 82.820 301.645 82.990 ;
        RECT 299.225 82.290 300.255 82.620 ;
        RECT 300.520 82.090 300.690 82.820 ;
        RECT 301.815 82.620 301.985 83.190 ;
        RECT 300.955 82.290 301.985 82.620 ;
        RECT 299.225 81.840 301.985 82.090 ;
        RECT 297.190 81.065 297.360 81.805 ;
        RECT 298.690 81.565 298.890 81.815 ;
        RECT 297.625 81.235 300.255 81.565 ;
        RECT 300.520 81.065 300.690 81.840 ;
        RECT 302.155 81.815 302.585 83.490 ;
        RECT 302.755 83.465 302.925 83.735 ;
        RECT 303.095 83.645 304.020 83.975 ;
        RECT 302.755 83.295 303.585 83.465 ;
        RECT 302.755 82.555 302.925 83.295 ;
        RECT 303.850 83.065 304.020 83.645 ;
        RECT 303.095 82.735 304.020 83.065 ;
        RECT 302.755 82.305 303.585 82.555 ;
        RECT 303.850 82.135 304.020 82.735 ;
        RECT 302.320 81.565 302.520 81.815 ;
        RECT 302.805 81.805 304.020 82.135 ;
        RECT 300.955 81.235 303.585 81.565 ;
        RECT 303.850 81.065 304.020 81.805 ;
        RECT 297.190 80.735 298.405 81.065 ;
        RECT 297.190 80.160 297.360 80.735 ;
        RECT 298.575 80.375 299.055 81.065 ;
        RECT 299.225 80.735 301.985 81.065 ;
        RECT 297.190 79.860 298.380 80.160 ;
        RECT 297.190 79.145 297.360 79.860 ;
        RECT 298.640 79.645 298.840 80.375 ;
        RECT 300.520 80.160 300.690 80.735 ;
        RECT 302.155 80.375 302.635 81.065 ;
        RECT 302.805 80.735 304.020 81.065 ;
        RECT 299.480 79.860 301.730 80.160 ;
        RECT 297.625 79.315 300.255 79.645 ;
        RECT 300.520 79.145 300.690 79.860 ;
        RECT 302.370 79.645 302.570 80.375 ;
        RECT 303.850 80.160 304.020 80.735 ;
        RECT 302.830 79.860 304.020 80.160 ;
        RECT 300.955 79.315 303.585 79.645 ;
        RECT 303.850 79.145 304.020 79.860 ;
        RECT 297.190 78.815 298.405 79.145 ;
        RECT 297.190 77.350 297.360 78.815 ;
        RECT 298.575 78.455 299.055 79.145 ;
        RECT 299.225 78.815 301.985 79.145 ;
        RECT 300.520 78.225 300.690 78.815 ;
        RECT 302.155 78.455 302.635 79.145 ;
        RECT 302.805 78.815 304.020 79.145 ;
        RECT 297.625 77.840 298.285 78.170 ;
        RECT 298.455 77.895 298.825 78.225 ;
        RECT 299.095 77.895 302.115 78.225 ;
        RECT 302.385 77.895 302.755 78.225 ;
        RECT 303.850 78.200 304.020 78.815 ;
        RECT 298.115 77.725 298.285 77.840 ;
        RECT 298.115 77.555 300.255 77.725 ;
        RECT 298.455 77.495 300.255 77.555 ;
        RECT 297.190 77.020 298.285 77.350 ;
        RECT 300.520 77.325 300.690 77.895 ;
        RECT 302.925 77.870 304.020 78.200 ;
        RECT 300.955 77.665 302.755 77.725 ;
        RECT 300.955 77.495 303.095 77.665 ;
        RECT 302.925 77.380 303.095 77.495 ;
        RECT 273.230 75.935 274.445 76.265 ;
        RECT 273.230 75.450 273.400 75.935 ;
        RECT 274.615 75.575 275.095 76.265 ;
        RECT 275.265 75.935 276.730 76.265 ;
        RECT 276.560 75.450 276.730 75.935 ;
        RECT 297.190 76.265 297.360 77.020 ;
        RECT 298.455 76.995 298.825 77.325 ;
        RECT 299.095 76.995 302.115 77.325 ;
        RECT 302.385 76.995 302.755 77.325 ;
        RECT 302.925 77.050 303.585 77.380 ;
        RECT 298.560 76.765 298.760 76.995 ;
        RECT 297.625 76.435 300.255 76.765 ;
        RECT 300.520 76.265 300.690 76.995 ;
        RECT 303.850 76.890 304.020 77.870 ;
        RECT 305.060 87.295 307.160 87.465 ;
        RECT 305.060 77.885 305.230 87.295 ;
        RECT 305.860 86.785 306.360 86.955 ;
        RECT 305.630 85.030 305.800 86.570 ;
        RECT 306.420 85.030 306.590 86.570 ;
        RECT 305.860 84.645 306.360 84.815 ;
        RECT 305.630 82.890 305.800 84.430 ;
        RECT 306.420 82.890 306.590 84.430 ;
        RECT 305.860 82.505 306.360 82.675 ;
        RECT 305.630 80.750 305.800 82.290 ;
        RECT 306.420 80.750 306.590 82.290 ;
        RECT 305.860 80.365 306.360 80.535 ;
        RECT 305.630 78.610 305.800 80.150 ;
        RECT 306.420 78.610 306.590 80.150 ;
        RECT 305.860 78.225 306.360 78.395 ;
        RECT 306.990 77.885 307.160 87.295 ;
        RECT 307.520 83.635 307.690 93.045 ;
        RECT 308.320 92.535 308.820 92.705 ;
        RECT 308.090 90.780 308.260 92.320 ;
        RECT 308.880 90.780 309.050 92.320 ;
        RECT 308.320 90.395 308.820 90.565 ;
        RECT 308.090 88.640 308.260 90.180 ;
        RECT 308.880 88.640 309.050 90.180 ;
        RECT 308.320 88.255 308.820 88.425 ;
        RECT 308.090 86.500 308.260 88.040 ;
        RECT 308.880 86.500 309.050 88.040 ;
        RECT 308.320 86.115 308.820 86.285 ;
        RECT 308.090 84.360 308.260 85.900 ;
        RECT 308.880 84.360 309.050 85.900 ;
        RECT 308.320 83.975 308.820 84.145 ;
        RECT 309.450 83.635 309.620 93.045 ;
        RECT 309.980 93.050 312.080 93.220 ;
        RECT 309.980 88.000 310.150 93.050 ;
        RECT 310.780 92.540 311.280 92.710 ;
        RECT 310.550 91.830 310.720 92.370 ;
        RECT 311.340 91.830 311.510 92.370 ;
        RECT 310.780 91.490 311.280 91.660 ;
        RECT 310.550 90.780 310.720 91.320 ;
        RECT 311.340 90.780 311.510 91.320 ;
        RECT 310.780 90.440 311.280 90.610 ;
        RECT 310.550 89.730 310.720 90.270 ;
        RECT 311.340 89.730 311.510 90.270 ;
        RECT 310.780 89.390 311.280 89.560 ;
        RECT 310.550 88.680 310.720 89.220 ;
        RECT 311.340 88.680 311.510 89.220 ;
        RECT 310.780 88.340 311.280 88.510 ;
        RECT 311.910 88.000 312.080 93.050 ;
        RECT 309.980 87.830 312.080 88.000 ;
        RECT 312.440 93.050 316.470 93.220 ;
        RECT 307.520 83.465 309.620 83.635 ;
        RECT 309.980 87.300 312.080 87.470 ;
        RECT 305.060 77.715 307.160 77.885 ;
        RECT 307.520 82.935 309.620 83.105 ;
        RECT 307.520 77.885 307.690 82.935 ;
        RECT 308.320 82.425 308.820 82.595 ;
        RECT 308.090 81.715 308.260 82.255 ;
        RECT 308.880 81.715 309.050 82.255 ;
        RECT 308.320 81.375 308.820 81.545 ;
        RECT 308.090 80.665 308.260 81.205 ;
        RECT 308.880 80.665 309.050 81.205 ;
        RECT 308.320 80.325 308.820 80.495 ;
        RECT 308.090 79.615 308.260 80.155 ;
        RECT 308.880 79.615 309.050 80.155 ;
        RECT 308.320 79.275 308.820 79.445 ;
        RECT 308.090 78.565 308.260 79.105 ;
        RECT 308.880 78.565 309.050 79.105 ;
        RECT 308.320 78.225 308.820 78.395 ;
        RECT 309.450 77.885 309.620 82.935 ;
        RECT 307.520 77.715 309.620 77.885 ;
        RECT 309.980 77.890 310.150 87.300 ;
        RECT 310.780 86.790 311.280 86.960 ;
        RECT 310.550 85.035 310.720 86.575 ;
        RECT 311.340 85.035 311.510 86.575 ;
        RECT 310.780 84.650 311.280 84.820 ;
        RECT 310.550 82.895 310.720 84.435 ;
        RECT 311.340 82.895 311.510 84.435 ;
        RECT 310.780 82.510 311.280 82.680 ;
        RECT 310.550 80.755 310.720 82.295 ;
        RECT 311.340 80.755 311.510 82.295 ;
        RECT 310.780 80.370 311.280 80.540 ;
        RECT 310.550 78.615 310.720 80.155 ;
        RECT 311.340 78.615 311.510 80.155 ;
        RECT 310.780 78.230 311.280 78.400 ;
        RECT 311.910 77.890 312.080 87.300 ;
        RECT 312.440 83.640 312.610 93.050 ;
        RECT 313.240 92.540 313.740 92.710 ;
        RECT 313.010 90.785 313.180 92.325 ;
        RECT 313.800 90.785 313.970 92.325 ;
        RECT 313.240 90.400 313.740 90.570 ;
        RECT 313.010 88.645 313.180 90.185 ;
        RECT 313.800 88.645 313.970 90.185 ;
        RECT 313.240 88.260 313.740 88.430 ;
        RECT 313.010 86.505 313.180 88.045 ;
        RECT 313.800 86.505 313.970 88.045 ;
        RECT 313.240 86.120 313.740 86.290 ;
        RECT 313.010 84.365 313.180 85.905 ;
        RECT 313.800 84.365 313.970 85.905 ;
        RECT 313.240 83.980 313.740 84.150 ;
        RECT 314.370 83.640 314.540 93.050 ;
        RECT 315.170 92.540 315.670 92.710 ;
        RECT 314.940 90.785 315.110 92.325 ;
        RECT 315.730 90.785 315.900 92.325 ;
        RECT 315.170 90.400 315.670 90.570 ;
        RECT 314.940 88.645 315.110 90.185 ;
        RECT 315.730 88.645 315.900 90.185 ;
        RECT 315.170 88.260 315.670 88.430 ;
        RECT 314.940 86.505 315.110 88.045 ;
        RECT 315.730 86.505 315.900 88.045 ;
        RECT 315.170 86.120 315.670 86.290 ;
        RECT 314.940 84.365 315.110 85.905 ;
        RECT 315.730 84.365 315.900 85.905 ;
        RECT 315.170 83.980 315.670 84.150 ;
        RECT 316.300 83.640 316.470 93.050 ;
        RECT 316.830 93.050 320.860 93.220 ;
        RECT 316.830 88.000 317.000 93.050 ;
        RECT 317.630 92.540 318.130 92.710 ;
        RECT 317.400 91.830 317.570 92.370 ;
        RECT 318.190 91.830 318.360 92.370 ;
        RECT 317.630 91.490 318.130 91.660 ;
        RECT 317.400 90.780 317.570 91.320 ;
        RECT 318.190 90.780 318.360 91.320 ;
        RECT 317.630 90.440 318.130 90.610 ;
        RECT 317.400 89.730 317.570 90.270 ;
        RECT 318.190 89.730 318.360 90.270 ;
        RECT 317.630 89.390 318.130 89.560 ;
        RECT 317.400 88.680 317.570 89.220 ;
        RECT 318.190 88.680 318.360 89.220 ;
        RECT 317.630 88.340 318.130 88.510 ;
        RECT 318.760 88.000 318.930 93.050 ;
        RECT 319.560 92.540 320.060 92.710 ;
        RECT 319.330 91.830 319.500 92.370 ;
        RECT 320.120 91.830 320.290 92.370 ;
        RECT 319.560 91.490 320.060 91.660 ;
        RECT 319.330 90.780 319.500 91.320 ;
        RECT 320.120 90.780 320.290 91.320 ;
        RECT 319.560 90.440 320.060 90.610 ;
        RECT 319.330 89.730 319.500 90.270 ;
        RECT 320.120 89.730 320.290 90.270 ;
        RECT 319.560 89.390 320.060 89.560 ;
        RECT 319.330 88.680 319.500 89.220 ;
        RECT 320.120 88.680 320.290 89.220 ;
        RECT 319.560 88.340 320.060 88.510 ;
        RECT 320.690 88.000 320.860 93.050 ;
        RECT 316.830 87.830 320.860 88.000 ;
        RECT 321.200 93.000 321.370 93.210 ;
        RECT 324.530 93.085 324.700 93.210 ;
        RECT 321.200 92.670 322.255 93.000 ;
        RECT 321.200 92.070 321.370 92.670 ;
        RECT 322.425 92.585 322.905 93.085 ;
        RECT 323.105 92.755 326.125 93.085 ;
        RECT 322.425 92.500 324.265 92.585 ;
        RECT 321.635 92.255 324.265 92.500 ;
        RECT 321.635 92.240 322.905 92.255 ;
        RECT 321.200 91.740 322.255 92.070 ;
        RECT 321.200 91.070 321.370 91.740 ;
        RECT 322.425 91.570 322.905 92.240 ;
        RECT 324.530 92.085 324.700 92.755 ;
        RECT 326.325 92.585 326.805 93.085 ;
        RECT 327.860 93.000 328.030 93.210 ;
        RECT 326.975 92.670 328.030 93.000 ;
        RECT 324.965 92.500 326.805 92.585 ;
        RECT 324.965 92.255 327.595 92.500 ;
        RECT 326.325 92.240 327.595 92.255 ;
        RECT 323.105 91.755 326.125 92.085 ;
        RECT 321.635 91.555 322.905 91.570 ;
        RECT 321.635 91.385 324.265 91.555 ;
        RECT 321.635 91.310 322.595 91.385 ;
        RECT 321.635 91.240 322.465 91.310 ;
        RECT 321.200 90.740 322.125 91.070 ;
        RECT 321.200 90.210 321.370 90.740 ;
        RECT 322.295 90.560 322.465 91.240 ;
        RECT 321.635 90.390 322.465 90.560 ;
        RECT 321.200 89.880 322.125 90.210 ;
        RECT 321.200 89.270 321.370 89.880 ;
        RECT 322.295 89.700 322.465 90.390 ;
        RECT 321.635 89.450 322.465 89.700 ;
        RECT 322.635 89.450 323.065 91.140 ;
        RECT 323.235 90.735 323.405 91.385 ;
        RECT 324.530 91.185 324.700 91.755 ;
        RECT 326.325 91.570 326.805 92.240 ;
        RECT 327.860 92.070 328.030 92.670 ;
        RECT 326.975 91.740 328.030 92.070 ;
        RECT 326.325 91.555 327.595 91.570 ;
        RECT 324.965 91.385 327.595 91.555 ;
        RECT 323.575 90.935 325.655 91.185 ;
        RECT 323.235 90.405 324.265 90.735 ;
        RECT 323.235 89.705 323.405 90.405 ;
        RECT 324.530 90.235 324.700 90.935 ;
        RECT 325.825 90.735 325.995 91.385 ;
        RECT 326.635 91.310 327.595 91.385 ;
        RECT 326.765 91.240 327.595 91.310 ;
        RECT 324.965 90.405 325.995 90.735 ;
        RECT 323.575 89.905 325.655 90.235 ;
        RECT 323.235 89.455 324.265 89.705 ;
        RECT 321.200 89.020 322.415 89.270 ;
        RECT 321.200 88.680 321.370 89.020 ;
        RECT 322.700 88.765 322.900 89.450 ;
        RECT 324.530 89.255 324.700 89.905 ;
        RECT 325.825 89.705 325.995 90.405 ;
        RECT 324.965 89.455 325.995 89.705 ;
        RECT 326.165 89.450 326.595 91.140 ;
        RECT 326.765 90.560 326.935 91.240 ;
        RECT 327.860 91.070 328.030 91.740 ;
        RECT 327.105 90.740 328.030 91.070 ;
        RECT 326.765 90.390 327.595 90.560 ;
        RECT 326.765 89.700 326.935 90.390 ;
        RECT 327.860 90.210 328.030 90.740 ;
        RECT 327.105 89.880 328.030 90.210 ;
        RECT 326.765 89.450 327.595 89.700 ;
        RECT 323.105 89.005 326.125 89.255 ;
        RECT 324.530 88.765 324.700 89.005 ;
        RECT 326.330 88.765 326.530 89.450 ;
        RECT 327.860 89.270 328.030 89.880 ;
        RECT 326.815 89.020 328.030 89.270 ;
        RECT 321.200 88.350 322.255 88.680 ;
        RECT 312.440 83.470 316.470 83.640 ;
        RECT 321.200 87.750 321.370 88.350 ;
        RECT 322.425 88.265 322.905 88.765 ;
        RECT 323.105 88.435 326.125 88.765 ;
        RECT 322.425 88.180 324.265 88.265 ;
        RECT 321.635 87.935 324.265 88.180 ;
        RECT 321.635 87.920 322.905 87.935 ;
        RECT 321.200 87.420 322.255 87.750 ;
        RECT 321.200 86.750 321.370 87.420 ;
        RECT 322.425 87.250 322.905 87.920 ;
        RECT 324.530 87.765 324.700 88.435 ;
        RECT 326.325 88.265 326.805 88.765 ;
        RECT 327.860 88.680 328.030 89.020 ;
        RECT 326.975 88.350 328.030 88.680 ;
        RECT 324.965 88.180 326.805 88.265 ;
        RECT 324.965 87.935 327.595 88.180 ;
        RECT 326.325 87.920 327.595 87.935 ;
        RECT 323.105 87.435 326.125 87.765 ;
        RECT 321.635 87.235 322.905 87.250 ;
        RECT 321.635 87.065 324.265 87.235 ;
        RECT 321.635 86.990 322.595 87.065 ;
        RECT 321.635 86.920 322.465 86.990 ;
        RECT 321.200 86.420 322.125 86.750 ;
        RECT 321.200 85.890 321.370 86.420 ;
        RECT 322.295 86.240 322.465 86.920 ;
        RECT 321.635 86.070 322.465 86.240 ;
        RECT 321.200 85.560 322.125 85.890 ;
        RECT 321.200 84.950 321.370 85.560 ;
        RECT 322.295 85.380 322.465 86.070 ;
        RECT 321.635 85.130 322.465 85.380 ;
        RECT 322.635 85.130 323.065 86.820 ;
        RECT 323.235 86.415 323.405 87.065 ;
        RECT 324.530 86.865 324.700 87.435 ;
        RECT 326.325 87.250 326.805 87.920 ;
        RECT 327.860 87.750 328.030 88.350 ;
        RECT 326.975 87.420 328.030 87.750 ;
        RECT 326.325 87.235 327.595 87.250 ;
        RECT 324.965 87.065 327.595 87.235 ;
        RECT 323.575 86.615 325.655 86.865 ;
        RECT 323.235 86.085 324.265 86.415 ;
        RECT 323.235 85.385 323.405 86.085 ;
        RECT 324.530 85.915 324.700 86.615 ;
        RECT 325.825 86.415 325.995 87.065 ;
        RECT 326.635 86.990 327.595 87.065 ;
        RECT 326.765 86.920 327.595 86.990 ;
        RECT 324.965 86.085 325.995 86.415 ;
        RECT 323.575 85.585 325.655 85.915 ;
        RECT 323.235 85.135 324.265 85.385 ;
        RECT 321.200 84.700 322.415 84.950 ;
        RECT 321.200 84.480 321.370 84.700 ;
        RECT 321.200 84.180 322.390 84.480 ;
        RECT 321.200 83.975 321.370 84.180 ;
        RECT 321.200 83.645 322.125 83.975 ;
        RECT 322.700 83.965 322.900 85.130 ;
        RECT 324.530 84.935 324.700 85.585 ;
        RECT 325.825 85.385 325.995 86.085 ;
        RECT 324.965 85.135 325.995 85.385 ;
        RECT 326.165 85.130 326.595 86.820 ;
        RECT 326.765 86.240 326.935 86.920 ;
        RECT 327.860 86.750 328.030 87.420 ;
        RECT 327.105 86.420 328.030 86.750 ;
        RECT 326.765 86.070 327.595 86.240 ;
        RECT 326.765 85.380 326.935 86.070 ;
        RECT 327.860 85.890 328.030 86.420 ;
        RECT 327.105 85.560 328.030 85.890 ;
        RECT 326.765 85.130 327.595 85.380 ;
        RECT 323.105 84.685 326.125 84.935 ;
        RECT 324.530 84.480 324.700 84.685 ;
        RECT 323.490 84.180 325.740 84.480 ;
        RECT 324.530 83.970 324.700 84.180 ;
        RECT 322.295 83.735 323.405 83.965 ;
        RECT 309.980 77.720 312.080 77.890 ;
        RECT 321.200 83.065 321.370 83.645 ;
        RECT 322.295 83.465 322.465 83.735 ;
        RECT 323.235 83.520 323.405 83.735 ;
        RECT 323.575 83.720 325.655 83.970 ;
        RECT 326.335 83.965 326.535 85.130 ;
        RECT 327.860 84.950 328.030 85.560 ;
        RECT 326.815 84.700 328.030 84.950 ;
        RECT 327.860 84.480 328.030 84.700 ;
        RECT 326.840 84.180 328.030 84.480 ;
        RECT 327.860 83.975 328.030 84.180 ;
        RECT 325.825 83.735 326.935 83.965 ;
        RECT 321.635 83.295 322.465 83.465 ;
        RECT 321.200 82.735 322.125 83.065 ;
        RECT 321.200 82.135 321.370 82.735 ;
        RECT 322.295 82.555 322.465 83.295 ;
        RECT 321.635 82.305 322.465 82.555 ;
        RECT 321.200 81.805 322.415 82.135 ;
        RECT 322.635 81.815 323.065 83.490 ;
        RECT 323.235 83.190 324.265 83.520 ;
        RECT 323.235 82.620 323.405 83.190 ;
        RECT 324.530 82.990 324.700 83.720 ;
        RECT 325.825 83.520 325.995 83.735 ;
        RECT 324.965 83.190 325.995 83.520 ;
        RECT 323.575 82.820 325.655 82.990 ;
        RECT 323.235 82.290 324.265 82.620 ;
        RECT 324.530 82.090 324.700 82.820 ;
        RECT 325.825 82.620 325.995 83.190 ;
        RECT 324.965 82.290 325.995 82.620 ;
        RECT 323.235 81.840 325.995 82.090 ;
        RECT 321.200 81.065 321.370 81.805 ;
        RECT 322.700 81.565 322.900 81.815 ;
        RECT 321.635 81.235 324.265 81.565 ;
        RECT 324.530 81.065 324.700 81.840 ;
        RECT 326.165 81.815 326.595 83.490 ;
        RECT 326.765 83.465 326.935 83.735 ;
        RECT 327.105 83.645 328.030 83.975 ;
        RECT 326.765 83.295 327.595 83.465 ;
        RECT 326.765 82.555 326.935 83.295 ;
        RECT 327.860 83.065 328.030 83.645 ;
        RECT 327.105 82.735 328.030 83.065 ;
        RECT 326.765 82.305 327.595 82.555 ;
        RECT 327.860 82.135 328.030 82.735 ;
        RECT 326.330 81.565 326.530 81.815 ;
        RECT 326.815 81.805 328.030 82.135 ;
        RECT 324.965 81.235 327.595 81.565 ;
        RECT 327.860 81.065 328.030 81.805 ;
        RECT 321.200 80.735 322.415 81.065 ;
        RECT 321.200 80.160 321.370 80.735 ;
        RECT 322.585 80.375 323.065 81.065 ;
        RECT 323.235 80.735 325.995 81.065 ;
        RECT 321.200 79.860 322.390 80.160 ;
        RECT 321.200 79.145 321.370 79.860 ;
        RECT 322.650 79.645 322.850 80.375 ;
        RECT 324.530 80.160 324.700 80.735 ;
        RECT 326.165 80.375 326.645 81.065 ;
        RECT 326.815 80.735 328.030 81.065 ;
        RECT 323.490 79.860 325.740 80.160 ;
        RECT 321.635 79.315 324.265 79.645 ;
        RECT 324.530 79.145 324.700 79.860 ;
        RECT 326.380 79.645 326.580 80.375 ;
        RECT 327.860 80.160 328.030 80.735 ;
        RECT 326.840 79.860 328.030 80.160 ;
        RECT 324.965 79.315 327.595 79.645 ;
        RECT 327.860 79.145 328.030 79.860 ;
        RECT 321.200 78.815 322.415 79.145 ;
        RECT 321.200 77.350 321.370 78.815 ;
        RECT 322.585 78.455 323.065 79.145 ;
        RECT 323.235 78.815 325.995 79.145 ;
        RECT 324.530 78.225 324.700 78.815 ;
        RECT 326.165 78.455 326.645 79.145 ;
        RECT 326.815 78.815 328.030 79.145 ;
        RECT 321.635 77.840 322.295 78.170 ;
        RECT 322.465 77.895 322.835 78.225 ;
        RECT 323.105 77.895 326.125 78.225 ;
        RECT 326.395 77.895 326.765 78.225 ;
        RECT 327.860 78.200 328.030 78.815 ;
        RECT 322.125 77.725 322.295 77.840 ;
        RECT 322.125 77.555 324.265 77.725 ;
        RECT 322.465 77.495 324.265 77.555 ;
        RECT 321.200 77.020 322.295 77.350 ;
        RECT 324.530 77.325 324.700 77.895 ;
        RECT 326.935 77.870 328.030 78.200 ;
        RECT 324.965 77.665 326.765 77.725 ;
        RECT 324.965 77.495 327.105 77.665 ;
        RECT 326.935 77.380 327.105 77.495 ;
        RECT 297.190 75.935 298.405 76.265 ;
        RECT 297.190 75.450 297.360 75.935 ;
        RECT 298.575 75.575 299.055 76.265 ;
        RECT 299.225 75.935 300.690 76.265 ;
        RECT 300.520 75.450 300.690 75.935 ;
        RECT 321.200 76.265 321.370 77.020 ;
        RECT 322.465 76.995 322.835 77.325 ;
        RECT 323.105 76.995 326.125 77.325 ;
        RECT 326.395 76.995 326.765 77.325 ;
        RECT 326.935 77.050 327.595 77.380 ;
        RECT 322.570 76.765 322.770 76.995 ;
        RECT 321.635 76.435 324.265 76.765 ;
        RECT 324.530 76.265 324.700 76.995 ;
        RECT 327.860 76.890 328.030 77.870 ;
        RECT 321.200 75.935 322.415 76.265 ;
        RECT 321.200 75.450 321.370 75.935 ;
        RECT 322.585 75.575 323.065 76.265 ;
        RECT 323.235 75.935 324.700 76.265 ;
        RECT 324.530 75.450 324.700 75.935 ;
        RECT 80.470 66.090 80.640 67.235 ;
        RECT 80.905 66.980 82.905 67.150 ;
        RECT 80.905 66.760 82.065 66.980 ;
        RECT 82.235 66.590 82.565 66.810 ;
        RECT 80.905 66.260 81.595 66.590 ;
        RECT 80.470 65.650 81.235 66.090 ;
        RECT 80.470 64.050 80.640 65.650 ;
        RECT 81.425 65.480 81.595 66.260 ;
        RECT 80.905 65.150 81.595 65.480 ;
        RECT 81.765 66.420 82.565 66.590 ;
        RECT 81.765 64.920 81.935 66.420 ;
        RECT 82.735 66.365 82.905 66.980 ;
        RECT 83.800 66.935 83.970 67.235 ;
        RECT 83.140 66.605 83.970 66.935 ;
        RECT 82.105 65.910 82.535 66.240 ;
        RECT 82.735 65.920 83.470 66.365 ;
        RECT 80.905 64.510 81.935 64.920 ;
        RECT 82.190 64.680 82.520 65.910 ;
        RECT 83.800 65.545 83.970 66.605 ;
        RECT 82.690 65.215 83.970 65.545 ;
        RECT 82.845 64.510 83.175 65.035 ;
        RECT 80.905 64.340 83.175 64.510 ;
        RECT 83.800 64.170 83.970 65.215 ;
        RECT 80.470 63.720 81.945 64.050 ;
        RECT 80.470 63.305 80.640 63.720 ;
        RECT 82.270 63.500 82.705 64.170 ;
        RECT 82.895 63.570 83.970 64.170 ;
        RECT 83.800 63.305 83.970 63.570 ;
        RECT 80.470 63.005 81.680 63.305 ;
        RECT 82.780 63.005 83.970 63.305 ;
        RECT 80.470 62.810 80.640 63.005 ;
        RECT 80.470 62.480 82.065 62.810 ;
        RECT 82.335 62.480 82.705 62.810 ;
        RECT 80.470 61.910 80.640 62.480 ;
        RECT 82.875 62.425 83.535 62.755 ;
        RECT 82.875 62.310 83.045 62.425 ;
        RECT 80.905 62.140 83.045 62.310 ;
        RECT 80.905 62.080 82.705 62.140 ;
        RECT 83.800 61.935 83.970 63.005 ;
        RECT 80.470 61.580 82.065 61.910 ;
        RECT 82.335 61.580 82.705 61.910 ;
        RECT 82.875 61.605 83.970 61.935 ;
        RECT 80.470 61.370 80.640 61.580 ;
        RECT 80.470 61.040 82.065 61.370 ;
        RECT 82.335 61.040 82.705 61.370 ;
        RECT 80.470 60.470 80.640 61.040 ;
        RECT 82.875 60.985 83.535 61.315 ;
        RECT 82.875 60.870 83.045 60.985 ;
        RECT 80.905 60.700 83.045 60.870 ;
        RECT 80.905 60.640 82.705 60.700 ;
        RECT 83.800 60.495 83.970 61.605 ;
        RECT 80.470 60.140 82.065 60.470 ;
        RECT 82.335 60.140 82.705 60.470 ;
        RECT 82.875 60.165 83.970 60.495 ;
        RECT 80.470 60.035 80.640 60.140 ;
        RECT 83.800 60.035 83.970 60.165 ;
        RECT 74.620 56.810 74.790 58.515 ;
        RECT 76.160 57.930 76.490 58.260 ;
        RECT 76.685 57.930 77.015 58.260 ;
        RECT 76.320 57.690 76.490 57.930 ;
        RECT 80.470 57.690 80.640 58.515 ;
        RECT 84.095 57.930 84.425 58.260 ;
        RECT 84.620 57.930 84.950 58.260 ;
        RECT 84.620 57.690 84.790 57.930 ;
        RECT 75.240 57.520 76.685 57.690 ;
        RECT 76.980 57.520 84.130 57.690 ;
        RECT 84.425 57.520 85.870 57.690 ;
        RECT 76.515 57.250 76.685 57.520 ;
        RECT 75.240 57.080 76.280 57.250 ;
        RECT 76.515 57.080 80.020 57.250 ;
        RECT 74.620 56.640 76.280 56.810 ;
        RECT 76.980 56.640 80.020 56.810 ;
        RECT 74.620 56.300 74.790 56.640 ;
        RECT 80.470 56.370 80.640 57.520 ;
        RECT 84.425 57.250 84.595 57.520 ;
        RECT 81.090 57.080 84.595 57.250 ;
        RECT 84.830 57.080 85.870 57.250 ;
        RECT 86.320 56.810 86.490 58.515 ;
        RECT 81.090 56.640 84.130 56.810 ;
        RECT 84.830 56.640 86.490 56.810 ;
        RECT 74.620 56.130 76.110 56.300 ;
        RECT 76.980 56.200 84.130 56.370 ;
        RECT 86.320 56.300 86.490 56.640 ;
        RECT 74.620 54.845 74.790 56.130 ;
        RECT 80.470 55.860 80.640 56.200 ;
        RECT 85.000 56.130 86.490 56.300 ;
        RECT 77.150 55.690 83.960 55.860 ;
        RECT 75.940 55.180 76.270 55.510 ;
        RECT 76.685 55.180 77.015 55.510 ;
        RECT 80.470 54.845 80.640 55.690 ;
        RECT 84.095 55.180 84.425 55.510 ;
        RECT 84.840 55.180 85.170 55.510 ;
        RECT 86.320 54.845 86.490 56.130 ;
        RECT 73.550 50.095 73.720 53.395 ;
        RECT 75.300 52.235 75.470 52.965 ;
        RECT 76.855 52.880 77.025 53.050 ;
        RECT 75.855 52.710 78.365 52.880 ;
        RECT 75.855 52.405 76.565 52.710 ;
        RECT 76.735 52.315 77.065 52.540 ;
        RECT 77.235 52.485 78.365 52.710 ;
        RECT 75.300 51.905 76.395 52.235 ;
        RECT 76.735 52.145 77.405 52.315 ;
        RECT 78.630 52.285 78.800 52.965 ;
        RECT 75.300 50.095 75.470 51.905 ;
        RECT 76.565 51.640 77.065 51.970 ;
        RECT 77.235 51.750 77.405 52.145 ;
        RECT 77.575 51.955 78.800 52.285 ;
        RECT 77.235 51.420 78.385 51.750 ;
        RECT 75.640 50.670 76.055 51.400 ;
        RECT 77.235 51.155 77.405 51.420 ;
        RECT 78.630 51.250 78.800 51.955 ;
        RECT 76.225 50.825 77.405 51.155 ;
        RECT 77.575 50.915 78.800 51.250 ;
        RECT 73.550 49.925 75.505 50.095 ;
        RECT 73.550 48.295 73.720 49.925 ;
        RECT 75.705 49.585 75.875 50.670 ;
        RECT 78.630 50.095 78.800 50.915 ;
        RECT 80.470 50.095 80.640 53.395 ;
        RECT 82.310 52.285 82.480 52.965 ;
        RECT 84.085 52.880 84.255 53.050 ;
        RECT 82.745 52.710 85.255 52.880 ;
        RECT 82.745 52.485 83.875 52.710 ;
        RECT 84.045 52.315 84.375 52.540 ;
        RECT 84.545 52.405 85.255 52.710 ;
        RECT 82.310 51.955 83.535 52.285 ;
        RECT 83.705 52.145 84.375 52.315 ;
        RECT 85.640 52.235 85.810 52.965 ;
        RECT 82.310 51.250 82.480 51.955 ;
        RECT 83.705 51.750 83.875 52.145 ;
        RECT 82.725 51.420 83.875 51.750 ;
        RECT 84.045 51.640 84.545 51.970 ;
        RECT 84.715 51.905 85.810 52.235 ;
        RECT 82.310 50.915 83.535 51.250 ;
        RECT 83.705 51.155 83.875 51.420 ;
        RECT 82.310 50.095 82.480 50.915 ;
        RECT 83.705 50.825 84.885 51.155 ;
        RECT 85.055 50.670 85.470 51.400 ;
        RECT 76.305 49.925 84.805 50.095 ;
        RECT 74.465 49.415 79.345 49.585 ;
        RECT 73.550 48.125 75.505 48.295 ;
        RECT 73.550 45.205 73.720 48.125 ;
        RECT 74.125 47.275 74.295 47.855 ;
        RECT 74.465 46.835 75.505 47.005 ;
        RECT 75.920 45.715 76.090 49.145 ;
        RECT 76.305 48.125 79.345 48.295 ;
        RECT 79.560 47.275 79.730 47.855 ;
        RECT 80.470 47.005 80.640 49.925 ;
        RECT 85.235 49.585 85.405 50.670 ;
        RECT 85.640 50.095 85.810 51.905 ;
        RECT 87.390 50.095 87.560 53.395 ;
        RECT 85.605 49.925 87.560 50.095 ;
        RECT 81.765 49.415 86.645 49.585 ;
        RECT 81.765 48.125 84.805 48.295 ;
        RECT 81.380 47.275 81.550 47.855 ;
        RECT 76.305 46.835 84.805 47.005 ;
        RECT 79.560 45.985 79.730 46.565 ;
        RECT 74.465 45.545 79.345 45.715 ;
        RECT 80.470 45.205 80.640 46.835 ;
        RECT 81.380 45.985 81.550 46.565 ;
        RECT 85.020 45.715 85.190 49.145 ;
        RECT 87.390 48.295 87.560 49.925 ;
        RECT 85.605 48.125 87.560 48.295 ;
        RECT 86.815 47.275 86.985 47.855 ;
        RECT 85.605 46.835 86.645 47.005 ;
        RECT 81.765 45.545 86.645 45.715 ;
        RECT 87.390 45.205 87.560 48.125 ;
        RECT 73.550 45.035 75.505 45.205 ;
        RECT 76.305 45.035 84.805 45.205 ;
        RECT 85.605 45.035 87.560 45.205 ;
        RECT 73.550 44.755 73.720 45.035 ;
        RECT 80.470 44.755 80.640 45.035 ;
        RECT 87.390 44.755 87.560 45.035 ;
        RECT 44.610 39.230 55.650 39.400 ;
        RECT 105.470 39.230 116.510 39.400 ;
        RECT 44.700 38.190 45.000 39.230 ;
        RECT 45.205 37.935 45.455 39.230 ;
        RECT 45.655 38.105 45.985 38.965 ;
        RECT 46.185 38.275 46.355 39.230 ;
        RECT 46.555 38.105 46.885 38.965 ;
        RECT 47.085 38.275 47.255 39.230 ;
        RECT 47.455 38.105 47.785 38.965 ;
        RECT 47.955 38.275 48.205 39.230 ;
        RECT 45.655 37.935 48.230 38.105 ;
        RECT 45.215 37.335 47.875 37.765 ;
        RECT 48.060 37.165 48.230 37.935 ;
        RECT 48.405 37.235 48.670 38.965 ;
        RECT 48.935 37.950 49.105 39.230 ;
        RECT 48.840 37.285 49.150 37.765 ;
        RECT 44.700 36.070 45.000 37.090 ;
        RECT 45.205 36.070 45.535 37.115 ;
        RECT 45.705 36.995 48.230 37.165 ;
        RECT 45.705 36.335 45.955 36.995 ;
        RECT 46.170 36.070 46.500 36.825 ;
        RECT 46.680 36.335 46.850 36.995 ;
        RECT 47.030 36.070 47.360 36.825 ;
        RECT 47.540 36.335 47.710 36.995 ;
        RECT 47.890 36.070 48.220 36.825 ;
        RECT 48.400 36.335 48.650 37.235 ;
        RECT 49.320 37.115 49.590 38.965 ;
        RECT 49.835 37.950 50.005 39.230 ;
        RECT 49.760 37.285 50.070 37.765 ;
        RECT 50.240 37.360 50.535 38.965 ;
        RECT 50.735 37.950 50.905 39.230 ;
        RECT 51.105 37.885 51.435 38.965 ;
        RECT 51.635 37.950 51.805 39.230 ;
        RECT 50.785 37.715 50.975 37.765 ;
        RECT 50.240 37.190 50.615 37.360 ;
        RECT 50.785 37.285 51.095 37.715 ;
        RECT 48.820 36.070 49.150 37.115 ;
        RECT 49.320 36.335 49.650 37.115 ;
        RECT 49.820 36.070 50.150 37.020 ;
        RECT 50.320 36.335 50.615 37.190 ;
        RECT 51.265 37.115 51.435 37.885 ;
        RECT 52.085 37.805 52.340 38.965 ;
        RECT 52.535 37.950 52.705 39.230 ;
        RECT 51.605 37.640 51.915 37.765 ;
        RECT 51.605 37.285 51.995 37.640 ;
        RECT 52.170 37.115 52.340 37.805 ;
        RECT 52.510 37.285 52.805 37.765 ;
        RECT 52.975 37.340 53.235 38.965 ;
        RECT 53.435 37.950 53.685 39.230 ;
        RECT 52.975 37.170 53.305 37.340 ;
        RECT 53.475 37.285 53.760 37.765 ;
        RECT 50.820 36.070 51.095 37.115 ;
        RECT 51.265 36.335 51.650 37.115 ;
        RECT 51.830 36.070 52.000 37.115 ;
        RECT 52.170 36.335 52.430 37.115 ;
        RECT 52.690 36.070 52.860 37.000 ;
        RECT 53.040 36.335 53.305 37.170 ;
        RECT 53.550 36.070 53.755 37.115 ;
        RECT 53.930 36.335 54.185 38.965 ;
        RECT 54.385 37.950 54.555 39.230 ;
        RECT 54.355 37.285 54.665 37.765 ;
        RECT 54.365 36.070 54.660 37.115 ;
        RECT 54.835 36.335 55.090 38.965 ;
        RECT 55.285 37.805 55.535 39.230 ;
        RECT 105.585 37.805 105.835 39.230 ;
        RECT 55.270 36.070 55.520 37.115 ;
        RECT 105.600 36.070 105.850 37.115 ;
        RECT 106.030 36.335 106.285 38.965 ;
        RECT 106.565 37.950 106.735 39.230 ;
        RECT 106.455 37.285 106.765 37.765 ;
        RECT 106.460 36.070 106.755 37.115 ;
        RECT 106.935 36.335 107.190 38.965 ;
        RECT 107.435 37.950 107.685 39.230 ;
        RECT 107.360 37.285 107.645 37.765 ;
        RECT 107.885 37.340 108.145 38.965 ;
        RECT 108.415 37.950 108.585 39.230 ;
        RECT 108.780 37.805 109.035 38.965 ;
        RECT 109.315 37.950 109.485 39.230 ;
        RECT 109.685 37.885 110.015 38.965 ;
        RECT 110.215 37.950 110.385 39.230 ;
        RECT 107.815 37.170 108.145 37.340 ;
        RECT 108.315 37.285 108.610 37.765 ;
        RECT 107.365 36.070 107.570 37.115 ;
        RECT 107.815 36.335 108.080 37.170 ;
        RECT 108.780 37.115 108.950 37.805 ;
        RECT 109.205 37.640 109.515 37.765 ;
        RECT 109.125 37.285 109.515 37.640 ;
        RECT 109.685 37.115 109.855 37.885 ;
        RECT 110.145 37.715 110.335 37.765 ;
        RECT 110.025 37.285 110.335 37.715 ;
        RECT 110.585 37.360 110.880 38.965 ;
        RECT 111.115 37.950 111.285 39.230 ;
        RECT 110.505 37.190 110.880 37.360 ;
        RECT 111.050 37.285 111.360 37.765 ;
        RECT 108.260 36.070 108.430 37.000 ;
        RECT 108.690 36.335 108.950 37.115 ;
        RECT 109.120 36.070 109.290 37.115 ;
        RECT 109.470 36.335 109.855 37.115 ;
        RECT 110.025 36.070 110.300 37.115 ;
        RECT 110.505 36.335 110.800 37.190 ;
        RECT 111.530 37.115 111.800 38.965 ;
        RECT 112.015 37.950 112.185 39.230 ;
        RECT 111.970 37.285 112.280 37.765 ;
        RECT 112.450 37.235 112.715 38.965 ;
        RECT 112.915 38.275 113.165 39.230 ;
        RECT 113.335 38.105 113.665 38.965 ;
        RECT 113.865 38.275 114.035 39.230 ;
        RECT 114.235 38.105 114.565 38.965 ;
        RECT 114.765 38.275 114.935 39.230 ;
        RECT 115.135 38.105 115.465 38.965 ;
        RECT 112.890 37.935 115.465 38.105 ;
        RECT 115.665 37.935 115.915 39.230 ;
        RECT 116.120 38.190 116.420 39.230 ;
        RECT 110.970 36.070 111.300 37.020 ;
        RECT 111.470 36.335 111.800 37.115 ;
        RECT 111.970 36.070 112.300 37.115 ;
        RECT 112.470 36.335 112.720 37.235 ;
        RECT 112.890 37.165 113.060 37.935 ;
        RECT 113.245 37.335 115.905 37.765 ;
        RECT 112.890 36.995 115.415 37.165 ;
        RECT 112.900 36.070 113.230 36.825 ;
        RECT 113.410 36.335 113.580 36.995 ;
        RECT 113.760 36.070 114.090 36.825 ;
        RECT 114.270 36.335 114.440 36.995 ;
        RECT 114.620 36.070 114.950 36.825 ;
        RECT 115.165 36.335 115.415 36.995 ;
        RECT 115.585 36.070 115.915 37.115 ;
        RECT 116.120 36.070 116.420 37.090 ;
        RECT 16.805 35.900 58.375 36.070 ;
        RECT 50.320 33.840 53.650 34.010 ;
        RECT 50.320 30.750 50.490 33.840 ;
        RECT 51.030 33.330 51.360 33.500 ;
        RECT 50.890 31.120 51.060 33.160 ;
        RECT 51.330 31.120 51.500 33.160 ;
        RECT 51.900 30.750 52.070 33.840 ;
        RECT 52.610 33.330 52.940 33.500 ;
        RECT 50.320 30.580 52.070 30.750 ;
        RECT 51.900 25.250 52.070 30.580 ;
        RECT 52.470 25.620 52.640 33.160 ;
        RECT 52.910 25.620 53.080 33.160 ;
        RECT 53.480 30.510 53.650 33.840 ;
        RECT 58.205 33.645 58.375 35.900 ;
        RECT 102.745 35.900 144.315 36.070 ;
        RECT 80.475 33.645 80.645 33.825 ;
        RECT 102.745 33.645 102.915 35.900 ;
        RECT 58.205 33.475 102.915 33.645 ;
        RECT 58.205 32.065 58.375 33.475 ;
        RECT 58.710 32.065 58.880 33.475 ;
        RECT 59.220 32.605 59.390 32.935 ;
        RECT 59.560 32.905 79.600 33.075 ;
        RECT 59.560 32.465 79.600 32.635 ;
        RECT 79.970 32.065 80.140 33.475 ;
        RECT 80.475 32.065 80.645 33.475 ;
        RECT 80.980 32.065 81.150 33.475 ;
        RECT 81.520 32.905 101.560 33.075 ;
        RECT 81.520 32.465 101.560 32.635 ;
        RECT 101.730 32.605 101.900 32.935 ;
        RECT 102.240 32.065 102.410 33.475 ;
        RECT 102.745 32.065 102.915 33.475 ;
        RECT 58.205 31.895 102.915 32.065 ;
        RECT 53.480 30.340 55.230 30.510 ;
        RECT 53.480 25.250 53.650 30.340 ;
        RECT 54.050 25.930 54.220 29.970 ;
        RECT 54.490 25.930 54.660 29.970 ;
        RECT 54.190 25.590 54.520 25.760 ;
        RECT 55.060 25.250 55.230 30.340 ;
        RECT 58.205 30.485 58.375 31.895 ;
        RECT 58.710 30.485 58.880 31.895 ;
        RECT 59.220 31.025 59.390 31.355 ;
        RECT 59.560 31.325 79.600 31.495 ;
        RECT 59.560 30.885 79.600 31.055 ;
        RECT 79.970 30.485 80.140 31.895 ;
        RECT 80.475 30.485 80.645 31.895 ;
        RECT 80.980 30.485 81.150 31.895 ;
        RECT 81.520 31.325 101.560 31.495 ;
        RECT 81.520 30.885 101.560 31.055 ;
        RECT 101.730 31.025 101.900 31.355 ;
        RECT 102.240 30.485 102.410 31.895 ;
        RECT 102.745 30.485 102.915 31.895 ;
        RECT 107.470 33.840 110.800 34.010 ;
        RECT 107.470 30.510 107.640 33.840 ;
        RECT 108.180 33.330 108.510 33.500 ;
        RECT 58.205 30.315 102.915 30.485 ;
        RECT 58.205 28.905 58.375 30.315 ;
        RECT 58.710 28.905 58.880 30.315 ;
        RECT 59.220 29.445 59.390 29.775 ;
        RECT 59.560 29.745 79.600 29.915 ;
        RECT 59.560 29.305 79.600 29.475 ;
        RECT 79.970 28.905 80.140 30.315 ;
        RECT 80.475 28.905 80.645 30.315 ;
        RECT 80.980 28.905 81.150 30.315 ;
        RECT 81.520 29.745 101.560 29.915 ;
        RECT 81.520 29.305 101.560 29.475 ;
        RECT 101.730 29.445 101.900 29.775 ;
        RECT 102.240 28.905 102.410 30.315 ;
        RECT 102.745 28.905 102.915 30.315 ;
        RECT 58.205 28.735 102.915 28.905 ;
        RECT 58.205 28.555 58.375 28.735 ;
        RECT 80.475 28.555 80.645 28.735 ;
        RECT 102.745 28.555 102.915 28.735 ;
        RECT 105.890 30.340 107.640 30.510 ;
        RECT 51.900 25.080 55.230 25.250 ;
        RECT 51.900 18.250 52.070 25.080 ;
        RECT 50.320 18.080 52.070 18.250 ;
        RECT 50.320 16.490 50.490 18.080 ;
        RECT 50.890 17.170 51.060 17.710 ;
        RECT 51.330 17.170 51.500 17.710 ;
        RECT 51.030 16.830 51.360 17.000 ;
        RECT 51.900 16.490 52.070 18.080 ;
        RECT 52.470 17.170 52.640 24.710 ;
        RECT 52.910 17.170 53.080 24.710 ;
        RECT 53.480 19.990 53.650 25.080 ;
        RECT 54.190 24.570 54.520 24.740 ;
        RECT 54.050 20.360 54.220 24.400 ;
        RECT 54.490 20.360 54.660 24.400 ;
        RECT 55.060 19.990 55.230 25.080 ;
        RECT 53.480 19.820 55.230 19.990 ;
        RECT 105.890 25.250 106.060 30.340 ;
        RECT 106.460 25.930 106.630 29.970 ;
        RECT 106.900 25.930 107.070 29.970 ;
        RECT 106.600 25.590 106.930 25.760 ;
        RECT 107.470 25.250 107.640 30.340 ;
        RECT 108.040 25.620 108.210 33.160 ;
        RECT 108.480 25.620 108.650 33.160 ;
        RECT 109.050 30.750 109.220 33.840 ;
        RECT 109.760 33.330 110.090 33.500 ;
        RECT 109.620 31.120 109.790 33.160 ;
        RECT 110.060 31.120 110.230 33.160 ;
        RECT 110.630 30.750 110.800 33.840 ;
        RECT 109.050 30.580 110.800 30.750 ;
        RECT 109.050 25.250 109.220 30.580 ;
        RECT 105.890 25.080 109.220 25.250 ;
        RECT 105.890 19.990 106.060 25.080 ;
        RECT 106.600 24.570 106.930 24.740 ;
        RECT 106.460 20.360 106.630 24.400 ;
        RECT 106.900 20.360 107.070 24.400 ;
        RECT 107.470 19.990 107.640 25.080 ;
        RECT 105.890 19.820 107.640 19.990 ;
        RECT 52.610 16.830 52.940 17.000 ;
        RECT 53.480 16.490 53.650 19.820 ;
        RECT 50.320 16.320 53.650 16.490 ;
        RECT 62.830 18.980 75.120 19.150 ;
        RECT 50.320 15.790 52.070 15.960 ;
        RECT 50.320 13.900 50.490 15.790 ;
        RECT 51.030 15.275 51.360 15.445 ;
        RECT 50.890 14.270 51.060 15.060 ;
        RECT 51.330 14.270 51.500 15.060 ;
        RECT 51.900 13.900 52.070 15.790 ;
        RECT 50.320 13.730 52.070 13.900 ;
        RECT 50.800 6.000 51.590 13.730 ;
        RECT 62.830 7.030 63.000 18.980 ;
        RECT 67.430 15.790 70.760 15.960 ;
        RECT 67.430 10.650 67.600 15.790 ;
        RECT 68.000 11.380 68.170 15.420 ;
        RECT 68.440 11.380 68.610 15.420 ;
        RECT 69.010 12.650 69.180 15.790 ;
        RECT 69.720 15.275 70.050 15.445 ;
        RECT 69.580 13.020 69.750 15.060 ;
        RECT 70.020 13.020 70.190 15.060 ;
        RECT 70.590 12.650 70.760 15.790 ;
        RECT 69.010 12.480 70.760 12.650 ;
        RECT 68.140 10.995 68.470 11.165 ;
        RECT 69.010 10.650 69.180 12.480 ;
        RECT 67.430 10.480 69.180 10.650 ;
        RECT 74.950 7.030 75.120 18.980 ;
        RECT 62.830 6.860 75.120 7.030 ;
        RECT 86.005 18.945 98.235 19.115 ;
        RECT 86.005 7.055 86.175 18.945 ;
        RECT 90.360 15.790 93.690 15.960 ;
        RECT 90.360 12.650 90.530 15.790 ;
        RECT 91.070 15.275 91.400 15.445 ;
        RECT 90.930 13.020 91.100 15.060 ;
        RECT 91.370 13.020 91.540 15.060 ;
        RECT 91.940 12.650 92.110 15.790 ;
        RECT 90.360 12.480 92.110 12.650 ;
        RECT 91.940 10.650 92.110 12.480 ;
        RECT 92.510 11.380 92.680 15.420 ;
        RECT 92.950 11.380 93.120 15.420 ;
        RECT 92.650 10.995 92.980 11.165 ;
        RECT 93.520 10.650 93.690 15.790 ;
        RECT 91.940 10.480 93.690 10.650 ;
        RECT 98.065 7.055 98.235 18.945 ;
        RECT 107.470 16.490 107.640 19.820 ;
        RECT 108.040 17.170 108.210 24.710 ;
        RECT 108.480 17.170 108.650 24.710 ;
        RECT 109.050 18.250 109.220 25.080 ;
        RECT 109.050 18.080 110.800 18.250 ;
        RECT 108.180 16.830 108.510 17.000 ;
        RECT 109.050 16.490 109.220 18.080 ;
        RECT 109.620 17.170 109.790 17.710 ;
        RECT 110.060 17.170 110.230 17.710 ;
        RECT 109.760 16.830 110.090 17.000 ;
        RECT 110.630 16.490 110.800 18.080 ;
        RECT 107.470 16.320 110.800 16.490 ;
        RECT 109.050 15.790 110.800 15.960 ;
        RECT 109.050 13.900 109.220 15.790 ;
        RECT 109.760 15.275 110.090 15.445 ;
        RECT 109.620 14.270 109.790 15.060 ;
        RECT 110.060 14.270 110.230 15.060 ;
        RECT 110.630 13.900 110.800 15.790 ;
        RECT 109.050 13.730 110.800 13.900 ;
        RECT 86.005 6.885 98.235 7.055 ;
        RECT 109.530 6.000 110.320 13.730 ;
        RECT 16.805 5.830 58.050 6.000 ;
        RECT 103.070 5.830 144.315 6.000 ;
      LAYER met1 ;
        RECT 134.530 232.470 135.110 232.950 ;
        RECT 241.475 214.400 249.115 214.880 ;
        RECT 241.475 203.600 249.115 204.080 ;
        RECT 241.475 200.000 249.115 200.480 ;
        RECT 248.535 195.860 254.135 196.340 ;
        RECT 241.475 194.060 252.535 194.540 ;
        RECT 241.475 192.260 253.335 192.740 ;
        RECT 248.535 190.460 252.535 190.940 ;
        RECT 241.475 189.200 249.115 189.680 ;
        RECT 241.475 182.000 249.115 182.480 ;
        RECT 241.475 171.200 249.115 171.680 ;
        RECT 112.800 162.680 330.185 163.200 ;
        RECT 112.800 161.640 330.185 162.160 ;
        RECT 112.800 160.600 330.185 161.120 ;
        RECT 112.800 159.560 330.185 160.080 ;
        RECT 112.800 158.520 330.185 159.040 ;
        RECT 112.800 157.480 330.185 158.000 ;
        RECT 112.800 156.440 330.185 156.960 ;
        RECT 112.800 155.400 330.185 155.920 ;
        RECT 112.800 154.360 330.185 154.880 ;
        RECT 111.750 153.320 330.185 153.840 ;
        RECT 10.200 143.375 69.720 143.865 ;
        RECT 62.120 143.135 62.440 143.195 ;
        RECT 48.290 142.995 62.440 143.135 ;
        RECT 32.450 142.625 41.230 142.765 ;
        RECT 13.640 142.395 13.960 142.455 ;
        RECT 15.095 142.395 15.385 142.440 ;
        RECT 13.640 142.255 15.385 142.395 ;
        RECT 13.640 142.195 13.960 142.255 ;
        RECT 15.095 142.210 15.385 142.255 ;
        RECT 20.840 142.195 21.160 142.455 ;
        RECT 24.215 142.395 24.505 142.440 ;
        RECT 32.450 142.395 32.590 142.625 ;
        RECT 24.215 142.255 32.590 142.395 ;
        RECT 35.240 142.395 35.560 142.455 ;
        RECT 41.090 142.440 41.230 142.625 ;
        RECT 38.135 142.395 38.425 142.440 ;
        RECT 35.240 142.255 38.425 142.395 ;
        RECT 24.215 142.210 24.505 142.255 ;
        RECT 35.240 142.195 35.560 142.255 ;
        RECT 38.135 142.210 38.425 142.255 ;
        RECT 41.015 142.210 41.305 142.440 ;
        RECT 43.880 142.195 44.200 142.455 ;
        RECT 48.290 142.440 48.430 142.995 ;
        RECT 62.120 142.935 62.440 142.995 ;
        RECT 65.495 142.765 65.785 142.810 ;
        RECT 61.250 142.625 65.785 142.765 ;
        RECT 48.215 142.210 48.505 142.440 ;
        RECT 50.120 142.195 50.440 142.455 ;
        RECT 51.080 142.395 51.400 142.455 ;
        RECT 61.250 142.440 61.390 142.625 ;
        RECT 65.495 142.580 65.785 142.625 ;
        RECT 55.415 142.395 55.705 142.440 ;
        RECT 51.080 142.255 55.705 142.395 ;
        RECT 51.080 142.195 51.400 142.255 ;
        RECT 55.415 142.210 55.705 142.255 ;
        RECT 61.175 142.210 61.465 142.440 ;
        RECT 63.095 142.395 63.385 142.440 ;
        RECT 65.960 142.395 66.280 142.455 ;
        RECT 61.730 142.255 63.385 142.395 ;
        RECT 17.975 141.840 18.265 142.070 ;
        RECT 18.935 142.025 19.225 142.070 ;
        RECT 18.935 141.885 24.430 142.025 ;
        RECT 18.935 141.840 19.225 141.885 ;
        RECT 13.160 141.455 13.480 141.715 ;
        RECT 13.655 141.655 13.945 141.700 ;
        RECT 18.050 141.655 18.190 141.840 ;
        RECT 24.290 141.715 24.430 141.885 ;
        RECT 32.360 141.825 32.680 142.085 ;
        RECT 32.840 142.025 33.160 142.085 ;
        RECT 59.720 142.025 60.040 142.085 ;
        RECT 61.730 142.025 61.870 142.255 ;
        RECT 63.095 142.210 63.385 142.255 ;
        RECT 63.650 142.255 66.280 142.395 ;
        RECT 32.840 141.885 41.710 142.025 ;
        RECT 32.840 141.825 33.160 141.885 ;
        RECT 13.655 141.515 18.190 141.655 ;
        RECT 13.655 141.470 13.945 141.515 ;
        RECT 14.120 141.285 14.440 141.345 ;
        RECT 15.575 141.285 15.865 141.330 ;
        RECT 14.120 141.145 15.865 141.285 ;
        RECT 18.050 141.285 18.190 141.515 ;
        RECT 21.320 141.455 21.640 141.715 ;
        RECT 24.200 141.455 24.520 141.715 ;
        RECT 24.680 141.655 25.000 141.715 ;
        RECT 41.570 141.700 41.710 141.885 ;
        RECT 59.720 141.885 61.870 142.025 ;
        RECT 59.720 141.825 60.040 141.885 ;
        RECT 26.615 141.655 26.905 141.700 ;
        RECT 29.495 141.655 29.785 141.700 ;
        RECT 33.335 141.655 33.625 141.700 ;
        RECT 24.680 141.515 33.625 141.655 ;
        RECT 24.680 141.455 25.000 141.515 ;
        RECT 26.615 141.470 26.905 141.515 ;
        RECT 29.495 141.470 29.785 141.515 ;
        RECT 33.335 141.470 33.625 141.515 ;
        RECT 34.295 141.655 34.585 141.700 ;
        RECT 34.295 141.515 40.510 141.655 ;
        RECT 34.295 141.470 34.585 141.515 ;
        RECT 37.160 141.285 37.480 141.345 ;
        RECT 38.615 141.285 38.905 141.330 ;
        RECT 18.050 141.145 33.070 141.285 ;
        RECT 14.120 141.085 14.440 141.145 ;
        RECT 15.575 141.100 15.865 141.145 ;
        RECT 32.930 140.975 33.070 141.145 ;
        RECT 37.160 141.145 38.905 141.285 ;
        RECT 37.160 141.085 37.480 141.145 ;
        RECT 38.615 141.100 38.905 141.145 ;
        RECT 32.840 140.715 33.160 140.975 ;
        RECT 40.370 140.915 40.510 141.515 ;
        RECT 41.495 141.470 41.785 141.700 ;
        RECT 44.360 141.455 44.680 141.715 ;
        RECT 60.695 141.655 60.985 141.700 ;
        RECT 63.650 141.655 63.790 142.255 ;
        RECT 65.960 142.195 66.280 142.255 ;
        RECT 64.520 142.025 64.840 142.085 ;
        RECT 66.455 142.025 66.745 142.070 ;
        RECT 64.520 141.885 66.745 142.025 ;
        RECT 64.520 141.825 64.840 141.885 ;
        RECT 66.455 141.840 66.745 141.885 ;
        RECT 60.695 141.515 63.790 141.655 ;
        RECT 60.695 141.470 60.985 141.515 ;
        RECT 46.775 141.285 47.065 141.330 ;
        RECT 47.720 141.285 48.040 141.345 ;
        RECT 46.775 141.145 48.040 141.285 ;
        RECT 46.775 141.100 47.065 141.145 ;
        RECT 47.720 141.085 48.040 141.145 ;
        RECT 48.680 141.285 49.000 141.345 ;
        RECT 50.615 141.285 50.905 141.330 ;
        RECT 48.680 141.145 50.905 141.285 ;
        RECT 48.680 141.085 49.000 141.145 ;
        RECT 50.615 141.100 50.905 141.145 ;
        RECT 54.440 141.285 54.760 141.345 ;
        RECT 55.895 141.285 56.185 141.330 ;
        RECT 54.440 141.145 56.185 141.285 ;
        RECT 54.440 141.085 54.760 141.145 ;
        RECT 55.895 141.100 56.185 141.145 ;
        RECT 61.640 141.285 61.960 141.345 ;
        RECT 63.575 141.285 63.865 141.330 ;
        RECT 61.640 141.145 63.865 141.285 ;
        RECT 61.640 141.085 61.960 141.145 ;
        RECT 63.575 141.100 63.865 141.145 ;
        RECT 52.520 140.915 52.840 140.975 ;
        RECT 40.370 140.775 52.840 140.915 ;
        RECT 52.520 140.715 52.840 140.775 ;
        RECT 10.200 140.045 69.720 140.535 ;
        RECT 13.175 139.805 13.465 139.850 ;
        RECT 20.840 139.805 21.160 139.865 ;
        RECT 13.175 139.665 21.160 139.805 ;
        RECT 13.175 139.620 13.465 139.665 ;
        RECT 20.840 139.605 21.160 139.665 ;
        RECT 25.640 139.805 25.960 139.865 ;
        RECT 27.095 139.805 27.385 139.850 ;
        RECT 25.640 139.665 27.385 139.805 ;
        RECT 25.640 139.605 25.960 139.665 ;
        RECT 27.095 139.620 27.385 139.665 ;
        RECT 43.415 139.805 43.705 139.850 ;
        RECT 43.880 139.805 44.200 139.865 ;
        RECT 43.415 139.665 44.200 139.805 ;
        RECT 43.415 139.620 43.705 139.665 ;
        RECT 43.880 139.605 44.200 139.665 ;
        RECT 46.775 139.805 47.065 139.850 ;
        RECT 47.240 139.805 47.560 139.865 ;
        RECT 46.775 139.665 47.560 139.805 ;
        RECT 46.775 139.620 47.065 139.665 ;
        RECT 47.240 139.605 47.560 139.665 ;
        RECT 59.720 139.605 60.040 139.865 ;
        RECT 32.360 139.435 32.680 139.495 ;
        RECT 31.490 139.295 45.550 139.435 ;
        RECT 15.095 139.065 15.385 139.110 ;
        RECT 17.975 139.065 18.265 139.110 ;
        RECT 21.815 139.065 22.105 139.110 ;
        RECT 24.680 139.065 25.000 139.125 ;
        RECT 15.095 138.925 25.000 139.065 ;
        RECT 15.095 138.880 15.385 138.925 ;
        RECT 17.975 138.880 18.265 138.925 ;
        RECT 21.815 138.880 22.105 138.925 ;
        RECT 24.680 138.865 25.000 138.925 ;
        RECT 20.855 138.695 21.145 138.740 ;
        RECT 22.280 138.695 22.600 138.755 ;
        RECT 20.855 138.555 22.600 138.695 ;
        RECT 20.855 138.510 21.145 138.555 ;
        RECT 22.280 138.495 22.600 138.555 ;
        RECT 25.640 138.495 25.960 138.755 ;
        RECT 22.775 138.140 23.065 138.370 ;
        RECT 24.200 138.325 24.520 138.385 ;
        RECT 25.730 138.325 25.870 138.495 ;
        RECT 24.200 138.185 25.870 138.325 ;
        RECT 22.850 137.955 22.990 138.140 ;
        RECT 24.200 138.125 24.520 138.185 ;
        RECT 26.600 138.125 26.920 138.385 ;
        RECT 31.490 138.325 31.630 139.295 ;
        RECT 32.360 139.235 32.680 139.295 ;
        RECT 32.840 139.065 33.160 139.125 ;
        RECT 45.410 139.110 45.550 139.295 ;
        RECT 50.630 139.110 50.890 139.155 ;
        RECT 34.295 139.065 34.585 139.110 ;
        RECT 38.135 139.065 38.425 139.110 ;
        RECT 41.015 139.065 41.305 139.110 ;
        RECT 32.840 138.925 41.305 139.065 ;
        RECT 32.840 138.865 33.160 138.925 ;
        RECT 34.295 138.880 34.585 138.925 ;
        RECT 38.135 138.880 38.425 138.925 ;
        RECT 41.015 138.880 41.305 138.925 ;
        RECT 45.335 138.880 45.625 139.110 ;
        RECT 50.615 139.065 50.905 139.110 ;
        RECT 54.455 139.065 54.745 139.110 ;
        RECT 57.335 139.065 57.625 139.110 ;
        RECT 50.615 138.925 57.625 139.065 ;
        RECT 50.615 138.880 50.905 138.925 ;
        RECT 54.455 138.880 54.745 138.925 ;
        RECT 57.335 138.880 57.625 138.925 ;
        RECT 31.880 138.740 32.200 138.755 ;
        RECT 31.880 138.695 32.265 138.740 ;
        RECT 35.255 138.695 35.545 138.740 ;
        RECT 31.880 138.555 35.545 138.695 ;
        RECT 45.410 138.695 45.550 138.880 ;
        RECT 50.630 138.835 50.890 138.880 ;
        RECT 51.575 138.695 51.865 138.740 ;
        RECT 45.410 138.555 53.710 138.695 ;
        RECT 31.880 138.510 32.265 138.555 ;
        RECT 35.255 138.510 35.545 138.555 ;
        RECT 51.575 138.510 51.865 138.555 ;
        RECT 31.880 138.495 32.200 138.510 ;
        RECT 32.375 138.325 32.665 138.370 ;
        RECT 31.490 138.185 32.665 138.325 ;
        RECT 32.375 138.140 32.665 138.185 ;
        RECT 33.320 138.125 33.640 138.385 ;
        RECT 43.400 138.325 43.720 138.385 ;
        RECT 44.855 138.325 45.145 138.370 ;
        RECT 43.400 138.185 45.145 138.325 ;
        RECT 43.400 138.125 43.720 138.185 ;
        RECT 44.855 138.140 45.145 138.185 ;
        RECT 48.215 138.140 48.505 138.370 ;
        RECT 49.160 138.325 49.480 138.385 ;
        RECT 49.655 138.325 49.945 138.370 ;
        RECT 49.160 138.185 49.945 138.325 ;
        RECT 47.720 137.955 48.040 138.015 ;
        RECT 22.850 137.815 48.040 137.955 ;
        RECT 48.290 137.955 48.430 138.140 ;
        RECT 49.160 138.125 49.480 138.185 ;
        RECT 49.655 138.140 49.945 138.185 ;
        RECT 48.290 137.815 51.790 137.955 ;
        RECT 47.720 137.755 48.040 137.815 ;
        RECT 51.650 137.645 51.790 137.815 ;
        RECT 53.570 137.645 53.710 138.555 ;
        RECT 64.055 138.325 64.345 138.370 ;
        RECT 66.440 138.325 66.760 138.385 ;
        RECT 64.055 138.185 66.760 138.325 ;
        RECT 64.055 138.140 64.345 138.185 ;
        RECT 66.440 138.125 66.760 138.185 ;
        RECT 66.935 138.325 67.225 138.370 ;
        RECT 68.360 138.325 68.680 138.385 ;
        RECT 66.935 138.185 68.680 138.325 ;
        RECT 66.935 138.140 67.225 138.185 ;
        RECT 68.360 138.125 68.680 138.185 ;
        RECT 51.560 137.385 51.880 137.645 ;
        RECT 53.480 137.385 53.800 137.645 ;
        RECT 62.615 137.585 62.905 137.630 ;
        RECT 63.560 137.585 63.880 137.645 ;
        RECT 62.615 137.445 63.880 137.585 ;
        RECT 62.615 137.400 62.905 137.445 ;
        RECT 63.560 137.385 63.880 137.445 ;
        RECT 65.495 137.585 65.785 137.630 ;
        RECT 66.440 137.585 66.760 137.645 ;
        RECT 65.495 137.445 66.760 137.585 ;
        RECT 65.495 137.400 65.785 137.445 ;
        RECT 66.440 137.385 66.760 137.445 ;
        RECT 10.200 136.715 69.720 137.205 ;
        RECT 13.160 136.475 13.480 136.535 ;
        RECT 13.655 136.475 13.945 136.520 ;
        RECT 13.160 136.335 13.945 136.475 ;
        RECT 13.160 136.275 13.480 136.335 ;
        RECT 13.655 136.290 13.945 136.335 ;
        RECT 14.615 136.475 14.905 136.520 ;
        RECT 26.600 136.475 26.920 136.535 ;
        RECT 14.615 136.335 26.920 136.475 ;
        RECT 14.615 136.290 14.905 136.335 ;
        RECT 26.600 136.275 26.920 136.335 ;
        RECT 35.240 136.275 35.560 136.535 ;
        RECT 44.855 136.475 45.145 136.520 ;
        RECT 51.080 136.475 51.400 136.535 ;
        RECT 44.855 136.335 51.400 136.475 ;
        RECT 44.855 136.290 45.145 136.335 ;
        RECT 51.080 136.275 51.400 136.335 ;
        RECT 56.855 136.475 57.145 136.520 ;
        RECT 57.800 136.475 58.120 136.535 ;
        RECT 62.615 136.475 62.905 136.520 ;
        RECT 56.855 136.335 58.120 136.475 ;
        RECT 56.855 136.290 57.145 136.335 ;
        RECT 57.800 136.275 58.120 136.335 ;
        RECT 58.370 136.335 62.905 136.475 ;
        RECT 46.760 136.105 47.080 136.165 ;
        RECT 24.770 135.965 47.080 136.105 ;
        RECT 24.770 135.780 24.910 135.965 ;
        RECT 46.760 135.905 47.080 135.965 ;
        RECT 47.720 136.105 48.040 136.165 ;
        RECT 54.440 136.105 54.760 136.165 ;
        RECT 58.370 136.105 58.510 136.335 ;
        RECT 62.615 136.290 62.905 136.335 ;
        RECT 64.520 136.275 64.840 136.535 ;
        RECT 65.960 136.275 66.280 136.535 ;
        RECT 47.720 135.965 54.760 136.105 ;
        RECT 47.720 135.905 48.040 135.965 ;
        RECT 54.440 135.905 54.760 135.965 ;
        RECT 57.890 135.965 58.510 136.105 ;
        RECT 59.735 136.105 60.025 136.150 ;
        RECT 66.050 136.105 66.190 136.275 ;
        RECT 59.735 135.965 66.190 136.105 ;
        RECT 57.890 135.795 58.030 135.965 ;
        RECT 59.735 135.920 60.025 135.965 ;
        RECT 24.695 135.550 24.985 135.780 ;
        RECT 31.880 135.735 32.200 135.795 ;
        RECT 25.250 135.595 32.200 135.735 ;
        RECT 8.360 135.365 8.680 135.425 ;
        RECT 12.215 135.365 12.505 135.410 ;
        RECT 8.360 135.225 12.505 135.365 ;
        RECT 8.360 135.165 8.680 135.225 ;
        RECT 12.215 135.180 12.505 135.225 ;
        RECT 22.280 135.365 22.600 135.425 ;
        RECT 22.775 135.365 23.065 135.410 ;
        RECT 25.250 135.365 25.390 135.595 ;
        RECT 26.600 135.365 26.920 135.425 ;
        RECT 27.170 135.410 27.310 135.595 ;
        RECT 31.880 135.535 32.200 135.595 ;
        RECT 53.480 135.735 53.800 135.795 ;
        RECT 53.480 135.595 56.110 135.735 ;
        RECT 53.480 135.535 53.800 135.595 ;
        RECT 22.280 135.225 25.390 135.365 ;
        RECT 25.730 135.225 26.920 135.365 ;
        RECT 22.280 135.165 22.600 135.225 ;
        RECT 22.775 135.180 23.065 135.225 ;
        RECT 17.015 134.995 17.305 135.040 ;
        RECT 19.895 134.995 20.185 135.040 ;
        RECT 23.735 134.995 24.025 135.040 ;
        RECT 17.015 134.855 24.025 134.995 ;
        RECT 17.015 134.810 17.305 134.855 ;
        RECT 19.895 134.810 20.185 134.855 ;
        RECT 23.735 134.810 24.025 134.855 ;
        RECT 25.175 134.995 25.465 135.040 ;
        RECT 25.730 134.995 25.870 135.225 ;
        RECT 26.600 135.165 26.920 135.225 ;
        RECT 27.095 135.180 27.385 135.410 ;
        RECT 53.015 135.365 53.305 135.410 ;
        RECT 53.570 135.365 53.710 135.535 ;
        RECT 53.015 135.225 53.710 135.365 ;
        RECT 54.935 135.365 55.225 135.410 ;
        RECT 55.400 135.365 55.720 135.425 ;
        RECT 54.935 135.225 55.720 135.365 ;
        RECT 55.970 135.365 56.110 135.595 ;
        RECT 57.800 135.535 58.120 135.795 ;
        RECT 58.280 135.535 58.600 135.795 ;
        RECT 61.175 135.735 61.465 135.780 ;
        RECT 61.640 135.735 61.960 135.795 ;
        RECT 61.175 135.595 61.960 135.735 ;
        RECT 61.175 135.550 61.465 135.595 ;
        RECT 61.640 135.535 61.960 135.595 ;
        RECT 63.575 135.550 63.865 135.780 ;
        RECT 63.650 135.365 63.790 135.550 ;
        RECT 65.480 135.535 65.800 135.795 ;
        RECT 55.970 135.225 63.790 135.365 ;
        RECT 53.015 135.180 53.305 135.225 ;
        RECT 54.935 135.180 55.225 135.225 ;
        RECT 55.400 135.165 55.720 135.225 ;
        RECT 25.175 134.855 25.870 134.995 ;
        RECT 26.135 134.995 26.425 135.040 ;
        RECT 29.975 134.995 30.265 135.040 ;
        RECT 32.855 134.995 33.145 135.040 ;
        RECT 26.135 134.855 33.145 134.995 ;
        RECT 25.175 134.810 25.465 134.855 ;
        RECT 26.135 134.810 26.425 134.855 ;
        RECT 29.975 134.810 30.265 134.855 ;
        RECT 32.855 134.810 33.145 134.855 ;
        RECT 47.255 134.995 47.545 135.040 ;
        RECT 48.200 134.995 48.520 135.055 ;
        RECT 50.135 134.995 50.425 135.040 ;
        RECT 53.975 134.995 54.265 135.040 ;
        RECT 47.255 134.855 54.265 134.995 ;
        RECT 47.255 134.810 47.545 134.855 ;
        RECT 23.810 134.625 23.950 134.810 ;
        RECT 24.680 134.625 25.000 134.685 ;
        RECT 26.210 134.625 26.350 134.810 ;
        RECT 48.200 134.795 48.520 134.855 ;
        RECT 50.135 134.810 50.425 134.855 ;
        RECT 53.975 134.810 54.265 134.855 ;
        RECT 23.810 134.485 26.350 134.625 ;
        RECT 48.290 134.625 48.430 134.795 ;
        RECT 50.600 134.625 50.920 134.685 ;
        RECT 48.290 134.485 50.920 134.625 ;
        RECT 24.680 134.425 25.000 134.485 ;
        RECT 50.600 134.425 50.920 134.485 ;
        RECT 66.920 134.055 67.240 134.315 ;
        RECT 10.200 133.385 69.720 133.875 ;
        RECT 13.175 133.145 13.465 133.190 ;
        RECT 13.640 133.145 13.960 133.205 ;
        RECT 13.175 133.005 13.960 133.145 ;
        RECT 13.175 132.960 13.465 133.005 ;
        RECT 13.640 132.945 13.960 133.005 ;
        RECT 39.095 133.145 39.385 133.190 ;
        RECT 50.120 133.145 50.440 133.205 ;
        RECT 39.095 133.005 50.440 133.145 ;
        RECT 39.095 132.960 39.385 133.005 ;
        RECT 50.120 132.945 50.440 133.005 ;
        RECT 53.960 133.145 54.280 133.205 ;
        RECT 55.415 133.145 55.705 133.190 ;
        RECT 53.960 133.005 55.705 133.145 ;
        RECT 53.960 132.945 54.280 133.005 ;
        RECT 55.415 132.960 55.705 133.005 ;
        RECT 48.200 132.775 48.520 132.835 ;
        RECT 41.090 132.635 48.520 132.775 ;
        RECT 15.095 132.405 15.385 132.450 ;
        RECT 17.975 132.405 18.265 132.450 ;
        RECT 21.815 132.405 22.105 132.450 ;
        RECT 25.640 132.405 25.960 132.465 ;
        RECT 41.090 132.450 41.230 132.635 ;
        RECT 48.200 132.575 48.520 132.635 ;
        RECT 57.830 132.450 58.090 132.495 ;
        RECT 41.015 132.405 41.305 132.450 ;
        RECT 43.895 132.405 44.185 132.450 ;
        RECT 47.735 132.405 48.025 132.450 ;
        RECT 15.095 132.265 48.025 132.405 ;
        RECT 15.095 132.220 15.385 132.265 ;
        RECT 17.975 132.220 18.265 132.265 ;
        RECT 21.815 132.220 22.105 132.265 ;
        RECT 25.640 132.205 25.960 132.265 ;
        RECT 41.015 132.220 41.305 132.265 ;
        RECT 43.895 132.220 44.185 132.265 ;
        RECT 47.735 132.220 48.025 132.265 ;
        RECT 57.815 132.405 58.105 132.450 ;
        RECT 61.655 132.405 61.945 132.450 ;
        RECT 64.535 132.405 64.825 132.450 ;
        RECT 57.815 132.265 64.825 132.405 ;
        RECT 57.815 132.220 58.105 132.265 ;
        RECT 61.655 132.220 61.945 132.265 ;
        RECT 64.535 132.220 64.825 132.265 ;
        RECT 57.830 132.175 58.090 132.220 ;
        RECT 20.855 132.035 21.145 132.080 ;
        RECT 22.280 132.035 22.600 132.095 ;
        RECT 20.855 131.895 22.600 132.035 ;
        RECT 20.855 131.850 21.145 131.895 ;
        RECT 22.280 131.835 22.600 131.895 ;
        RECT 40.520 132.035 40.840 132.095 ;
        RECT 43.400 132.035 43.720 132.095 ;
        RECT 46.775 132.035 47.065 132.080 ;
        RECT 40.520 131.895 47.065 132.035 ;
        RECT 40.520 131.835 40.840 131.895 ;
        RECT 43.400 131.835 43.720 131.895 ;
        RECT 46.775 131.850 47.065 131.895 ;
        RECT 58.760 131.835 59.080 132.095 ;
        RECT 22.775 131.665 23.065 131.710 ;
        RECT 37.160 131.665 37.480 131.725 ;
        RECT 22.775 131.525 37.480 131.665 ;
        RECT 22.775 131.480 23.065 131.525 ;
        RECT 37.160 131.465 37.480 131.525 ;
        RECT 48.695 131.665 48.985 131.710 ;
        RECT 49.160 131.665 49.480 131.725 ;
        RECT 48.695 131.525 49.480 131.665 ;
        RECT 48.695 131.480 48.985 131.525 ;
        RECT 49.160 131.465 49.480 131.525 ;
        RECT 55.895 131.480 56.185 131.710 ;
        RECT 55.970 131.295 56.110 131.480 ;
        RECT 56.840 131.465 57.160 131.725 ;
        RECT 66.935 131.295 67.225 131.340 ;
        RECT 55.970 131.155 67.225 131.295 ;
        RECT 66.935 131.110 67.225 131.155 ;
        RECT 10.200 130.055 69.720 130.545 ;
        RECT 51.560 129.615 51.880 129.875 ;
        RECT 56.840 129.075 57.160 129.135 ;
        RECT 61.655 129.075 61.945 129.120 ;
        RECT 56.840 128.935 61.945 129.075 ;
        RECT 56.840 128.875 57.160 128.935 ;
        RECT 61.655 128.890 61.945 128.935 ;
        RECT 65.495 128.890 65.785 129.120 ;
        RECT 17.480 128.505 17.800 128.765 ;
        RECT 18.440 128.705 18.760 128.765 ;
        RECT 26.135 128.705 26.425 128.750 ;
        RECT 18.440 128.565 26.425 128.705 ;
        RECT 18.440 128.505 18.760 128.565 ;
        RECT 26.135 128.520 26.425 128.565 ;
        RECT 59.240 128.705 59.560 128.765 ;
        RECT 59.735 128.705 60.025 128.750 ;
        RECT 65.570 128.705 65.710 128.890 ;
        RECT 59.240 128.565 65.710 128.705 ;
        RECT 59.240 128.505 59.560 128.565 ;
        RECT 59.735 128.520 60.025 128.565 ;
        RECT 13.160 128.335 13.480 128.395 ;
        RECT 16.535 128.335 16.825 128.380 ;
        RECT 13.160 128.195 16.825 128.335 ;
        RECT 13.160 128.135 13.480 128.195 ;
        RECT 16.535 128.150 16.825 128.195 ;
        RECT 24.215 128.335 24.505 128.380 ;
        RECT 27.560 128.335 27.880 128.395 ;
        RECT 24.215 128.195 27.880 128.335 ;
        RECT 24.215 128.150 24.505 128.195 ;
        RECT 27.560 128.135 27.880 128.195 ;
        RECT 53.975 128.335 54.265 128.380 ;
        RECT 56.855 128.335 57.145 128.380 ;
        RECT 60.695 128.335 60.985 128.380 ;
        RECT 53.975 128.195 60.985 128.335 ;
        RECT 53.975 128.150 54.265 128.195 ;
        RECT 56.855 128.150 57.145 128.195 ;
        RECT 60.695 128.150 60.985 128.195 ;
        RECT 54.050 127.965 54.190 128.150 ;
        RECT 66.920 128.135 67.240 128.395 ;
        RECT 57.800 127.965 58.120 128.025 ;
        RECT 54.050 127.825 58.120 127.965 ;
        RECT 17.960 127.595 18.280 127.655 ;
        RECT 18.455 127.595 18.745 127.640 ;
        RECT 17.960 127.455 18.745 127.595 ;
        RECT 17.960 127.395 18.280 127.455 ;
        RECT 18.455 127.410 18.745 127.455 ;
        RECT 46.760 127.595 47.080 127.655 ;
        RECT 54.050 127.595 54.190 127.825 ;
        RECT 57.800 127.765 58.120 127.825 ;
        RECT 46.760 127.455 54.190 127.595 ;
        RECT 46.760 127.395 47.080 127.455 ;
        RECT 111.750 127.400 112.250 153.320 ;
        RECT 116.800 150.215 117.310 150.815 ;
        RECT 119.260 150.215 119.770 150.815 ;
        RECT 113.800 149.765 114.260 149.815 ;
        RECT 116.260 149.765 116.720 149.815 ;
        RECT 112.800 132.850 113.180 149.765 ;
        RECT 113.780 148.875 114.280 149.765 ;
        RECT 114.510 148.670 114.680 149.765 ;
        RECT 113.380 147.170 113.750 148.670 ;
        RECT 114.310 147.170 114.680 148.670 ;
        RECT 113.380 146.530 113.550 147.170 ;
        RECT 113.800 146.735 114.260 146.965 ;
        RECT 114.510 146.530 114.680 147.170 ;
        RECT 113.380 145.030 113.750 146.530 ;
        RECT 114.310 145.030 114.680 146.530 ;
        RECT 113.380 144.390 113.550 145.030 ;
        RECT 113.800 144.595 114.260 144.825 ;
        RECT 114.510 144.390 114.680 145.030 ;
        RECT 113.380 142.890 113.750 144.390 ;
        RECT 114.310 142.890 114.680 144.390 ;
        RECT 113.380 142.250 113.550 142.890 ;
        RECT 113.800 142.455 114.260 142.685 ;
        RECT 114.510 142.250 114.680 142.890 ;
        RECT 113.380 140.750 113.750 142.250 ;
        RECT 114.310 140.750 114.680 142.250 ;
        RECT 113.380 139.740 113.550 140.750 ;
        RECT 113.800 140.315 114.260 140.545 ;
        RECT 114.510 139.740 114.680 140.750 ;
        RECT 113.380 139.570 114.680 139.740 ;
        RECT 113.380 138.605 113.550 139.570 ;
        RECT 113.800 138.765 114.260 138.995 ;
        RECT 114.510 138.605 114.680 139.570 ;
        RECT 113.380 138.105 113.750 138.605 ;
        RECT 114.310 138.105 114.680 138.605 ;
        RECT 113.380 137.555 113.550 138.105 ;
        RECT 113.800 137.715 114.260 137.945 ;
        RECT 114.510 137.555 114.680 138.105 ;
        RECT 113.380 137.055 113.750 137.555 ;
        RECT 114.310 137.055 114.680 137.555 ;
        RECT 113.380 136.505 113.550 137.055 ;
        RECT 113.800 136.665 114.260 136.895 ;
        RECT 114.510 136.505 114.680 137.055 ;
        RECT 113.380 136.005 113.750 136.505 ;
        RECT 114.310 136.005 114.680 136.505 ;
        RECT 113.380 135.455 113.550 136.005 ;
        RECT 113.800 135.615 114.260 135.845 ;
        RECT 114.510 135.455 114.680 136.005 ;
        RECT 113.380 134.955 113.750 135.455 ;
        RECT 114.310 134.955 114.680 135.455 ;
        RECT 113.380 127.450 113.550 134.955 ;
        RECT 113.780 133.905 114.280 134.795 ;
        RECT 114.510 133.905 114.680 134.955 ;
        RECT 113.800 133.855 114.260 133.905 ;
        RECT 114.880 131.850 115.640 149.765 ;
        RECT 115.840 148.715 116.010 149.765 ;
        RECT 116.240 148.875 116.740 149.765 ;
        RECT 116.970 148.715 117.140 150.215 ;
        RECT 115.840 148.215 116.210 148.715 ;
        RECT 116.770 148.215 117.140 148.715 ;
        RECT 115.840 147.665 116.010 148.215 ;
        RECT 116.260 147.825 116.720 148.055 ;
        RECT 116.970 147.665 117.140 148.215 ;
        RECT 115.840 147.165 116.210 147.665 ;
        RECT 116.770 147.165 117.140 147.665 ;
        RECT 115.840 146.615 116.010 147.165 ;
        RECT 116.260 146.775 116.720 147.005 ;
        RECT 116.970 146.615 117.140 147.165 ;
        RECT 115.840 146.115 116.210 146.615 ;
        RECT 116.770 146.115 117.140 146.615 ;
        RECT 115.840 145.565 116.010 146.115 ;
        RECT 116.260 145.725 116.720 145.955 ;
        RECT 116.970 145.565 117.140 146.115 ;
        RECT 115.840 145.065 116.210 145.565 ;
        RECT 116.770 145.065 117.140 145.565 ;
        RECT 115.840 142.920 116.010 145.065 ;
        RECT 116.260 144.675 116.720 144.905 ;
        RECT 116.260 143.125 116.720 143.355 ;
        RECT 116.970 142.920 117.140 145.065 ;
        RECT 115.840 141.420 116.210 142.920 ;
        RECT 116.770 141.420 117.140 142.920 ;
        RECT 115.840 140.780 116.010 141.420 ;
        RECT 116.260 140.985 116.720 141.215 ;
        RECT 116.970 140.780 117.140 141.420 ;
        RECT 115.840 139.280 116.210 140.780 ;
        RECT 116.770 139.280 117.140 140.780 ;
        RECT 115.840 138.640 116.010 139.280 ;
        RECT 116.260 138.845 116.720 139.075 ;
        RECT 116.970 138.640 117.140 139.280 ;
        RECT 115.840 137.140 116.210 138.640 ;
        RECT 116.770 137.140 117.140 138.640 ;
        RECT 115.840 136.500 116.010 137.140 ;
        RECT 116.260 136.705 116.720 136.935 ;
        RECT 116.970 136.500 117.140 137.140 ;
        RECT 115.840 135.000 116.210 136.500 ;
        RECT 116.770 135.000 117.140 136.500 ;
        RECT 117.340 149.760 117.720 149.765 ;
        RECT 118.720 149.760 119.180 149.815 ;
        RECT 115.840 127.450 116.010 135.000 ;
        RECT 116.240 133.905 116.740 134.795 ;
        RECT 116.260 127.850 116.720 133.905 ;
        RECT 117.340 132.850 118.100 149.760 ;
        RECT 118.700 148.870 119.200 149.760 ;
        RECT 119.430 148.665 119.600 150.215 ;
        RECT 118.300 147.165 118.670 148.665 ;
        RECT 119.230 147.165 119.600 148.665 ;
        RECT 118.300 146.525 118.470 147.165 ;
        RECT 118.720 146.730 119.180 146.960 ;
        RECT 119.430 146.525 119.600 147.165 ;
        RECT 118.300 145.025 118.670 146.525 ;
        RECT 119.230 145.025 119.600 146.525 ;
        RECT 118.300 144.385 118.470 145.025 ;
        RECT 118.720 144.590 119.180 144.820 ;
        RECT 119.430 144.385 119.600 145.025 ;
        RECT 118.300 142.885 118.670 144.385 ;
        RECT 119.230 142.885 119.600 144.385 ;
        RECT 118.300 142.245 118.470 142.885 ;
        RECT 118.720 142.450 119.180 142.680 ;
        RECT 119.430 142.245 119.600 142.885 ;
        RECT 118.300 140.745 118.670 142.245 ;
        RECT 119.230 140.745 119.600 142.245 ;
        RECT 118.300 139.735 118.470 140.745 ;
        RECT 118.720 140.310 119.180 140.540 ;
        RECT 119.430 139.735 119.600 140.745 ;
        RECT 118.300 139.565 119.600 139.735 ;
        RECT 118.300 138.600 118.470 139.565 ;
        RECT 118.720 138.760 119.180 138.990 ;
        RECT 119.430 138.600 119.600 139.565 ;
        RECT 118.300 138.100 118.670 138.600 ;
        RECT 119.230 138.100 119.600 138.600 ;
        RECT 118.300 137.550 118.470 138.100 ;
        RECT 118.720 137.710 119.180 137.940 ;
        RECT 119.430 137.550 119.600 138.100 ;
        RECT 118.300 137.050 118.670 137.550 ;
        RECT 119.230 137.050 119.600 137.550 ;
        RECT 118.300 136.500 118.470 137.050 ;
        RECT 118.720 136.660 119.180 136.890 ;
        RECT 119.430 136.500 119.600 137.050 ;
        RECT 118.300 136.000 118.670 136.500 ;
        RECT 119.230 136.000 119.600 136.500 ;
        RECT 118.300 135.450 118.470 136.000 ;
        RECT 118.720 135.610 119.180 135.840 ;
        RECT 119.430 135.450 119.600 136.000 ;
        RECT 118.300 134.950 118.670 135.450 ;
        RECT 119.230 134.950 119.600 135.450 ;
        RECT 118.300 133.900 118.470 134.950 ;
        RECT 118.700 133.900 119.200 134.790 ;
        RECT 119.430 133.900 119.600 134.950 ;
        RECT 119.800 144.010 120.180 149.760 ;
        RECT 119.800 142.915 120.560 144.010 ;
        RECT 121.180 143.120 121.640 143.350 ;
        RECT 123.110 143.120 123.570 143.350 ;
        RECT 123.820 142.915 125.320 150.815 ;
        RECT 119.800 141.415 121.130 142.915 ;
        RECT 121.690 141.415 123.060 142.915 ;
        RECT 123.620 141.855 125.320 142.915 ;
        RECT 123.620 141.685 125.370 141.855 ;
        RECT 123.620 141.415 125.315 141.685 ;
        RECT 119.800 140.775 120.930 141.415 ;
        RECT 121.180 140.980 121.640 141.210 ;
        RECT 121.890 140.775 122.860 141.415 ;
        RECT 123.110 140.980 123.570 141.210 ;
        RECT 123.820 140.775 125.315 141.415 ;
        RECT 119.800 139.275 121.130 140.775 ;
        RECT 121.690 139.275 123.060 140.775 ;
        RECT 123.620 139.275 125.315 140.775 ;
        RECT 128.960 139.600 129.450 151.850 ;
        RECT 130.495 151.330 130.855 151.750 ;
        RECT 130.415 149.030 130.775 149.450 ;
        RECT 130.490 148.110 130.850 148.530 ;
        RECT 131.455 148.120 131.755 149.850 ;
        RECT 130.540 144.785 130.900 145.205 ;
        RECT 119.800 138.635 120.930 139.275 ;
        RECT 121.180 138.840 121.640 139.070 ;
        RECT 121.890 138.635 122.860 139.275 ;
        RECT 123.110 138.840 123.570 139.070 ;
        RECT 123.820 138.635 125.315 139.275 ;
        RECT 125.570 138.760 126.030 138.990 ;
        RECT 127.500 138.760 127.960 138.990 ;
        RECT 119.800 137.135 121.130 138.635 ;
        RECT 121.690 137.135 123.060 138.635 ;
        RECT 123.620 138.600 125.315 138.635 ;
        RECT 128.580 138.600 129.450 139.600 ;
        RECT 123.620 138.100 125.520 138.600 ;
        RECT 126.080 138.100 127.450 138.600 ;
        RECT 128.010 138.100 129.450 138.600 ;
        RECT 123.620 137.550 125.315 138.100 ;
        RECT 125.570 137.710 126.030 137.940 ;
        RECT 126.280 137.550 127.250 138.100 ;
        RECT 127.500 137.710 127.960 137.940 ;
        RECT 128.210 137.550 129.450 138.100 ;
        RECT 123.620 137.135 125.520 137.550 ;
        RECT 119.800 136.495 120.930 137.135 ;
        RECT 121.180 136.700 121.640 136.930 ;
        RECT 121.890 136.495 122.860 137.135 ;
        RECT 123.820 137.050 125.520 137.135 ;
        RECT 126.080 137.050 127.450 137.550 ;
        RECT 128.010 137.050 129.450 137.550 ;
        RECT 123.110 136.700 123.570 136.930 ;
        RECT 123.820 136.500 125.315 137.050 ;
        RECT 125.570 136.660 126.030 136.890 ;
        RECT 126.280 136.500 127.250 137.050 ;
        RECT 127.500 136.660 127.960 136.890 ;
        RECT 128.210 136.500 129.450 137.050 ;
        RECT 123.820 136.495 125.520 136.500 ;
        RECT 119.800 134.995 121.130 136.495 ;
        RECT 121.690 134.995 123.060 136.495 ;
        RECT 123.620 136.000 125.520 136.495 ;
        RECT 126.080 136.000 127.450 136.500 ;
        RECT 128.010 136.000 129.450 136.500 ;
        RECT 123.620 135.450 125.315 136.000 ;
        RECT 125.570 135.610 126.030 135.840 ;
        RECT 126.280 135.450 127.250 136.000 ;
        RECT 127.500 135.610 127.960 135.840 ;
        RECT 128.210 135.450 129.450 136.000 ;
        RECT 123.620 134.995 125.520 135.450 ;
        RECT 118.720 133.855 119.180 133.900 ;
        RECT 10.200 126.725 69.720 127.215 ;
        RECT 111.700 126.900 112.300 127.400 ;
        RECT 14.135 126.485 14.425 126.530 ;
        RECT 17.480 126.485 17.800 126.545 ;
        RECT 14.135 126.345 17.800 126.485 ;
        RECT 14.135 126.300 14.425 126.345 ;
        RECT 17.480 126.285 17.800 126.345 ;
        RECT 27.560 126.285 27.880 126.545 ;
        RECT 40.520 126.285 40.840 126.545 ;
        RECT 66.935 126.485 67.225 126.530 ;
        RECT 69.320 126.485 69.640 126.545 ;
        RECT 66.935 126.345 69.640 126.485 ;
        RECT 66.935 126.300 67.225 126.345 ;
        RECT 69.320 126.285 69.640 126.345 ;
        RECT 59.240 126.115 59.560 126.175 ;
        RECT 46.370 125.975 59.560 126.115 ;
        RECT 25.160 125.745 25.480 125.805 ;
        RECT 12.770 125.605 25.480 125.745 ;
        RECT 12.770 125.050 12.910 125.605 ;
        RECT 25.160 125.545 25.480 125.605 ;
        RECT 31.415 125.745 31.705 125.790 ;
        RECT 35.255 125.745 35.545 125.790 ;
        RECT 38.135 125.745 38.425 125.790 ;
        RECT 40.520 125.745 40.840 125.805 ;
        RECT 31.415 125.605 40.840 125.745 ;
        RECT 31.415 125.560 31.705 125.605 ;
        RECT 35.255 125.560 35.545 125.605 ;
        RECT 38.135 125.560 38.425 125.605 ;
        RECT 40.520 125.545 40.840 125.605 ;
        RECT 16.055 125.190 16.345 125.420 ;
        RECT 17.960 125.375 18.280 125.435 ;
        RECT 20.855 125.375 21.145 125.420 ;
        RECT 17.960 125.235 21.145 125.375 ;
        RECT 12.695 124.820 12.985 125.050 ;
        RECT 13.655 125.005 13.945 125.050 ;
        RECT 13.250 124.865 13.945 125.005 ;
        RECT 13.250 124.265 13.390 124.865 ;
        RECT 13.655 124.820 13.945 124.865 ;
        RECT 13.655 124.635 13.945 124.680 ;
        RECT 16.130 124.635 16.270 125.190 ;
        RECT 17.960 125.175 18.280 125.235 ;
        RECT 20.855 125.190 21.145 125.235 ;
        RECT 21.320 125.375 21.640 125.435 ;
        RECT 26.615 125.375 26.905 125.420 ;
        RECT 21.320 125.235 26.905 125.375 ;
        RECT 21.320 125.175 21.640 125.235 ;
        RECT 26.615 125.190 26.905 125.235 ;
        RECT 28.520 125.175 28.840 125.435 ;
        RECT 31.880 125.375 32.200 125.435 ;
        RECT 32.375 125.375 32.665 125.420 ;
        RECT 46.370 125.375 46.510 125.975 ;
        RECT 59.240 125.915 59.560 125.975 ;
        RECT 46.760 125.745 47.080 125.805 ;
        RECT 50.615 125.745 50.905 125.790 ;
        RECT 54.455 125.745 54.745 125.790 ;
        RECT 57.335 125.745 57.625 125.790 ;
        RECT 46.760 125.605 57.625 125.745 ;
        RECT 46.760 125.545 47.080 125.605 ;
        RECT 50.615 125.560 50.905 125.605 ;
        RECT 54.455 125.560 54.745 125.605 ;
        RECT 57.335 125.560 57.625 125.605 ;
        RECT 31.880 125.235 32.665 125.375 ;
        RECT 31.880 125.175 32.200 125.235 ;
        RECT 32.375 125.190 32.665 125.235 ;
        RECT 33.410 125.235 46.510 125.375 ;
        RECT 33.410 125.065 33.550 125.235 ;
        RECT 47.720 125.175 48.040 125.435 ;
        RECT 51.575 125.375 51.865 125.420 ;
        RECT 48.290 125.235 51.865 125.375 ;
        RECT 17.495 125.005 17.785 125.050 ;
        RECT 25.655 125.005 25.945 125.050 ;
        RECT 17.495 124.865 25.945 125.005 ;
        RECT 17.495 124.820 17.785 124.865 ;
        RECT 25.655 124.820 25.945 124.865 ;
        RECT 30.455 125.005 30.745 125.050 ;
        RECT 33.320 125.005 33.640 125.065 ;
        RECT 30.455 124.865 33.640 125.005 ;
        RECT 30.455 124.820 30.745 124.865 ;
        RECT 33.320 124.805 33.640 124.865 ;
        RECT 46.760 124.805 47.080 125.065 ;
        RECT 13.655 124.495 23.950 124.635 ;
        RECT 13.655 124.450 13.945 124.495 ;
        RECT 23.810 124.325 23.950 124.495 ;
        RECT 19.895 124.265 20.185 124.310 ;
        RECT 22.280 124.265 22.600 124.325 ;
        RECT 13.250 124.125 22.600 124.265 ;
        RECT 19.895 124.080 20.185 124.125 ;
        RECT 22.280 124.065 22.600 124.125 ;
        RECT 23.720 124.065 24.040 124.325 ;
        RECT 41.960 124.265 42.280 124.325 ;
        RECT 48.290 124.265 48.430 125.235 ;
        RECT 51.575 125.190 51.865 125.235 ;
        RECT 49.640 125.005 49.960 125.065 ;
        RECT 58.760 125.005 59.080 125.065 ;
        RECT 62.615 125.005 62.905 125.050 ;
        RECT 49.640 124.865 62.905 125.005 ;
        RECT 49.640 124.805 49.960 124.865 ;
        RECT 58.760 124.805 59.080 124.865 ;
        RECT 62.615 124.820 62.905 124.865 ;
        RECT 63.080 125.005 63.400 125.065 ;
        RECT 65.495 125.005 65.785 125.050 ;
        RECT 63.080 124.865 65.785 125.005 ;
        RECT 63.080 124.805 63.400 124.865 ;
        RECT 65.495 124.820 65.785 124.865 ;
        RECT 41.960 124.125 48.430 124.265 ;
        RECT 41.960 124.065 42.280 124.125 ;
        RECT 64.040 124.065 64.360 124.325 ;
        RECT 10.200 123.395 69.720 123.885 ;
        RECT 23.255 123.155 23.545 123.200 ;
        RECT 24.680 123.155 25.000 123.215 ;
        RECT 23.255 123.015 25.000 123.155 ;
        RECT 23.255 122.970 23.545 123.015 ;
        RECT 24.680 122.955 25.000 123.015 ;
        RECT 28.520 122.955 28.840 123.215 ;
        RECT 33.320 122.955 33.640 123.215 ;
        RECT 14.135 122.045 14.425 122.090 ;
        RECT 18.440 122.045 18.760 122.105 ;
        RECT 14.135 121.905 18.760 122.045 ;
        RECT 14.135 121.860 14.425 121.905 ;
        RECT 18.440 121.845 18.760 121.905 ;
        RECT 23.240 121.845 23.560 122.105 ;
        RECT 23.720 121.845 24.040 122.105 ;
        RECT 28.610 122.045 28.750 122.955 ;
        RECT 24.770 121.905 28.750 122.045 ;
        RECT 33.410 122.045 33.550 122.955 ;
        RECT 40.040 122.785 40.360 122.845 ;
        RECT 50.120 122.785 50.440 122.845 ;
        RECT 40.040 122.645 50.440 122.785 ;
        RECT 40.040 122.585 40.360 122.645 ;
        RECT 50.120 122.585 50.440 122.645 ;
        RECT 54.920 122.415 55.240 122.475 ;
        RECT 34.850 122.275 37.870 122.415 ;
        RECT 33.815 122.045 34.105 122.090 ;
        RECT 33.410 121.905 34.105 122.045 ;
        RECT 16.055 121.675 16.345 121.720 ;
        RECT 16.520 121.675 16.840 121.735 ;
        RECT 24.770 121.720 24.910 121.905 ;
        RECT 33.815 121.860 34.105 121.905 ;
        RECT 34.850 121.720 34.990 122.275 ;
        RECT 36.695 122.045 36.985 122.090 ;
        RECT 35.330 121.905 36.985 122.045 ;
        RECT 16.055 121.535 16.840 121.675 ;
        RECT 16.055 121.490 16.345 121.535 ;
        RECT 16.520 121.475 16.840 121.535 ;
        RECT 24.695 121.490 24.985 121.720 ;
        RECT 28.055 121.675 28.345 121.720 ;
        RECT 30.935 121.675 31.225 121.720 ;
        RECT 34.775 121.675 35.065 121.720 ;
        RECT 28.055 121.535 35.065 121.675 ;
        RECT 28.055 121.490 28.345 121.535 ;
        RECT 30.935 121.490 31.225 121.535 ;
        RECT 34.775 121.490 35.065 121.535 ;
        RECT 32.840 121.305 33.160 121.365 ;
        RECT 35.330 121.305 35.470 121.905 ;
        RECT 36.695 121.860 36.985 121.905 ;
        RECT 37.730 121.720 37.870 122.275 ;
        RECT 45.890 122.275 55.240 122.415 ;
        RECT 45.890 122.090 46.030 122.275 ;
        RECT 54.920 122.215 55.240 122.275 ;
        RECT 59.240 122.415 59.560 122.475 ;
        RECT 65.495 122.415 65.785 122.460 ;
        RECT 59.240 122.275 65.785 122.415 ;
        RECT 59.240 122.215 59.560 122.275 ;
        RECT 65.495 122.230 65.785 122.275 ;
        RECT 45.815 121.860 46.105 122.090 ;
        RECT 48.215 122.045 48.505 122.090 ;
        RECT 49.640 122.045 49.960 122.105 ;
        RECT 48.215 121.905 49.960 122.045 ;
        RECT 48.215 121.860 48.505 121.905 ;
        RECT 49.640 121.845 49.960 121.905 ;
        RECT 35.735 121.490 36.025 121.720 ;
        RECT 37.655 121.675 37.945 121.720 ;
        RECT 40.520 121.675 40.840 121.735 ;
        RECT 46.295 121.675 46.585 121.720 ;
        RECT 37.655 121.535 40.840 121.675 ;
        RECT 37.655 121.490 37.945 121.535 ;
        RECT 32.840 121.165 35.470 121.305 ;
        RECT 35.810 121.305 35.950 121.490 ;
        RECT 40.520 121.475 40.840 121.535 ;
        RECT 44.450 121.535 46.585 121.675 ;
        RECT 35.810 121.165 41.230 121.305 ;
        RECT 32.840 121.105 33.160 121.165 ;
        RECT 41.090 120.995 41.230 121.165 ;
        RECT 21.320 120.935 21.640 120.995 ;
        RECT 21.815 120.935 22.105 120.980 ;
        RECT 21.320 120.795 22.105 120.935 ;
        RECT 21.320 120.735 21.640 120.795 ;
        RECT 21.815 120.750 22.105 120.795 ;
        RECT 25.655 120.935 25.945 120.980 ;
        RECT 40.040 120.935 40.360 120.995 ;
        RECT 25.655 120.795 40.360 120.935 ;
        RECT 25.655 120.750 25.945 120.795 ;
        RECT 40.040 120.735 40.360 120.795 ;
        RECT 41.000 120.935 41.320 120.995 ;
        RECT 44.450 120.980 44.590 121.535 ;
        RECT 46.295 121.490 46.585 121.535 ;
        RECT 47.255 121.675 47.545 121.720 ;
        RECT 51.095 121.675 51.385 121.720 ;
        RECT 52.040 121.675 52.360 121.735 ;
        RECT 53.975 121.675 54.265 121.720 ;
        RECT 47.255 121.535 54.265 121.675 ;
        RECT 47.255 121.490 47.545 121.535 ;
        RECT 51.095 121.490 51.385 121.535 ;
        RECT 52.040 121.475 52.360 121.535 ;
        RECT 53.975 121.490 54.265 121.535 ;
        RECT 50.120 121.305 50.440 121.365 ;
        RECT 55.880 121.305 56.200 121.365 ;
        RECT 50.120 121.165 56.200 121.305 ;
        RECT 50.120 121.105 50.440 121.165 ;
        RECT 55.880 121.105 56.200 121.165 ;
        RECT 44.375 120.935 44.665 120.980 ;
        RECT 41.000 120.795 44.665 120.935 ;
        RECT 41.000 120.735 41.320 120.795 ;
        RECT 44.375 120.750 44.665 120.795 ;
        RECT 55.400 120.935 55.720 120.995 ;
        RECT 56.375 120.935 56.665 120.980 ;
        RECT 57.320 120.935 57.640 120.995 ;
        RECT 55.400 120.795 57.640 120.935 ;
        RECT 55.400 120.735 55.720 120.795 ;
        RECT 56.375 120.750 56.665 120.795 ;
        RECT 57.320 120.735 57.640 120.795 ;
        RECT 66.920 120.735 67.240 120.995 ;
        RECT 10.200 120.065 69.720 120.555 ;
        RECT 23.240 119.825 23.560 119.885 ;
        RECT 23.735 119.825 24.025 119.870 ;
        RECT 23.240 119.685 24.025 119.825 ;
        RECT 23.240 119.625 23.560 119.685 ;
        RECT 23.735 119.640 24.025 119.685 ;
        RECT 48.215 119.825 48.505 119.870 ;
        RECT 49.640 119.825 49.960 119.885 ;
        RECT 48.215 119.685 49.960 119.825 ;
        RECT 48.215 119.640 48.505 119.685 ;
        RECT 49.640 119.625 49.960 119.685 ;
        RECT 62.120 119.825 62.440 119.885 ;
        RECT 66.455 119.825 66.745 119.870 ;
        RECT 62.120 119.685 66.745 119.825 ;
        RECT 62.120 119.625 62.440 119.685 ;
        RECT 66.455 119.640 66.745 119.685 ;
        RECT 40.520 119.455 40.840 119.515 ;
        RECT 36.770 119.315 47.470 119.455 ;
        RECT 18.440 119.130 18.760 119.145 ;
        RECT 36.770 119.130 36.910 119.315 ;
        RECT 40.520 119.255 40.840 119.315 ;
        RECT 12.630 118.900 19.330 119.130 ;
        RECT 29.975 119.085 30.265 119.130 ;
        RECT 32.855 119.085 33.145 119.130 ;
        RECT 36.695 119.085 36.985 119.130 ;
        RECT 29.975 118.945 36.985 119.085 ;
        RECT 29.975 118.900 30.265 118.945 ;
        RECT 32.855 118.900 33.145 118.945 ;
        RECT 36.695 118.900 36.985 118.945 ;
        RECT 39.095 119.085 39.385 119.130 ;
        RECT 42.935 119.085 43.225 119.130 ;
        RECT 45.815 119.085 46.105 119.130 ;
        RECT 46.760 119.085 47.080 119.145 ;
        RECT 39.095 118.945 47.080 119.085 ;
        RECT 39.095 118.900 39.385 118.945 ;
        RECT 42.935 118.900 43.225 118.945 ;
        RECT 45.815 118.900 46.105 118.945 ;
        RECT 18.440 118.885 18.760 118.900 ;
        RECT 46.760 118.885 47.080 118.945 ;
        RECT 47.330 118.775 47.470 119.315 ;
        RECT 47.720 119.085 48.040 119.145 ;
        RECT 52.040 119.085 52.360 119.145 ;
        RECT 57.830 119.130 58.090 119.175 ;
        RECT 57.815 119.085 58.105 119.130 ;
        RECT 61.655 119.085 61.945 119.130 ;
        RECT 64.535 119.085 64.825 119.130 ;
        RECT 47.720 118.945 64.825 119.085 ;
        RECT 47.720 118.885 48.040 118.945 ;
        RECT 52.040 118.885 52.360 118.945 ;
        RECT 57.815 118.900 58.105 118.945 ;
        RECT 61.655 118.900 61.945 118.945 ;
        RECT 64.535 118.900 64.825 118.945 ;
        RECT 57.830 118.855 58.090 118.900 ;
        RECT 21.335 118.715 21.625 118.760 ;
        RECT 21.800 118.715 22.120 118.775 ;
        RECT 21.335 118.575 22.120 118.715 ;
        RECT 21.335 118.530 21.625 118.575 ;
        RECT 21.800 118.515 22.120 118.575 ;
        RECT 22.280 118.715 22.600 118.775 ;
        RECT 24.695 118.715 24.985 118.760 ;
        RECT 22.280 118.575 24.985 118.715 ;
        RECT 22.280 118.515 22.600 118.575 ;
        RECT 24.695 118.530 24.985 118.575 ;
        RECT 27.080 118.715 27.400 118.775 ;
        RECT 35.735 118.715 36.025 118.760 ;
        RECT 40.055 118.715 40.345 118.760 ;
        RECT 41.960 118.715 42.280 118.775 ;
        RECT 27.080 118.575 42.280 118.715 ;
        RECT 27.080 118.515 27.400 118.575 ;
        RECT 35.735 118.530 36.025 118.575 ;
        RECT 40.055 118.530 40.345 118.575 ;
        RECT 41.960 118.515 42.280 118.575 ;
        RECT 47.240 118.715 47.560 118.775 ;
        RECT 51.095 118.715 51.385 118.760 ;
        RECT 47.240 118.575 51.385 118.715 ;
        RECT 47.240 118.515 47.560 118.575 ;
        RECT 51.095 118.530 51.385 118.575 ;
        RECT 53.495 118.530 53.785 118.760 ;
        RECT 58.775 118.715 59.065 118.760 ;
        RECT 59.240 118.715 59.560 118.775 ;
        RECT 58.775 118.575 59.560 118.715 ;
        RECT 58.775 118.530 59.065 118.575 ;
        RECT 13.080 118.160 19.780 118.390 ;
        RECT 25.160 118.345 25.480 118.405 ;
        RECT 25.655 118.345 25.945 118.390 ;
        RECT 33.320 118.345 33.640 118.405 ;
        RECT 25.160 118.205 33.640 118.345 ;
        RECT 25.160 118.145 25.480 118.205 ;
        RECT 25.655 118.160 25.945 118.205 ;
        RECT 33.320 118.145 33.640 118.205 ;
        RECT 37.640 118.145 37.960 118.405 ;
        RECT 38.135 118.345 38.425 118.390 ;
        RECT 48.200 118.345 48.520 118.405 ;
        RECT 53.570 118.345 53.710 118.530 ;
        RECT 59.240 118.515 59.560 118.575 ;
        RECT 56.840 118.345 57.160 118.405 ;
        RECT 38.135 118.205 41.710 118.345 ;
        RECT 38.135 118.160 38.425 118.205 ;
        RECT 27.575 117.975 27.865 118.020 ;
        RECT 38.210 117.975 38.350 118.160 ;
        RECT 27.575 117.835 38.350 117.975 ;
        RECT 27.575 117.790 27.865 117.835 ;
        RECT 41.570 117.665 41.710 118.205 ;
        RECT 48.200 118.205 53.710 118.345 ;
        RECT 55.010 118.205 57.160 118.345 ;
        RECT 48.200 118.145 48.520 118.205 ;
        RECT 55.010 117.665 55.150 118.205 ;
        RECT 56.840 118.145 57.160 118.205 ;
        RECT 41.480 117.405 41.800 117.665 ;
        RECT 54.920 117.405 55.240 117.665 ;
        RECT 10.200 116.735 69.720 117.225 ;
        RECT 17.015 116.495 17.305 116.540 ;
        RECT 27.560 116.495 27.880 116.555 ;
        RECT 17.015 116.355 27.880 116.495 ;
        RECT 17.015 116.310 17.305 116.355 ;
        RECT 27.560 116.295 27.880 116.355 ;
        RECT 58.760 116.295 59.080 116.555 ;
        RECT 61.160 116.295 61.480 116.555 ;
        RECT 66.920 116.295 67.240 116.555 ;
        RECT 17.960 116.125 18.280 116.185 ;
        RECT 41.480 116.125 41.800 116.185 ;
        RECT 58.850 116.125 58.990 116.295 ;
        RECT 16.130 115.985 37.390 116.125 ;
        RECT 16.130 115.430 16.270 115.985 ;
        RECT 17.960 115.925 18.280 115.985 ;
        RECT 22.200 115.570 28.900 115.800 ;
        RECT 31.400 115.755 31.720 115.815 ;
        RECT 32.375 115.755 32.665 115.800 ;
        RECT 29.090 115.615 32.665 115.755 ;
        RECT 15.575 115.200 15.865 115.430 ;
        RECT 16.055 115.200 16.345 115.430 ;
        RECT 18.935 115.200 19.225 115.430 ;
        RECT 13.640 114.275 13.960 114.335 ;
        RECT 14.135 114.275 14.425 114.320 ;
        RECT 13.640 114.135 14.425 114.275 ;
        RECT 15.650 114.275 15.790 115.200 ;
        RECT 19.010 114.645 19.150 115.200 ;
        RECT 19.400 115.185 19.720 115.445 ;
        RECT 20.375 115.385 20.665 115.430 ;
        RECT 29.090 115.385 29.230 115.615 ;
        RECT 31.400 115.555 31.720 115.615 ;
        RECT 32.375 115.570 32.665 115.615 ;
        RECT 33.320 115.755 33.640 115.815 ;
        RECT 37.250 115.800 37.390 115.985 ;
        RECT 41.480 115.985 58.990 116.125 ;
        RECT 41.480 115.925 41.800 115.985 ;
        RECT 35.735 115.755 36.025 115.800 ;
        RECT 33.320 115.615 36.025 115.755 ;
        RECT 33.320 115.555 33.640 115.615 ;
        RECT 35.735 115.570 36.025 115.615 ;
        RECT 37.175 115.570 37.465 115.800 ;
        RECT 37.655 115.570 37.945 115.800 ;
        RECT 38.135 115.570 38.425 115.800 ;
        RECT 20.375 115.245 29.230 115.385 ;
        RECT 20.375 115.200 20.665 115.245 ;
        RECT 30.440 115.185 30.760 115.445 ;
        RECT 30.920 115.185 31.240 115.445 ;
        RECT 31.895 115.385 32.185 115.430 ;
        RECT 33.410 115.385 33.550 115.555 ;
        RECT 31.895 115.245 33.550 115.385 ;
        RECT 35.810 115.385 35.950 115.570 ;
        RECT 37.730 115.385 37.870 115.570 ;
        RECT 35.810 115.245 37.870 115.385 ;
        RECT 31.895 115.200 32.185 115.245 ;
        RECT 21.800 115.060 22.120 115.075 ;
        RECT 21.750 114.830 28.450 115.060 ;
        RECT 38.210 115.015 38.350 115.570 ;
        RECT 41.570 115.430 41.710 115.925 ;
        RECT 51.095 115.755 51.385 115.800 ;
        RECT 54.920 115.755 55.240 115.815 ;
        RECT 51.095 115.615 55.240 115.755 ;
        RECT 51.095 115.570 51.385 115.615 ;
        RECT 54.920 115.555 55.240 115.615 ;
        RECT 59.240 115.755 59.560 115.815 ;
        RECT 65.495 115.755 65.785 115.800 ;
        RECT 59.240 115.615 65.785 115.755 ;
        RECT 59.240 115.555 59.560 115.615 ;
        RECT 65.495 115.570 65.785 115.615 ;
        RECT 41.495 115.200 41.785 115.430 ;
        RECT 53.015 115.385 53.305 115.430 ;
        RECT 53.480 115.385 53.800 115.445 ;
        RECT 53.015 115.245 53.800 115.385 ;
        RECT 53.015 115.200 53.305 115.245 ;
        RECT 53.480 115.185 53.800 115.245 ;
        RECT 28.610 114.875 38.350 115.015 ;
        RECT 39.575 115.015 39.865 115.060 ;
        RECT 40.040 115.015 40.360 115.075 ;
        RECT 47.270 115.060 47.530 115.105 ;
        RECT 39.575 114.875 40.360 115.015 ;
        RECT 21.800 114.815 22.120 114.830 ;
        RECT 21.320 114.645 21.640 114.705 ;
        RECT 28.610 114.645 28.750 114.875 ;
        RECT 39.575 114.830 39.865 114.875 ;
        RECT 40.040 114.815 40.360 114.875 ;
        RECT 40.535 115.015 40.825 115.060 ;
        RECT 44.375 115.015 44.665 115.060 ;
        RECT 47.255 115.015 47.545 115.060 ;
        RECT 40.535 114.875 47.545 115.015 ;
        RECT 40.535 114.830 40.825 114.875 ;
        RECT 44.375 114.830 44.665 114.875 ;
        RECT 47.255 114.830 47.545 114.875 ;
        RECT 52.055 115.015 52.345 115.060 ;
        RECT 55.895 115.015 56.185 115.060 ;
        RECT 57.800 115.015 58.120 115.075 ;
        RECT 58.775 115.015 59.065 115.060 ;
        RECT 52.055 114.875 59.065 115.015 ;
        RECT 52.055 114.830 52.345 114.875 ;
        RECT 55.895 114.830 56.185 114.875 ;
        RECT 47.270 114.785 47.530 114.830 ;
        RECT 57.800 114.815 58.120 114.875 ;
        RECT 58.775 114.830 59.065 114.875 ;
        RECT 19.010 114.505 28.750 114.645 ;
        RECT 32.360 114.645 32.680 114.705 ;
        RECT 36.695 114.645 36.985 114.690 ;
        RECT 32.360 114.505 36.985 114.645 ;
        RECT 21.320 114.445 21.640 114.505 ;
        RECT 32.360 114.445 32.680 114.505 ;
        RECT 36.695 114.460 36.985 114.505 ;
        RECT 26.120 114.275 26.440 114.335 ;
        RECT 15.650 114.135 26.440 114.275 ;
        RECT 13.640 114.075 13.960 114.135 ;
        RECT 14.135 114.090 14.425 114.135 ;
        RECT 26.120 114.075 26.440 114.135 ;
        RECT 31.415 114.275 31.705 114.320 ;
        RECT 33.320 114.275 33.640 114.335 ;
        RECT 31.415 114.135 33.640 114.275 ;
        RECT 31.415 114.090 31.705 114.135 ;
        RECT 33.320 114.075 33.640 114.135 ;
        RECT 49.640 114.075 49.960 114.335 ;
        RECT 10.200 113.405 69.720 113.895 ;
        RECT 13.640 112.965 13.960 113.225 ;
        RECT 31.400 112.965 31.720 113.225 ;
        RECT 58.280 113.165 58.600 113.225 ;
        RECT 66.455 113.165 66.745 113.210 ;
        RECT 58.280 113.025 66.745 113.165 ;
        RECT 58.280 112.965 58.600 113.025 ;
        RECT 66.455 112.980 66.745 113.025 ;
        RECT 13.730 112.425 13.870 112.965 ;
        RECT 37.640 112.795 37.960 112.855 ;
        RECT 37.640 112.655 54.190 112.795 ;
        RECT 37.640 112.595 37.960 112.655 ;
        RECT 38.150 112.470 38.410 112.515 ;
        RECT 35.255 112.425 35.545 112.470 ;
        RECT 38.135 112.425 38.425 112.470 ;
        RECT 41.975 112.425 42.265 112.470 ;
        RECT 13.730 112.285 14.830 112.425 ;
        RECT 12.215 111.870 12.505 112.100 ;
        RECT 12.290 111.685 12.430 111.870 ;
        RECT 13.160 111.855 13.480 112.115 ;
        RECT 14.690 112.100 14.830 112.285 ;
        RECT 35.255 112.285 42.265 112.425 ;
        RECT 35.255 112.240 35.545 112.285 ;
        RECT 38.135 112.240 38.425 112.285 ;
        RECT 41.975 112.240 42.265 112.285 ;
        RECT 38.150 112.195 38.410 112.240 ;
        RECT 13.655 111.870 13.945 112.100 ;
        RECT 14.615 111.870 14.905 112.100 ;
        RECT 15.095 112.055 15.385 112.100 ;
        RECT 16.520 112.055 16.840 112.115 ;
        RECT 15.095 111.915 16.840 112.055 ;
        RECT 15.095 111.870 15.385 111.915 ;
        RECT 13.730 111.685 13.870 111.870 ;
        RECT 16.520 111.855 16.840 111.915 ;
        RECT 18.440 112.055 18.760 112.115 ;
        RECT 23.735 112.055 24.025 112.100 ;
        RECT 18.440 111.915 24.025 112.055 ;
        RECT 18.440 111.855 18.760 111.915 ;
        RECT 23.735 111.870 24.025 111.915 ;
        RECT 41.015 112.055 41.305 112.100 ;
        RECT 43.400 112.055 43.720 112.115 ;
        RECT 53.480 112.055 53.800 112.115 ;
        RECT 41.015 111.915 53.800 112.055 ;
        RECT 54.050 112.055 54.190 112.655 ;
        RECT 57.830 112.470 58.090 112.515 ;
        RECT 57.815 112.425 58.105 112.470 ;
        RECT 61.655 112.425 61.945 112.470 ;
        RECT 64.535 112.425 64.825 112.470 ;
        RECT 57.815 112.285 64.825 112.425 ;
        RECT 57.815 112.240 58.105 112.285 ;
        RECT 61.655 112.240 61.945 112.285 ;
        RECT 64.535 112.240 64.825 112.285 ;
        RECT 57.830 112.195 58.090 112.240 ;
        RECT 58.775 112.055 59.065 112.100 ;
        RECT 59.240 112.055 59.560 112.115 ;
        RECT 54.050 111.915 59.560 112.055 ;
        RECT 41.015 111.870 41.305 111.915 ;
        RECT 43.400 111.855 43.720 111.915 ;
        RECT 53.480 111.855 53.800 111.915 ;
        RECT 58.775 111.870 59.065 111.915 ;
        RECT 59.240 111.855 59.560 111.915 ;
        RECT 12.290 111.545 13.870 111.685 ;
        RECT 13.730 111.315 13.870 111.545 ;
        RECT 17.000 111.485 17.320 111.745 ;
        RECT 25.640 111.485 25.960 111.745 ;
        RECT 42.920 111.485 43.240 111.745 ;
        RECT 56.840 111.485 57.160 111.745 ;
        RECT 30.920 111.315 31.240 111.375 ;
        RECT 13.730 111.175 31.240 111.315 ;
        RECT 30.920 111.115 31.240 111.175 ;
        RECT 12.680 110.745 13.000 111.005 ;
        RECT 14.120 110.745 14.440 111.005 ;
        RECT 22.760 110.745 23.080 111.005 ;
        RECT 26.600 110.945 26.920 111.005 ;
        RECT 32.855 110.945 33.145 110.990 ;
        RECT 57.800 110.945 58.120 111.005 ;
        RECT 26.600 110.805 58.120 110.945 ;
        RECT 26.600 110.745 26.920 110.805 ;
        RECT 32.855 110.760 33.145 110.805 ;
        RECT 57.800 110.745 58.120 110.805 ;
        RECT 10.200 110.075 69.720 110.565 ;
        RECT 12.680 109.635 13.000 109.895 ;
        RECT 14.120 109.635 14.440 109.895 ;
        RECT 16.040 109.835 16.360 109.895 ;
        RECT 16.535 109.835 16.825 109.880 ;
        RECT 16.040 109.695 16.825 109.835 ;
        RECT 16.040 109.635 16.360 109.695 ;
        RECT 16.535 109.650 16.825 109.695 ;
        RECT 17.000 109.835 17.320 109.895 ;
        RECT 20.855 109.835 21.145 109.880 ;
        RECT 17.000 109.695 21.145 109.835 ;
        RECT 17.000 109.635 17.320 109.695 ;
        RECT 20.855 109.650 21.145 109.695 ;
        RECT 22.760 109.635 23.080 109.895 ;
        RECT 25.640 109.835 25.960 109.895 ;
        RECT 31.895 109.835 32.185 109.880 ;
        RECT 25.640 109.695 32.185 109.835 ;
        RECT 25.640 109.635 25.960 109.695 ;
        RECT 31.895 109.650 32.185 109.695 ;
        RECT 66.935 109.835 67.225 109.880 ;
        RECT 68.840 109.835 69.160 109.895 ;
        RECT 66.935 109.695 69.160 109.835 ;
        RECT 66.935 109.650 67.225 109.695 ;
        RECT 68.840 109.635 69.160 109.695 ;
        RECT 12.770 108.725 12.910 109.635 ;
        RECT 14.210 109.095 14.350 109.635 ;
        RECT 14.210 108.955 18.910 109.095 ;
        RECT 15.095 108.725 15.385 108.770 ;
        RECT 12.770 108.585 15.385 108.725 ;
        RECT 18.770 108.725 18.910 108.955 ;
        RECT 21.815 108.725 22.105 108.770 ;
        RECT 18.770 108.585 22.105 108.725 ;
        RECT 22.850 108.725 22.990 109.635 ;
        RECT 28.520 109.265 28.840 109.525 ;
        RECT 29.495 109.465 29.785 109.510 ;
        RECT 31.400 109.465 31.720 109.525 ;
        RECT 29.495 109.325 31.720 109.465 ;
        RECT 29.495 109.280 29.785 109.325 ;
        RECT 31.400 109.265 31.720 109.325 ;
        RECT 53.480 109.465 53.800 109.525 ;
        RECT 54.935 109.465 55.225 109.510 ;
        RECT 53.480 109.325 65.710 109.465 ;
        RECT 53.480 109.265 53.800 109.325 ;
        RECT 54.935 109.280 55.225 109.325 ;
        RECT 24.695 108.725 24.985 108.770 ;
        RECT 22.850 108.585 24.985 108.725 ;
        RECT 15.095 108.540 15.385 108.585 ;
        RECT 21.815 108.540 22.105 108.585 ;
        RECT 24.695 108.540 24.985 108.585 ;
        RECT 27.560 108.525 27.880 108.785 ;
        RECT 28.610 108.770 28.750 109.265 ;
        RECT 38.120 108.895 38.440 109.155 ;
        RECT 56.360 109.095 56.680 109.155 ;
        RECT 65.570 109.140 65.710 109.325 ;
        RECT 59.735 109.095 60.025 109.140 ;
        RECT 56.360 108.955 60.025 109.095 ;
        RECT 56.360 108.895 56.680 108.955 ;
        RECT 59.735 108.910 60.025 108.955 ;
        RECT 65.495 108.910 65.785 109.140 ;
        RECT 28.535 108.725 28.825 108.770 ;
        RECT 29.480 108.725 29.800 108.785 ;
        RECT 28.535 108.585 29.800 108.725 ;
        RECT 28.535 108.540 28.825 108.585 ;
        RECT 29.480 108.525 29.800 108.585 ;
        RECT 33.320 108.525 33.640 108.785 ;
        RECT 37.175 108.725 37.465 108.770 ;
        RECT 40.040 108.725 40.360 108.785 ;
        RECT 37.175 108.585 40.360 108.725 ;
        RECT 37.175 108.540 37.465 108.585 ;
        RECT 40.040 108.525 40.360 108.585 ;
        RECT 41.960 108.725 42.280 108.785 ;
        RECT 46.775 108.725 47.065 108.770 ;
        RECT 41.960 108.585 47.065 108.725 ;
        RECT 41.960 108.525 42.280 108.585 ;
        RECT 46.775 108.540 47.065 108.585 ;
        RECT 19.400 108.355 19.720 108.415 ;
        RECT 23.720 108.355 24.040 108.415 ;
        RECT 19.400 108.215 24.040 108.355 ;
        RECT 19.400 108.155 19.720 108.215 ;
        RECT 23.720 108.155 24.040 108.215 ;
        RECT 43.880 108.355 44.200 108.415 ;
        RECT 44.855 108.355 45.145 108.400 ;
        RECT 43.880 108.215 45.145 108.355 ;
        RECT 43.880 108.155 44.200 108.215 ;
        RECT 44.855 108.170 45.145 108.215 ;
        RECT 45.815 108.355 46.105 108.400 ;
        RECT 49.655 108.355 49.945 108.400 ;
        RECT 51.560 108.355 51.880 108.415 ;
        RECT 52.535 108.355 52.825 108.400 ;
        RECT 45.815 108.215 52.825 108.355 ;
        RECT 45.815 108.170 46.105 108.215 ;
        RECT 49.655 108.170 49.945 108.215 ;
        RECT 51.560 108.155 51.880 108.215 ;
        RECT 52.535 108.170 52.825 108.215 ;
        RECT 61.175 108.355 61.465 108.400 ;
        RECT 65.960 108.355 66.280 108.415 ;
        RECT 61.175 108.215 66.280 108.355 ;
        RECT 61.175 108.170 61.465 108.215 ;
        RECT 65.960 108.155 66.280 108.215 ;
        RECT 10.200 106.745 69.720 107.235 ;
        RECT 37.640 106.505 37.960 106.565 ;
        RECT 33.890 106.365 37.960 106.505 ;
        RECT 26.120 106.135 26.440 106.195 ;
        RECT 33.890 106.180 34.030 106.365 ;
        RECT 37.640 106.305 37.960 106.365 ;
        RECT 27.095 106.135 27.385 106.180 ;
        RECT 26.120 105.995 27.385 106.135 ;
        RECT 26.120 105.935 26.440 105.995 ;
        RECT 27.095 105.950 27.385 105.995 ;
        RECT 33.815 105.950 34.105 106.180 ;
        RECT 51.560 106.135 51.880 106.195 ;
        RECT 47.810 105.995 51.880 106.135 ;
        RECT 16.520 105.810 16.840 105.825 ;
        RECT 12.630 105.580 19.330 105.810 ;
        RECT 35.735 105.765 36.025 105.810 ;
        RECT 38.120 105.765 38.440 105.825 ;
        RECT 38.615 105.765 38.905 105.810 ;
        RECT 42.455 105.765 42.745 105.810 ;
        RECT 26.210 105.625 32.590 105.765 ;
        RECT 16.520 105.565 16.840 105.580 ;
        RECT 21.335 105.395 21.625 105.440 ;
        RECT 21.800 105.395 22.120 105.455 ;
        RECT 26.210 105.440 26.350 105.625 ;
        RECT 32.450 105.455 32.590 105.625 ;
        RECT 35.735 105.625 42.745 105.765 ;
        RECT 35.735 105.580 36.025 105.625 ;
        RECT 38.120 105.565 38.440 105.625 ;
        RECT 38.615 105.580 38.905 105.625 ;
        RECT 42.455 105.580 42.745 105.625 ;
        RECT 43.400 105.565 43.720 105.825 ;
        RECT 47.810 105.810 47.950 105.995 ;
        RECT 51.560 105.935 51.880 105.995 ;
        RECT 43.970 105.625 47.470 105.765 ;
        RECT 21.335 105.255 22.120 105.395 ;
        RECT 21.335 105.210 21.625 105.255 ;
        RECT 21.800 105.195 22.120 105.255 ;
        RECT 26.135 105.210 26.425 105.440 ;
        RECT 26.600 105.395 26.920 105.455 ;
        RECT 28.535 105.395 28.825 105.440 ;
        RECT 31.895 105.395 32.185 105.440 ;
        RECT 26.600 105.255 28.825 105.395 ;
        RECT 26.600 105.195 26.920 105.255 ;
        RECT 28.535 105.210 28.825 105.255 ;
        RECT 29.090 105.255 32.185 105.395 ;
        RECT 13.080 104.840 19.780 105.070 ;
        RECT 23.720 104.825 24.040 105.085 ;
        RECT 24.200 105.025 24.520 105.085 ;
        RECT 29.090 105.025 29.230 105.255 ;
        RECT 31.895 105.210 32.185 105.255 ;
        RECT 32.360 105.195 32.680 105.455 ;
        RECT 41.495 105.395 41.785 105.440 ;
        RECT 43.970 105.395 44.110 105.625 ;
        RECT 47.330 105.455 47.470 105.625 ;
        RECT 47.735 105.580 48.025 105.810 ;
        RECT 50.615 105.765 50.905 105.810 ;
        RECT 51.650 105.765 51.790 105.935 ;
        RECT 54.455 105.765 54.745 105.810 ;
        RECT 57.335 105.765 57.625 105.810 ;
        RECT 50.615 105.625 57.625 105.765 ;
        RECT 50.615 105.580 50.905 105.625 ;
        RECT 54.455 105.580 54.745 105.625 ;
        RECT 57.335 105.580 57.625 105.625 ;
        RECT 66.920 105.565 67.240 105.825 ;
        RECT 41.495 105.255 44.110 105.395 ;
        RECT 41.495 105.210 41.785 105.255 ;
        RECT 46.775 105.210 47.065 105.440 ;
        RECT 47.240 105.395 47.560 105.455 ;
        RECT 51.575 105.395 51.865 105.440 ;
        RECT 47.240 105.255 51.865 105.395 ;
        RECT 24.200 104.885 29.230 105.025 ;
        RECT 29.480 105.025 29.800 105.085 ;
        RECT 30.455 105.025 30.745 105.070 ;
        RECT 29.480 104.885 30.745 105.025 ;
        RECT 24.200 104.825 24.520 104.885 ;
        RECT 29.480 104.825 29.800 104.885 ;
        RECT 30.455 104.840 30.745 104.885 ;
        RECT 40.040 105.025 40.360 105.085 ;
        RECT 46.850 105.025 46.990 105.210 ;
        RECT 47.240 105.195 47.560 105.255 ;
        RECT 51.575 105.210 51.865 105.255 ;
        RECT 49.655 105.025 49.945 105.070 ;
        RECT 56.360 105.025 56.680 105.085 ;
        RECT 40.040 104.885 47.470 105.025 ;
        RECT 40.040 104.825 40.360 104.885 ;
        RECT 26.120 104.655 26.440 104.715 ;
        RECT 29.570 104.655 29.710 104.825 ;
        RECT 47.330 104.715 47.470 104.885 ;
        RECT 49.655 104.885 56.680 105.025 ;
        RECT 49.655 104.840 49.945 104.885 ;
        RECT 56.360 104.825 56.680 104.885 ;
        RECT 62.600 104.825 62.920 105.085 ;
        RECT 65.495 104.840 65.785 105.070 ;
        RECT 26.120 104.515 29.710 104.655 ;
        RECT 26.120 104.455 26.440 104.515 ;
        RECT 47.240 104.455 47.560 104.715 ;
        RECT 64.040 104.455 64.360 104.715 ;
        RECT 27.560 104.085 27.880 104.345 ;
        RECT 28.520 104.285 28.840 104.345 ;
        RECT 30.935 104.285 31.225 104.330 ;
        RECT 28.520 104.145 31.225 104.285 ;
        RECT 28.520 104.085 28.840 104.145 ;
        RECT 30.935 104.100 31.225 104.145 ;
        RECT 43.880 104.285 44.200 104.345 ;
        RECT 58.760 104.285 59.080 104.345 ;
        RECT 59.735 104.285 60.025 104.330 ;
        RECT 65.570 104.285 65.710 104.840 ;
        RECT 43.880 104.145 65.710 104.285 ;
        RECT 43.880 104.085 44.200 104.145 ;
        RECT 58.760 104.085 59.080 104.145 ;
        RECT 59.735 104.100 60.025 104.145 ;
        RECT 10.200 103.415 69.720 103.905 ;
        RECT 22.775 102.990 23.065 103.220 ;
        RECT 22.850 102.805 22.990 102.990 ;
        RECT 24.200 102.975 24.520 103.235 ;
        RECT 26.120 102.975 26.440 103.235 ;
        RECT 28.520 103.175 28.840 103.235 ;
        RECT 26.690 103.035 28.840 103.175 ;
        RECT 26.210 102.805 26.350 102.975 ;
        RECT 22.850 102.665 26.350 102.805 ;
        RECT 23.255 102.435 23.545 102.480 ;
        RECT 26.120 102.435 26.440 102.495 ;
        RECT 26.690 102.480 26.830 103.035 ;
        RECT 28.520 102.975 28.840 103.035 ;
        RECT 52.520 103.175 52.840 103.235 ;
        RECT 53.495 103.175 53.785 103.220 ;
        RECT 52.520 103.035 53.785 103.175 ;
        RECT 52.520 102.975 52.840 103.035 ;
        RECT 53.495 102.990 53.785 103.035 ;
        RECT 23.255 102.295 26.440 102.435 ;
        RECT 23.255 102.250 23.545 102.295 ;
        RECT 26.120 102.235 26.440 102.295 ;
        RECT 26.615 102.250 26.905 102.480 ;
        RECT 42.920 102.435 43.240 102.495 ;
        RECT 43.415 102.435 43.705 102.480 ;
        RECT 42.920 102.295 43.705 102.435 ;
        RECT 42.920 102.235 43.240 102.295 ;
        RECT 43.415 102.250 43.705 102.295 ;
        RECT 55.880 102.435 56.200 102.495 ;
        RECT 59.735 102.435 60.025 102.480 ;
        RECT 55.880 102.295 60.025 102.435 ;
        RECT 55.880 102.235 56.200 102.295 ;
        RECT 59.735 102.250 60.025 102.295 ;
        RECT 65.495 102.250 65.785 102.480 ;
        RECT 13.655 102.065 13.945 102.110 ;
        RECT 16.520 102.065 16.840 102.125 ;
        RECT 24.695 102.065 24.985 102.110 ;
        RECT 13.655 101.925 24.985 102.065 ;
        RECT 13.655 101.880 13.945 101.925 ;
        RECT 16.520 101.865 16.840 101.925 ;
        RECT 24.695 101.880 24.985 101.925 ;
        RECT 43.880 102.065 44.200 102.125 ;
        RECT 45.335 102.065 45.625 102.110 ;
        RECT 43.880 101.925 45.625 102.065 ;
        RECT 43.880 101.865 44.200 101.925 ;
        RECT 45.335 101.880 45.625 101.925 ;
        RECT 47.240 102.065 47.560 102.125 ;
        RECT 64.055 102.065 64.345 102.110 ;
        RECT 47.240 101.925 64.345 102.065 ;
        RECT 47.240 101.865 47.560 101.925 ;
        RECT 64.055 101.880 64.345 101.925 ;
        RECT 15.575 101.695 15.865 101.740 ;
        RECT 44.375 101.695 44.665 101.740 ;
        RECT 48.215 101.695 48.505 101.740 ;
        RECT 51.095 101.695 51.385 101.740 ;
        RECT 51.560 101.695 51.880 101.755 ;
        RECT 65.570 101.695 65.710 102.250 ;
        RECT 15.575 101.555 16.750 101.695 ;
        RECT 15.575 101.510 15.865 101.555 ;
        RECT 16.610 101.385 16.750 101.555 ;
        RECT 44.375 101.555 51.880 101.695 ;
        RECT 44.375 101.510 44.665 101.555 ;
        RECT 48.215 101.510 48.505 101.555 ;
        RECT 51.095 101.510 51.385 101.555 ;
        RECT 51.560 101.495 51.880 101.555 ;
        RECT 52.130 101.555 65.710 101.695 ;
        RECT 16.520 101.125 16.840 101.385 ;
        RECT 47.240 101.325 47.560 101.385 ;
        RECT 52.130 101.325 52.270 101.555 ;
        RECT 66.920 101.495 67.240 101.755 ;
        RECT 63.095 101.325 63.385 101.370 ;
        RECT 47.240 101.185 52.270 101.325 ;
        RECT 58.370 101.185 63.385 101.325 ;
        RECT 47.240 101.125 47.560 101.185 ;
        RECT 58.370 101.015 58.510 101.185 ;
        RECT 63.095 101.140 63.385 101.185 ;
        RECT 21.320 100.755 21.640 101.015 ;
        RECT 32.360 100.755 32.680 101.015 ;
        RECT 58.280 100.755 58.600 101.015 ;
        RECT 61.160 100.755 61.480 101.015 ;
        RECT 10.200 100.085 69.720 100.575 ;
        RECT 111.750 100.400 112.250 126.900 ;
        RECT 113.210 126.850 113.720 127.450 ;
        RECT 115.670 126.850 116.180 127.450 ;
        RECT 112.800 117.900 113.300 126.450 ;
        RECT 113.800 124.200 114.300 125.450 ;
        RECT 112.750 117.400 113.350 117.900 ;
        RECT 112.800 100.850 113.300 117.400 ;
        RECT 113.750 108.400 114.350 108.900 ;
        RECT 113.800 101.850 114.300 108.400 ;
        RECT 15.575 99.845 15.865 99.890 ;
        RECT 16.520 99.845 16.840 99.905 ;
        RECT 15.575 99.705 16.840 99.845 ;
        RECT 15.575 99.660 15.865 99.705 ;
        RECT 16.520 99.645 16.840 99.705 ;
        RECT 26.120 99.845 26.440 99.905 ;
        RECT 111.700 99.900 112.300 100.400 ;
        RECT 27.575 99.845 27.865 99.890 ;
        RECT 26.120 99.705 27.865 99.845 ;
        RECT 26.120 99.645 26.440 99.705 ;
        RECT 27.575 99.660 27.865 99.705 ;
        RECT 27.560 99.105 27.880 99.165 ;
        RECT 17.090 98.965 27.880 99.105 ;
        RECT 17.090 98.780 17.230 98.965 ;
        RECT 27.560 98.905 27.880 98.965 ;
        RECT 34.775 99.105 35.065 99.150 ;
        RECT 37.655 99.105 37.945 99.150 ;
        RECT 38.120 99.105 38.440 99.165 ;
        RECT 41.495 99.105 41.785 99.150 ;
        RECT 34.775 98.965 41.785 99.105 ;
        RECT 34.775 98.920 35.065 98.965 ;
        RECT 37.655 98.920 37.945 98.965 ;
        RECT 38.120 98.905 38.440 98.965 ;
        RECT 41.495 98.920 41.785 98.965 ;
        RECT 56.840 98.905 57.160 99.165 ;
        RECT 57.815 99.105 58.105 99.150 ;
        RECT 58.280 99.105 58.600 99.165 ;
        RECT 61.655 99.105 61.945 99.150 ;
        RECT 64.535 99.105 64.825 99.150 ;
        RECT 57.815 98.965 64.825 99.105 ;
        RECT 57.815 98.920 58.105 98.965 ;
        RECT 58.280 98.905 58.600 98.965 ;
        RECT 61.655 98.920 61.945 98.965 ;
        RECT 64.535 98.920 64.825 98.965 ;
        RECT 66.935 99.105 67.225 99.150 ;
        RECT 67.400 99.105 67.720 99.165 ;
        RECT 66.935 98.965 67.720 99.105 ;
        RECT 66.935 98.920 67.225 98.965 ;
        RECT 67.400 98.905 67.720 98.965 ;
        RECT 17.015 98.550 17.305 98.780 ;
        RECT 19.415 98.550 19.705 98.780 ;
        RECT 21.320 98.735 21.640 98.795 ;
        RECT 26.615 98.735 26.905 98.780 ;
        RECT 21.320 98.595 26.905 98.735 ;
        RECT 19.490 97.995 19.630 98.550 ;
        RECT 21.320 98.535 21.640 98.595 ;
        RECT 26.615 98.550 26.905 98.595 ;
        RECT 28.040 98.735 28.360 98.795 ;
        RECT 28.535 98.735 28.825 98.780 ;
        RECT 28.040 98.595 28.825 98.735 ;
        RECT 28.040 98.535 28.360 98.595 ;
        RECT 28.535 98.550 28.825 98.595 ;
        RECT 20.855 98.365 21.145 98.410 ;
        RECT 25.655 98.365 25.945 98.410 ;
        RECT 20.855 98.225 25.945 98.365 ;
        RECT 20.855 98.180 21.145 98.225 ;
        RECT 25.655 98.180 25.945 98.225 ;
        RECT 30.935 98.365 31.225 98.410 ;
        RECT 38.210 98.365 38.350 98.905 ;
        RECT 40.535 98.550 40.825 98.780 ;
        RECT 41.000 98.735 41.320 98.795 ;
        RECT 42.455 98.735 42.745 98.780 ;
        RECT 41.000 98.595 42.745 98.735 ;
        RECT 30.935 98.225 38.350 98.365 ;
        RECT 30.935 98.180 31.225 98.225 ;
        RECT 19.490 97.855 21.070 97.995 ;
        RECT 20.930 97.685 21.070 97.855 ;
        RECT 21.335 97.810 21.625 98.040 ;
        RECT 22.775 97.995 23.065 98.040 ;
        RECT 26.600 97.995 26.920 98.055 ;
        RECT 22.775 97.855 26.920 97.995 ;
        RECT 22.775 97.810 23.065 97.855 ;
        RECT 20.840 97.425 21.160 97.685 ;
        RECT 21.410 97.625 21.550 97.810 ;
        RECT 26.600 97.795 26.920 97.855 ;
        RECT 37.640 97.995 37.960 98.055 ;
        RECT 40.610 97.995 40.750 98.550 ;
        RECT 41.000 98.535 41.320 98.595 ;
        RECT 42.455 98.550 42.745 98.595 ;
        RECT 58.760 98.535 59.080 98.795 ;
        RECT 50.615 98.365 50.905 98.410 ;
        RECT 51.560 98.365 51.880 98.425 ;
        RECT 50.615 98.225 51.880 98.365 ;
        RECT 50.615 98.180 50.905 98.225 ;
        RECT 51.560 98.165 51.880 98.225 ;
        RECT 54.440 98.165 54.760 98.425 ;
        RECT 37.640 97.855 40.750 97.995 ;
        RECT 43.970 97.855 65.710 97.995 ;
        RECT 37.640 97.795 37.960 97.855 ;
        RECT 25.160 97.625 25.480 97.685 ;
        RECT 21.410 97.485 25.480 97.625 ;
        RECT 25.160 97.425 25.480 97.485 ;
        RECT 32.375 97.625 32.665 97.670 ;
        RECT 33.320 97.625 33.640 97.685 ;
        RECT 43.970 97.625 44.110 97.855 ;
        RECT 65.570 97.685 65.710 97.855 ;
        RECT 111.750 97.750 112.250 99.900 ;
        RECT 113.210 99.850 113.720 100.450 ;
        RECT 115.670 99.850 116.180 100.450 ;
        RECT 32.375 97.485 44.110 97.625 ;
        RECT 32.375 97.440 32.665 97.485 ;
        RECT 33.320 97.425 33.640 97.485 ;
        RECT 52.040 97.425 52.360 97.685 ;
        RECT 55.880 97.425 56.200 97.685 ;
        RECT 65.480 97.425 65.800 97.685 ;
        RECT 10.200 96.755 69.720 97.245 ;
        RECT 109.400 96.850 112.250 97.750 ;
        RECT 20.840 96.515 21.160 96.575 ;
        RECT 28.040 96.515 28.360 96.575 ;
        RECT 20.840 96.375 28.360 96.515 ;
        RECT 20.840 96.315 21.160 96.375 ;
        RECT 28.040 96.315 28.360 96.375 ;
        RECT 30.920 96.515 31.240 96.575 ;
        RECT 32.840 96.515 33.160 96.575 ;
        RECT 30.920 96.375 33.160 96.515 ;
        RECT 30.920 96.315 31.240 96.375 ;
        RECT 32.840 96.315 33.160 96.375 ;
        RECT 40.040 96.315 40.360 96.575 ;
        RECT 46.280 96.515 46.600 96.575 ;
        RECT 49.655 96.515 49.945 96.560 ;
        RECT 46.280 96.375 49.945 96.515 ;
        RECT 46.280 96.315 46.600 96.375 ;
        RECT 49.655 96.330 49.945 96.375 ;
        RECT 66.920 96.315 67.240 96.575 ;
        RECT 30.455 96.145 30.745 96.190 ;
        RECT 40.130 96.145 40.270 96.315 ;
        RECT 30.455 96.005 40.270 96.145 ;
        RECT 48.215 96.145 48.505 96.190 ;
        RECT 63.080 96.145 63.400 96.205 ;
        RECT 48.215 96.005 63.400 96.145 ;
        RECT 30.455 95.960 30.745 96.005 ;
        RECT 28.040 95.775 28.360 95.835 ;
        RECT 31.880 95.775 32.200 95.835 ;
        RECT 28.040 95.635 32.200 95.775 ;
        RECT 28.040 95.575 28.360 95.635 ;
        RECT 31.880 95.575 32.200 95.635 ;
        RECT 29.495 95.405 29.785 95.450 ;
        RECT 30.920 95.405 31.240 95.465 ;
        RECT 29.495 95.265 31.240 95.405 ;
        RECT 29.495 95.220 29.785 95.265 ;
        RECT 30.920 95.205 31.240 95.265 ;
        RECT 32.360 95.205 32.680 95.465 ;
        RECT 32.930 95.450 33.070 96.005 ;
        RECT 48.215 95.960 48.505 96.005 ;
        RECT 63.080 95.945 63.400 96.005 ;
        RECT 33.815 95.775 34.105 95.820 ;
        RECT 57.320 95.775 57.640 95.835 ;
        RECT 65.495 95.775 65.785 95.820 ;
        RECT 33.815 95.635 40.750 95.775 ;
        RECT 33.815 95.590 34.105 95.635 ;
        RECT 40.610 95.465 40.750 95.635 ;
        RECT 57.320 95.635 65.785 95.775 ;
        RECT 57.320 95.575 57.640 95.635 ;
        RECT 65.495 95.590 65.785 95.635 ;
        RECT 32.855 95.220 33.145 95.450 ;
        RECT 40.040 95.205 40.360 95.465 ;
        RECT 40.520 95.205 40.840 95.465 ;
        RECT 56.360 95.405 56.680 95.465 ;
        RECT 57.815 95.405 58.105 95.450 ;
        RECT 56.360 95.265 58.105 95.405 ;
        RECT 56.360 95.205 56.680 95.265 ;
        RECT 57.815 95.220 58.105 95.265 ;
        RECT 27.080 95.035 27.400 95.095 ;
        RECT 27.575 95.035 27.865 95.080 ;
        RECT 27.080 94.895 27.865 95.035 ;
        RECT 27.080 94.835 27.400 94.895 ;
        RECT 27.575 94.850 27.865 94.895 ;
        RECT 38.120 94.835 38.440 95.095 ;
        RECT 39.095 95.035 39.385 95.080 ;
        RECT 42.935 95.035 43.225 95.080 ;
        RECT 45.815 95.035 46.105 95.080 ;
        RECT 47.720 95.035 48.040 95.095 ;
        RECT 52.070 95.080 52.330 95.125 ;
        RECT 52.055 95.035 52.345 95.080 ;
        RECT 54.935 95.035 55.225 95.080 ;
        RECT 58.775 95.035 59.065 95.080 ;
        RECT 39.095 94.895 59.065 95.035 ;
        RECT 39.095 94.850 39.385 94.895 ;
        RECT 42.935 94.850 43.225 94.895 ;
        RECT 45.815 94.850 46.105 94.895 ;
        RECT 47.720 94.835 48.040 94.895 ;
        RECT 52.055 94.850 52.345 94.895 ;
        RECT 54.935 94.850 55.225 94.895 ;
        RECT 58.775 94.850 59.065 94.895 ;
        RECT 59.735 94.850 60.025 95.080 ;
        RECT 52.070 94.805 52.330 94.850 ;
        RECT 59.810 94.665 59.950 94.850 ;
        RECT 57.410 94.525 59.950 94.665 ;
        RECT 57.410 94.355 57.550 94.525 ;
        RECT 57.320 94.095 57.640 94.355 ;
        RECT 10.200 93.425 69.720 93.915 ;
        RECT 47.720 93.185 48.040 93.245 ;
        RECT 34.850 93.045 48.040 93.185 ;
        RECT 28.535 92.445 28.825 92.490 ;
        RECT 31.415 92.445 31.705 92.490 ;
        RECT 34.850 92.445 34.990 93.045 ;
        RECT 47.720 92.985 48.040 93.045 ;
        RECT 47.240 92.615 47.560 92.875 ;
        RECT 35.255 92.445 35.545 92.490 ;
        RECT 28.535 92.305 35.545 92.445 ;
        RECT 28.535 92.260 28.825 92.305 ;
        RECT 31.415 92.260 31.705 92.305 ;
        RECT 35.255 92.260 35.545 92.305 ;
        RECT 39.575 92.445 39.865 92.490 ;
        RECT 40.520 92.445 40.840 92.505 ;
        RECT 42.455 92.445 42.745 92.490 ;
        RECT 46.295 92.445 46.585 92.490 ;
        RECT 39.575 92.305 46.585 92.445 ;
        RECT 39.575 92.260 39.865 92.305 ;
        RECT 40.520 92.245 40.840 92.305 ;
        RECT 42.455 92.260 42.745 92.305 ;
        RECT 46.295 92.260 46.585 92.305 ;
        RECT 34.295 92.075 34.585 92.120 ;
        RECT 45.335 92.075 45.625 92.120 ;
        RECT 46.760 92.075 47.080 92.135 ;
        RECT 34.295 91.935 35.950 92.075 ;
        RECT 34.295 91.890 34.585 91.935 ;
        RECT 24.695 91.705 24.985 91.750 ;
        RECT 27.080 91.705 27.400 91.765 ;
        RECT 24.695 91.565 27.400 91.705 ;
        RECT 24.695 91.520 24.985 91.565 ;
        RECT 27.080 91.505 27.400 91.565 ;
        RECT 24.215 90.965 24.505 91.010 ;
        RECT 25.640 90.965 25.960 91.025 ;
        RECT 24.215 90.825 25.960 90.965 ;
        RECT 24.215 90.780 24.505 90.825 ;
        RECT 25.640 90.765 25.960 90.825 ;
        RECT 26.135 90.965 26.425 91.010 ;
        RECT 26.600 90.965 26.920 91.025 ;
        RECT 26.135 90.825 26.920 90.965 ;
        RECT 35.810 90.965 35.950 91.935 ;
        RECT 45.335 91.935 47.080 92.075 ;
        RECT 45.335 91.890 45.625 91.935 ;
        RECT 46.760 91.875 47.080 91.935 ;
        RECT 36.215 91.520 36.505 91.750 ;
        RECT 40.040 91.705 40.360 91.765 ;
        RECT 43.880 91.705 44.200 91.765 ;
        RECT 47.330 91.750 47.470 92.615 ;
        RECT 56.840 92.445 57.160 92.505 ;
        RECT 55.010 92.305 57.160 92.445 ;
        RECT 55.010 92.075 55.150 92.305 ;
        RECT 56.840 92.245 57.160 92.305 ;
        RECT 57.815 92.445 58.105 92.490 ;
        RECT 58.280 92.445 58.600 92.505 ;
        RECT 61.655 92.445 61.945 92.490 ;
        RECT 64.535 92.445 64.825 92.490 ;
        RECT 57.815 92.305 64.825 92.445 ;
        RECT 57.815 92.260 58.105 92.305 ;
        RECT 58.280 92.245 58.600 92.305 ;
        RECT 61.655 92.260 61.945 92.305 ;
        RECT 64.535 92.260 64.825 92.305 ;
        RECT 52.130 91.935 55.150 92.075 ;
        RECT 56.360 92.075 56.680 92.135 ;
        RECT 58.775 92.075 59.065 92.120 ;
        RECT 56.360 91.935 59.065 92.075 ;
        RECT 47.255 91.705 47.545 91.750 ;
        RECT 40.040 91.565 47.545 91.705 ;
        RECT 36.290 91.335 36.430 91.520 ;
        RECT 40.040 91.505 40.360 91.565 ;
        RECT 43.880 91.505 44.200 91.565 ;
        RECT 47.255 91.520 47.545 91.565 ;
        RECT 51.560 91.505 51.880 91.765 ;
        RECT 38.120 91.335 38.440 91.395 ;
        RECT 52.130 91.335 52.270 91.935 ;
        RECT 56.360 91.875 56.680 91.935 ;
        RECT 58.775 91.890 59.065 91.935 ;
        RECT 52.520 91.705 52.840 91.765 ;
        RECT 54.455 91.705 54.745 91.750 ;
        RECT 52.520 91.565 54.745 91.705 ;
        RECT 52.520 91.505 52.840 91.565 ;
        RECT 54.455 91.520 54.745 91.565 ;
        RECT 66.935 91.705 67.225 91.750 ;
        RECT 68.360 91.705 68.680 91.765 ;
        RECT 66.935 91.565 68.680 91.705 ;
        RECT 66.935 91.520 67.225 91.565 ;
        RECT 68.360 91.505 68.680 91.565 ;
        RECT 67.880 91.335 68.200 91.395 ;
        RECT 36.290 91.195 52.270 91.335 ;
        RECT 53.090 91.195 68.200 91.335 ;
        RECT 38.120 91.135 38.440 91.195 ;
        RECT 37.175 90.965 37.465 91.010 ;
        RECT 37.640 90.965 37.960 91.025 ;
        RECT 35.810 90.825 37.960 90.965 ;
        RECT 26.135 90.780 26.425 90.825 ;
        RECT 26.600 90.765 26.920 90.825 ;
        RECT 37.175 90.780 37.465 90.825 ;
        RECT 37.640 90.765 37.960 90.825 ;
        RECT 39.560 90.965 39.880 91.025 ;
        RECT 48.200 90.965 48.520 91.025 ;
        RECT 53.090 91.010 53.230 91.195 ;
        RECT 67.880 91.135 68.200 91.195 ;
        RECT 39.560 90.825 48.520 90.965 ;
        RECT 39.560 90.765 39.880 90.825 ;
        RECT 48.200 90.765 48.520 90.825 ;
        RECT 53.015 90.780 53.305 91.010 ;
        RECT 55.895 90.965 56.185 91.010 ;
        RECT 61.640 90.965 61.960 91.025 ;
        RECT 55.895 90.825 61.960 90.965 ;
        RECT 55.895 90.780 56.185 90.825 ;
        RECT 61.640 90.765 61.960 90.825 ;
        RECT 10.200 90.095 69.720 90.585 ;
        RECT 36.695 89.855 36.985 89.900 ;
        RECT 38.120 89.855 38.440 89.915 ;
        RECT 36.695 89.715 38.440 89.855 ;
        RECT 36.695 89.670 36.985 89.715 ;
        RECT 38.120 89.655 38.440 89.715 ;
        RECT 40.040 89.655 40.360 89.915 ;
        RECT 42.920 89.855 43.240 89.915 ;
        RECT 55.895 89.855 56.185 89.900 ;
        RECT 56.360 89.855 56.680 89.915 ;
        RECT 42.920 89.715 51.790 89.855 ;
        RECT 42.920 89.655 43.240 89.715 ;
        RECT 35.255 89.485 35.545 89.530 ;
        RECT 40.130 89.485 40.270 89.655 ;
        RECT 35.255 89.345 40.270 89.485 ;
        RECT 40.610 89.345 46.510 89.485 ;
        RECT 35.255 89.300 35.545 89.345 ;
        RECT 25.160 89.115 25.480 89.175 ;
        RECT 39.560 89.115 39.880 89.175 ;
        RECT 25.160 88.975 33.070 89.115 ;
        RECT 25.160 88.915 25.480 88.975 ;
        RECT 25.640 88.745 25.960 88.805 ;
        RECT 27.095 88.745 27.385 88.790 ;
        RECT 25.640 88.605 27.385 88.745 ;
        RECT 25.640 88.545 25.960 88.605 ;
        RECT 27.095 88.560 27.385 88.605 ;
        RECT 25.730 88.005 25.870 88.545 ;
        RECT 32.930 88.420 33.070 88.975 ;
        RECT 38.210 88.975 39.880 89.115 ;
        RECT 35.720 88.745 36.040 88.805 ;
        RECT 38.210 88.790 38.350 88.975 ;
        RECT 39.560 88.915 39.880 88.975 ;
        RECT 40.040 88.915 40.360 89.175 ;
        RECT 40.610 89.160 40.750 89.345 ;
        RECT 46.370 89.175 46.510 89.345 ;
        RECT 47.720 89.285 48.040 89.545 ;
        RECT 51.650 89.485 51.790 89.715 ;
        RECT 55.895 89.715 56.680 89.855 ;
        RECT 55.895 89.670 56.185 89.715 ;
        RECT 56.360 89.655 56.680 89.715 ;
        RECT 66.935 89.855 67.225 89.900 ;
        RECT 68.840 89.855 69.160 89.915 ;
        RECT 66.935 89.715 69.160 89.855 ;
        RECT 66.935 89.670 67.225 89.715 ;
        RECT 68.840 89.655 69.160 89.715 ;
        RECT 56.855 89.485 57.145 89.530 ;
        RECT 57.320 89.485 57.640 89.545 ;
        RECT 51.650 89.345 57.640 89.485 ;
        RECT 56.855 89.300 57.145 89.345 ;
        RECT 57.320 89.285 57.640 89.345 ;
        RECT 57.890 89.345 65.710 89.485 ;
        RECT 40.535 88.930 40.825 89.160 ;
        RECT 43.415 89.115 43.705 89.160 ;
        RECT 41.090 88.975 43.705 89.115 ;
        RECT 38.135 88.745 38.425 88.790 ;
        RECT 35.720 88.605 38.425 88.745 ;
        RECT 40.130 88.745 40.270 88.915 ;
        RECT 41.090 88.745 41.230 88.975 ;
        RECT 43.415 88.930 43.705 88.975 ;
        RECT 46.280 88.915 46.600 89.175 ;
        RECT 47.810 88.790 47.950 89.285 ;
        RECT 49.640 89.115 49.960 89.175 ;
        RECT 57.890 89.115 58.030 89.345 ;
        RECT 49.640 88.975 58.030 89.115 ;
        RECT 58.280 89.115 58.600 89.175 ;
        RECT 65.570 89.160 65.710 89.345 ;
        RECT 59.735 89.115 60.025 89.160 ;
        RECT 58.280 88.975 60.025 89.115 ;
        RECT 49.640 88.915 49.960 88.975 ;
        RECT 58.280 88.915 58.600 88.975 ;
        RECT 59.735 88.930 60.025 88.975 ;
        RECT 65.495 88.930 65.785 89.160 ;
        RECT 47.735 88.745 48.025 88.790 ;
        RECT 40.130 88.605 41.230 88.745 ;
        RECT 42.050 88.605 48.025 88.745 ;
        RECT 35.720 88.545 36.040 88.605 ;
        RECT 38.135 88.560 38.425 88.605 ;
        RECT 26.135 88.375 26.425 88.420 ;
        RECT 29.975 88.375 30.265 88.420 ;
        RECT 32.855 88.375 33.145 88.420 ;
        RECT 40.520 88.375 40.840 88.435 ;
        RECT 42.050 88.375 42.190 88.605 ;
        RECT 47.735 88.560 48.025 88.605 ;
        RECT 55.400 88.745 55.720 88.805 ;
        RECT 57.815 88.745 58.105 88.790 ;
        RECT 60.680 88.745 61.000 88.805 ;
        RECT 55.400 88.605 61.000 88.745 ;
        RECT 55.400 88.545 55.720 88.605 ;
        RECT 57.815 88.560 58.105 88.605 ;
        RECT 60.680 88.545 61.000 88.605 ;
        RECT 26.135 88.235 40.840 88.375 ;
        RECT 26.135 88.190 26.425 88.235 ;
        RECT 29.975 88.190 30.265 88.235 ;
        RECT 32.855 88.190 33.145 88.235 ;
        RECT 40.520 88.175 40.840 88.235 ;
        RECT 41.570 88.235 42.190 88.375 ;
        RECT 45.815 88.375 46.105 88.420 ;
        RECT 46.280 88.375 46.600 88.435 ;
        RECT 45.815 88.235 46.600 88.375 ;
        RECT 41.570 88.005 41.710 88.235 ;
        RECT 45.815 88.190 46.105 88.235 ;
        RECT 46.280 88.175 46.600 88.235 ;
        RECT 46.775 88.375 47.065 88.420 ;
        RECT 50.615 88.375 50.905 88.420 ;
        RECT 52.520 88.375 52.840 88.435 ;
        RECT 53.495 88.375 53.785 88.420 ;
        RECT 46.775 88.235 53.785 88.375 ;
        RECT 46.775 88.190 47.065 88.235 ;
        RECT 50.615 88.190 50.905 88.235 ;
        RECT 52.520 88.175 52.840 88.235 ;
        RECT 53.495 88.190 53.785 88.235 ;
        RECT 61.175 88.375 61.465 88.420 ;
        RECT 65.960 88.375 66.280 88.435 ;
        RECT 61.175 88.235 66.280 88.375 ;
        RECT 61.175 88.190 61.465 88.235 ;
        RECT 65.960 88.175 66.280 88.235 ;
        RECT 54.440 88.005 54.760 88.065 ;
        RECT 25.730 87.865 41.710 88.005 ;
        RECT 42.050 87.865 54.760 88.005 ;
        RECT 37.160 87.635 37.480 87.695 ;
        RECT 40.040 87.635 40.360 87.695 ;
        RECT 42.050 87.680 42.190 87.865 ;
        RECT 54.440 87.805 54.760 87.865 ;
        RECT 55.400 88.005 55.720 88.065 ;
        RECT 65.000 88.005 65.320 88.065 ;
        RECT 55.400 87.865 65.320 88.005 ;
        RECT 55.400 87.805 55.720 87.865 ;
        RECT 65.000 87.805 65.320 87.865 ;
        RECT 37.160 87.495 40.360 87.635 ;
        RECT 37.160 87.435 37.480 87.495 ;
        RECT 40.040 87.435 40.360 87.495 ;
        RECT 41.975 87.450 42.265 87.680 ;
        RECT 44.855 87.635 45.145 87.680 ;
        RECT 53.480 87.635 53.800 87.695 ;
        RECT 44.855 87.495 53.800 87.635 ;
        RECT 44.855 87.450 45.145 87.495 ;
        RECT 53.480 87.435 53.800 87.495 ;
        RECT 10.200 86.765 69.720 87.255 ;
        RECT 28.040 86.325 28.360 86.585 ;
        RECT 35.720 86.325 36.040 86.585 ;
        RECT 37.160 86.325 37.480 86.585 ;
        RECT 37.640 86.525 37.960 86.585 ;
        RECT 46.760 86.525 47.080 86.585 ;
        RECT 37.640 86.385 47.080 86.525 ;
        RECT 37.640 86.325 37.960 86.385 ;
        RECT 46.760 86.325 47.080 86.385 ;
        RECT 50.615 86.525 50.905 86.570 ;
        RECT 53.960 86.525 54.280 86.585 ;
        RECT 50.615 86.385 54.280 86.525 ;
        RECT 50.615 86.340 50.905 86.385 ;
        RECT 53.960 86.325 54.280 86.385 ;
        RECT 55.400 86.325 55.720 86.585 ;
        RECT 57.320 86.325 57.640 86.585 ;
        RECT 58.280 86.525 58.600 86.585 ;
        RECT 62.600 86.525 62.920 86.585 ;
        RECT 58.280 86.385 62.920 86.525 ;
        RECT 58.280 86.325 58.600 86.385 ;
        RECT 62.600 86.325 62.920 86.385 ;
        RECT 66.920 86.325 67.240 86.585 ;
        RECT 26.600 86.155 26.920 86.215 ;
        RECT 55.490 86.155 55.630 86.325 ;
        RECT 26.600 86.015 55.630 86.155 ;
        RECT 57.410 86.155 57.550 86.325 ;
        RECT 57.410 86.015 60.430 86.155 ;
        RECT 26.600 85.955 26.920 86.015 ;
        RECT 39.575 85.785 39.865 85.830 ;
        RECT 40.520 85.785 40.840 85.845 ;
        RECT 52.550 85.830 52.810 85.875 ;
        RECT 60.290 85.830 60.430 86.015 ;
        RECT 60.680 85.955 61.000 86.215 ;
        RECT 42.455 85.785 42.745 85.830 ;
        RECT 46.295 85.785 46.585 85.830 ;
        RECT 39.575 85.645 46.585 85.785 ;
        RECT 39.575 85.600 39.865 85.645 ;
        RECT 40.520 85.585 40.840 85.645 ;
        RECT 42.455 85.600 42.745 85.645 ;
        RECT 46.295 85.600 46.585 85.645 ;
        RECT 52.535 85.785 52.825 85.830 ;
        RECT 55.415 85.785 55.705 85.830 ;
        RECT 59.255 85.785 59.545 85.830 ;
        RECT 52.535 85.645 59.545 85.785 ;
        RECT 52.535 85.600 52.825 85.645 ;
        RECT 55.415 85.600 55.705 85.645 ;
        RECT 59.255 85.600 59.545 85.645 ;
        RECT 60.215 85.600 60.505 85.830 ;
        RECT 60.770 85.785 60.910 85.955 ;
        RECT 62.615 85.785 62.905 85.830 ;
        RECT 60.770 85.645 62.905 85.785 ;
        RECT 62.615 85.600 62.905 85.645 ;
        RECT 52.550 85.555 52.810 85.600 ;
        RECT 26.600 85.215 26.920 85.475 ;
        RECT 34.775 85.415 35.065 85.460 ;
        RECT 40.040 85.415 40.360 85.475 ;
        RECT 34.775 85.275 40.360 85.415 ;
        RECT 34.775 85.230 35.065 85.275 ;
        RECT 40.040 85.215 40.360 85.275 ;
        RECT 42.920 85.215 43.240 85.475 ;
        RECT 43.880 85.415 44.200 85.475 ;
        RECT 45.335 85.415 45.625 85.460 ;
        RECT 43.880 85.275 45.625 85.415 ;
        RECT 43.880 85.215 44.200 85.275 ;
        RECT 45.335 85.230 45.625 85.275 ;
        RECT 46.760 85.415 47.080 85.475 ;
        RECT 58.280 85.415 58.600 85.475 ;
        RECT 63.575 85.415 63.865 85.460 ;
        RECT 46.760 85.275 58.600 85.415 ;
        RECT 46.760 85.215 47.080 85.275 ;
        RECT 58.280 85.215 58.600 85.275 ;
        RECT 58.850 85.275 63.865 85.415 ;
        RECT 14.615 85.045 14.905 85.090 ;
        RECT 21.320 85.045 21.640 85.105 ;
        RECT 14.615 84.905 21.640 85.045 ;
        RECT 43.010 85.045 43.150 85.215 ;
        RECT 47.255 85.045 47.545 85.090 ;
        RECT 43.010 84.905 47.545 85.045 ;
        RECT 14.615 84.860 14.905 84.905 ;
        RECT 21.320 84.845 21.640 84.905 ;
        RECT 47.255 84.860 47.545 84.905 ;
        RECT 53.960 85.045 54.280 85.105 ;
        RECT 58.850 85.045 58.990 85.275 ;
        RECT 63.575 85.230 63.865 85.275 ;
        RECT 53.960 84.905 58.990 85.045 ;
        RECT 53.960 84.845 54.280 84.905 ;
        RECT 65.480 84.845 65.800 85.105 ;
        RECT 13.160 84.105 13.480 84.365 ;
        RECT 10.200 83.435 69.720 83.925 ;
        RECT 111.750 73.980 112.250 96.850 ;
        RECT 112.800 77.535 113.180 94.450 ;
        RECT 113.380 92.345 113.550 99.850 ;
        RECT 113.800 93.395 114.260 93.445 ;
        RECT 113.780 92.505 114.280 93.395 ;
        RECT 114.510 92.345 114.680 93.395 ;
        RECT 113.380 91.845 113.750 92.345 ;
        RECT 114.310 91.845 114.680 92.345 ;
        RECT 113.380 91.295 113.550 91.845 ;
        RECT 113.800 91.455 114.260 91.685 ;
        RECT 114.510 91.295 114.680 91.845 ;
        RECT 113.380 90.795 113.750 91.295 ;
        RECT 114.310 90.795 114.680 91.295 ;
        RECT 113.380 90.245 113.550 90.795 ;
        RECT 113.800 90.405 114.260 90.635 ;
        RECT 114.510 90.245 114.680 90.795 ;
        RECT 113.380 89.745 113.750 90.245 ;
        RECT 114.310 89.745 114.680 90.245 ;
        RECT 113.380 89.195 113.550 89.745 ;
        RECT 113.800 89.355 114.260 89.585 ;
        RECT 114.510 89.195 114.680 89.745 ;
        RECT 113.380 88.695 113.750 89.195 ;
        RECT 114.310 88.695 114.680 89.195 ;
        RECT 113.380 87.730 113.550 88.695 ;
        RECT 113.800 88.305 114.260 88.535 ;
        RECT 114.510 87.730 114.680 88.695 ;
        RECT 113.380 87.560 114.680 87.730 ;
        RECT 113.380 86.550 113.550 87.560 ;
        RECT 113.800 86.755 114.260 86.985 ;
        RECT 114.510 86.550 114.680 87.560 ;
        RECT 113.380 85.050 113.750 86.550 ;
        RECT 114.310 85.050 114.680 86.550 ;
        RECT 113.380 84.410 113.550 85.050 ;
        RECT 113.800 84.615 114.260 84.845 ;
        RECT 114.510 84.410 114.680 85.050 ;
        RECT 113.380 82.910 113.750 84.410 ;
        RECT 114.310 82.910 114.680 84.410 ;
        RECT 113.380 82.270 113.550 82.910 ;
        RECT 113.800 82.475 114.260 82.705 ;
        RECT 114.510 82.270 114.680 82.910 ;
        RECT 113.380 80.770 113.750 82.270 ;
        RECT 114.310 80.770 114.680 82.270 ;
        RECT 113.380 80.130 113.550 80.770 ;
        RECT 113.800 80.335 114.260 80.565 ;
        RECT 114.510 80.130 114.680 80.770 ;
        RECT 113.380 78.630 113.750 80.130 ;
        RECT 114.310 78.630 114.680 80.130 ;
        RECT 113.780 77.535 114.280 78.425 ;
        RECT 114.510 77.535 114.680 78.630 ;
        RECT 114.880 77.535 115.640 95.450 ;
        RECT 115.840 92.300 116.010 99.850 ;
        RECT 116.260 93.395 116.720 99.450 ;
        RECT 116.240 92.505 116.740 93.395 ;
        RECT 115.840 90.800 116.210 92.300 ;
        RECT 116.770 90.800 117.140 92.300 ;
        RECT 115.840 90.160 116.010 90.800 ;
        RECT 116.260 90.365 116.720 90.595 ;
        RECT 116.970 90.160 117.140 90.800 ;
        RECT 115.840 88.660 116.210 90.160 ;
        RECT 116.770 88.660 117.140 90.160 ;
        RECT 115.840 88.020 116.010 88.660 ;
        RECT 116.260 88.225 116.720 88.455 ;
        RECT 116.970 88.020 117.140 88.660 ;
        RECT 115.840 86.520 116.210 88.020 ;
        RECT 116.770 86.520 117.140 88.020 ;
        RECT 115.840 85.880 116.010 86.520 ;
        RECT 116.260 86.085 116.720 86.315 ;
        RECT 116.970 85.880 117.140 86.520 ;
        RECT 115.840 84.380 116.210 85.880 ;
        RECT 116.770 84.380 117.140 85.880 ;
        RECT 115.840 82.235 116.010 84.380 ;
        RECT 116.260 83.945 116.720 84.175 ;
        RECT 116.260 82.395 116.720 82.625 ;
        RECT 116.970 82.235 117.140 84.380 ;
        RECT 115.840 81.735 116.210 82.235 ;
        RECT 116.770 81.735 117.140 82.235 ;
        RECT 115.840 81.185 116.010 81.735 ;
        RECT 116.260 81.345 116.720 81.575 ;
        RECT 116.970 81.185 117.140 81.735 ;
        RECT 115.840 80.685 116.210 81.185 ;
        RECT 116.770 80.685 117.140 81.185 ;
        RECT 115.840 80.135 116.010 80.685 ;
        RECT 116.260 80.295 116.720 80.525 ;
        RECT 116.970 80.135 117.140 80.685 ;
        RECT 115.840 79.635 116.210 80.135 ;
        RECT 116.770 79.635 117.140 80.135 ;
        RECT 115.840 79.085 116.010 79.635 ;
        RECT 116.260 79.245 116.720 79.475 ;
        RECT 116.970 79.085 117.140 79.635 ;
        RECT 115.840 78.585 116.210 79.085 ;
        RECT 116.770 78.585 117.140 79.085 ;
        RECT 115.840 77.535 116.010 78.585 ;
        RECT 116.240 77.535 116.740 78.425 ;
        RECT 113.800 77.485 114.260 77.535 ;
        RECT 116.260 77.485 116.720 77.535 ;
        RECT 116.970 77.085 117.140 78.585 ;
        RECT 117.340 77.540 118.100 94.450 ;
        RECT 118.720 93.400 119.180 93.445 ;
        RECT 118.300 92.350 118.470 93.400 ;
        RECT 118.700 92.510 119.200 93.400 ;
        RECT 119.430 92.350 119.600 93.400 ;
        RECT 118.300 91.850 118.670 92.350 ;
        RECT 119.230 91.850 119.600 92.350 ;
        RECT 118.300 91.300 118.470 91.850 ;
        RECT 118.720 91.460 119.180 91.690 ;
        RECT 119.430 91.300 119.600 91.850 ;
        RECT 118.300 90.800 118.670 91.300 ;
        RECT 119.230 90.800 119.600 91.300 ;
        RECT 118.300 90.250 118.470 90.800 ;
        RECT 118.720 90.410 119.180 90.640 ;
        RECT 119.430 90.250 119.600 90.800 ;
        RECT 118.300 89.750 118.670 90.250 ;
        RECT 119.230 89.750 119.600 90.250 ;
        RECT 118.300 89.200 118.470 89.750 ;
        RECT 118.720 89.360 119.180 89.590 ;
        RECT 119.430 89.200 119.600 89.750 ;
        RECT 118.300 88.700 118.670 89.200 ;
        RECT 119.230 88.700 119.600 89.200 ;
        RECT 118.300 87.735 118.470 88.700 ;
        RECT 118.720 88.310 119.180 88.540 ;
        RECT 119.430 87.735 119.600 88.700 ;
        RECT 118.300 87.565 119.600 87.735 ;
        RECT 118.300 86.555 118.470 87.565 ;
        RECT 118.720 86.760 119.180 86.990 ;
        RECT 119.430 86.555 119.600 87.565 ;
        RECT 118.300 85.055 118.670 86.555 ;
        RECT 119.230 85.055 119.600 86.555 ;
        RECT 118.300 84.415 118.470 85.055 ;
        RECT 118.720 84.620 119.180 84.850 ;
        RECT 119.430 84.415 119.600 85.055 ;
        RECT 118.300 82.915 118.670 84.415 ;
        RECT 119.230 82.915 119.600 84.415 ;
        RECT 118.300 82.275 118.470 82.915 ;
        RECT 118.720 82.480 119.180 82.710 ;
        RECT 119.430 82.275 119.600 82.915 ;
        RECT 118.300 80.775 118.670 82.275 ;
        RECT 119.230 80.775 119.600 82.275 ;
        RECT 118.300 80.135 118.470 80.775 ;
        RECT 118.720 80.340 119.180 80.570 ;
        RECT 119.430 80.135 119.600 80.775 ;
        RECT 118.300 78.635 118.670 80.135 ;
        RECT 119.230 78.635 119.600 80.135 ;
        RECT 118.700 77.540 119.200 78.430 ;
        RECT 117.340 77.535 117.720 77.540 ;
        RECT 118.720 77.485 119.180 77.540 ;
        RECT 119.430 77.085 119.600 78.635 ;
        RECT 119.800 92.305 120.560 134.995 ;
        RECT 123.820 134.950 125.520 134.995 ;
        RECT 126.080 134.950 127.450 135.450 ;
        RECT 128.010 134.950 129.450 135.450 ;
        RECT 121.180 134.785 121.640 134.790 ;
        RECT 121.160 124.850 121.660 134.785 ;
        RECT 123.090 129.850 123.590 134.790 ;
        RECT 123.820 133.900 125.315 134.950 ;
        RECT 125.550 130.850 126.050 134.790 ;
        RECT 127.480 134.200 127.980 134.790 ;
        RECT 121.160 92.515 121.660 102.450 ;
        RECT 121.180 92.510 121.640 92.515 ;
        RECT 123.090 92.510 123.590 97.450 ;
        RECT 123.820 92.350 125.315 93.400 ;
        RECT 125.550 92.510 126.050 96.450 ;
        RECT 127.480 92.510 127.980 93.100 ;
        RECT 128.580 92.350 129.450 134.950 ;
        RECT 129.800 127.850 130.100 136.510 ;
        RECT 130.525 136.100 130.885 136.520 ;
        RECT 130.575 128.850 130.875 134.475 ;
        RECT 132.290 131.850 132.780 151.850 ;
        RECT 134.330 150.350 134.630 151.740 ;
        RECT 134.300 149.930 134.660 150.350 ;
        RECT 133.315 148.120 133.615 149.850 ;
        RECT 134.305 149.030 134.665 149.450 ;
        RECT 134.250 148.120 134.550 148.520 ;
        RECT 135.000 144.795 135.300 149.440 ;
        RECT 134.165 143.765 134.525 144.185 ;
        RECT 133.315 129.850 133.615 136.510 ;
        RECT 134.185 136.100 134.545 136.520 ;
        RECT 134.950 135.145 135.350 135.645 ;
        RECT 134.195 130.850 134.495 134.475 ;
        RECT 134.950 125.850 135.250 135.145 ;
        RECT 135.620 132.850 136.110 150.410 ;
        RECT 140.810 150.215 141.320 150.815 ;
        RECT 143.270 150.215 143.780 150.815 ;
        RECT 137.810 149.765 138.270 149.815 ;
        RECT 140.270 149.765 140.730 149.815 ;
        RECT 136.810 132.850 137.190 149.765 ;
        RECT 137.790 148.875 138.290 149.765 ;
        RECT 138.520 148.670 138.690 149.765 ;
        RECT 137.390 147.170 137.760 148.670 ;
        RECT 138.320 147.170 138.690 148.670 ;
        RECT 137.390 146.530 137.560 147.170 ;
        RECT 137.810 146.735 138.270 146.965 ;
        RECT 138.520 146.530 138.690 147.170 ;
        RECT 137.390 145.030 137.760 146.530 ;
        RECT 138.320 145.030 138.690 146.530 ;
        RECT 137.390 144.390 137.560 145.030 ;
        RECT 137.810 144.595 138.270 144.825 ;
        RECT 138.520 144.390 138.690 145.030 ;
        RECT 137.390 142.890 137.760 144.390 ;
        RECT 138.320 142.890 138.690 144.390 ;
        RECT 137.390 142.250 137.560 142.890 ;
        RECT 137.810 142.455 138.270 142.685 ;
        RECT 138.520 142.250 138.690 142.890 ;
        RECT 137.390 140.750 137.760 142.250 ;
        RECT 138.320 140.750 138.690 142.250 ;
        RECT 137.390 139.740 137.560 140.750 ;
        RECT 137.810 140.315 138.270 140.545 ;
        RECT 138.520 139.740 138.690 140.750 ;
        RECT 137.390 139.570 138.690 139.740 ;
        RECT 137.390 138.605 137.560 139.570 ;
        RECT 137.810 138.765 138.270 138.995 ;
        RECT 138.520 138.605 138.690 139.570 ;
        RECT 137.390 138.105 137.760 138.605 ;
        RECT 138.320 138.105 138.690 138.605 ;
        RECT 137.390 137.555 137.560 138.105 ;
        RECT 137.810 137.715 138.270 137.945 ;
        RECT 138.520 137.555 138.690 138.105 ;
        RECT 137.390 137.055 137.760 137.555 ;
        RECT 138.320 137.055 138.690 137.555 ;
        RECT 137.390 136.505 137.560 137.055 ;
        RECT 137.810 136.665 138.270 136.895 ;
        RECT 138.520 136.505 138.690 137.055 ;
        RECT 137.390 136.005 137.760 136.505 ;
        RECT 138.320 136.005 138.690 136.505 ;
        RECT 137.390 135.455 137.560 136.005 ;
        RECT 137.810 135.615 138.270 135.845 ;
        RECT 138.520 135.455 138.690 136.005 ;
        RECT 137.390 134.955 137.760 135.455 ;
        RECT 138.320 134.955 138.690 135.455 ;
        RECT 137.390 127.450 137.560 134.955 ;
        RECT 137.790 133.905 138.290 134.795 ;
        RECT 138.520 133.905 138.690 134.955 ;
        RECT 137.810 133.855 138.270 133.905 ;
        RECT 138.890 131.850 139.650 149.765 ;
        RECT 139.850 148.715 140.020 149.765 ;
        RECT 140.250 148.875 140.750 149.765 ;
        RECT 140.980 148.715 141.150 150.215 ;
        RECT 139.850 148.215 140.220 148.715 ;
        RECT 140.780 148.215 141.150 148.715 ;
        RECT 139.850 147.665 140.020 148.215 ;
        RECT 140.270 147.825 140.730 148.055 ;
        RECT 140.980 147.665 141.150 148.215 ;
        RECT 139.850 147.165 140.220 147.665 ;
        RECT 140.780 147.165 141.150 147.665 ;
        RECT 139.850 146.615 140.020 147.165 ;
        RECT 140.270 146.775 140.730 147.005 ;
        RECT 140.980 146.615 141.150 147.165 ;
        RECT 139.850 146.115 140.220 146.615 ;
        RECT 140.780 146.115 141.150 146.615 ;
        RECT 139.850 145.565 140.020 146.115 ;
        RECT 140.270 145.725 140.730 145.955 ;
        RECT 140.980 145.565 141.150 146.115 ;
        RECT 139.850 145.065 140.220 145.565 ;
        RECT 140.780 145.065 141.150 145.565 ;
        RECT 139.850 142.920 140.020 145.065 ;
        RECT 140.270 144.675 140.730 144.905 ;
        RECT 140.270 143.125 140.730 143.355 ;
        RECT 140.980 142.920 141.150 145.065 ;
        RECT 139.850 141.420 140.220 142.920 ;
        RECT 140.780 141.420 141.150 142.920 ;
        RECT 139.850 140.780 140.020 141.420 ;
        RECT 140.270 140.985 140.730 141.215 ;
        RECT 140.980 140.780 141.150 141.420 ;
        RECT 139.850 139.280 140.220 140.780 ;
        RECT 140.780 139.280 141.150 140.780 ;
        RECT 139.850 138.640 140.020 139.280 ;
        RECT 140.270 138.845 140.730 139.075 ;
        RECT 140.980 138.640 141.150 139.280 ;
        RECT 139.850 137.140 140.220 138.640 ;
        RECT 140.780 137.140 141.150 138.640 ;
        RECT 139.850 136.500 140.020 137.140 ;
        RECT 140.270 136.705 140.730 136.935 ;
        RECT 140.980 136.500 141.150 137.140 ;
        RECT 139.850 135.000 140.220 136.500 ;
        RECT 140.780 135.000 141.150 136.500 ;
        RECT 141.350 149.760 141.730 149.765 ;
        RECT 142.730 149.760 143.190 149.815 ;
        RECT 139.850 127.450 140.020 135.000 ;
        RECT 140.250 133.905 140.750 134.795 ;
        RECT 140.270 127.850 140.730 133.905 ;
        RECT 141.350 132.850 142.110 149.760 ;
        RECT 142.710 148.870 143.210 149.760 ;
        RECT 143.440 148.665 143.610 150.215 ;
        RECT 142.310 147.165 142.680 148.665 ;
        RECT 143.240 147.165 143.610 148.665 ;
        RECT 142.310 146.525 142.480 147.165 ;
        RECT 142.730 146.730 143.190 146.960 ;
        RECT 143.440 146.525 143.610 147.165 ;
        RECT 142.310 145.025 142.680 146.525 ;
        RECT 143.240 145.025 143.610 146.525 ;
        RECT 142.310 144.385 142.480 145.025 ;
        RECT 142.730 144.590 143.190 144.820 ;
        RECT 143.440 144.385 143.610 145.025 ;
        RECT 142.310 142.885 142.680 144.385 ;
        RECT 143.240 142.885 143.610 144.385 ;
        RECT 142.310 142.245 142.480 142.885 ;
        RECT 142.730 142.450 143.190 142.680 ;
        RECT 143.440 142.245 143.610 142.885 ;
        RECT 142.310 140.745 142.680 142.245 ;
        RECT 143.240 140.745 143.610 142.245 ;
        RECT 142.310 139.735 142.480 140.745 ;
        RECT 142.730 140.310 143.190 140.540 ;
        RECT 143.440 139.735 143.610 140.745 ;
        RECT 142.310 139.565 143.610 139.735 ;
        RECT 142.310 138.600 142.480 139.565 ;
        RECT 142.730 138.760 143.190 138.990 ;
        RECT 143.440 138.600 143.610 139.565 ;
        RECT 142.310 138.100 142.680 138.600 ;
        RECT 143.240 138.100 143.610 138.600 ;
        RECT 142.310 137.550 142.480 138.100 ;
        RECT 142.730 137.710 143.190 137.940 ;
        RECT 143.440 137.550 143.610 138.100 ;
        RECT 142.310 137.050 142.680 137.550 ;
        RECT 143.240 137.050 143.610 137.550 ;
        RECT 142.310 136.500 142.480 137.050 ;
        RECT 142.730 136.660 143.190 136.890 ;
        RECT 143.440 136.500 143.610 137.050 ;
        RECT 142.310 136.000 142.680 136.500 ;
        RECT 143.240 136.000 143.610 136.500 ;
        RECT 142.310 135.450 142.480 136.000 ;
        RECT 142.730 135.610 143.190 135.840 ;
        RECT 143.440 135.450 143.610 136.000 ;
        RECT 142.310 134.950 142.680 135.450 ;
        RECT 143.240 134.950 143.610 135.450 ;
        RECT 142.310 133.900 142.480 134.950 ;
        RECT 142.710 133.900 143.210 134.790 ;
        RECT 143.440 133.900 143.610 134.950 ;
        RECT 143.810 144.010 144.190 149.760 ;
        RECT 143.810 142.915 144.570 144.010 ;
        RECT 145.190 143.120 145.650 143.350 ;
        RECT 147.120 143.120 147.580 143.350 ;
        RECT 147.830 142.915 149.330 150.815 ;
        RECT 143.810 141.415 145.140 142.915 ;
        RECT 145.700 141.415 147.070 142.915 ;
        RECT 147.630 141.855 149.330 142.915 ;
        RECT 147.630 141.415 149.380 141.855 ;
        RECT 143.810 140.775 144.940 141.415 ;
        RECT 145.190 140.980 145.650 141.210 ;
        RECT 145.900 140.775 146.870 141.415 ;
        RECT 147.120 140.980 147.580 141.210 ;
        RECT 147.830 140.775 149.380 141.415 ;
        RECT 143.810 139.275 145.140 140.775 ;
        RECT 145.700 139.275 147.070 140.775 ;
        RECT 147.630 139.275 149.380 140.775 ;
        RECT 152.970 139.600 153.460 151.850 ;
        RECT 154.505 151.330 154.865 151.750 ;
        RECT 154.425 149.030 154.785 149.450 ;
        RECT 154.500 148.110 154.860 148.530 ;
        RECT 155.465 148.120 155.765 149.850 ;
        RECT 154.550 144.785 154.910 145.205 ;
        RECT 143.810 138.635 144.940 139.275 ;
        RECT 145.190 138.840 145.650 139.070 ;
        RECT 145.900 138.635 146.870 139.275 ;
        RECT 147.120 138.840 147.580 139.070 ;
        RECT 147.830 138.635 149.380 139.275 ;
        RECT 149.580 138.760 150.040 138.990 ;
        RECT 151.510 138.760 151.970 138.990 ;
        RECT 143.810 137.135 145.140 138.635 ;
        RECT 145.700 137.135 147.070 138.635 ;
        RECT 147.630 138.600 149.380 138.635 ;
        RECT 152.590 138.600 153.460 139.600 ;
        RECT 147.630 138.100 149.530 138.600 ;
        RECT 150.090 138.100 151.460 138.600 ;
        RECT 152.020 138.100 153.460 138.600 ;
        RECT 147.630 137.550 149.380 138.100 ;
        RECT 149.580 137.710 150.040 137.940 ;
        RECT 150.290 137.550 151.260 138.100 ;
        RECT 151.510 137.710 151.970 137.940 ;
        RECT 152.220 137.550 153.460 138.100 ;
        RECT 147.630 137.135 149.530 137.550 ;
        RECT 143.810 136.495 144.940 137.135 ;
        RECT 145.190 136.700 145.650 136.930 ;
        RECT 145.900 136.495 146.870 137.135 ;
        RECT 147.830 137.050 149.530 137.135 ;
        RECT 150.090 137.050 151.460 137.550 ;
        RECT 152.020 137.050 153.460 137.550 ;
        RECT 147.120 136.700 147.580 136.930 ;
        RECT 147.830 136.500 149.380 137.050 ;
        RECT 149.580 136.660 150.040 136.890 ;
        RECT 150.290 136.500 151.260 137.050 ;
        RECT 151.510 136.660 151.970 136.890 ;
        RECT 152.220 136.500 153.460 137.050 ;
        RECT 147.830 136.495 149.530 136.500 ;
        RECT 143.810 134.995 145.140 136.495 ;
        RECT 145.700 134.995 147.070 136.495 ;
        RECT 147.630 136.000 149.530 136.495 ;
        RECT 150.090 136.000 151.460 136.500 ;
        RECT 152.020 136.000 153.460 136.500 ;
        RECT 147.630 135.450 149.380 136.000 ;
        RECT 149.580 135.610 150.040 135.840 ;
        RECT 150.290 135.450 151.260 136.000 ;
        RECT 151.510 135.610 151.970 135.840 ;
        RECT 152.220 135.450 153.460 136.000 ;
        RECT 147.630 134.995 149.530 135.450 ;
        RECT 142.730 133.855 143.190 133.900 ;
        RECT 137.220 126.850 137.730 127.450 ;
        RECT 139.680 126.850 140.190 127.450 ;
        RECT 136.810 116.900 137.310 126.450 ;
        RECT 137.810 124.200 138.310 125.450 ;
        RECT 136.760 116.400 137.360 116.900 ;
        RECT 123.820 92.305 125.520 92.350 ;
        RECT 119.800 90.805 121.130 92.305 ;
        RECT 121.690 90.805 123.060 92.305 ;
        RECT 123.620 91.850 125.520 92.305 ;
        RECT 126.080 91.850 127.450 92.350 ;
        RECT 128.010 91.850 129.450 92.350 ;
        RECT 123.620 91.300 125.315 91.850 ;
        RECT 125.570 91.460 126.030 91.690 ;
        RECT 126.280 91.300 127.250 91.850 ;
        RECT 127.500 91.460 127.960 91.690 ;
        RECT 128.210 91.300 129.450 91.850 ;
        RECT 123.620 90.805 125.520 91.300 ;
        RECT 119.800 90.165 120.930 90.805 ;
        RECT 121.180 90.370 121.640 90.600 ;
        RECT 121.890 90.165 122.860 90.805 ;
        RECT 123.820 90.800 125.520 90.805 ;
        RECT 126.080 90.800 127.450 91.300 ;
        RECT 128.010 90.800 129.450 91.300 ;
        RECT 123.110 90.370 123.570 90.600 ;
        RECT 123.820 90.250 125.315 90.800 ;
        RECT 125.570 90.410 126.030 90.640 ;
        RECT 126.280 90.250 127.250 90.800 ;
        RECT 127.500 90.410 127.960 90.640 ;
        RECT 128.210 90.250 129.450 90.800 ;
        RECT 129.800 90.790 130.100 99.450 ;
        RECT 130.575 92.825 130.875 98.450 ;
        RECT 130.525 90.780 130.885 91.200 ;
        RECT 123.820 90.165 125.520 90.250 ;
        RECT 119.800 88.665 121.130 90.165 ;
        RECT 121.690 88.665 123.060 90.165 ;
        RECT 123.620 89.750 125.520 90.165 ;
        RECT 126.080 89.750 127.450 90.250 ;
        RECT 128.010 89.750 129.450 90.250 ;
        RECT 123.620 89.200 125.315 89.750 ;
        RECT 125.570 89.360 126.030 89.590 ;
        RECT 126.280 89.200 127.250 89.750 ;
        RECT 127.500 89.360 127.960 89.590 ;
        RECT 128.210 89.200 129.450 89.750 ;
        RECT 123.620 88.700 125.520 89.200 ;
        RECT 126.080 88.700 127.450 89.200 ;
        RECT 128.010 88.700 129.450 89.200 ;
        RECT 123.620 88.665 125.315 88.700 ;
        RECT 119.800 88.025 120.930 88.665 ;
        RECT 121.180 88.230 121.640 88.460 ;
        RECT 121.890 88.025 122.860 88.665 ;
        RECT 123.110 88.230 123.570 88.460 ;
        RECT 123.820 88.025 125.315 88.665 ;
        RECT 125.570 88.310 126.030 88.540 ;
        RECT 127.500 88.310 127.960 88.540 ;
        RECT 119.800 86.525 121.130 88.025 ;
        RECT 121.690 86.525 123.060 88.025 ;
        RECT 123.620 86.525 125.315 88.025 ;
        RECT 128.580 87.700 129.450 88.700 ;
        RECT 119.800 85.885 120.930 86.525 ;
        RECT 121.180 86.090 121.640 86.320 ;
        RECT 121.890 85.885 122.860 86.525 ;
        RECT 123.110 86.090 123.570 86.320 ;
        RECT 123.820 85.885 125.315 86.525 ;
        RECT 119.800 84.385 121.130 85.885 ;
        RECT 121.690 84.385 123.060 85.885 ;
        RECT 123.620 85.615 125.315 85.885 ;
        RECT 123.620 85.445 125.370 85.615 ;
        RECT 123.620 84.385 125.320 85.445 ;
        RECT 119.800 83.290 120.560 84.385 ;
        RECT 121.180 83.950 121.640 84.180 ;
        RECT 123.110 83.950 123.570 84.180 ;
        RECT 119.800 77.540 120.180 83.290 ;
        RECT 116.800 76.485 117.310 77.085 ;
        RECT 119.260 76.485 119.770 77.085 ;
        RECT 123.820 76.485 125.320 84.385 ;
        RECT 128.960 75.450 129.450 87.700 ;
        RECT 130.540 82.095 130.900 82.515 ;
        RECT 130.490 78.770 130.850 79.190 ;
        RECT 130.415 77.850 130.775 78.270 ;
        RECT 131.455 77.450 131.755 79.180 ;
        RECT 130.495 75.550 130.855 75.970 ;
        RECT 132.290 75.450 132.780 95.450 ;
        RECT 133.315 90.790 133.615 97.450 ;
        RECT 134.195 92.825 134.495 96.450 ;
        RECT 134.950 92.155 135.250 101.450 ;
        RECT 136.810 100.850 137.310 116.400 ;
        RECT 137.760 107.400 138.360 107.900 ;
        RECT 137.810 101.850 138.310 107.400 ;
        RECT 137.220 99.850 137.730 100.450 ;
        RECT 139.680 99.850 140.190 100.450 ;
        RECT 134.950 91.655 135.350 92.155 ;
        RECT 134.185 90.780 134.545 91.200 ;
        RECT 134.165 83.115 134.525 83.535 ;
        RECT 133.315 77.450 133.615 79.180 ;
        RECT 134.250 78.780 134.550 79.180 ;
        RECT 134.305 77.850 134.665 78.270 ;
        RECT 135.000 77.860 135.300 82.505 ;
        RECT 134.300 76.950 134.660 77.370 ;
        RECT 134.330 75.560 134.630 76.950 ;
        RECT 135.620 76.890 136.110 94.450 ;
        RECT 136.810 77.535 137.190 94.450 ;
        RECT 137.390 92.345 137.560 99.850 ;
        RECT 137.810 93.395 138.270 93.445 ;
        RECT 137.790 92.505 138.290 93.395 ;
        RECT 138.520 92.345 138.690 93.395 ;
        RECT 137.390 91.845 137.760 92.345 ;
        RECT 138.320 91.845 138.690 92.345 ;
        RECT 137.390 91.295 137.560 91.845 ;
        RECT 137.810 91.455 138.270 91.685 ;
        RECT 138.520 91.295 138.690 91.845 ;
        RECT 137.390 90.795 137.760 91.295 ;
        RECT 138.320 90.795 138.690 91.295 ;
        RECT 137.390 90.245 137.560 90.795 ;
        RECT 137.810 90.405 138.270 90.635 ;
        RECT 138.520 90.245 138.690 90.795 ;
        RECT 137.390 89.745 137.760 90.245 ;
        RECT 138.320 89.745 138.690 90.245 ;
        RECT 137.390 89.195 137.560 89.745 ;
        RECT 137.810 89.355 138.270 89.585 ;
        RECT 138.520 89.195 138.690 89.745 ;
        RECT 137.390 88.695 137.760 89.195 ;
        RECT 138.320 88.695 138.690 89.195 ;
        RECT 137.390 87.730 137.560 88.695 ;
        RECT 137.810 88.305 138.270 88.535 ;
        RECT 138.520 87.730 138.690 88.695 ;
        RECT 137.390 87.560 138.690 87.730 ;
        RECT 137.390 86.550 137.560 87.560 ;
        RECT 137.810 86.755 138.270 86.985 ;
        RECT 138.520 86.550 138.690 87.560 ;
        RECT 137.390 85.050 137.760 86.550 ;
        RECT 138.320 85.050 138.690 86.550 ;
        RECT 137.390 84.410 137.560 85.050 ;
        RECT 137.810 84.615 138.270 84.845 ;
        RECT 138.520 84.410 138.690 85.050 ;
        RECT 137.390 82.910 137.760 84.410 ;
        RECT 138.320 82.910 138.690 84.410 ;
        RECT 137.390 82.270 137.560 82.910 ;
        RECT 137.810 82.475 138.270 82.705 ;
        RECT 138.520 82.270 138.690 82.910 ;
        RECT 137.390 80.770 137.760 82.270 ;
        RECT 138.320 80.770 138.690 82.270 ;
        RECT 137.390 80.130 137.560 80.770 ;
        RECT 137.810 80.335 138.270 80.565 ;
        RECT 138.520 80.130 138.690 80.770 ;
        RECT 137.390 78.630 137.760 80.130 ;
        RECT 138.320 78.630 138.690 80.130 ;
        RECT 137.790 77.535 138.290 78.425 ;
        RECT 138.520 77.535 138.690 78.630 ;
        RECT 138.890 77.535 139.650 95.450 ;
        RECT 139.850 92.300 140.020 99.850 ;
        RECT 140.270 93.395 140.730 99.450 ;
        RECT 140.250 92.505 140.750 93.395 ;
        RECT 139.850 90.800 140.220 92.300 ;
        RECT 140.780 90.800 141.150 92.300 ;
        RECT 139.850 90.160 140.020 90.800 ;
        RECT 140.270 90.365 140.730 90.595 ;
        RECT 140.980 90.160 141.150 90.800 ;
        RECT 139.850 88.660 140.220 90.160 ;
        RECT 140.780 88.660 141.150 90.160 ;
        RECT 139.850 88.020 140.020 88.660 ;
        RECT 140.270 88.225 140.730 88.455 ;
        RECT 140.980 88.020 141.150 88.660 ;
        RECT 139.850 86.520 140.220 88.020 ;
        RECT 140.780 86.520 141.150 88.020 ;
        RECT 139.850 85.880 140.020 86.520 ;
        RECT 140.270 86.085 140.730 86.315 ;
        RECT 140.980 85.880 141.150 86.520 ;
        RECT 139.850 84.380 140.220 85.880 ;
        RECT 140.780 84.380 141.150 85.880 ;
        RECT 139.850 82.235 140.020 84.380 ;
        RECT 140.270 83.945 140.730 84.175 ;
        RECT 140.270 82.395 140.730 82.625 ;
        RECT 140.980 82.235 141.150 84.380 ;
        RECT 139.850 81.735 140.220 82.235 ;
        RECT 140.780 81.735 141.150 82.235 ;
        RECT 139.850 81.185 140.020 81.735 ;
        RECT 140.270 81.345 140.730 81.575 ;
        RECT 140.980 81.185 141.150 81.735 ;
        RECT 139.850 80.685 140.220 81.185 ;
        RECT 140.780 80.685 141.150 81.185 ;
        RECT 139.850 80.135 140.020 80.685 ;
        RECT 140.270 80.295 140.730 80.525 ;
        RECT 140.980 80.135 141.150 80.685 ;
        RECT 139.850 79.635 140.220 80.135 ;
        RECT 140.780 79.635 141.150 80.135 ;
        RECT 139.850 79.085 140.020 79.635 ;
        RECT 140.270 79.245 140.730 79.475 ;
        RECT 140.980 79.085 141.150 79.635 ;
        RECT 139.850 78.585 140.220 79.085 ;
        RECT 140.780 78.585 141.150 79.085 ;
        RECT 139.850 77.535 140.020 78.585 ;
        RECT 140.250 77.535 140.750 78.425 ;
        RECT 137.810 77.485 138.270 77.535 ;
        RECT 140.270 77.485 140.730 77.535 ;
        RECT 140.980 77.085 141.150 78.585 ;
        RECT 141.350 77.540 142.110 94.450 ;
        RECT 142.730 93.400 143.190 93.445 ;
        RECT 142.310 92.350 142.480 93.400 ;
        RECT 142.710 92.510 143.210 93.400 ;
        RECT 143.440 92.350 143.610 93.400 ;
        RECT 142.310 91.850 142.680 92.350 ;
        RECT 143.240 91.850 143.610 92.350 ;
        RECT 142.310 91.300 142.480 91.850 ;
        RECT 142.730 91.460 143.190 91.690 ;
        RECT 143.440 91.300 143.610 91.850 ;
        RECT 142.310 90.800 142.680 91.300 ;
        RECT 143.240 90.800 143.610 91.300 ;
        RECT 142.310 90.250 142.480 90.800 ;
        RECT 142.730 90.410 143.190 90.640 ;
        RECT 143.440 90.250 143.610 90.800 ;
        RECT 142.310 89.750 142.680 90.250 ;
        RECT 143.240 89.750 143.610 90.250 ;
        RECT 142.310 89.200 142.480 89.750 ;
        RECT 142.730 89.360 143.190 89.590 ;
        RECT 143.440 89.200 143.610 89.750 ;
        RECT 142.310 88.700 142.680 89.200 ;
        RECT 143.240 88.700 143.610 89.200 ;
        RECT 142.310 87.735 142.480 88.700 ;
        RECT 142.730 88.310 143.190 88.540 ;
        RECT 143.440 87.735 143.610 88.700 ;
        RECT 142.310 87.565 143.610 87.735 ;
        RECT 142.310 86.555 142.480 87.565 ;
        RECT 142.730 86.760 143.190 86.990 ;
        RECT 143.440 86.555 143.610 87.565 ;
        RECT 142.310 85.055 142.680 86.555 ;
        RECT 143.240 85.055 143.610 86.555 ;
        RECT 142.310 84.415 142.480 85.055 ;
        RECT 142.730 84.620 143.190 84.850 ;
        RECT 143.440 84.415 143.610 85.055 ;
        RECT 142.310 82.915 142.680 84.415 ;
        RECT 143.240 82.915 143.610 84.415 ;
        RECT 142.310 82.275 142.480 82.915 ;
        RECT 142.730 82.480 143.190 82.710 ;
        RECT 143.440 82.275 143.610 82.915 ;
        RECT 142.310 80.775 142.680 82.275 ;
        RECT 143.240 80.775 143.610 82.275 ;
        RECT 142.310 80.135 142.480 80.775 ;
        RECT 142.730 80.340 143.190 80.570 ;
        RECT 143.440 80.135 143.610 80.775 ;
        RECT 142.310 78.635 142.680 80.135 ;
        RECT 143.240 78.635 143.610 80.135 ;
        RECT 142.710 77.540 143.210 78.430 ;
        RECT 141.350 77.535 141.730 77.540 ;
        RECT 142.730 77.485 143.190 77.540 ;
        RECT 143.440 77.085 143.610 78.635 ;
        RECT 143.810 92.305 144.570 134.995 ;
        RECT 147.830 134.950 149.530 134.995 ;
        RECT 150.090 134.950 151.460 135.450 ;
        RECT 152.020 134.950 153.460 135.450 ;
        RECT 145.190 134.785 145.650 134.790 ;
        RECT 145.170 124.850 145.670 134.785 ;
        RECT 147.100 129.850 147.600 134.790 ;
        RECT 147.830 133.900 149.380 134.950 ;
        RECT 149.560 130.850 150.060 134.790 ;
        RECT 151.490 134.200 151.990 134.790 ;
        RECT 145.170 92.515 145.670 102.450 ;
        RECT 145.190 92.510 145.650 92.515 ;
        RECT 147.100 92.510 147.600 97.450 ;
        RECT 147.830 92.350 149.380 93.400 ;
        RECT 149.560 92.510 150.060 96.450 ;
        RECT 151.490 92.510 151.990 93.100 ;
        RECT 152.590 92.350 153.460 134.950 ;
        RECT 153.810 127.850 154.110 136.510 ;
        RECT 154.535 136.100 154.895 136.520 ;
        RECT 154.585 128.850 154.885 134.475 ;
        RECT 156.300 131.850 156.790 151.850 ;
        RECT 158.340 150.350 158.640 151.740 ;
        RECT 158.310 149.930 158.670 150.350 ;
        RECT 157.325 148.120 157.625 149.850 ;
        RECT 158.315 149.030 158.675 149.450 ;
        RECT 158.260 148.120 158.560 148.520 ;
        RECT 159.010 144.795 159.310 149.440 ;
        RECT 158.175 143.765 158.535 144.185 ;
        RECT 157.325 129.850 157.625 136.510 ;
        RECT 158.195 136.100 158.555 136.520 ;
        RECT 158.960 135.145 159.360 135.645 ;
        RECT 158.205 130.850 158.505 134.475 ;
        RECT 158.960 125.850 159.260 135.145 ;
        RECT 159.630 132.850 160.120 150.410 ;
        RECT 164.820 150.215 165.330 150.815 ;
        RECT 167.280 150.215 167.790 150.815 ;
        RECT 161.820 149.765 162.280 149.815 ;
        RECT 164.280 149.765 164.740 149.815 ;
        RECT 160.820 132.850 161.200 149.765 ;
        RECT 161.800 148.875 162.300 149.765 ;
        RECT 162.530 148.670 162.700 149.765 ;
        RECT 161.400 147.170 161.770 148.670 ;
        RECT 162.330 147.170 162.700 148.670 ;
        RECT 161.400 146.530 161.570 147.170 ;
        RECT 161.820 146.735 162.280 146.965 ;
        RECT 162.530 146.530 162.700 147.170 ;
        RECT 161.400 145.030 161.770 146.530 ;
        RECT 162.330 145.030 162.700 146.530 ;
        RECT 161.400 144.390 161.570 145.030 ;
        RECT 161.820 144.595 162.280 144.825 ;
        RECT 162.530 144.390 162.700 145.030 ;
        RECT 161.400 142.890 161.770 144.390 ;
        RECT 162.330 142.890 162.700 144.390 ;
        RECT 161.400 142.250 161.570 142.890 ;
        RECT 161.820 142.455 162.280 142.685 ;
        RECT 162.530 142.250 162.700 142.890 ;
        RECT 161.400 140.750 161.770 142.250 ;
        RECT 162.330 140.750 162.700 142.250 ;
        RECT 161.400 139.740 161.570 140.750 ;
        RECT 161.820 140.315 162.280 140.545 ;
        RECT 162.530 139.740 162.700 140.750 ;
        RECT 161.400 139.570 162.700 139.740 ;
        RECT 161.400 138.605 161.570 139.570 ;
        RECT 161.820 138.765 162.280 138.995 ;
        RECT 162.530 138.605 162.700 139.570 ;
        RECT 161.400 138.105 161.770 138.605 ;
        RECT 162.330 138.105 162.700 138.605 ;
        RECT 161.400 137.555 161.570 138.105 ;
        RECT 161.820 137.715 162.280 137.945 ;
        RECT 162.530 137.555 162.700 138.105 ;
        RECT 161.400 137.055 161.770 137.555 ;
        RECT 162.330 137.055 162.700 137.555 ;
        RECT 161.400 136.505 161.570 137.055 ;
        RECT 161.820 136.665 162.280 136.895 ;
        RECT 162.530 136.505 162.700 137.055 ;
        RECT 161.400 136.005 161.770 136.505 ;
        RECT 162.330 136.005 162.700 136.505 ;
        RECT 161.400 135.455 161.570 136.005 ;
        RECT 161.820 135.615 162.280 135.845 ;
        RECT 162.530 135.455 162.700 136.005 ;
        RECT 161.400 134.955 161.770 135.455 ;
        RECT 162.330 134.955 162.700 135.455 ;
        RECT 161.400 127.450 161.570 134.955 ;
        RECT 161.800 133.905 162.300 134.795 ;
        RECT 162.530 133.905 162.700 134.955 ;
        RECT 161.820 133.855 162.280 133.905 ;
        RECT 162.900 131.850 163.660 149.765 ;
        RECT 163.860 148.715 164.030 149.765 ;
        RECT 164.260 148.875 164.760 149.765 ;
        RECT 164.990 148.715 165.160 150.215 ;
        RECT 163.860 148.215 164.230 148.715 ;
        RECT 164.790 148.215 165.160 148.715 ;
        RECT 163.860 147.665 164.030 148.215 ;
        RECT 164.280 147.825 164.740 148.055 ;
        RECT 164.990 147.665 165.160 148.215 ;
        RECT 163.860 147.165 164.230 147.665 ;
        RECT 164.790 147.165 165.160 147.665 ;
        RECT 163.860 146.615 164.030 147.165 ;
        RECT 164.280 146.775 164.740 147.005 ;
        RECT 164.990 146.615 165.160 147.165 ;
        RECT 163.860 146.115 164.230 146.615 ;
        RECT 164.790 146.115 165.160 146.615 ;
        RECT 163.860 145.565 164.030 146.115 ;
        RECT 164.280 145.725 164.740 145.955 ;
        RECT 164.990 145.565 165.160 146.115 ;
        RECT 163.860 145.065 164.230 145.565 ;
        RECT 164.790 145.065 165.160 145.565 ;
        RECT 163.860 142.920 164.030 145.065 ;
        RECT 164.280 144.675 164.740 144.905 ;
        RECT 164.280 143.125 164.740 143.355 ;
        RECT 164.990 142.920 165.160 145.065 ;
        RECT 163.860 141.420 164.230 142.920 ;
        RECT 164.790 141.420 165.160 142.920 ;
        RECT 163.860 140.780 164.030 141.420 ;
        RECT 164.280 140.985 164.740 141.215 ;
        RECT 164.990 140.780 165.160 141.420 ;
        RECT 163.860 139.280 164.230 140.780 ;
        RECT 164.790 139.280 165.160 140.780 ;
        RECT 163.860 138.640 164.030 139.280 ;
        RECT 164.280 138.845 164.740 139.075 ;
        RECT 164.990 138.640 165.160 139.280 ;
        RECT 163.860 137.140 164.230 138.640 ;
        RECT 164.790 137.140 165.160 138.640 ;
        RECT 163.860 136.500 164.030 137.140 ;
        RECT 164.280 136.705 164.740 136.935 ;
        RECT 164.990 136.500 165.160 137.140 ;
        RECT 163.860 135.000 164.230 136.500 ;
        RECT 164.790 135.000 165.160 136.500 ;
        RECT 165.360 149.760 165.740 149.765 ;
        RECT 166.740 149.760 167.200 149.815 ;
        RECT 163.860 127.450 164.030 135.000 ;
        RECT 164.260 133.905 164.760 134.795 ;
        RECT 164.280 127.850 164.740 133.905 ;
        RECT 165.360 132.850 166.120 149.760 ;
        RECT 166.720 148.870 167.220 149.760 ;
        RECT 167.450 148.665 167.620 150.215 ;
        RECT 166.320 147.165 166.690 148.665 ;
        RECT 167.250 147.165 167.620 148.665 ;
        RECT 166.320 146.525 166.490 147.165 ;
        RECT 166.740 146.730 167.200 146.960 ;
        RECT 167.450 146.525 167.620 147.165 ;
        RECT 166.320 145.025 166.690 146.525 ;
        RECT 167.250 145.025 167.620 146.525 ;
        RECT 166.320 144.385 166.490 145.025 ;
        RECT 166.740 144.590 167.200 144.820 ;
        RECT 167.450 144.385 167.620 145.025 ;
        RECT 166.320 142.885 166.690 144.385 ;
        RECT 167.250 142.885 167.620 144.385 ;
        RECT 166.320 142.245 166.490 142.885 ;
        RECT 166.740 142.450 167.200 142.680 ;
        RECT 167.450 142.245 167.620 142.885 ;
        RECT 166.320 140.745 166.690 142.245 ;
        RECT 167.250 140.745 167.620 142.245 ;
        RECT 166.320 139.735 166.490 140.745 ;
        RECT 166.740 140.310 167.200 140.540 ;
        RECT 167.450 139.735 167.620 140.745 ;
        RECT 166.320 139.565 167.620 139.735 ;
        RECT 166.320 138.600 166.490 139.565 ;
        RECT 166.740 138.760 167.200 138.990 ;
        RECT 167.450 138.600 167.620 139.565 ;
        RECT 166.320 138.100 166.690 138.600 ;
        RECT 167.250 138.100 167.620 138.600 ;
        RECT 166.320 137.550 166.490 138.100 ;
        RECT 166.740 137.710 167.200 137.940 ;
        RECT 167.450 137.550 167.620 138.100 ;
        RECT 166.320 137.050 166.690 137.550 ;
        RECT 167.250 137.050 167.620 137.550 ;
        RECT 166.320 136.500 166.490 137.050 ;
        RECT 166.740 136.660 167.200 136.890 ;
        RECT 167.450 136.500 167.620 137.050 ;
        RECT 166.320 136.000 166.690 136.500 ;
        RECT 167.250 136.000 167.620 136.500 ;
        RECT 166.320 135.450 166.490 136.000 ;
        RECT 166.740 135.610 167.200 135.840 ;
        RECT 167.450 135.450 167.620 136.000 ;
        RECT 166.320 134.950 166.690 135.450 ;
        RECT 167.250 134.950 167.620 135.450 ;
        RECT 166.320 133.900 166.490 134.950 ;
        RECT 166.720 133.900 167.220 134.790 ;
        RECT 167.450 133.900 167.620 134.950 ;
        RECT 167.820 144.010 168.200 149.760 ;
        RECT 167.820 142.915 168.580 144.010 ;
        RECT 169.200 143.120 169.660 143.350 ;
        RECT 171.130 143.120 171.590 143.350 ;
        RECT 171.840 142.915 173.340 150.815 ;
        RECT 167.820 141.415 169.150 142.915 ;
        RECT 169.710 141.415 171.080 142.915 ;
        RECT 171.640 141.685 173.340 142.915 ;
        RECT 171.640 141.415 173.335 141.685 ;
        RECT 167.820 140.775 168.950 141.415 ;
        RECT 169.200 140.980 169.660 141.210 ;
        RECT 169.910 140.775 170.880 141.415 ;
        RECT 171.130 140.980 171.590 141.210 ;
        RECT 171.840 140.775 173.335 141.415 ;
        RECT 167.820 139.275 169.150 140.775 ;
        RECT 169.710 139.275 171.080 140.775 ;
        RECT 171.640 139.275 173.335 140.775 ;
        RECT 176.980 139.600 177.470 151.850 ;
        RECT 178.515 151.330 178.875 151.750 ;
        RECT 178.435 149.030 178.795 149.450 ;
        RECT 178.510 148.110 178.870 148.530 ;
        RECT 179.475 148.120 179.775 149.850 ;
        RECT 178.560 144.785 178.920 145.205 ;
        RECT 167.820 138.635 168.950 139.275 ;
        RECT 169.200 138.840 169.660 139.070 ;
        RECT 169.910 138.635 170.880 139.275 ;
        RECT 171.130 138.840 171.590 139.070 ;
        RECT 171.840 138.635 173.335 139.275 ;
        RECT 173.590 138.760 174.050 138.990 ;
        RECT 175.520 138.760 175.980 138.990 ;
        RECT 167.820 137.135 169.150 138.635 ;
        RECT 169.710 137.135 171.080 138.635 ;
        RECT 171.640 138.600 173.335 138.635 ;
        RECT 176.600 138.600 177.470 139.600 ;
        RECT 171.640 138.100 173.540 138.600 ;
        RECT 174.100 138.100 175.470 138.600 ;
        RECT 176.030 138.100 177.470 138.600 ;
        RECT 171.640 137.550 173.335 138.100 ;
        RECT 173.590 137.710 174.050 137.940 ;
        RECT 174.300 137.550 175.270 138.100 ;
        RECT 175.520 137.710 175.980 137.940 ;
        RECT 176.230 137.550 177.470 138.100 ;
        RECT 171.640 137.135 173.540 137.550 ;
        RECT 167.820 136.495 168.950 137.135 ;
        RECT 169.200 136.700 169.660 136.930 ;
        RECT 169.910 136.495 170.880 137.135 ;
        RECT 171.840 137.050 173.540 137.135 ;
        RECT 174.100 137.050 175.470 137.550 ;
        RECT 176.030 137.050 177.470 137.550 ;
        RECT 171.130 136.700 171.590 136.930 ;
        RECT 171.840 136.500 173.335 137.050 ;
        RECT 173.590 136.660 174.050 136.890 ;
        RECT 174.300 136.500 175.270 137.050 ;
        RECT 175.520 136.660 175.980 136.890 ;
        RECT 176.230 136.500 177.470 137.050 ;
        RECT 171.840 136.495 173.540 136.500 ;
        RECT 167.820 134.995 169.150 136.495 ;
        RECT 169.710 134.995 171.080 136.495 ;
        RECT 171.640 136.000 173.540 136.495 ;
        RECT 174.100 136.000 175.470 136.500 ;
        RECT 176.030 136.000 177.470 136.500 ;
        RECT 171.640 135.450 173.335 136.000 ;
        RECT 173.590 135.610 174.050 135.840 ;
        RECT 174.300 135.450 175.270 136.000 ;
        RECT 175.520 135.610 175.980 135.840 ;
        RECT 176.230 135.450 177.470 136.000 ;
        RECT 171.640 134.995 173.540 135.450 ;
        RECT 166.740 133.855 167.200 133.900 ;
        RECT 161.230 126.850 161.740 127.450 ;
        RECT 163.690 126.850 164.200 127.450 ;
        RECT 160.820 115.900 161.320 126.450 ;
        RECT 161.815 125.400 162.315 125.450 ;
        RECT 161.815 124.850 162.320 125.400 ;
        RECT 161.820 124.200 162.320 124.850 ;
        RECT 160.770 115.400 161.370 115.900 ;
        RECT 147.830 92.305 149.530 92.350 ;
        RECT 143.810 90.805 145.140 92.305 ;
        RECT 145.700 90.805 147.070 92.305 ;
        RECT 147.630 91.850 149.530 92.305 ;
        RECT 150.090 91.850 151.460 92.350 ;
        RECT 152.020 91.850 153.460 92.350 ;
        RECT 147.630 91.300 149.380 91.850 ;
        RECT 149.580 91.460 150.040 91.690 ;
        RECT 150.290 91.300 151.260 91.850 ;
        RECT 151.510 91.460 151.970 91.690 ;
        RECT 152.220 91.300 153.460 91.850 ;
        RECT 147.630 90.805 149.530 91.300 ;
        RECT 143.810 90.165 144.940 90.805 ;
        RECT 145.190 90.370 145.650 90.600 ;
        RECT 145.900 90.165 146.870 90.805 ;
        RECT 147.830 90.800 149.530 90.805 ;
        RECT 150.090 90.800 151.460 91.300 ;
        RECT 152.020 90.800 153.460 91.300 ;
        RECT 147.120 90.370 147.580 90.600 ;
        RECT 147.830 90.250 149.380 90.800 ;
        RECT 149.580 90.410 150.040 90.640 ;
        RECT 150.290 90.250 151.260 90.800 ;
        RECT 151.510 90.410 151.970 90.640 ;
        RECT 152.220 90.250 153.460 90.800 ;
        RECT 153.810 90.790 154.110 99.450 ;
        RECT 154.585 92.825 154.885 98.450 ;
        RECT 154.535 90.780 154.895 91.200 ;
        RECT 147.830 90.165 149.530 90.250 ;
        RECT 143.810 88.665 145.140 90.165 ;
        RECT 145.700 88.665 147.070 90.165 ;
        RECT 147.630 89.750 149.530 90.165 ;
        RECT 150.090 89.750 151.460 90.250 ;
        RECT 152.020 89.750 153.460 90.250 ;
        RECT 147.630 89.200 149.380 89.750 ;
        RECT 149.580 89.360 150.040 89.590 ;
        RECT 150.290 89.200 151.260 89.750 ;
        RECT 151.510 89.360 151.970 89.590 ;
        RECT 152.220 89.200 153.460 89.750 ;
        RECT 147.630 88.700 149.530 89.200 ;
        RECT 150.090 88.700 151.460 89.200 ;
        RECT 152.020 88.700 153.460 89.200 ;
        RECT 147.630 88.665 149.380 88.700 ;
        RECT 143.810 88.025 144.940 88.665 ;
        RECT 145.190 88.230 145.650 88.460 ;
        RECT 145.900 88.025 146.870 88.665 ;
        RECT 147.120 88.230 147.580 88.460 ;
        RECT 147.830 88.025 149.380 88.665 ;
        RECT 149.580 88.310 150.040 88.540 ;
        RECT 151.510 88.310 151.970 88.540 ;
        RECT 143.810 86.525 145.140 88.025 ;
        RECT 145.700 86.525 147.070 88.025 ;
        RECT 147.630 86.525 149.380 88.025 ;
        RECT 152.590 87.700 153.460 88.700 ;
        RECT 143.810 85.885 144.940 86.525 ;
        RECT 145.190 86.090 145.650 86.320 ;
        RECT 145.900 85.885 146.870 86.525 ;
        RECT 147.120 86.090 147.580 86.320 ;
        RECT 147.830 85.885 149.380 86.525 ;
        RECT 143.810 84.385 145.140 85.885 ;
        RECT 145.700 84.385 147.070 85.885 ;
        RECT 147.630 85.445 149.380 85.885 ;
        RECT 147.630 84.385 149.330 85.445 ;
        RECT 143.810 83.290 144.570 84.385 ;
        RECT 145.190 83.950 145.650 84.180 ;
        RECT 147.120 83.950 147.580 84.180 ;
        RECT 143.810 77.540 144.190 83.290 ;
        RECT 140.810 76.485 141.320 77.085 ;
        RECT 143.270 76.485 143.780 77.085 ;
        RECT 147.830 76.485 149.330 84.385 ;
        RECT 152.970 75.450 153.460 87.700 ;
        RECT 154.550 82.095 154.910 82.515 ;
        RECT 154.500 78.770 154.860 79.190 ;
        RECT 154.425 77.850 154.785 78.270 ;
        RECT 155.465 77.450 155.765 79.180 ;
        RECT 154.505 75.550 154.865 75.970 ;
        RECT 156.300 75.450 156.790 95.450 ;
        RECT 157.325 90.790 157.625 97.450 ;
        RECT 158.205 92.825 158.505 96.450 ;
        RECT 158.960 92.155 159.260 101.450 ;
        RECT 160.820 100.850 161.320 115.400 ;
        RECT 161.770 106.400 162.370 106.900 ;
        RECT 161.820 102.450 162.320 106.400 ;
        RECT 161.815 101.900 162.320 102.450 ;
        RECT 161.815 101.850 162.315 101.900 ;
        RECT 161.230 99.850 161.740 100.450 ;
        RECT 163.690 99.850 164.200 100.450 ;
        RECT 158.960 91.655 159.360 92.155 ;
        RECT 158.195 90.780 158.555 91.200 ;
        RECT 158.175 83.115 158.535 83.535 ;
        RECT 157.325 77.450 157.625 79.180 ;
        RECT 158.260 78.780 158.560 79.180 ;
        RECT 158.315 77.850 158.675 78.270 ;
        RECT 159.010 77.860 159.310 82.505 ;
        RECT 158.310 76.950 158.670 77.370 ;
        RECT 158.340 75.560 158.640 76.950 ;
        RECT 159.630 76.890 160.120 94.450 ;
        RECT 160.820 77.535 161.200 94.450 ;
        RECT 161.400 92.345 161.570 99.850 ;
        RECT 161.820 93.395 162.280 93.445 ;
        RECT 161.800 92.505 162.300 93.395 ;
        RECT 162.530 92.345 162.700 93.395 ;
        RECT 161.400 91.845 161.770 92.345 ;
        RECT 162.330 91.845 162.700 92.345 ;
        RECT 161.400 91.295 161.570 91.845 ;
        RECT 161.820 91.455 162.280 91.685 ;
        RECT 162.530 91.295 162.700 91.845 ;
        RECT 161.400 90.795 161.770 91.295 ;
        RECT 162.330 90.795 162.700 91.295 ;
        RECT 161.400 90.245 161.570 90.795 ;
        RECT 161.820 90.405 162.280 90.635 ;
        RECT 162.530 90.245 162.700 90.795 ;
        RECT 161.400 89.745 161.770 90.245 ;
        RECT 162.330 89.745 162.700 90.245 ;
        RECT 161.400 89.195 161.570 89.745 ;
        RECT 161.820 89.355 162.280 89.585 ;
        RECT 162.530 89.195 162.700 89.745 ;
        RECT 161.400 88.695 161.770 89.195 ;
        RECT 162.330 88.695 162.700 89.195 ;
        RECT 161.400 87.730 161.570 88.695 ;
        RECT 161.820 88.305 162.280 88.535 ;
        RECT 162.530 87.730 162.700 88.695 ;
        RECT 161.400 87.560 162.700 87.730 ;
        RECT 161.400 86.550 161.570 87.560 ;
        RECT 161.820 86.755 162.280 86.985 ;
        RECT 162.530 86.550 162.700 87.560 ;
        RECT 161.400 85.050 161.770 86.550 ;
        RECT 162.330 85.050 162.700 86.550 ;
        RECT 161.400 84.410 161.570 85.050 ;
        RECT 161.820 84.615 162.280 84.845 ;
        RECT 162.530 84.410 162.700 85.050 ;
        RECT 161.400 82.910 161.770 84.410 ;
        RECT 162.330 82.910 162.700 84.410 ;
        RECT 161.400 82.270 161.570 82.910 ;
        RECT 161.820 82.475 162.280 82.705 ;
        RECT 162.530 82.270 162.700 82.910 ;
        RECT 161.400 80.770 161.770 82.270 ;
        RECT 162.330 80.770 162.700 82.270 ;
        RECT 161.400 80.130 161.570 80.770 ;
        RECT 161.820 80.335 162.280 80.565 ;
        RECT 162.530 80.130 162.700 80.770 ;
        RECT 161.400 78.630 161.770 80.130 ;
        RECT 162.330 78.630 162.700 80.130 ;
        RECT 161.800 77.535 162.300 78.425 ;
        RECT 162.530 77.535 162.700 78.630 ;
        RECT 162.900 77.535 163.660 95.450 ;
        RECT 163.860 92.300 164.030 99.850 ;
        RECT 164.280 93.395 164.740 99.450 ;
        RECT 164.260 92.505 164.760 93.395 ;
        RECT 163.860 90.800 164.230 92.300 ;
        RECT 164.790 90.800 165.160 92.300 ;
        RECT 163.860 90.160 164.030 90.800 ;
        RECT 164.280 90.365 164.740 90.595 ;
        RECT 164.990 90.160 165.160 90.800 ;
        RECT 163.860 88.660 164.230 90.160 ;
        RECT 164.790 88.660 165.160 90.160 ;
        RECT 163.860 88.020 164.030 88.660 ;
        RECT 164.280 88.225 164.740 88.455 ;
        RECT 164.990 88.020 165.160 88.660 ;
        RECT 163.860 86.520 164.230 88.020 ;
        RECT 164.790 86.520 165.160 88.020 ;
        RECT 163.860 85.880 164.030 86.520 ;
        RECT 164.280 86.085 164.740 86.315 ;
        RECT 164.990 85.880 165.160 86.520 ;
        RECT 163.860 84.380 164.230 85.880 ;
        RECT 164.790 84.380 165.160 85.880 ;
        RECT 163.860 82.235 164.030 84.380 ;
        RECT 164.280 83.945 164.740 84.175 ;
        RECT 164.280 82.395 164.740 82.625 ;
        RECT 164.990 82.235 165.160 84.380 ;
        RECT 163.860 81.735 164.230 82.235 ;
        RECT 164.790 81.735 165.160 82.235 ;
        RECT 163.860 81.185 164.030 81.735 ;
        RECT 164.280 81.345 164.740 81.575 ;
        RECT 164.990 81.185 165.160 81.735 ;
        RECT 163.860 80.685 164.230 81.185 ;
        RECT 164.790 80.685 165.160 81.185 ;
        RECT 163.860 80.135 164.030 80.685 ;
        RECT 164.280 80.295 164.740 80.525 ;
        RECT 164.990 80.135 165.160 80.685 ;
        RECT 163.860 79.635 164.230 80.135 ;
        RECT 164.790 79.635 165.160 80.135 ;
        RECT 163.860 79.085 164.030 79.635 ;
        RECT 164.280 79.245 164.740 79.475 ;
        RECT 164.990 79.085 165.160 79.635 ;
        RECT 163.860 78.585 164.230 79.085 ;
        RECT 164.790 78.585 165.160 79.085 ;
        RECT 163.860 77.535 164.030 78.585 ;
        RECT 164.260 77.535 164.760 78.425 ;
        RECT 161.820 77.485 162.280 77.535 ;
        RECT 164.280 77.485 164.740 77.535 ;
        RECT 164.990 77.085 165.160 78.585 ;
        RECT 165.360 77.540 166.120 94.450 ;
        RECT 166.740 93.400 167.200 93.445 ;
        RECT 166.320 92.350 166.490 93.400 ;
        RECT 166.720 92.510 167.220 93.400 ;
        RECT 167.450 92.350 167.620 93.400 ;
        RECT 166.320 91.850 166.690 92.350 ;
        RECT 167.250 91.850 167.620 92.350 ;
        RECT 166.320 91.300 166.490 91.850 ;
        RECT 166.740 91.460 167.200 91.690 ;
        RECT 167.450 91.300 167.620 91.850 ;
        RECT 166.320 90.800 166.690 91.300 ;
        RECT 167.250 90.800 167.620 91.300 ;
        RECT 166.320 90.250 166.490 90.800 ;
        RECT 166.740 90.410 167.200 90.640 ;
        RECT 167.450 90.250 167.620 90.800 ;
        RECT 166.320 89.750 166.690 90.250 ;
        RECT 167.250 89.750 167.620 90.250 ;
        RECT 166.320 89.200 166.490 89.750 ;
        RECT 166.740 89.360 167.200 89.590 ;
        RECT 167.450 89.200 167.620 89.750 ;
        RECT 166.320 88.700 166.690 89.200 ;
        RECT 167.250 88.700 167.620 89.200 ;
        RECT 166.320 87.735 166.490 88.700 ;
        RECT 166.740 88.310 167.200 88.540 ;
        RECT 167.450 87.735 167.620 88.700 ;
        RECT 166.320 87.565 167.620 87.735 ;
        RECT 166.320 86.555 166.490 87.565 ;
        RECT 166.740 86.760 167.200 86.990 ;
        RECT 167.450 86.555 167.620 87.565 ;
        RECT 166.320 85.055 166.690 86.555 ;
        RECT 167.250 85.055 167.620 86.555 ;
        RECT 166.320 84.415 166.490 85.055 ;
        RECT 166.740 84.620 167.200 84.850 ;
        RECT 167.450 84.415 167.620 85.055 ;
        RECT 166.320 82.915 166.690 84.415 ;
        RECT 167.250 82.915 167.620 84.415 ;
        RECT 166.320 82.275 166.490 82.915 ;
        RECT 166.740 82.480 167.200 82.710 ;
        RECT 167.450 82.275 167.620 82.915 ;
        RECT 166.320 80.775 166.690 82.275 ;
        RECT 167.250 80.775 167.620 82.275 ;
        RECT 166.320 80.135 166.490 80.775 ;
        RECT 166.740 80.340 167.200 80.570 ;
        RECT 167.450 80.135 167.620 80.775 ;
        RECT 166.320 78.635 166.690 80.135 ;
        RECT 167.250 78.635 167.620 80.135 ;
        RECT 166.720 77.540 167.220 78.430 ;
        RECT 165.360 77.535 165.740 77.540 ;
        RECT 166.740 77.485 167.200 77.540 ;
        RECT 167.450 77.085 167.620 78.635 ;
        RECT 167.820 92.305 168.580 134.995 ;
        RECT 171.840 134.950 173.540 134.995 ;
        RECT 174.100 134.950 175.470 135.450 ;
        RECT 176.030 134.950 177.470 135.450 ;
        RECT 169.200 134.785 169.660 134.790 ;
        RECT 169.180 124.850 169.680 134.785 ;
        RECT 171.110 129.850 171.610 134.790 ;
        RECT 171.840 133.900 173.335 134.950 ;
        RECT 173.570 130.850 174.070 134.790 ;
        RECT 175.500 134.200 176.000 134.790 ;
        RECT 169.180 92.515 169.680 102.450 ;
        RECT 169.200 92.510 169.660 92.515 ;
        RECT 171.110 92.510 171.610 97.450 ;
        RECT 171.840 92.350 173.335 93.400 ;
        RECT 173.570 92.510 174.070 96.450 ;
        RECT 175.500 92.510 176.000 93.100 ;
        RECT 176.600 92.350 177.470 134.950 ;
        RECT 177.820 127.850 178.120 136.510 ;
        RECT 178.545 136.100 178.905 136.520 ;
        RECT 178.595 128.850 178.895 134.475 ;
        RECT 180.310 131.850 180.800 151.850 ;
        RECT 182.350 150.350 182.650 151.740 ;
        RECT 182.320 149.930 182.680 150.350 ;
        RECT 181.335 148.120 181.635 149.850 ;
        RECT 182.325 149.030 182.685 149.450 ;
        RECT 182.270 148.120 182.570 148.520 ;
        RECT 183.020 144.795 183.320 149.440 ;
        RECT 182.185 143.765 182.545 144.185 ;
        RECT 181.335 129.850 181.635 136.510 ;
        RECT 182.205 136.100 182.565 136.520 ;
        RECT 182.970 135.145 183.370 135.645 ;
        RECT 182.215 130.850 182.515 134.475 ;
        RECT 182.970 125.850 183.270 135.145 ;
        RECT 183.640 132.850 184.130 150.410 ;
        RECT 188.830 150.215 189.340 150.815 ;
        RECT 191.290 150.215 191.800 150.815 ;
        RECT 185.830 149.765 186.290 149.815 ;
        RECT 188.290 149.765 188.750 149.815 ;
        RECT 184.830 132.850 185.210 149.765 ;
        RECT 185.810 148.875 186.310 149.765 ;
        RECT 186.540 148.670 186.710 149.765 ;
        RECT 185.410 147.170 185.780 148.670 ;
        RECT 186.340 147.170 186.710 148.670 ;
        RECT 185.410 146.530 185.580 147.170 ;
        RECT 185.830 146.735 186.290 146.965 ;
        RECT 186.540 146.530 186.710 147.170 ;
        RECT 185.410 145.030 185.780 146.530 ;
        RECT 186.340 145.030 186.710 146.530 ;
        RECT 185.410 144.390 185.580 145.030 ;
        RECT 185.830 144.595 186.290 144.825 ;
        RECT 186.540 144.390 186.710 145.030 ;
        RECT 185.410 142.890 185.780 144.390 ;
        RECT 186.340 142.890 186.710 144.390 ;
        RECT 185.410 142.250 185.580 142.890 ;
        RECT 185.830 142.455 186.290 142.685 ;
        RECT 186.540 142.250 186.710 142.890 ;
        RECT 185.410 140.750 185.780 142.250 ;
        RECT 186.340 140.750 186.710 142.250 ;
        RECT 185.410 139.740 185.580 140.750 ;
        RECT 185.830 140.315 186.290 140.545 ;
        RECT 186.540 139.740 186.710 140.750 ;
        RECT 185.410 139.570 186.710 139.740 ;
        RECT 185.410 138.605 185.580 139.570 ;
        RECT 185.830 138.765 186.290 138.995 ;
        RECT 186.540 138.605 186.710 139.570 ;
        RECT 185.410 138.105 185.780 138.605 ;
        RECT 186.340 138.105 186.710 138.605 ;
        RECT 185.410 137.555 185.580 138.105 ;
        RECT 185.830 137.715 186.290 137.945 ;
        RECT 186.540 137.555 186.710 138.105 ;
        RECT 185.410 137.055 185.780 137.555 ;
        RECT 186.340 137.055 186.710 137.555 ;
        RECT 185.410 136.505 185.580 137.055 ;
        RECT 185.830 136.665 186.290 136.895 ;
        RECT 186.540 136.505 186.710 137.055 ;
        RECT 185.410 136.005 185.780 136.505 ;
        RECT 186.340 136.005 186.710 136.505 ;
        RECT 185.410 135.455 185.580 136.005 ;
        RECT 185.830 135.615 186.290 135.845 ;
        RECT 186.540 135.455 186.710 136.005 ;
        RECT 185.410 134.955 185.780 135.455 ;
        RECT 186.340 134.955 186.710 135.455 ;
        RECT 185.410 127.450 185.580 134.955 ;
        RECT 185.810 133.905 186.310 134.795 ;
        RECT 186.540 133.905 186.710 134.955 ;
        RECT 185.830 133.855 186.290 133.905 ;
        RECT 186.910 131.850 187.670 149.765 ;
        RECT 187.870 148.715 188.040 149.765 ;
        RECT 188.270 148.875 188.770 149.765 ;
        RECT 189.000 148.715 189.170 150.215 ;
        RECT 187.870 148.215 188.240 148.715 ;
        RECT 188.800 148.215 189.170 148.715 ;
        RECT 187.870 147.665 188.040 148.215 ;
        RECT 188.290 147.825 188.750 148.055 ;
        RECT 189.000 147.665 189.170 148.215 ;
        RECT 187.870 147.165 188.240 147.665 ;
        RECT 188.800 147.165 189.170 147.665 ;
        RECT 187.870 146.615 188.040 147.165 ;
        RECT 188.290 146.775 188.750 147.005 ;
        RECT 189.000 146.615 189.170 147.165 ;
        RECT 187.870 146.115 188.240 146.615 ;
        RECT 188.800 146.115 189.170 146.615 ;
        RECT 187.870 145.565 188.040 146.115 ;
        RECT 188.290 145.725 188.750 145.955 ;
        RECT 189.000 145.565 189.170 146.115 ;
        RECT 187.870 145.065 188.240 145.565 ;
        RECT 188.800 145.065 189.170 145.565 ;
        RECT 187.870 142.920 188.040 145.065 ;
        RECT 188.290 144.675 188.750 144.905 ;
        RECT 188.290 143.125 188.750 143.355 ;
        RECT 189.000 142.920 189.170 145.065 ;
        RECT 187.870 141.420 188.240 142.920 ;
        RECT 188.800 141.420 189.170 142.920 ;
        RECT 187.870 140.780 188.040 141.420 ;
        RECT 188.290 140.985 188.750 141.215 ;
        RECT 189.000 140.780 189.170 141.420 ;
        RECT 187.870 139.280 188.240 140.780 ;
        RECT 188.800 139.280 189.170 140.780 ;
        RECT 187.870 138.640 188.040 139.280 ;
        RECT 188.290 138.845 188.750 139.075 ;
        RECT 189.000 138.640 189.170 139.280 ;
        RECT 187.870 137.140 188.240 138.640 ;
        RECT 188.800 137.140 189.170 138.640 ;
        RECT 187.870 136.500 188.040 137.140 ;
        RECT 188.290 136.705 188.750 136.935 ;
        RECT 189.000 136.500 189.170 137.140 ;
        RECT 187.870 135.000 188.240 136.500 ;
        RECT 188.800 135.000 189.170 136.500 ;
        RECT 189.370 149.760 189.750 149.765 ;
        RECT 190.750 149.760 191.210 149.815 ;
        RECT 187.870 127.450 188.040 135.000 ;
        RECT 188.270 133.905 188.770 134.795 ;
        RECT 188.290 127.850 188.750 133.905 ;
        RECT 189.370 132.850 190.130 149.760 ;
        RECT 190.730 148.870 191.230 149.760 ;
        RECT 191.460 148.665 191.630 150.215 ;
        RECT 190.330 147.165 190.700 148.665 ;
        RECT 191.260 147.165 191.630 148.665 ;
        RECT 190.330 146.525 190.500 147.165 ;
        RECT 190.750 146.730 191.210 146.960 ;
        RECT 191.460 146.525 191.630 147.165 ;
        RECT 190.330 145.025 190.700 146.525 ;
        RECT 191.260 145.025 191.630 146.525 ;
        RECT 190.330 144.385 190.500 145.025 ;
        RECT 190.750 144.590 191.210 144.820 ;
        RECT 191.460 144.385 191.630 145.025 ;
        RECT 190.330 142.885 190.700 144.385 ;
        RECT 191.260 142.885 191.630 144.385 ;
        RECT 190.330 142.245 190.500 142.885 ;
        RECT 190.750 142.450 191.210 142.680 ;
        RECT 191.460 142.245 191.630 142.885 ;
        RECT 190.330 140.745 190.700 142.245 ;
        RECT 191.260 140.745 191.630 142.245 ;
        RECT 190.330 139.735 190.500 140.745 ;
        RECT 190.750 140.310 191.210 140.540 ;
        RECT 191.460 139.735 191.630 140.745 ;
        RECT 190.330 139.565 191.630 139.735 ;
        RECT 190.330 138.600 190.500 139.565 ;
        RECT 190.750 138.760 191.210 138.990 ;
        RECT 191.460 138.600 191.630 139.565 ;
        RECT 190.330 138.100 190.700 138.600 ;
        RECT 191.260 138.100 191.630 138.600 ;
        RECT 190.330 137.550 190.500 138.100 ;
        RECT 190.750 137.710 191.210 137.940 ;
        RECT 191.460 137.550 191.630 138.100 ;
        RECT 190.330 137.050 190.700 137.550 ;
        RECT 191.260 137.050 191.630 137.550 ;
        RECT 190.330 136.500 190.500 137.050 ;
        RECT 190.750 136.660 191.210 136.890 ;
        RECT 191.460 136.500 191.630 137.050 ;
        RECT 190.330 136.000 190.700 136.500 ;
        RECT 191.260 136.000 191.630 136.500 ;
        RECT 190.330 135.450 190.500 136.000 ;
        RECT 190.750 135.610 191.210 135.840 ;
        RECT 191.460 135.450 191.630 136.000 ;
        RECT 190.330 134.950 190.700 135.450 ;
        RECT 191.260 134.950 191.630 135.450 ;
        RECT 190.330 133.900 190.500 134.950 ;
        RECT 190.730 133.900 191.230 134.790 ;
        RECT 191.460 133.900 191.630 134.950 ;
        RECT 191.830 144.010 192.210 149.760 ;
        RECT 191.830 142.915 192.590 144.010 ;
        RECT 193.210 143.120 193.670 143.350 ;
        RECT 195.140 143.120 195.600 143.350 ;
        RECT 195.850 142.915 197.350 150.815 ;
        RECT 191.830 141.415 193.160 142.915 ;
        RECT 193.720 141.415 195.090 142.915 ;
        RECT 195.650 141.855 197.350 142.915 ;
        RECT 195.650 141.415 197.400 141.855 ;
        RECT 191.830 140.775 192.960 141.415 ;
        RECT 193.210 140.980 193.670 141.210 ;
        RECT 193.920 140.775 194.890 141.415 ;
        RECT 195.140 140.980 195.600 141.210 ;
        RECT 195.850 140.775 197.400 141.415 ;
        RECT 191.830 139.275 193.160 140.775 ;
        RECT 193.720 139.275 195.090 140.775 ;
        RECT 195.650 139.275 197.400 140.775 ;
        RECT 200.990 139.600 201.480 151.850 ;
        RECT 202.525 151.330 202.885 151.750 ;
        RECT 202.445 149.030 202.805 149.450 ;
        RECT 202.520 148.110 202.880 148.530 ;
        RECT 203.485 148.120 203.785 149.850 ;
        RECT 202.570 144.785 202.930 145.205 ;
        RECT 191.830 138.635 192.960 139.275 ;
        RECT 193.210 138.840 193.670 139.070 ;
        RECT 193.920 138.635 194.890 139.275 ;
        RECT 195.140 138.840 195.600 139.070 ;
        RECT 195.850 138.635 197.400 139.275 ;
        RECT 197.600 138.760 198.060 138.990 ;
        RECT 199.530 138.760 199.990 138.990 ;
        RECT 191.830 137.135 193.160 138.635 ;
        RECT 193.720 137.135 195.090 138.635 ;
        RECT 195.650 138.600 197.400 138.635 ;
        RECT 200.610 138.600 201.480 139.600 ;
        RECT 195.650 138.100 197.550 138.600 ;
        RECT 198.110 138.100 199.480 138.600 ;
        RECT 200.040 138.100 201.480 138.600 ;
        RECT 195.650 137.550 197.400 138.100 ;
        RECT 197.600 137.710 198.060 137.940 ;
        RECT 198.310 137.550 199.280 138.100 ;
        RECT 199.530 137.710 199.990 137.940 ;
        RECT 200.240 137.550 201.480 138.100 ;
        RECT 195.650 137.135 197.550 137.550 ;
        RECT 191.830 136.495 192.960 137.135 ;
        RECT 193.210 136.700 193.670 136.930 ;
        RECT 193.920 136.495 194.890 137.135 ;
        RECT 195.850 137.050 197.550 137.135 ;
        RECT 198.110 137.050 199.480 137.550 ;
        RECT 200.040 137.050 201.480 137.550 ;
        RECT 195.140 136.700 195.600 136.930 ;
        RECT 195.850 136.500 197.400 137.050 ;
        RECT 197.600 136.660 198.060 136.890 ;
        RECT 198.310 136.500 199.280 137.050 ;
        RECT 199.530 136.660 199.990 136.890 ;
        RECT 200.240 136.500 201.480 137.050 ;
        RECT 195.850 136.495 197.550 136.500 ;
        RECT 191.830 134.995 193.160 136.495 ;
        RECT 193.720 134.995 195.090 136.495 ;
        RECT 195.650 136.000 197.550 136.495 ;
        RECT 198.110 136.000 199.480 136.500 ;
        RECT 200.040 136.000 201.480 136.500 ;
        RECT 195.650 135.450 197.400 136.000 ;
        RECT 197.600 135.610 198.060 135.840 ;
        RECT 198.310 135.450 199.280 136.000 ;
        RECT 199.530 135.610 199.990 135.840 ;
        RECT 200.240 135.450 201.480 136.000 ;
        RECT 195.650 134.995 197.550 135.450 ;
        RECT 190.750 133.855 191.210 133.900 ;
        RECT 185.240 126.850 185.750 127.450 ;
        RECT 187.700 126.850 188.210 127.450 ;
        RECT 184.830 114.900 185.330 126.450 ;
        RECT 185.830 123.900 186.330 125.450 ;
        RECT 185.780 123.400 186.380 123.900 ;
        RECT 184.780 114.400 185.380 114.900 ;
        RECT 171.840 92.305 173.540 92.350 ;
        RECT 167.820 90.805 169.150 92.305 ;
        RECT 169.710 90.805 171.080 92.305 ;
        RECT 171.640 91.850 173.540 92.305 ;
        RECT 174.100 91.850 175.470 92.350 ;
        RECT 176.030 91.850 177.470 92.350 ;
        RECT 171.640 91.300 173.335 91.850 ;
        RECT 173.590 91.460 174.050 91.690 ;
        RECT 174.300 91.300 175.270 91.850 ;
        RECT 175.520 91.460 175.980 91.690 ;
        RECT 176.230 91.300 177.470 91.850 ;
        RECT 171.640 90.805 173.540 91.300 ;
        RECT 167.820 90.165 168.950 90.805 ;
        RECT 169.200 90.370 169.660 90.600 ;
        RECT 169.910 90.165 170.880 90.805 ;
        RECT 171.840 90.800 173.540 90.805 ;
        RECT 174.100 90.800 175.470 91.300 ;
        RECT 176.030 90.800 177.470 91.300 ;
        RECT 171.130 90.370 171.590 90.600 ;
        RECT 171.840 90.250 173.335 90.800 ;
        RECT 173.590 90.410 174.050 90.640 ;
        RECT 174.300 90.250 175.270 90.800 ;
        RECT 175.520 90.410 175.980 90.640 ;
        RECT 176.230 90.250 177.470 90.800 ;
        RECT 177.820 90.790 178.120 99.450 ;
        RECT 178.595 92.825 178.895 98.450 ;
        RECT 178.545 90.780 178.905 91.200 ;
        RECT 171.840 90.165 173.540 90.250 ;
        RECT 167.820 88.665 169.150 90.165 ;
        RECT 169.710 88.665 171.080 90.165 ;
        RECT 171.640 89.750 173.540 90.165 ;
        RECT 174.100 89.750 175.470 90.250 ;
        RECT 176.030 89.750 177.470 90.250 ;
        RECT 171.640 89.200 173.335 89.750 ;
        RECT 173.590 89.360 174.050 89.590 ;
        RECT 174.300 89.200 175.270 89.750 ;
        RECT 175.520 89.360 175.980 89.590 ;
        RECT 176.230 89.200 177.470 89.750 ;
        RECT 171.640 88.700 173.540 89.200 ;
        RECT 174.100 88.700 175.470 89.200 ;
        RECT 176.030 88.700 177.470 89.200 ;
        RECT 171.640 88.665 173.335 88.700 ;
        RECT 167.820 88.025 168.950 88.665 ;
        RECT 169.200 88.230 169.660 88.460 ;
        RECT 169.910 88.025 170.880 88.665 ;
        RECT 171.130 88.230 171.590 88.460 ;
        RECT 171.840 88.025 173.335 88.665 ;
        RECT 173.590 88.310 174.050 88.540 ;
        RECT 175.520 88.310 175.980 88.540 ;
        RECT 167.820 86.525 169.150 88.025 ;
        RECT 169.710 86.525 171.080 88.025 ;
        RECT 171.640 86.525 173.335 88.025 ;
        RECT 176.600 87.700 177.470 88.700 ;
        RECT 167.820 85.885 168.950 86.525 ;
        RECT 169.200 86.090 169.660 86.320 ;
        RECT 169.910 85.885 170.880 86.525 ;
        RECT 171.130 86.090 171.590 86.320 ;
        RECT 171.840 85.885 173.335 86.525 ;
        RECT 167.820 84.385 169.150 85.885 ;
        RECT 169.710 84.385 171.080 85.885 ;
        RECT 171.640 85.615 173.335 85.885 ;
        RECT 171.640 84.385 173.340 85.615 ;
        RECT 167.820 83.290 168.580 84.385 ;
        RECT 169.200 83.950 169.660 84.180 ;
        RECT 171.130 83.950 171.590 84.180 ;
        RECT 167.820 77.540 168.200 83.290 ;
        RECT 164.820 76.485 165.330 77.085 ;
        RECT 167.280 76.485 167.790 77.085 ;
        RECT 171.840 76.485 173.340 84.385 ;
        RECT 176.980 75.450 177.470 87.700 ;
        RECT 178.560 82.095 178.920 82.515 ;
        RECT 178.510 78.770 178.870 79.190 ;
        RECT 178.435 77.850 178.795 78.270 ;
        RECT 179.475 77.450 179.775 79.180 ;
        RECT 178.515 75.550 178.875 75.970 ;
        RECT 180.310 75.450 180.800 95.450 ;
        RECT 181.335 90.790 181.635 97.450 ;
        RECT 182.215 92.825 182.515 96.450 ;
        RECT 182.970 92.155 183.270 101.450 ;
        RECT 184.830 100.850 185.330 114.400 ;
        RECT 185.780 105.400 186.380 105.900 ;
        RECT 185.830 101.850 186.330 105.400 ;
        RECT 185.240 99.850 185.750 100.450 ;
        RECT 187.700 99.850 188.210 100.450 ;
        RECT 182.970 91.655 183.370 92.155 ;
        RECT 182.205 90.780 182.565 91.200 ;
        RECT 182.185 83.115 182.545 83.535 ;
        RECT 181.335 77.450 181.635 79.180 ;
        RECT 182.270 78.780 182.570 79.180 ;
        RECT 182.325 77.850 182.685 78.270 ;
        RECT 183.020 77.860 183.320 82.505 ;
        RECT 182.320 76.950 182.680 77.370 ;
        RECT 182.350 75.560 182.650 76.950 ;
        RECT 183.640 76.890 184.130 94.450 ;
        RECT 184.830 77.535 185.210 94.450 ;
        RECT 185.410 92.345 185.580 99.850 ;
        RECT 185.830 93.395 186.290 93.445 ;
        RECT 185.810 92.505 186.310 93.395 ;
        RECT 186.540 92.345 186.710 93.395 ;
        RECT 185.410 91.845 185.780 92.345 ;
        RECT 186.340 91.845 186.710 92.345 ;
        RECT 185.410 91.295 185.580 91.845 ;
        RECT 185.830 91.455 186.290 91.685 ;
        RECT 186.540 91.295 186.710 91.845 ;
        RECT 185.410 90.795 185.780 91.295 ;
        RECT 186.340 90.795 186.710 91.295 ;
        RECT 185.410 90.245 185.580 90.795 ;
        RECT 185.830 90.405 186.290 90.635 ;
        RECT 186.540 90.245 186.710 90.795 ;
        RECT 185.410 89.745 185.780 90.245 ;
        RECT 186.340 89.745 186.710 90.245 ;
        RECT 185.410 89.195 185.580 89.745 ;
        RECT 185.830 89.355 186.290 89.585 ;
        RECT 186.540 89.195 186.710 89.745 ;
        RECT 185.410 88.695 185.780 89.195 ;
        RECT 186.340 88.695 186.710 89.195 ;
        RECT 185.410 87.730 185.580 88.695 ;
        RECT 185.830 88.305 186.290 88.535 ;
        RECT 186.540 87.730 186.710 88.695 ;
        RECT 185.410 87.560 186.710 87.730 ;
        RECT 185.410 86.550 185.580 87.560 ;
        RECT 185.830 86.755 186.290 86.985 ;
        RECT 186.540 86.550 186.710 87.560 ;
        RECT 185.410 85.050 185.780 86.550 ;
        RECT 186.340 85.050 186.710 86.550 ;
        RECT 185.410 84.410 185.580 85.050 ;
        RECT 185.830 84.615 186.290 84.845 ;
        RECT 186.540 84.410 186.710 85.050 ;
        RECT 185.410 82.910 185.780 84.410 ;
        RECT 186.340 82.910 186.710 84.410 ;
        RECT 185.410 82.270 185.580 82.910 ;
        RECT 185.830 82.475 186.290 82.705 ;
        RECT 186.540 82.270 186.710 82.910 ;
        RECT 185.410 80.770 185.780 82.270 ;
        RECT 186.340 80.770 186.710 82.270 ;
        RECT 185.410 80.130 185.580 80.770 ;
        RECT 185.830 80.335 186.290 80.565 ;
        RECT 186.540 80.130 186.710 80.770 ;
        RECT 185.410 78.630 185.780 80.130 ;
        RECT 186.340 78.630 186.710 80.130 ;
        RECT 185.810 77.535 186.310 78.425 ;
        RECT 186.540 77.535 186.710 78.630 ;
        RECT 186.910 77.535 187.670 95.450 ;
        RECT 187.870 92.300 188.040 99.850 ;
        RECT 188.290 93.395 188.750 99.450 ;
        RECT 188.270 92.505 188.770 93.395 ;
        RECT 187.870 90.800 188.240 92.300 ;
        RECT 188.800 90.800 189.170 92.300 ;
        RECT 187.870 90.160 188.040 90.800 ;
        RECT 188.290 90.365 188.750 90.595 ;
        RECT 189.000 90.160 189.170 90.800 ;
        RECT 187.870 88.660 188.240 90.160 ;
        RECT 188.800 88.660 189.170 90.160 ;
        RECT 187.870 88.020 188.040 88.660 ;
        RECT 188.290 88.225 188.750 88.455 ;
        RECT 189.000 88.020 189.170 88.660 ;
        RECT 187.870 86.520 188.240 88.020 ;
        RECT 188.800 86.520 189.170 88.020 ;
        RECT 187.870 85.880 188.040 86.520 ;
        RECT 188.290 86.085 188.750 86.315 ;
        RECT 189.000 85.880 189.170 86.520 ;
        RECT 187.870 84.380 188.240 85.880 ;
        RECT 188.800 84.380 189.170 85.880 ;
        RECT 187.870 82.235 188.040 84.380 ;
        RECT 188.290 83.945 188.750 84.175 ;
        RECT 188.290 82.395 188.750 82.625 ;
        RECT 189.000 82.235 189.170 84.380 ;
        RECT 187.870 81.735 188.240 82.235 ;
        RECT 188.800 81.735 189.170 82.235 ;
        RECT 187.870 81.185 188.040 81.735 ;
        RECT 188.290 81.345 188.750 81.575 ;
        RECT 189.000 81.185 189.170 81.735 ;
        RECT 187.870 80.685 188.240 81.185 ;
        RECT 188.800 80.685 189.170 81.185 ;
        RECT 187.870 80.135 188.040 80.685 ;
        RECT 188.290 80.295 188.750 80.525 ;
        RECT 189.000 80.135 189.170 80.685 ;
        RECT 187.870 79.635 188.240 80.135 ;
        RECT 188.800 79.635 189.170 80.135 ;
        RECT 187.870 79.085 188.040 79.635 ;
        RECT 188.290 79.245 188.750 79.475 ;
        RECT 189.000 79.085 189.170 79.635 ;
        RECT 187.870 78.585 188.240 79.085 ;
        RECT 188.800 78.585 189.170 79.085 ;
        RECT 187.870 77.535 188.040 78.585 ;
        RECT 188.270 77.535 188.770 78.425 ;
        RECT 185.830 77.485 186.290 77.535 ;
        RECT 188.290 77.485 188.750 77.535 ;
        RECT 189.000 77.085 189.170 78.585 ;
        RECT 189.370 77.540 190.130 94.450 ;
        RECT 190.750 93.400 191.210 93.445 ;
        RECT 190.330 92.350 190.500 93.400 ;
        RECT 190.730 92.510 191.230 93.400 ;
        RECT 191.460 92.350 191.630 93.400 ;
        RECT 190.330 91.850 190.700 92.350 ;
        RECT 191.260 91.850 191.630 92.350 ;
        RECT 190.330 91.300 190.500 91.850 ;
        RECT 190.750 91.460 191.210 91.690 ;
        RECT 191.460 91.300 191.630 91.850 ;
        RECT 190.330 90.800 190.700 91.300 ;
        RECT 191.260 90.800 191.630 91.300 ;
        RECT 190.330 90.250 190.500 90.800 ;
        RECT 190.750 90.410 191.210 90.640 ;
        RECT 191.460 90.250 191.630 90.800 ;
        RECT 190.330 89.750 190.700 90.250 ;
        RECT 191.260 89.750 191.630 90.250 ;
        RECT 190.330 89.200 190.500 89.750 ;
        RECT 190.750 89.360 191.210 89.590 ;
        RECT 191.460 89.200 191.630 89.750 ;
        RECT 190.330 88.700 190.700 89.200 ;
        RECT 191.260 88.700 191.630 89.200 ;
        RECT 190.330 87.735 190.500 88.700 ;
        RECT 190.750 88.310 191.210 88.540 ;
        RECT 191.460 87.735 191.630 88.700 ;
        RECT 190.330 87.565 191.630 87.735 ;
        RECT 190.330 86.555 190.500 87.565 ;
        RECT 190.750 86.760 191.210 86.990 ;
        RECT 191.460 86.555 191.630 87.565 ;
        RECT 190.330 85.055 190.700 86.555 ;
        RECT 191.260 85.055 191.630 86.555 ;
        RECT 190.330 84.415 190.500 85.055 ;
        RECT 190.750 84.620 191.210 84.850 ;
        RECT 191.460 84.415 191.630 85.055 ;
        RECT 190.330 82.915 190.700 84.415 ;
        RECT 191.260 82.915 191.630 84.415 ;
        RECT 190.330 82.275 190.500 82.915 ;
        RECT 190.750 82.480 191.210 82.710 ;
        RECT 191.460 82.275 191.630 82.915 ;
        RECT 190.330 80.775 190.700 82.275 ;
        RECT 191.260 80.775 191.630 82.275 ;
        RECT 190.330 80.135 190.500 80.775 ;
        RECT 190.750 80.340 191.210 80.570 ;
        RECT 191.460 80.135 191.630 80.775 ;
        RECT 190.330 78.635 190.700 80.135 ;
        RECT 191.260 78.635 191.630 80.135 ;
        RECT 190.730 77.540 191.230 78.430 ;
        RECT 189.370 77.535 189.750 77.540 ;
        RECT 190.750 77.485 191.210 77.540 ;
        RECT 191.460 77.085 191.630 78.635 ;
        RECT 191.830 92.305 192.590 134.995 ;
        RECT 195.850 134.950 197.550 134.995 ;
        RECT 198.110 134.950 199.480 135.450 ;
        RECT 200.040 134.950 201.480 135.450 ;
        RECT 193.210 134.785 193.670 134.790 ;
        RECT 193.190 124.850 193.690 134.785 ;
        RECT 195.120 129.850 195.620 134.790 ;
        RECT 195.850 133.900 197.345 134.950 ;
        RECT 197.580 130.850 198.080 134.790 ;
        RECT 199.510 134.200 200.010 134.790 ;
        RECT 193.190 92.515 193.690 102.450 ;
        RECT 193.210 92.510 193.670 92.515 ;
        RECT 195.120 92.510 195.620 97.450 ;
        RECT 195.850 92.350 197.345 93.400 ;
        RECT 197.580 92.510 198.080 96.450 ;
        RECT 199.510 92.510 200.010 93.100 ;
        RECT 200.610 92.350 201.480 134.950 ;
        RECT 201.830 127.850 202.130 136.510 ;
        RECT 202.555 136.100 202.915 136.520 ;
        RECT 202.605 128.850 202.905 134.475 ;
        RECT 204.320 131.850 204.810 151.850 ;
        RECT 206.360 150.350 206.660 151.740 ;
        RECT 206.330 149.930 206.690 150.350 ;
        RECT 205.345 148.120 205.645 149.850 ;
        RECT 206.335 149.030 206.695 149.450 ;
        RECT 206.280 148.120 206.580 148.520 ;
        RECT 207.030 144.795 207.330 149.440 ;
        RECT 206.195 143.765 206.555 144.185 ;
        RECT 205.345 129.850 205.645 136.510 ;
        RECT 206.215 136.100 206.575 136.520 ;
        RECT 206.980 135.145 207.380 135.645 ;
        RECT 206.225 130.850 206.525 134.475 ;
        RECT 206.980 125.850 207.280 135.145 ;
        RECT 207.650 132.850 208.140 150.410 ;
        RECT 212.840 150.215 213.350 150.815 ;
        RECT 215.300 150.215 215.810 150.815 ;
        RECT 209.840 149.765 210.300 149.815 ;
        RECT 212.300 149.765 212.760 149.815 ;
        RECT 208.840 132.850 209.220 149.765 ;
        RECT 209.820 148.875 210.320 149.765 ;
        RECT 210.550 148.670 210.720 149.765 ;
        RECT 209.420 147.170 209.790 148.670 ;
        RECT 210.350 147.170 210.720 148.670 ;
        RECT 209.420 146.530 209.590 147.170 ;
        RECT 209.840 146.735 210.300 146.965 ;
        RECT 210.550 146.530 210.720 147.170 ;
        RECT 209.420 145.030 209.790 146.530 ;
        RECT 210.350 145.030 210.720 146.530 ;
        RECT 209.420 144.390 209.590 145.030 ;
        RECT 209.840 144.595 210.300 144.825 ;
        RECT 210.550 144.390 210.720 145.030 ;
        RECT 209.420 142.890 209.790 144.390 ;
        RECT 210.350 142.890 210.720 144.390 ;
        RECT 209.420 142.250 209.590 142.890 ;
        RECT 209.840 142.455 210.300 142.685 ;
        RECT 210.550 142.250 210.720 142.890 ;
        RECT 209.420 140.750 209.790 142.250 ;
        RECT 210.350 140.750 210.720 142.250 ;
        RECT 209.420 139.740 209.590 140.750 ;
        RECT 209.840 140.315 210.300 140.545 ;
        RECT 210.550 139.740 210.720 140.750 ;
        RECT 209.420 139.570 210.720 139.740 ;
        RECT 209.420 138.605 209.590 139.570 ;
        RECT 209.840 138.765 210.300 138.995 ;
        RECT 210.550 138.605 210.720 139.570 ;
        RECT 209.420 138.105 209.790 138.605 ;
        RECT 210.350 138.105 210.720 138.605 ;
        RECT 209.420 137.555 209.590 138.105 ;
        RECT 209.840 137.715 210.300 137.945 ;
        RECT 210.550 137.555 210.720 138.105 ;
        RECT 209.420 137.055 209.790 137.555 ;
        RECT 210.350 137.055 210.720 137.555 ;
        RECT 209.420 136.505 209.590 137.055 ;
        RECT 209.840 136.665 210.300 136.895 ;
        RECT 210.550 136.505 210.720 137.055 ;
        RECT 209.420 136.005 209.790 136.505 ;
        RECT 210.350 136.005 210.720 136.505 ;
        RECT 209.420 135.455 209.590 136.005 ;
        RECT 209.840 135.615 210.300 135.845 ;
        RECT 210.550 135.455 210.720 136.005 ;
        RECT 209.420 134.955 209.790 135.455 ;
        RECT 210.350 134.955 210.720 135.455 ;
        RECT 209.420 127.450 209.590 134.955 ;
        RECT 209.820 133.905 210.320 134.795 ;
        RECT 210.550 133.905 210.720 134.955 ;
        RECT 209.840 133.855 210.300 133.905 ;
        RECT 210.920 131.850 211.680 149.765 ;
        RECT 211.880 148.715 212.050 149.765 ;
        RECT 212.280 148.875 212.780 149.765 ;
        RECT 213.010 148.715 213.180 150.215 ;
        RECT 211.880 148.215 212.250 148.715 ;
        RECT 212.810 148.215 213.180 148.715 ;
        RECT 211.880 147.665 212.050 148.215 ;
        RECT 212.300 147.825 212.760 148.055 ;
        RECT 213.010 147.665 213.180 148.215 ;
        RECT 211.880 147.165 212.250 147.665 ;
        RECT 212.810 147.165 213.180 147.665 ;
        RECT 211.880 146.615 212.050 147.165 ;
        RECT 212.300 146.775 212.760 147.005 ;
        RECT 213.010 146.615 213.180 147.165 ;
        RECT 211.880 146.115 212.250 146.615 ;
        RECT 212.810 146.115 213.180 146.615 ;
        RECT 211.880 145.565 212.050 146.115 ;
        RECT 212.300 145.725 212.760 145.955 ;
        RECT 213.010 145.565 213.180 146.115 ;
        RECT 211.880 145.065 212.250 145.565 ;
        RECT 212.810 145.065 213.180 145.565 ;
        RECT 211.880 142.920 212.050 145.065 ;
        RECT 212.300 144.675 212.760 144.905 ;
        RECT 212.300 143.125 212.760 143.355 ;
        RECT 213.010 142.920 213.180 145.065 ;
        RECT 211.880 141.420 212.250 142.920 ;
        RECT 212.810 141.420 213.180 142.920 ;
        RECT 211.880 140.780 212.050 141.420 ;
        RECT 212.300 140.985 212.760 141.215 ;
        RECT 213.010 140.780 213.180 141.420 ;
        RECT 211.880 139.280 212.250 140.780 ;
        RECT 212.810 139.280 213.180 140.780 ;
        RECT 211.880 138.640 212.050 139.280 ;
        RECT 212.300 138.845 212.760 139.075 ;
        RECT 213.010 138.640 213.180 139.280 ;
        RECT 211.880 137.140 212.250 138.640 ;
        RECT 212.810 137.140 213.180 138.640 ;
        RECT 211.880 136.500 212.050 137.140 ;
        RECT 212.300 136.705 212.760 136.935 ;
        RECT 213.010 136.500 213.180 137.140 ;
        RECT 211.880 135.000 212.250 136.500 ;
        RECT 212.810 135.000 213.180 136.500 ;
        RECT 213.380 149.760 213.760 149.765 ;
        RECT 214.760 149.760 215.220 149.815 ;
        RECT 211.880 127.450 212.050 135.000 ;
        RECT 212.280 133.905 212.780 134.795 ;
        RECT 212.300 127.850 212.760 133.905 ;
        RECT 213.380 132.850 214.140 149.760 ;
        RECT 214.740 148.870 215.240 149.760 ;
        RECT 215.470 148.665 215.640 150.215 ;
        RECT 214.340 147.165 214.710 148.665 ;
        RECT 215.270 147.165 215.640 148.665 ;
        RECT 214.340 146.525 214.510 147.165 ;
        RECT 214.760 146.730 215.220 146.960 ;
        RECT 215.470 146.525 215.640 147.165 ;
        RECT 214.340 145.025 214.710 146.525 ;
        RECT 215.270 145.025 215.640 146.525 ;
        RECT 214.340 144.385 214.510 145.025 ;
        RECT 214.760 144.590 215.220 144.820 ;
        RECT 215.470 144.385 215.640 145.025 ;
        RECT 214.340 142.885 214.710 144.385 ;
        RECT 215.270 142.885 215.640 144.385 ;
        RECT 214.340 142.245 214.510 142.885 ;
        RECT 214.760 142.450 215.220 142.680 ;
        RECT 215.470 142.245 215.640 142.885 ;
        RECT 214.340 140.745 214.710 142.245 ;
        RECT 215.270 140.745 215.640 142.245 ;
        RECT 214.340 139.735 214.510 140.745 ;
        RECT 214.760 140.310 215.220 140.540 ;
        RECT 215.470 139.735 215.640 140.745 ;
        RECT 214.340 139.565 215.640 139.735 ;
        RECT 214.340 138.600 214.510 139.565 ;
        RECT 214.760 138.760 215.220 138.990 ;
        RECT 215.470 138.600 215.640 139.565 ;
        RECT 214.340 138.100 214.710 138.600 ;
        RECT 215.270 138.100 215.640 138.600 ;
        RECT 214.340 137.550 214.510 138.100 ;
        RECT 214.760 137.710 215.220 137.940 ;
        RECT 215.470 137.550 215.640 138.100 ;
        RECT 214.340 137.050 214.710 137.550 ;
        RECT 215.270 137.050 215.640 137.550 ;
        RECT 214.340 136.500 214.510 137.050 ;
        RECT 214.760 136.660 215.220 136.890 ;
        RECT 215.470 136.500 215.640 137.050 ;
        RECT 214.340 136.000 214.710 136.500 ;
        RECT 215.270 136.000 215.640 136.500 ;
        RECT 214.340 135.450 214.510 136.000 ;
        RECT 214.760 135.610 215.220 135.840 ;
        RECT 215.470 135.450 215.640 136.000 ;
        RECT 214.340 134.950 214.710 135.450 ;
        RECT 215.270 134.950 215.640 135.450 ;
        RECT 214.340 133.900 214.510 134.950 ;
        RECT 214.740 133.900 215.240 134.790 ;
        RECT 215.470 133.900 215.640 134.950 ;
        RECT 215.840 144.010 216.220 149.760 ;
        RECT 215.840 142.915 216.600 144.010 ;
        RECT 217.220 143.120 217.680 143.350 ;
        RECT 219.150 143.120 219.610 143.350 ;
        RECT 219.860 142.915 221.360 150.815 ;
        RECT 215.840 141.415 217.170 142.915 ;
        RECT 217.730 141.415 219.100 142.915 ;
        RECT 219.660 141.855 221.360 142.915 ;
        RECT 219.660 141.415 221.410 141.855 ;
        RECT 215.840 140.775 216.970 141.415 ;
        RECT 217.220 140.980 217.680 141.210 ;
        RECT 217.930 140.775 218.900 141.415 ;
        RECT 219.150 140.980 219.610 141.210 ;
        RECT 219.860 140.775 221.410 141.415 ;
        RECT 215.840 139.275 217.170 140.775 ;
        RECT 217.730 139.275 219.100 140.775 ;
        RECT 219.660 139.275 221.410 140.775 ;
        RECT 225.000 139.600 225.490 151.850 ;
        RECT 226.535 151.330 226.895 151.750 ;
        RECT 226.455 149.030 226.815 149.450 ;
        RECT 226.530 148.110 226.890 148.530 ;
        RECT 227.495 148.120 227.795 149.850 ;
        RECT 226.580 144.785 226.940 145.205 ;
        RECT 215.840 138.635 216.970 139.275 ;
        RECT 217.220 138.840 217.680 139.070 ;
        RECT 217.930 138.635 218.900 139.275 ;
        RECT 219.150 138.840 219.610 139.070 ;
        RECT 219.860 138.635 221.410 139.275 ;
        RECT 221.610 138.760 222.070 138.990 ;
        RECT 223.540 138.760 224.000 138.990 ;
        RECT 215.840 137.135 217.170 138.635 ;
        RECT 217.730 137.135 219.100 138.635 ;
        RECT 219.660 138.600 221.410 138.635 ;
        RECT 224.620 138.600 225.490 139.600 ;
        RECT 219.660 138.100 221.560 138.600 ;
        RECT 222.120 138.100 223.490 138.600 ;
        RECT 224.050 138.100 225.490 138.600 ;
        RECT 219.660 137.550 221.410 138.100 ;
        RECT 221.610 137.710 222.070 137.940 ;
        RECT 222.320 137.550 223.290 138.100 ;
        RECT 223.540 137.710 224.000 137.940 ;
        RECT 224.250 137.550 225.490 138.100 ;
        RECT 219.660 137.135 221.560 137.550 ;
        RECT 215.840 136.495 216.970 137.135 ;
        RECT 217.220 136.700 217.680 136.930 ;
        RECT 217.930 136.495 218.900 137.135 ;
        RECT 219.860 137.050 221.560 137.135 ;
        RECT 222.120 137.050 223.490 137.550 ;
        RECT 224.050 137.050 225.490 137.550 ;
        RECT 219.150 136.700 219.610 136.930 ;
        RECT 219.860 136.500 221.410 137.050 ;
        RECT 221.610 136.660 222.070 136.890 ;
        RECT 222.320 136.500 223.290 137.050 ;
        RECT 223.540 136.660 224.000 136.890 ;
        RECT 224.250 136.500 225.490 137.050 ;
        RECT 219.860 136.495 221.560 136.500 ;
        RECT 215.840 134.995 217.170 136.495 ;
        RECT 217.730 134.995 219.100 136.495 ;
        RECT 219.660 136.000 221.560 136.495 ;
        RECT 222.120 136.000 223.490 136.500 ;
        RECT 224.050 136.000 225.490 136.500 ;
        RECT 219.660 135.450 221.410 136.000 ;
        RECT 221.610 135.610 222.070 135.840 ;
        RECT 222.320 135.450 223.290 136.000 ;
        RECT 223.540 135.610 224.000 135.840 ;
        RECT 224.250 135.450 225.490 136.000 ;
        RECT 219.660 134.995 221.560 135.450 ;
        RECT 214.760 133.855 215.220 133.900 ;
        RECT 209.250 126.850 209.760 127.450 ;
        RECT 211.710 126.850 212.220 127.450 ;
        RECT 208.840 113.900 209.340 126.450 ;
        RECT 209.840 122.900 210.340 125.450 ;
        RECT 209.790 122.400 210.390 122.900 ;
        RECT 208.790 113.400 209.390 113.900 ;
        RECT 195.850 92.305 197.550 92.350 ;
        RECT 191.830 90.805 193.160 92.305 ;
        RECT 193.720 90.805 195.090 92.305 ;
        RECT 195.650 91.850 197.550 92.305 ;
        RECT 198.110 91.850 199.480 92.350 ;
        RECT 200.040 91.850 201.480 92.350 ;
        RECT 195.650 91.300 197.400 91.850 ;
        RECT 197.600 91.460 198.060 91.690 ;
        RECT 198.310 91.300 199.280 91.850 ;
        RECT 199.530 91.460 199.990 91.690 ;
        RECT 200.240 91.300 201.480 91.850 ;
        RECT 195.650 90.805 197.550 91.300 ;
        RECT 191.830 90.165 192.960 90.805 ;
        RECT 193.210 90.370 193.670 90.600 ;
        RECT 193.920 90.165 194.890 90.805 ;
        RECT 195.850 90.800 197.550 90.805 ;
        RECT 198.110 90.800 199.480 91.300 ;
        RECT 200.040 90.800 201.480 91.300 ;
        RECT 195.140 90.370 195.600 90.600 ;
        RECT 195.850 90.250 197.400 90.800 ;
        RECT 197.600 90.410 198.060 90.640 ;
        RECT 198.310 90.250 199.280 90.800 ;
        RECT 199.530 90.410 199.990 90.640 ;
        RECT 200.240 90.250 201.480 90.800 ;
        RECT 201.830 90.790 202.130 99.450 ;
        RECT 202.605 92.825 202.905 98.450 ;
        RECT 202.555 90.780 202.915 91.200 ;
        RECT 195.850 90.165 197.550 90.250 ;
        RECT 191.830 88.665 193.160 90.165 ;
        RECT 193.720 88.665 195.090 90.165 ;
        RECT 195.650 89.750 197.550 90.165 ;
        RECT 198.110 89.750 199.480 90.250 ;
        RECT 200.040 89.750 201.480 90.250 ;
        RECT 195.650 89.200 197.400 89.750 ;
        RECT 197.600 89.360 198.060 89.590 ;
        RECT 198.310 89.200 199.280 89.750 ;
        RECT 199.530 89.360 199.990 89.590 ;
        RECT 200.240 89.200 201.480 89.750 ;
        RECT 195.650 88.700 197.550 89.200 ;
        RECT 198.110 88.700 199.480 89.200 ;
        RECT 200.040 88.700 201.480 89.200 ;
        RECT 195.650 88.665 197.400 88.700 ;
        RECT 191.830 88.025 192.960 88.665 ;
        RECT 193.210 88.230 193.670 88.460 ;
        RECT 193.920 88.025 194.890 88.665 ;
        RECT 195.140 88.230 195.600 88.460 ;
        RECT 195.850 88.025 197.400 88.665 ;
        RECT 197.600 88.310 198.060 88.540 ;
        RECT 199.530 88.310 199.990 88.540 ;
        RECT 191.830 86.525 193.160 88.025 ;
        RECT 193.720 86.525 195.090 88.025 ;
        RECT 195.650 86.525 197.400 88.025 ;
        RECT 200.610 87.700 201.480 88.700 ;
        RECT 191.830 85.885 192.960 86.525 ;
        RECT 193.210 86.090 193.670 86.320 ;
        RECT 193.920 85.885 194.890 86.525 ;
        RECT 195.140 86.090 195.600 86.320 ;
        RECT 195.850 85.885 197.400 86.525 ;
        RECT 191.830 84.385 193.160 85.885 ;
        RECT 193.720 84.385 195.090 85.885 ;
        RECT 195.650 85.445 197.400 85.885 ;
        RECT 195.650 84.385 197.350 85.445 ;
        RECT 191.830 83.290 192.590 84.385 ;
        RECT 193.210 83.950 193.670 84.180 ;
        RECT 195.140 83.950 195.600 84.180 ;
        RECT 191.830 77.540 192.210 83.290 ;
        RECT 188.830 76.485 189.340 77.085 ;
        RECT 191.290 76.485 191.800 77.085 ;
        RECT 195.850 76.485 197.350 84.385 ;
        RECT 200.990 75.450 201.480 87.700 ;
        RECT 202.570 82.095 202.930 82.515 ;
        RECT 202.520 78.770 202.880 79.190 ;
        RECT 202.445 77.850 202.805 78.270 ;
        RECT 203.485 77.450 203.785 79.180 ;
        RECT 202.525 75.550 202.885 75.970 ;
        RECT 204.320 75.450 204.810 95.450 ;
        RECT 205.345 90.790 205.645 97.450 ;
        RECT 206.225 92.825 206.525 96.450 ;
        RECT 206.980 92.155 207.280 101.450 ;
        RECT 208.840 100.850 209.340 113.400 ;
        RECT 209.790 104.400 210.390 104.900 ;
        RECT 209.840 101.850 210.340 104.400 ;
        RECT 209.250 99.850 209.760 100.450 ;
        RECT 211.710 99.850 212.220 100.450 ;
        RECT 206.980 91.655 207.380 92.155 ;
        RECT 206.215 90.780 206.575 91.200 ;
        RECT 206.195 83.115 206.555 83.535 ;
        RECT 205.345 77.450 205.645 79.180 ;
        RECT 206.280 78.780 206.580 79.180 ;
        RECT 206.335 77.850 206.695 78.270 ;
        RECT 207.030 77.860 207.330 82.505 ;
        RECT 206.330 76.950 206.690 77.370 ;
        RECT 206.360 75.560 206.660 76.950 ;
        RECT 207.650 76.890 208.140 94.450 ;
        RECT 208.840 77.535 209.220 94.450 ;
        RECT 209.420 92.345 209.590 99.850 ;
        RECT 209.840 93.395 210.300 93.445 ;
        RECT 209.820 92.505 210.320 93.395 ;
        RECT 210.550 92.345 210.720 93.395 ;
        RECT 209.420 91.845 209.790 92.345 ;
        RECT 210.350 91.845 210.720 92.345 ;
        RECT 209.420 91.295 209.590 91.845 ;
        RECT 209.840 91.455 210.300 91.685 ;
        RECT 210.550 91.295 210.720 91.845 ;
        RECT 209.420 90.795 209.790 91.295 ;
        RECT 210.350 90.795 210.720 91.295 ;
        RECT 209.420 90.245 209.590 90.795 ;
        RECT 209.840 90.405 210.300 90.635 ;
        RECT 210.550 90.245 210.720 90.795 ;
        RECT 209.420 89.745 209.790 90.245 ;
        RECT 210.350 89.745 210.720 90.245 ;
        RECT 209.420 89.195 209.590 89.745 ;
        RECT 209.840 89.355 210.300 89.585 ;
        RECT 210.550 89.195 210.720 89.745 ;
        RECT 209.420 88.695 209.790 89.195 ;
        RECT 210.350 88.695 210.720 89.195 ;
        RECT 209.420 87.730 209.590 88.695 ;
        RECT 209.840 88.305 210.300 88.535 ;
        RECT 210.550 87.730 210.720 88.695 ;
        RECT 209.420 87.560 210.720 87.730 ;
        RECT 209.420 86.550 209.590 87.560 ;
        RECT 209.840 86.755 210.300 86.985 ;
        RECT 210.550 86.550 210.720 87.560 ;
        RECT 209.420 85.050 209.790 86.550 ;
        RECT 210.350 85.050 210.720 86.550 ;
        RECT 209.420 84.410 209.590 85.050 ;
        RECT 209.840 84.615 210.300 84.845 ;
        RECT 210.550 84.410 210.720 85.050 ;
        RECT 209.420 82.910 209.790 84.410 ;
        RECT 210.350 82.910 210.720 84.410 ;
        RECT 209.420 82.270 209.590 82.910 ;
        RECT 209.840 82.475 210.300 82.705 ;
        RECT 210.550 82.270 210.720 82.910 ;
        RECT 209.420 80.770 209.790 82.270 ;
        RECT 210.350 80.770 210.720 82.270 ;
        RECT 209.420 80.130 209.590 80.770 ;
        RECT 209.840 80.335 210.300 80.565 ;
        RECT 210.550 80.130 210.720 80.770 ;
        RECT 209.420 78.630 209.790 80.130 ;
        RECT 210.350 78.630 210.720 80.130 ;
        RECT 209.820 77.535 210.320 78.425 ;
        RECT 210.550 77.535 210.720 78.630 ;
        RECT 210.920 77.535 211.680 95.450 ;
        RECT 211.880 92.300 212.050 99.850 ;
        RECT 212.300 93.395 212.760 99.450 ;
        RECT 212.280 92.505 212.780 93.395 ;
        RECT 211.880 90.800 212.250 92.300 ;
        RECT 212.810 90.800 213.180 92.300 ;
        RECT 211.880 90.160 212.050 90.800 ;
        RECT 212.300 90.365 212.760 90.595 ;
        RECT 213.010 90.160 213.180 90.800 ;
        RECT 211.880 88.660 212.250 90.160 ;
        RECT 212.810 88.660 213.180 90.160 ;
        RECT 211.880 88.020 212.050 88.660 ;
        RECT 212.300 88.225 212.760 88.455 ;
        RECT 213.010 88.020 213.180 88.660 ;
        RECT 211.880 86.520 212.250 88.020 ;
        RECT 212.810 86.520 213.180 88.020 ;
        RECT 211.880 85.880 212.050 86.520 ;
        RECT 212.300 86.085 212.760 86.315 ;
        RECT 213.010 85.880 213.180 86.520 ;
        RECT 211.880 84.380 212.250 85.880 ;
        RECT 212.810 84.380 213.180 85.880 ;
        RECT 211.880 82.235 212.050 84.380 ;
        RECT 212.300 83.945 212.760 84.175 ;
        RECT 212.300 82.395 212.760 82.625 ;
        RECT 213.010 82.235 213.180 84.380 ;
        RECT 211.880 81.735 212.250 82.235 ;
        RECT 212.810 81.735 213.180 82.235 ;
        RECT 211.880 81.185 212.050 81.735 ;
        RECT 212.300 81.345 212.760 81.575 ;
        RECT 213.010 81.185 213.180 81.735 ;
        RECT 211.880 80.685 212.250 81.185 ;
        RECT 212.810 80.685 213.180 81.185 ;
        RECT 211.880 80.135 212.050 80.685 ;
        RECT 212.300 80.295 212.760 80.525 ;
        RECT 213.010 80.135 213.180 80.685 ;
        RECT 211.880 79.635 212.250 80.135 ;
        RECT 212.810 79.635 213.180 80.135 ;
        RECT 211.880 79.085 212.050 79.635 ;
        RECT 212.300 79.245 212.760 79.475 ;
        RECT 213.010 79.085 213.180 79.635 ;
        RECT 211.880 78.585 212.250 79.085 ;
        RECT 212.810 78.585 213.180 79.085 ;
        RECT 211.880 77.535 212.050 78.585 ;
        RECT 212.280 77.535 212.780 78.425 ;
        RECT 209.840 77.485 210.300 77.535 ;
        RECT 212.300 77.485 212.760 77.535 ;
        RECT 213.010 77.085 213.180 78.585 ;
        RECT 213.380 77.540 214.140 94.450 ;
        RECT 214.760 93.400 215.220 93.445 ;
        RECT 214.340 92.350 214.510 93.400 ;
        RECT 214.740 92.510 215.240 93.400 ;
        RECT 215.470 92.350 215.640 93.400 ;
        RECT 214.340 91.850 214.710 92.350 ;
        RECT 215.270 91.850 215.640 92.350 ;
        RECT 214.340 91.300 214.510 91.850 ;
        RECT 214.760 91.460 215.220 91.690 ;
        RECT 215.470 91.300 215.640 91.850 ;
        RECT 214.340 90.800 214.710 91.300 ;
        RECT 215.270 90.800 215.640 91.300 ;
        RECT 214.340 90.250 214.510 90.800 ;
        RECT 214.760 90.410 215.220 90.640 ;
        RECT 215.470 90.250 215.640 90.800 ;
        RECT 214.340 89.750 214.710 90.250 ;
        RECT 215.270 89.750 215.640 90.250 ;
        RECT 214.340 89.200 214.510 89.750 ;
        RECT 214.760 89.360 215.220 89.590 ;
        RECT 215.470 89.200 215.640 89.750 ;
        RECT 214.340 88.700 214.710 89.200 ;
        RECT 215.270 88.700 215.640 89.200 ;
        RECT 214.340 87.735 214.510 88.700 ;
        RECT 214.760 88.310 215.220 88.540 ;
        RECT 215.470 87.735 215.640 88.700 ;
        RECT 214.340 87.565 215.640 87.735 ;
        RECT 214.340 86.555 214.510 87.565 ;
        RECT 214.760 86.760 215.220 86.990 ;
        RECT 215.470 86.555 215.640 87.565 ;
        RECT 214.340 85.055 214.710 86.555 ;
        RECT 215.270 85.055 215.640 86.555 ;
        RECT 214.340 84.415 214.510 85.055 ;
        RECT 214.760 84.620 215.220 84.850 ;
        RECT 215.470 84.415 215.640 85.055 ;
        RECT 214.340 82.915 214.710 84.415 ;
        RECT 215.270 82.915 215.640 84.415 ;
        RECT 214.340 82.275 214.510 82.915 ;
        RECT 214.760 82.480 215.220 82.710 ;
        RECT 215.470 82.275 215.640 82.915 ;
        RECT 214.340 80.775 214.710 82.275 ;
        RECT 215.270 80.775 215.640 82.275 ;
        RECT 214.340 80.135 214.510 80.775 ;
        RECT 214.760 80.340 215.220 80.570 ;
        RECT 215.470 80.135 215.640 80.775 ;
        RECT 214.340 78.635 214.710 80.135 ;
        RECT 215.270 78.635 215.640 80.135 ;
        RECT 214.740 77.540 215.240 78.430 ;
        RECT 213.380 77.535 213.760 77.540 ;
        RECT 214.760 77.485 215.220 77.540 ;
        RECT 215.470 77.085 215.640 78.635 ;
        RECT 215.840 92.305 216.600 134.995 ;
        RECT 219.860 134.950 221.560 134.995 ;
        RECT 222.120 134.950 223.490 135.450 ;
        RECT 224.050 134.950 225.490 135.450 ;
        RECT 217.220 134.785 217.680 134.790 ;
        RECT 217.200 124.850 217.700 134.785 ;
        RECT 219.130 129.850 219.630 134.790 ;
        RECT 219.860 133.900 221.410 134.950 ;
        RECT 221.590 130.850 222.090 134.790 ;
        RECT 223.520 134.200 224.020 134.790 ;
        RECT 217.200 92.515 217.700 102.450 ;
        RECT 217.220 92.510 217.680 92.515 ;
        RECT 219.130 92.510 219.630 97.450 ;
        RECT 219.860 92.350 221.410 93.400 ;
        RECT 221.590 92.510 222.090 96.450 ;
        RECT 223.520 92.510 224.020 93.100 ;
        RECT 224.620 92.350 225.490 134.950 ;
        RECT 225.840 127.850 226.140 136.510 ;
        RECT 226.565 136.100 226.925 136.520 ;
        RECT 226.615 128.850 226.915 134.475 ;
        RECT 228.330 131.850 228.820 151.850 ;
        RECT 230.370 150.350 230.670 151.740 ;
        RECT 230.340 149.930 230.700 150.350 ;
        RECT 229.355 148.120 229.655 149.850 ;
        RECT 230.345 149.030 230.705 149.450 ;
        RECT 230.290 148.120 230.590 148.520 ;
        RECT 231.040 144.795 231.340 149.440 ;
        RECT 230.205 143.765 230.565 144.185 ;
        RECT 229.355 129.850 229.655 136.510 ;
        RECT 230.225 136.100 230.585 136.520 ;
        RECT 230.990 135.145 231.390 135.645 ;
        RECT 230.235 130.850 230.535 134.475 ;
        RECT 230.990 125.850 231.290 135.145 ;
        RECT 231.660 132.850 232.150 150.410 ;
        RECT 236.855 150.215 237.365 150.815 ;
        RECT 239.315 150.215 239.825 150.815 ;
        RECT 233.855 149.765 234.315 149.815 ;
        RECT 236.315 149.765 236.775 149.815 ;
        RECT 232.855 132.850 233.235 149.765 ;
        RECT 233.835 148.875 234.335 149.765 ;
        RECT 234.565 148.670 234.735 149.765 ;
        RECT 233.435 147.170 233.805 148.670 ;
        RECT 234.365 147.170 234.735 148.670 ;
        RECT 233.435 146.530 233.605 147.170 ;
        RECT 233.855 146.735 234.315 146.965 ;
        RECT 234.565 146.530 234.735 147.170 ;
        RECT 233.435 145.030 233.805 146.530 ;
        RECT 234.365 145.030 234.735 146.530 ;
        RECT 233.435 144.390 233.605 145.030 ;
        RECT 233.855 144.595 234.315 144.825 ;
        RECT 234.565 144.390 234.735 145.030 ;
        RECT 233.435 142.890 233.805 144.390 ;
        RECT 234.365 142.890 234.735 144.390 ;
        RECT 233.435 142.250 233.605 142.890 ;
        RECT 233.855 142.455 234.315 142.685 ;
        RECT 234.565 142.250 234.735 142.890 ;
        RECT 233.435 140.750 233.805 142.250 ;
        RECT 234.365 140.750 234.735 142.250 ;
        RECT 233.435 139.740 233.605 140.750 ;
        RECT 233.855 140.315 234.315 140.545 ;
        RECT 234.565 139.740 234.735 140.750 ;
        RECT 233.435 139.570 234.735 139.740 ;
        RECT 233.435 138.605 233.605 139.570 ;
        RECT 233.855 138.765 234.315 138.995 ;
        RECT 234.565 138.605 234.735 139.570 ;
        RECT 233.435 138.105 233.805 138.605 ;
        RECT 234.365 138.105 234.735 138.605 ;
        RECT 233.435 137.555 233.605 138.105 ;
        RECT 233.855 137.715 234.315 137.945 ;
        RECT 234.565 137.555 234.735 138.105 ;
        RECT 233.435 137.055 233.805 137.555 ;
        RECT 234.365 137.055 234.735 137.555 ;
        RECT 233.435 136.505 233.605 137.055 ;
        RECT 233.855 136.665 234.315 136.895 ;
        RECT 234.565 136.505 234.735 137.055 ;
        RECT 233.435 136.005 233.805 136.505 ;
        RECT 234.365 136.005 234.735 136.505 ;
        RECT 233.435 135.455 233.605 136.005 ;
        RECT 233.855 135.615 234.315 135.845 ;
        RECT 234.565 135.455 234.735 136.005 ;
        RECT 233.435 134.955 233.805 135.455 ;
        RECT 234.365 134.955 234.735 135.455 ;
        RECT 233.435 127.450 233.605 134.955 ;
        RECT 233.835 133.905 234.335 134.795 ;
        RECT 234.565 133.905 234.735 134.955 ;
        RECT 233.855 133.855 234.315 133.905 ;
        RECT 234.935 131.850 235.695 149.765 ;
        RECT 235.895 148.715 236.065 149.765 ;
        RECT 236.295 148.875 236.795 149.765 ;
        RECT 237.025 148.715 237.195 150.215 ;
        RECT 235.895 148.215 236.265 148.715 ;
        RECT 236.825 148.215 237.195 148.715 ;
        RECT 235.895 147.665 236.065 148.215 ;
        RECT 236.315 147.825 236.775 148.055 ;
        RECT 237.025 147.665 237.195 148.215 ;
        RECT 235.895 147.165 236.265 147.665 ;
        RECT 236.825 147.165 237.195 147.665 ;
        RECT 235.895 146.615 236.065 147.165 ;
        RECT 236.315 146.775 236.775 147.005 ;
        RECT 237.025 146.615 237.195 147.165 ;
        RECT 235.895 146.115 236.265 146.615 ;
        RECT 236.825 146.115 237.195 146.615 ;
        RECT 235.895 145.565 236.065 146.115 ;
        RECT 236.315 145.725 236.775 145.955 ;
        RECT 237.025 145.565 237.195 146.115 ;
        RECT 235.895 145.065 236.265 145.565 ;
        RECT 236.825 145.065 237.195 145.565 ;
        RECT 235.895 142.920 236.065 145.065 ;
        RECT 236.315 144.675 236.775 144.905 ;
        RECT 236.315 143.125 236.775 143.355 ;
        RECT 237.025 142.920 237.195 145.065 ;
        RECT 235.895 141.420 236.265 142.920 ;
        RECT 236.825 141.420 237.195 142.920 ;
        RECT 235.895 140.780 236.065 141.420 ;
        RECT 236.315 140.985 236.775 141.215 ;
        RECT 237.025 140.780 237.195 141.420 ;
        RECT 235.895 139.280 236.265 140.780 ;
        RECT 236.825 139.280 237.195 140.780 ;
        RECT 235.895 138.640 236.065 139.280 ;
        RECT 236.315 138.845 236.775 139.075 ;
        RECT 237.025 138.640 237.195 139.280 ;
        RECT 235.895 137.140 236.265 138.640 ;
        RECT 236.825 137.140 237.195 138.640 ;
        RECT 235.895 136.500 236.065 137.140 ;
        RECT 236.315 136.705 236.775 136.935 ;
        RECT 237.025 136.500 237.195 137.140 ;
        RECT 235.895 135.000 236.265 136.500 ;
        RECT 236.825 135.000 237.195 136.500 ;
        RECT 237.395 149.760 237.775 149.765 ;
        RECT 238.775 149.760 239.235 149.815 ;
        RECT 235.895 127.450 236.065 135.000 ;
        RECT 236.295 133.905 236.795 134.795 ;
        RECT 236.315 127.850 236.775 133.905 ;
        RECT 237.395 132.850 238.155 149.760 ;
        RECT 238.755 148.870 239.255 149.760 ;
        RECT 239.485 148.665 239.655 150.215 ;
        RECT 238.355 147.165 238.725 148.665 ;
        RECT 239.285 147.165 239.655 148.665 ;
        RECT 238.355 146.525 238.525 147.165 ;
        RECT 238.775 146.730 239.235 146.960 ;
        RECT 239.485 146.525 239.655 147.165 ;
        RECT 238.355 145.025 238.725 146.525 ;
        RECT 239.285 145.025 239.655 146.525 ;
        RECT 238.355 144.385 238.525 145.025 ;
        RECT 238.775 144.590 239.235 144.820 ;
        RECT 239.485 144.385 239.655 145.025 ;
        RECT 238.355 142.885 238.725 144.385 ;
        RECT 239.285 142.885 239.655 144.385 ;
        RECT 238.355 142.245 238.525 142.885 ;
        RECT 238.775 142.450 239.235 142.680 ;
        RECT 239.485 142.245 239.655 142.885 ;
        RECT 238.355 140.745 238.725 142.245 ;
        RECT 239.285 140.745 239.655 142.245 ;
        RECT 238.355 139.735 238.525 140.745 ;
        RECT 238.775 140.310 239.235 140.540 ;
        RECT 239.485 139.735 239.655 140.745 ;
        RECT 238.355 139.565 239.655 139.735 ;
        RECT 238.355 138.600 238.525 139.565 ;
        RECT 238.775 138.760 239.235 138.990 ;
        RECT 239.485 138.600 239.655 139.565 ;
        RECT 238.355 138.100 238.725 138.600 ;
        RECT 239.285 138.100 239.655 138.600 ;
        RECT 238.355 137.550 238.525 138.100 ;
        RECT 238.775 137.710 239.235 137.940 ;
        RECT 239.485 137.550 239.655 138.100 ;
        RECT 238.355 137.050 238.725 137.550 ;
        RECT 239.285 137.050 239.655 137.550 ;
        RECT 238.355 136.500 238.525 137.050 ;
        RECT 238.775 136.660 239.235 136.890 ;
        RECT 239.485 136.500 239.655 137.050 ;
        RECT 238.355 136.000 238.725 136.500 ;
        RECT 239.285 136.000 239.655 136.500 ;
        RECT 238.355 135.450 238.525 136.000 ;
        RECT 238.775 135.610 239.235 135.840 ;
        RECT 239.485 135.450 239.655 136.000 ;
        RECT 238.355 134.950 238.725 135.450 ;
        RECT 239.285 134.950 239.655 135.450 ;
        RECT 238.355 133.900 238.525 134.950 ;
        RECT 238.755 133.900 239.255 134.790 ;
        RECT 239.485 133.900 239.655 134.950 ;
        RECT 239.855 144.010 240.235 149.760 ;
        RECT 239.855 142.915 240.615 144.010 ;
        RECT 241.235 143.120 241.695 143.350 ;
        RECT 243.165 143.120 243.625 143.350 ;
        RECT 243.875 142.915 245.375 150.815 ;
        RECT 239.855 141.415 241.185 142.915 ;
        RECT 241.745 141.415 243.115 142.915 ;
        RECT 243.675 141.855 245.375 142.915 ;
        RECT 243.675 141.415 245.420 141.855 ;
        RECT 239.855 140.775 240.985 141.415 ;
        RECT 241.235 140.980 241.695 141.210 ;
        RECT 241.945 140.775 242.915 141.415 ;
        RECT 243.165 140.980 243.625 141.210 ;
        RECT 243.875 140.775 245.420 141.415 ;
        RECT 239.855 139.275 241.185 140.775 ;
        RECT 241.745 139.275 243.115 140.775 ;
        RECT 243.675 139.275 245.420 140.775 ;
        RECT 249.015 139.600 249.505 151.850 ;
        RECT 250.550 151.330 250.910 151.750 ;
        RECT 250.470 149.030 250.830 149.450 ;
        RECT 250.545 148.110 250.905 148.530 ;
        RECT 251.510 148.120 251.810 149.850 ;
        RECT 250.595 144.785 250.955 145.205 ;
        RECT 239.855 138.635 240.985 139.275 ;
        RECT 241.235 138.840 241.695 139.070 ;
        RECT 241.945 138.635 242.915 139.275 ;
        RECT 243.165 138.840 243.625 139.070 ;
        RECT 243.875 138.635 245.420 139.275 ;
        RECT 245.625 138.760 246.085 138.990 ;
        RECT 247.555 138.760 248.015 138.990 ;
        RECT 239.855 137.135 241.185 138.635 ;
        RECT 241.745 137.135 243.115 138.635 ;
        RECT 243.675 138.600 245.420 138.635 ;
        RECT 248.635 138.600 249.505 139.600 ;
        RECT 243.675 138.100 245.575 138.600 ;
        RECT 246.135 138.100 247.505 138.600 ;
        RECT 248.065 138.100 249.505 138.600 ;
        RECT 243.675 137.550 245.420 138.100 ;
        RECT 245.625 137.710 246.085 137.940 ;
        RECT 246.335 137.550 247.305 138.100 ;
        RECT 247.555 137.710 248.015 137.940 ;
        RECT 248.265 137.550 249.505 138.100 ;
        RECT 243.675 137.135 245.575 137.550 ;
        RECT 239.855 136.495 240.985 137.135 ;
        RECT 241.235 136.700 241.695 136.930 ;
        RECT 241.945 136.495 242.915 137.135 ;
        RECT 243.875 137.050 245.575 137.135 ;
        RECT 246.135 137.050 247.505 137.550 ;
        RECT 248.065 137.050 249.505 137.550 ;
        RECT 243.165 136.700 243.625 136.930 ;
        RECT 243.875 136.500 245.420 137.050 ;
        RECT 245.625 136.660 246.085 136.890 ;
        RECT 246.335 136.500 247.305 137.050 ;
        RECT 247.555 136.660 248.015 136.890 ;
        RECT 248.265 136.500 249.505 137.050 ;
        RECT 243.875 136.495 245.575 136.500 ;
        RECT 239.855 134.995 241.185 136.495 ;
        RECT 241.745 134.995 243.115 136.495 ;
        RECT 243.675 136.000 245.575 136.495 ;
        RECT 246.135 136.000 247.505 136.500 ;
        RECT 248.065 136.000 249.505 136.500 ;
        RECT 243.675 135.450 245.420 136.000 ;
        RECT 245.625 135.610 246.085 135.840 ;
        RECT 246.335 135.450 247.305 136.000 ;
        RECT 247.555 135.610 248.015 135.840 ;
        RECT 248.265 135.450 249.505 136.000 ;
        RECT 243.675 134.995 245.575 135.450 ;
        RECT 238.775 133.855 239.235 133.900 ;
        RECT 233.265 126.850 233.775 127.450 ;
        RECT 235.725 126.850 236.235 127.450 ;
        RECT 232.855 126.400 233.355 126.450 ;
        RECT 232.850 125.850 233.355 126.400 ;
        RECT 232.850 112.900 233.350 125.850 ;
        RECT 233.850 121.900 234.350 125.450 ;
        RECT 233.800 121.400 234.400 121.900 ;
        RECT 232.800 112.400 233.400 112.900 ;
        RECT 232.850 101.450 233.350 112.400 ;
        RECT 233.790 103.370 234.410 103.930 ;
        RECT 233.850 101.850 234.350 103.370 ;
        RECT 219.860 92.305 221.560 92.350 ;
        RECT 215.840 90.805 217.170 92.305 ;
        RECT 217.730 90.805 219.100 92.305 ;
        RECT 219.660 91.850 221.560 92.305 ;
        RECT 222.120 91.850 223.490 92.350 ;
        RECT 224.050 91.850 225.490 92.350 ;
        RECT 219.660 91.300 221.410 91.850 ;
        RECT 221.610 91.460 222.070 91.690 ;
        RECT 222.320 91.300 223.290 91.850 ;
        RECT 223.540 91.460 224.000 91.690 ;
        RECT 224.250 91.300 225.490 91.850 ;
        RECT 219.660 90.805 221.560 91.300 ;
        RECT 215.840 90.165 216.970 90.805 ;
        RECT 217.220 90.370 217.680 90.600 ;
        RECT 217.930 90.165 218.900 90.805 ;
        RECT 219.860 90.800 221.560 90.805 ;
        RECT 222.120 90.800 223.490 91.300 ;
        RECT 224.050 90.800 225.490 91.300 ;
        RECT 219.150 90.370 219.610 90.600 ;
        RECT 219.860 90.250 221.410 90.800 ;
        RECT 221.610 90.410 222.070 90.640 ;
        RECT 222.320 90.250 223.290 90.800 ;
        RECT 223.540 90.410 224.000 90.640 ;
        RECT 224.250 90.250 225.490 90.800 ;
        RECT 225.840 90.790 226.140 99.450 ;
        RECT 226.615 92.825 226.915 98.450 ;
        RECT 226.565 90.780 226.925 91.200 ;
        RECT 219.860 90.165 221.560 90.250 ;
        RECT 215.840 88.665 217.170 90.165 ;
        RECT 217.730 88.665 219.100 90.165 ;
        RECT 219.660 89.750 221.560 90.165 ;
        RECT 222.120 89.750 223.490 90.250 ;
        RECT 224.050 89.750 225.490 90.250 ;
        RECT 219.660 89.200 221.410 89.750 ;
        RECT 221.610 89.360 222.070 89.590 ;
        RECT 222.320 89.200 223.290 89.750 ;
        RECT 223.540 89.360 224.000 89.590 ;
        RECT 224.250 89.200 225.490 89.750 ;
        RECT 219.660 88.700 221.560 89.200 ;
        RECT 222.120 88.700 223.490 89.200 ;
        RECT 224.050 88.700 225.490 89.200 ;
        RECT 219.660 88.665 221.410 88.700 ;
        RECT 215.840 88.025 216.970 88.665 ;
        RECT 217.220 88.230 217.680 88.460 ;
        RECT 217.930 88.025 218.900 88.665 ;
        RECT 219.150 88.230 219.610 88.460 ;
        RECT 219.860 88.025 221.410 88.665 ;
        RECT 221.610 88.310 222.070 88.540 ;
        RECT 223.540 88.310 224.000 88.540 ;
        RECT 215.840 86.525 217.170 88.025 ;
        RECT 217.730 86.525 219.100 88.025 ;
        RECT 219.660 86.525 221.410 88.025 ;
        RECT 224.620 87.700 225.490 88.700 ;
        RECT 215.840 85.885 216.970 86.525 ;
        RECT 217.220 86.090 217.680 86.320 ;
        RECT 217.930 85.885 218.900 86.525 ;
        RECT 219.150 86.090 219.610 86.320 ;
        RECT 219.860 85.885 221.410 86.525 ;
        RECT 215.840 84.385 217.170 85.885 ;
        RECT 217.730 84.385 219.100 85.885 ;
        RECT 219.660 85.445 221.410 85.885 ;
        RECT 219.660 84.385 221.360 85.445 ;
        RECT 215.840 83.290 216.600 84.385 ;
        RECT 217.220 83.950 217.680 84.180 ;
        RECT 219.150 83.950 219.610 84.180 ;
        RECT 215.840 77.540 216.220 83.290 ;
        RECT 212.840 76.485 213.350 77.085 ;
        RECT 215.300 76.485 215.810 77.085 ;
        RECT 219.860 76.485 221.360 84.385 ;
        RECT 225.000 75.450 225.490 87.700 ;
        RECT 226.580 82.095 226.940 82.515 ;
        RECT 226.530 78.770 226.890 79.190 ;
        RECT 226.455 77.850 226.815 78.270 ;
        RECT 227.495 77.450 227.795 79.180 ;
        RECT 226.535 75.550 226.895 75.970 ;
        RECT 228.330 75.450 228.820 95.450 ;
        RECT 229.355 90.790 229.655 97.450 ;
        RECT 230.235 92.825 230.535 96.450 ;
        RECT 230.990 92.155 231.290 101.450 ;
        RECT 232.850 100.900 233.355 101.450 ;
        RECT 232.855 100.850 233.355 100.900 ;
        RECT 233.265 99.850 233.775 100.450 ;
        RECT 235.725 99.850 236.235 100.450 ;
        RECT 230.990 91.655 231.390 92.155 ;
        RECT 230.225 90.780 230.585 91.200 ;
        RECT 230.205 83.115 230.565 83.535 ;
        RECT 229.355 77.450 229.655 79.180 ;
        RECT 230.290 78.780 230.590 79.180 ;
        RECT 230.345 77.850 230.705 78.270 ;
        RECT 231.040 77.860 231.340 82.505 ;
        RECT 230.340 76.950 230.700 77.370 ;
        RECT 230.370 75.560 230.670 76.950 ;
        RECT 231.660 76.890 232.150 94.450 ;
        RECT 232.855 77.535 233.235 94.450 ;
        RECT 233.435 92.345 233.605 99.850 ;
        RECT 233.855 93.395 234.315 93.445 ;
        RECT 233.835 92.505 234.335 93.395 ;
        RECT 234.565 92.345 234.735 93.395 ;
        RECT 233.435 91.845 233.805 92.345 ;
        RECT 234.365 91.845 234.735 92.345 ;
        RECT 233.435 91.295 233.605 91.845 ;
        RECT 233.855 91.455 234.315 91.685 ;
        RECT 234.565 91.295 234.735 91.845 ;
        RECT 233.435 90.795 233.805 91.295 ;
        RECT 234.365 90.795 234.735 91.295 ;
        RECT 233.435 90.245 233.605 90.795 ;
        RECT 233.855 90.405 234.315 90.635 ;
        RECT 234.565 90.245 234.735 90.795 ;
        RECT 233.435 89.745 233.805 90.245 ;
        RECT 234.365 89.745 234.735 90.245 ;
        RECT 233.435 89.195 233.605 89.745 ;
        RECT 233.855 89.355 234.315 89.585 ;
        RECT 234.565 89.195 234.735 89.745 ;
        RECT 233.435 88.695 233.805 89.195 ;
        RECT 234.365 88.695 234.735 89.195 ;
        RECT 233.435 87.730 233.605 88.695 ;
        RECT 233.855 88.305 234.315 88.535 ;
        RECT 234.565 87.730 234.735 88.695 ;
        RECT 233.435 87.560 234.735 87.730 ;
        RECT 233.435 86.550 233.605 87.560 ;
        RECT 233.855 86.755 234.315 86.985 ;
        RECT 234.565 86.550 234.735 87.560 ;
        RECT 233.435 85.050 233.805 86.550 ;
        RECT 234.365 85.050 234.735 86.550 ;
        RECT 233.435 84.410 233.605 85.050 ;
        RECT 233.855 84.615 234.315 84.845 ;
        RECT 234.565 84.410 234.735 85.050 ;
        RECT 233.435 82.910 233.805 84.410 ;
        RECT 234.365 82.910 234.735 84.410 ;
        RECT 233.435 82.270 233.605 82.910 ;
        RECT 233.855 82.475 234.315 82.705 ;
        RECT 234.565 82.270 234.735 82.910 ;
        RECT 233.435 80.770 233.805 82.270 ;
        RECT 234.365 80.770 234.735 82.270 ;
        RECT 233.435 80.130 233.605 80.770 ;
        RECT 233.855 80.335 234.315 80.565 ;
        RECT 234.565 80.130 234.735 80.770 ;
        RECT 233.435 78.630 233.805 80.130 ;
        RECT 234.365 78.630 234.735 80.130 ;
        RECT 233.835 77.535 234.335 78.425 ;
        RECT 234.565 77.535 234.735 78.630 ;
        RECT 234.935 77.535 235.695 95.450 ;
        RECT 235.895 92.300 236.065 99.850 ;
        RECT 236.315 93.395 236.775 99.450 ;
        RECT 236.295 92.505 236.795 93.395 ;
        RECT 235.895 90.800 236.265 92.300 ;
        RECT 236.825 90.800 237.195 92.300 ;
        RECT 235.895 90.160 236.065 90.800 ;
        RECT 236.315 90.365 236.775 90.595 ;
        RECT 237.025 90.160 237.195 90.800 ;
        RECT 235.895 88.660 236.265 90.160 ;
        RECT 236.825 88.660 237.195 90.160 ;
        RECT 235.895 88.020 236.065 88.660 ;
        RECT 236.315 88.225 236.775 88.455 ;
        RECT 237.025 88.020 237.195 88.660 ;
        RECT 235.895 86.520 236.265 88.020 ;
        RECT 236.825 86.520 237.195 88.020 ;
        RECT 235.895 85.880 236.065 86.520 ;
        RECT 236.315 86.085 236.775 86.315 ;
        RECT 237.025 85.880 237.195 86.520 ;
        RECT 235.895 84.380 236.265 85.880 ;
        RECT 236.825 84.380 237.195 85.880 ;
        RECT 235.895 82.235 236.065 84.380 ;
        RECT 236.315 83.945 236.775 84.175 ;
        RECT 236.315 82.395 236.775 82.625 ;
        RECT 237.025 82.235 237.195 84.380 ;
        RECT 235.895 81.735 236.265 82.235 ;
        RECT 236.825 81.735 237.195 82.235 ;
        RECT 235.895 81.185 236.065 81.735 ;
        RECT 236.315 81.345 236.775 81.575 ;
        RECT 237.025 81.185 237.195 81.735 ;
        RECT 235.895 80.685 236.265 81.185 ;
        RECT 236.825 80.685 237.195 81.185 ;
        RECT 235.895 80.135 236.065 80.685 ;
        RECT 236.315 80.295 236.775 80.525 ;
        RECT 237.025 80.135 237.195 80.685 ;
        RECT 235.895 79.635 236.265 80.135 ;
        RECT 236.825 79.635 237.195 80.135 ;
        RECT 235.895 79.085 236.065 79.635 ;
        RECT 236.315 79.245 236.775 79.475 ;
        RECT 237.025 79.085 237.195 79.635 ;
        RECT 235.895 78.585 236.265 79.085 ;
        RECT 236.825 78.585 237.195 79.085 ;
        RECT 235.895 77.535 236.065 78.585 ;
        RECT 236.295 77.535 236.795 78.425 ;
        RECT 233.855 77.485 234.315 77.535 ;
        RECT 236.315 77.485 236.775 77.535 ;
        RECT 237.025 77.085 237.195 78.585 ;
        RECT 237.395 77.540 238.155 94.450 ;
        RECT 238.775 93.400 239.235 93.445 ;
        RECT 238.355 92.350 238.525 93.400 ;
        RECT 238.755 92.510 239.255 93.400 ;
        RECT 239.485 92.350 239.655 93.400 ;
        RECT 238.355 91.850 238.725 92.350 ;
        RECT 239.285 91.850 239.655 92.350 ;
        RECT 238.355 91.300 238.525 91.850 ;
        RECT 238.775 91.460 239.235 91.690 ;
        RECT 239.485 91.300 239.655 91.850 ;
        RECT 238.355 90.800 238.725 91.300 ;
        RECT 239.285 90.800 239.655 91.300 ;
        RECT 238.355 90.250 238.525 90.800 ;
        RECT 238.775 90.410 239.235 90.640 ;
        RECT 239.485 90.250 239.655 90.800 ;
        RECT 238.355 89.750 238.725 90.250 ;
        RECT 239.285 89.750 239.655 90.250 ;
        RECT 238.355 89.200 238.525 89.750 ;
        RECT 238.775 89.360 239.235 89.590 ;
        RECT 239.485 89.200 239.655 89.750 ;
        RECT 238.355 88.700 238.725 89.200 ;
        RECT 239.285 88.700 239.655 89.200 ;
        RECT 238.355 87.735 238.525 88.700 ;
        RECT 238.775 88.310 239.235 88.540 ;
        RECT 239.485 87.735 239.655 88.700 ;
        RECT 238.355 87.565 239.655 87.735 ;
        RECT 238.355 86.555 238.525 87.565 ;
        RECT 238.775 86.760 239.235 86.990 ;
        RECT 239.485 86.555 239.655 87.565 ;
        RECT 238.355 85.055 238.725 86.555 ;
        RECT 239.285 85.055 239.655 86.555 ;
        RECT 238.355 84.415 238.525 85.055 ;
        RECT 238.775 84.620 239.235 84.850 ;
        RECT 239.485 84.415 239.655 85.055 ;
        RECT 238.355 82.915 238.725 84.415 ;
        RECT 239.285 82.915 239.655 84.415 ;
        RECT 238.355 82.275 238.525 82.915 ;
        RECT 238.775 82.480 239.235 82.710 ;
        RECT 239.485 82.275 239.655 82.915 ;
        RECT 238.355 80.775 238.725 82.275 ;
        RECT 239.285 80.775 239.655 82.275 ;
        RECT 238.355 80.135 238.525 80.775 ;
        RECT 238.775 80.340 239.235 80.570 ;
        RECT 239.485 80.135 239.655 80.775 ;
        RECT 238.355 78.635 238.725 80.135 ;
        RECT 239.285 78.635 239.655 80.135 ;
        RECT 238.755 77.540 239.255 78.430 ;
        RECT 237.395 77.535 237.775 77.540 ;
        RECT 238.775 77.485 239.235 77.540 ;
        RECT 239.485 77.085 239.655 78.635 ;
        RECT 239.855 92.305 240.615 134.995 ;
        RECT 243.875 134.950 245.575 134.995 ;
        RECT 246.135 134.950 247.505 135.450 ;
        RECT 248.065 134.950 249.505 135.450 ;
        RECT 241.235 134.785 241.695 134.790 ;
        RECT 241.215 124.850 241.715 134.785 ;
        RECT 243.145 129.850 243.645 134.790 ;
        RECT 243.875 133.900 245.420 134.950 ;
        RECT 245.605 130.850 246.105 134.790 ;
        RECT 247.535 134.200 248.035 134.790 ;
        RECT 241.215 92.515 241.715 102.450 ;
        RECT 241.235 92.510 241.695 92.515 ;
        RECT 243.145 92.510 243.645 97.450 ;
        RECT 243.875 92.350 245.420 93.400 ;
        RECT 245.605 92.510 246.105 96.450 ;
        RECT 247.535 92.510 248.035 93.100 ;
        RECT 248.635 92.350 249.505 134.950 ;
        RECT 249.855 127.850 250.155 136.510 ;
        RECT 250.580 136.100 250.940 136.520 ;
        RECT 250.630 128.850 250.930 134.475 ;
        RECT 252.345 131.850 252.835 151.850 ;
        RECT 254.385 150.350 254.685 151.740 ;
        RECT 254.355 149.930 254.715 150.350 ;
        RECT 253.370 148.120 253.670 149.850 ;
        RECT 254.360 149.030 254.720 149.450 ;
        RECT 254.305 148.120 254.605 148.520 ;
        RECT 255.055 144.795 255.355 149.440 ;
        RECT 254.220 143.765 254.580 144.185 ;
        RECT 253.370 129.850 253.670 136.510 ;
        RECT 254.240 136.100 254.600 136.520 ;
        RECT 255.005 135.145 255.405 135.645 ;
        RECT 254.250 130.850 254.550 134.475 ;
        RECT 255.005 125.850 255.305 135.145 ;
        RECT 255.675 132.850 256.165 150.410 ;
        RECT 260.910 150.215 261.420 150.815 ;
        RECT 263.370 150.215 263.880 150.815 ;
        RECT 257.910 149.765 258.370 149.815 ;
        RECT 260.370 149.765 260.830 149.815 ;
        RECT 256.910 132.850 257.290 149.765 ;
        RECT 257.890 148.875 258.390 149.765 ;
        RECT 258.620 148.670 258.790 149.765 ;
        RECT 257.490 147.170 257.860 148.670 ;
        RECT 258.420 147.170 258.790 148.670 ;
        RECT 257.490 146.530 257.660 147.170 ;
        RECT 257.910 146.735 258.370 146.965 ;
        RECT 258.620 146.530 258.790 147.170 ;
        RECT 257.490 145.030 257.860 146.530 ;
        RECT 258.420 145.030 258.790 146.530 ;
        RECT 257.490 144.390 257.660 145.030 ;
        RECT 257.910 144.595 258.370 144.825 ;
        RECT 258.620 144.390 258.790 145.030 ;
        RECT 257.490 142.890 257.860 144.390 ;
        RECT 258.420 142.890 258.790 144.390 ;
        RECT 257.490 142.250 257.660 142.890 ;
        RECT 257.910 142.455 258.370 142.685 ;
        RECT 258.620 142.250 258.790 142.890 ;
        RECT 257.490 140.750 257.860 142.250 ;
        RECT 258.420 140.750 258.790 142.250 ;
        RECT 257.490 139.740 257.660 140.750 ;
        RECT 257.910 140.315 258.370 140.545 ;
        RECT 258.620 139.740 258.790 140.750 ;
        RECT 257.490 139.570 258.790 139.740 ;
        RECT 257.490 138.605 257.660 139.570 ;
        RECT 257.910 138.765 258.370 138.995 ;
        RECT 258.620 138.605 258.790 139.570 ;
        RECT 257.490 138.105 257.860 138.605 ;
        RECT 258.420 138.105 258.790 138.605 ;
        RECT 257.490 137.555 257.660 138.105 ;
        RECT 257.910 137.715 258.370 137.945 ;
        RECT 258.620 137.555 258.790 138.105 ;
        RECT 257.490 137.055 257.860 137.555 ;
        RECT 258.420 137.055 258.790 137.555 ;
        RECT 257.490 136.505 257.660 137.055 ;
        RECT 257.910 136.665 258.370 136.895 ;
        RECT 258.620 136.505 258.790 137.055 ;
        RECT 257.490 136.005 257.860 136.505 ;
        RECT 258.420 136.005 258.790 136.505 ;
        RECT 257.490 135.455 257.660 136.005 ;
        RECT 257.910 135.615 258.370 135.845 ;
        RECT 258.620 135.455 258.790 136.005 ;
        RECT 257.490 134.955 257.860 135.455 ;
        RECT 258.420 134.955 258.790 135.455 ;
        RECT 257.490 127.450 257.660 134.955 ;
        RECT 257.890 133.905 258.390 134.795 ;
        RECT 258.620 133.905 258.790 134.955 ;
        RECT 257.910 133.855 258.370 133.905 ;
        RECT 258.990 131.850 259.750 149.765 ;
        RECT 259.950 148.715 260.120 149.765 ;
        RECT 260.350 148.875 260.850 149.765 ;
        RECT 261.080 148.715 261.250 150.215 ;
        RECT 259.950 148.215 260.320 148.715 ;
        RECT 260.880 148.215 261.250 148.715 ;
        RECT 259.950 147.665 260.120 148.215 ;
        RECT 260.370 147.825 260.830 148.055 ;
        RECT 261.080 147.665 261.250 148.215 ;
        RECT 259.950 147.165 260.320 147.665 ;
        RECT 260.880 147.165 261.250 147.665 ;
        RECT 259.950 146.615 260.120 147.165 ;
        RECT 260.370 146.775 260.830 147.005 ;
        RECT 261.080 146.615 261.250 147.165 ;
        RECT 259.950 146.115 260.320 146.615 ;
        RECT 260.880 146.115 261.250 146.615 ;
        RECT 259.950 145.565 260.120 146.115 ;
        RECT 260.370 145.725 260.830 145.955 ;
        RECT 261.080 145.565 261.250 146.115 ;
        RECT 259.950 145.065 260.320 145.565 ;
        RECT 260.880 145.065 261.250 145.565 ;
        RECT 259.950 142.920 260.120 145.065 ;
        RECT 260.370 144.675 260.830 144.905 ;
        RECT 260.370 143.125 260.830 143.355 ;
        RECT 261.080 142.920 261.250 145.065 ;
        RECT 259.950 141.420 260.320 142.920 ;
        RECT 260.880 141.420 261.250 142.920 ;
        RECT 259.950 140.780 260.120 141.420 ;
        RECT 260.370 140.985 260.830 141.215 ;
        RECT 261.080 140.780 261.250 141.420 ;
        RECT 259.950 139.280 260.320 140.780 ;
        RECT 260.880 139.280 261.250 140.780 ;
        RECT 259.950 138.640 260.120 139.280 ;
        RECT 260.370 138.845 260.830 139.075 ;
        RECT 261.080 138.640 261.250 139.280 ;
        RECT 259.950 137.140 260.320 138.640 ;
        RECT 260.880 137.140 261.250 138.640 ;
        RECT 259.950 136.500 260.120 137.140 ;
        RECT 260.370 136.705 260.830 136.935 ;
        RECT 261.080 136.500 261.250 137.140 ;
        RECT 259.950 135.000 260.320 136.500 ;
        RECT 260.880 135.000 261.250 136.500 ;
        RECT 261.450 149.760 261.830 149.765 ;
        RECT 262.830 149.760 263.290 149.815 ;
        RECT 259.950 127.450 260.120 135.000 ;
        RECT 260.350 133.905 260.850 134.795 ;
        RECT 260.370 127.850 260.830 133.905 ;
        RECT 261.450 132.850 262.210 149.760 ;
        RECT 262.810 148.870 263.310 149.760 ;
        RECT 263.540 148.665 263.710 150.215 ;
        RECT 262.410 147.165 262.780 148.665 ;
        RECT 263.340 147.165 263.710 148.665 ;
        RECT 262.410 146.525 262.580 147.165 ;
        RECT 262.830 146.730 263.290 146.960 ;
        RECT 263.540 146.525 263.710 147.165 ;
        RECT 262.410 145.025 262.780 146.525 ;
        RECT 263.340 145.025 263.710 146.525 ;
        RECT 262.410 144.385 262.580 145.025 ;
        RECT 262.830 144.590 263.290 144.820 ;
        RECT 263.540 144.385 263.710 145.025 ;
        RECT 262.410 142.885 262.780 144.385 ;
        RECT 263.340 142.885 263.710 144.385 ;
        RECT 262.410 142.245 262.580 142.885 ;
        RECT 262.830 142.450 263.290 142.680 ;
        RECT 263.540 142.245 263.710 142.885 ;
        RECT 262.410 140.745 262.780 142.245 ;
        RECT 263.340 140.745 263.710 142.245 ;
        RECT 262.410 139.735 262.580 140.745 ;
        RECT 262.830 140.310 263.290 140.540 ;
        RECT 263.540 139.735 263.710 140.745 ;
        RECT 262.410 139.565 263.710 139.735 ;
        RECT 262.410 138.600 262.580 139.565 ;
        RECT 262.830 138.760 263.290 138.990 ;
        RECT 263.540 138.600 263.710 139.565 ;
        RECT 262.410 138.100 262.780 138.600 ;
        RECT 263.340 138.100 263.710 138.600 ;
        RECT 262.410 137.550 262.580 138.100 ;
        RECT 262.830 137.710 263.290 137.940 ;
        RECT 263.540 137.550 263.710 138.100 ;
        RECT 262.410 137.050 262.780 137.550 ;
        RECT 263.340 137.050 263.710 137.550 ;
        RECT 262.410 136.500 262.580 137.050 ;
        RECT 262.830 136.660 263.290 136.890 ;
        RECT 263.540 136.500 263.710 137.050 ;
        RECT 262.410 136.000 262.780 136.500 ;
        RECT 263.340 136.000 263.710 136.500 ;
        RECT 262.410 135.450 262.580 136.000 ;
        RECT 262.830 135.610 263.290 135.840 ;
        RECT 263.540 135.450 263.710 136.000 ;
        RECT 262.410 134.950 262.780 135.450 ;
        RECT 263.340 134.950 263.710 135.450 ;
        RECT 262.410 133.900 262.580 134.950 ;
        RECT 262.810 133.900 263.310 134.790 ;
        RECT 263.540 133.900 263.710 134.950 ;
        RECT 263.910 144.010 264.290 149.760 ;
        RECT 263.910 142.915 264.670 144.010 ;
        RECT 265.290 143.120 265.750 143.350 ;
        RECT 267.220 143.120 267.680 143.350 ;
        RECT 267.930 142.915 269.430 150.815 ;
        RECT 263.910 141.415 265.240 142.915 ;
        RECT 265.800 141.415 267.170 142.915 ;
        RECT 267.730 141.415 269.430 142.915 ;
        RECT 263.910 140.775 265.040 141.415 ;
        RECT 265.290 140.980 265.750 141.210 ;
        RECT 266.000 140.775 266.970 141.415 ;
        RECT 267.220 140.980 267.680 141.210 ;
        RECT 267.930 140.775 269.430 141.415 ;
        RECT 263.910 139.275 265.240 140.775 ;
        RECT 265.800 139.275 267.170 140.775 ;
        RECT 267.730 139.275 269.430 140.775 ;
        RECT 273.070 139.600 273.560 151.850 ;
        RECT 274.605 151.330 274.965 151.750 ;
        RECT 274.525 149.030 274.885 149.450 ;
        RECT 274.600 148.110 274.960 148.530 ;
        RECT 275.565 148.120 275.865 149.850 ;
        RECT 274.650 144.785 275.010 145.205 ;
        RECT 263.910 138.635 265.040 139.275 ;
        RECT 265.290 138.840 265.750 139.070 ;
        RECT 266.000 138.635 266.970 139.275 ;
        RECT 267.220 138.840 267.680 139.070 ;
        RECT 267.930 138.635 269.430 139.275 ;
        RECT 269.680 138.760 270.140 138.990 ;
        RECT 271.610 138.760 272.070 138.990 ;
        RECT 263.910 137.135 265.240 138.635 ;
        RECT 265.800 137.135 267.170 138.635 ;
        RECT 267.730 138.600 269.430 138.635 ;
        RECT 272.690 138.600 273.560 139.600 ;
        RECT 267.730 138.100 269.630 138.600 ;
        RECT 270.190 138.100 271.560 138.600 ;
        RECT 272.120 138.100 273.560 138.600 ;
        RECT 267.730 137.550 269.430 138.100 ;
        RECT 269.680 137.710 270.140 137.940 ;
        RECT 270.390 137.550 271.360 138.100 ;
        RECT 271.610 137.710 272.070 137.940 ;
        RECT 272.320 137.550 273.560 138.100 ;
        RECT 267.730 137.135 269.630 137.550 ;
        RECT 263.910 136.495 265.040 137.135 ;
        RECT 265.290 136.700 265.750 136.930 ;
        RECT 266.000 136.495 266.970 137.135 ;
        RECT 267.930 137.050 269.630 137.135 ;
        RECT 270.190 137.050 271.560 137.550 ;
        RECT 272.120 137.050 273.560 137.550 ;
        RECT 267.220 136.700 267.680 136.930 ;
        RECT 267.930 136.500 269.430 137.050 ;
        RECT 269.680 136.660 270.140 136.890 ;
        RECT 270.390 136.500 271.360 137.050 ;
        RECT 271.610 136.660 272.070 136.890 ;
        RECT 272.320 136.500 273.560 137.050 ;
        RECT 267.930 136.495 269.630 136.500 ;
        RECT 263.910 134.995 265.240 136.495 ;
        RECT 265.800 134.995 267.170 136.495 ;
        RECT 267.730 136.000 269.630 136.495 ;
        RECT 270.190 136.000 271.560 136.500 ;
        RECT 272.120 136.000 273.560 136.500 ;
        RECT 267.730 135.450 269.430 136.000 ;
        RECT 269.680 135.610 270.140 135.840 ;
        RECT 270.390 135.450 271.360 136.000 ;
        RECT 271.610 135.610 272.070 135.840 ;
        RECT 272.320 135.450 273.560 136.000 ;
        RECT 267.730 134.995 269.630 135.450 ;
        RECT 262.830 133.855 263.290 133.900 ;
        RECT 257.320 126.850 257.830 127.450 ;
        RECT 259.780 126.850 260.290 127.450 ;
        RECT 256.860 111.900 257.360 126.450 ;
        RECT 257.860 120.900 258.360 125.430 ;
        RECT 257.810 120.400 258.410 120.900 ;
        RECT 256.810 111.400 257.410 111.900 ;
        RECT 243.875 92.305 245.575 92.350 ;
        RECT 239.855 90.805 241.185 92.305 ;
        RECT 241.745 90.805 243.115 92.305 ;
        RECT 243.675 91.850 245.575 92.305 ;
        RECT 246.135 91.850 247.505 92.350 ;
        RECT 248.065 91.850 249.505 92.350 ;
        RECT 243.675 91.300 245.420 91.850 ;
        RECT 245.625 91.460 246.085 91.690 ;
        RECT 246.335 91.300 247.305 91.850 ;
        RECT 247.555 91.460 248.015 91.690 ;
        RECT 248.265 91.300 249.505 91.850 ;
        RECT 243.675 90.805 245.575 91.300 ;
        RECT 239.855 90.165 240.985 90.805 ;
        RECT 241.235 90.370 241.695 90.600 ;
        RECT 241.945 90.165 242.915 90.805 ;
        RECT 243.875 90.800 245.575 90.805 ;
        RECT 246.135 90.800 247.505 91.300 ;
        RECT 248.065 90.800 249.505 91.300 ;
        RECT 243.165 90.370 243.625 90.600 ;
        RECT 243.875 90.250 245.420 90.800 ;
        RECT 245.625 90.410 246.085 90.640 ;
        RECT 246.335 90.250 247.305 90.800 ;
        RECT 247.555 90.410 248.015 90.640 ;
        RECT 248.265 90.250 249.505 90.800 ;
        RECT 249.855 90.790 250.155 99.450 ;
        RECT 250.630 92.825 250.930 98.450 ;
        RECT 250.580 90.780 250.940 91.200 ;
        RECT 243.875 90.165 245.575 90.250 ;
        RECT 239.855 88.665 241.185 90.165 ;
        RECT 241.745 88.665 243.115 90.165 ;
        RECT 243.675 89.750 245.575 90.165 ;
        RECT 246.135 89.750 247.505 90.250 ;
        RECT 248.065 89.750 249.505 90.250 ;
        RECT 243.675 89.200 245.420 89.750 ;
        RECT 245.625 89.360 246.085 89.590 ;
        RECT 246.335 89.200 247.305 89.750 ;
        RECT 247.555 89.360 248.015 89.590 ;
        RECT 248.265 89.200 249.505 89.750 ;
        RECT 243.675 88.700 245.575 89.200 ;
        RECT 246.135 88.700 247.505 89.200 ;
        RECT 248.065 88.700 249.505 89.200 ;
        RECT 243.675 88.665 245.420 88.700 ;
        RECT 239.855 88.025 240.985 88.665 ;
        RECT 241.235 88.230 241.695 88.460 ;
        RECT 241.945 88.025 242.915 88.665 ;
        RECT 243.165 88.230 243.625 88.460 ;
        RECT 243.875 88.025 245.420 88.665 ;
        RECT 245.625 88.310 246.085 88.540 ;
        RECT 247.555 88.310 248.015 88.540 ;
        RECT 239.855 86.525 241.185 88.025 ;
        RECT 241.745 86.525 243.115 88.025 ;
        RECT 243.675 86.525 245.420 88.025 ;
        RECT 248.635 87.700 249.505 88.700 ;
        RECT 239.855 85.885 240.985 86.525 ;
        RECT 241.235 86.090 241.695 86.320 ;
        RECT 241.945 85.885 242.915 86.525 ;
        RECT 243.165 86.090 243.625 86.320 ;
        RECT 243.875 85.885 245.420 86.525 ;
        RECT 239.855 84.385 241.185 85.885 ;
        RECT 241.745 84.385 243.115 85.885 ;
        RECT 243.675 85.445 245.420 85.885 ;
        RECT 243.675 84.385 245.375 85.445 ;
        RECT 239.855 83.290 240.615 84.385 ;
        RECT 241.235 83.950 241.695 84.180 ;
        RECT 243.165 83.950 243.625 84.180 ;
        RECT 239.855 77.540 240.235 83.290 ;
        RECT 236.855 76.485 237.365 77.085 ;
        RECT 239.315 76.485 239.825 77.085 ;
        RECT 243.875 76.485 245.375 84.385 ;
        RECT 249.015 75.450 249.505 87.700 ;
        RECT 250.595 82.095 250.955 82.515 ;
        RECT 250.545 78.770 250.905 79.190 ;
        RECT 250.470 77.850 250.830 78.270 ;
        RECT 251.510 77.450 251.810 79.180 ;
        RECT 250.550 75.550 250.910 75.970 ;
        RECT 252.345 75.450 252.835 95.450 ;
        RECT 253.370 90.790 253.670 97.450 ;
        RECT 254.250 92.825 254.550 96.450 ;
        RECT 255.005 92.155 255.305 101.450 ;
        RECT 256.860 100.850 257.360 111.400 ;
        RECT 257.860 102.900 258.360 103.100 ;
        RECT 257.810 102.400 258.410 102.900 ;
        RECT 257.860 101.870 258.360 102.400 ;
        RECT 257.320 99.850 257.830 100.450 ;
        RECT 259.780 99.850 260.290 100.450 ;
        RECT 255.005 91.655 255.405 92.155 ;
        RECT 254.240 90.780 254.600 91.200 ;
        RECT 254.220 83.115 254.580 83.535 ;
        RECT 253.370 77.450 253.670 79.180 ;
        RECT 254.305 78.780 254.605 79.180 ;
        RECT 254.360 77.850 254.720 78.270 ;
        RECT 255.055 77.860 255.355 82.505 ;
        RECT 254.355 76.950 254.715 77.370 ;
        RECT 254.385 75.560 254.685 76.950 ;
        RECT 255.675 76.890 256.165 94.450 ;
        RECT 256.910 77.535 257.290 94.450 ;
        RECT 257.490 92.345 257.660 99.850 ;
        RECT 257.910 93.395 258.370 93.445 ;
        RECT 257.890 92.505 258.390 93.395 ;
        RECT 258.620 92.345 258.790 93.395 ;
        RECT 257.490 91.845 257.860 92.345 ;
        RECT 258.420 91.845 258.790 92.345 ;
        RECT 257.490 91.295 257.660 91.845 ;
        RECT 257.910 91.455 258.370 91.685 ;
        RECT 258.620 91.295 258.790 91.845 ;
        RECT 257.490 90.795 257.860 91.295 ;
        RECT 258.420 90.795 258.790 91.295 ;
        RECT 257.490 90.245 257.660 90.795 ;
        RECT 257.910 90.405 258.370 90.635 ;
        RECT 258.620 90.245 258.790 90.795 ;
        RECT 257.490 89.745 257.860 90.245 ;
        RECT 258.420 89.745 258.790 90.245 ;
        RECT 257.490 89.195 257.660 89.745 ;
        RECT 257.910 89.355 258.370 89.585 ;
        RECT 258.620 89.195 258.790 89.745 ;
        RECT 257.490 88.695 257.860 89.195 ;
        RECT 258.420 88.695 258.790 89.195 ;
        RECT 257.490 87.730 257.660 88.695 ;
        RECT 257.910 88.305 258.370 88.535 ;
        RECT 258.620 87.730 258.790 88.695 ;
        RECT 257.490 87.560 258.790 87.730 ;
        RECT 257.490 86.550 257.660 87.560 ;
        RECT 257.910 86.755 258.370 86.985 ;
        RECT 258.620 86.550 258.790 87.560 ;
        RECT 257.490 85.050 257.860 86.550 ;
        RECT 258.420 85.050 258.790 86.550 ;
        RECT 257.490 84.410 257.660 85.050 ;
        RECT 257.910 84.615 258.370 84.845 ;
        RECT 258.620 84.410 258.790 85.050 ;
        RECT 257.490 82.910 257.860 84.410 ;
        RECT 258.420 82.910 258.790 84.410 ;
        RECT 257.490 82.270 257.660 82.910 ;
        RECT 257.910 82.475 258.370 82.705 ;
        RECT 258.620 82.270 258.790 82.910 ;
        RECT 257.490 80.770 257.860 82.270 ;
        RECT 258.420 80.770 258.790 82.270 ;
        RECT 257.490 80.130 257.660 80.770 ;
        RECT 257.910 80.335 258.370 80.565 ;
        RECT 258.620 80.130 258.790 80.770 ;
        RECT 257.490 78.630 257.860 80.130 ;
        RECT 258.420 78.630 258.790 80.130 ;
        RECT 257.890 77.535 258.390 78.425 ;
        RECT 258.620 77.535 258.790 78.630 ;
        RECT 258.990 77.535 259.750 95.450 ;
        RECT 259.950 92.300 260.120 99.850 ;
        RECT 260.370 93.395 260.830 99.450 ;
        RECT 260.350 92.505 260.850 93.395 ;
        RECT 259.950 90.800 260.320 92.300 ;
        RECT 260.880 90.800 261.250 92.300 ;
        RECT 259.950 90.160 260.120 90.800 ;
        RECT 260.370 90.365 260.830 90.595 ;
        RECT 261.080 90.160 261.250 90.800 ;
        RECT 259.950 88.660 260.320 90.160 ;
        RECT 260.880 88.660 261.250 90.160 ;
        RECT 259.950 88.020 260.120 88.660 ;
        RECT 260.370 88.225 260.830 88.455 ;
        RECT 261.080 88.020 261.250 88.660 ;
        RECT 259.950 86.520 260.320 88.020 ;
        RECT 260.880 86.520 261.250 88.020 ;
        RECT 259.950 85.880 260.120 86.520 ;
        RECT 260.370 86.085 260.830 86.315 ;
        RECT 261.080 85.880 261.250 86.520 ;
        RECT 259.950 84.380 260.320 85.880 ;
        RECT 260.880 84.380 261.250 85.880 ;
        RECT 259.950 82.235 260.120 84.380 ;
        RECT 260.370 83.945 260.830 84.175 ;
        RECT 260.370 82.395 260.830 82.625 ;
        RECT 261.080 82.235 261.250 84.380 ;
        RECT 259.950 81.735 260.320 82.235 ;
        RECT 260.880 81.735 261.250 82.235 ;
        RECT 259.950 81.185 260.120 81.735 ;
        RECT 260.370 81.345 260.830 81.575 ;
        RECT 261.080 81.185 261.250 81.735 ;
        RECT 259.950 80.685 260.320 81.185 ;
        RECT 260.880 80.685 261.250 81.185 ;
        RECT 259.950 80.135 260.120 80.685 ;
        RECT 260.370 80.295 260.830 80.525 ;
        RECT 261.080 80.135 261.250 80.685 ;
        RECT 259.950 79.635 260.320 80.135 ;
        RECT 260.880 79.635 261.250 80.135 ;
        RECT 259.950 79.085 260.120 79.635 ;
        RECT 260.370 79.245 260.830 79.475 ;
        RECT 261.080 79.085 261.250 79.635 ;
        RECT 259.950 78.585 260.320 79.085 ;
        RECT 260.880 78.585 261.250 79.085 ;
        RECT 259.950 77.535 260.120 78.585 ;
        RECT 260.350 77.535 260.850 78.425 ;
        RECT 257.910 77.485 258.370 77.535 ;
        RECT 260.370 77.485 260.830 77.535 ;
        RECT 261.080 77.085 261.250 78.585 ;
        RECT 261.450 77.540 262.210 94.450 ;
        RECT 262.830 93.400 263.290 93.445 ;
        RECT 262.410 92.350 262.580 93.400 ;
        RECT 262.810 92.510 263.310 93.400 ;
        RECT 263.540 92.350 263.710 93.400 ;
        RECT 262.410 91.850 262.780 92.350 ;
        RECT 263.340 91.850 263.710 92.350 ;
        RECT 262.410 91.300 262.580 91.850 ;
        RECT 262.830 91.460 263.290 91.690 ;
        RECT 263.540 91.300 263.710 91.850 ;
        RECT 262.410 90.800 262.780 91.300 ;
        RECT 263.340 90.800 263.710 91.300 ;
        RECT 262.410 90.250 262.580 90.800 ;
        RECT 262.830 90.410 263.290 90.640 ;
        RECT 263.540 90.250 263.710 90.800 ;
        RECT 262.410 89.750 262.780 90.250 ;
        RECT 263.340 89.750 263.710 90.250 ;
        RECT 262.410 89.200 262.580 89.750 ;
        RECT 262.830 89.360 263.290 89.590 ;
        RECT 263.540 89.200 263.710 89.750 ;
        RECT 262.410 88.700 262.780 89.200 ;
        RECT 263.340 88.700 263.710 89.200 ;
        RECT 262.410 87.735 262.580 88.700 ;
        RECT 262.830 88.310 263.290 88.540 ;
        RECT 263.540 87.735 263.710 88.700 ;
        RECT 262.410 87.565 263.710 87.735 ;
        RECT 262.410 86.555 262.580 87.565 ;
        RECT 262.830 86.760 263.290 86.990 ;
        RECT 263.540 86.555 263.710 87.565 ;
        RECT 262.410 85.055 262.780 86.555 ;
        RECT 263.340 85.055 263.710 86.555 ;
        RECT 262.410 84.415 262.580 85.055 ;
        RECT 262.830 84.620 263.290 84.850 ;
        RECT 263.540 84.415 263.710 85.055 ;
        RECT 262.410 82.915 262.780 84.415 ;
        RECT 263.340 82.915 263.710 84.415 ;
        RECT 262.410 82.275 262.580 82.915 ;
        RECT 262.830 82.480 263.290 82.710 ;
        RECT 263.540 82.275 263.710 82.915 ;
        RECT 262.410 80.775 262.780 82.275 ;
        RECT 263.340 80.775 263.710 82.275 ;
        RECT 262.410 80.135 262.580 80.775 ;
        RECT 262.830 80.340 263.290 80.570 ;
        RECT 263.540 80.135 263.710 80.775 ;
        RECT 262.410 78.635 262.780 80.135 ;
        RECT 263.340 78.635 263.710 80.135 ;
        RECT 262.810 77.540 263.310 78.430 ;
        RECT 261.450 77.535 261.830 77.540 ;
        RECT 262.830 77.485 263.290 77.540 ;
        RECT 263.540 77.085 263.710 78.635 ;
        RECT 263.910 92.305 264.670 134.995 ;
        RECT 267.930 134.950 269.630 134.995 ;
        RECT 270.190 134.950 271.560 135.450 ;
        RECT 272.120 134.950 273.560 135.450 ;
        RECT 265.290 134.785 265.750 134.790 ;
        RECT 265.270 124.850 265.770 134.785 ;
        RECT 267.200 129.850 267.700 134.790 ;
        RECT 267.930 133.900 269.430 134.950 ;
        RECT 269.660 130.850 270.160 134.790 ;
        RECT 271.590 134.200 272.090 134.790 ;
        RECT 265.270 92.515 265.770 102.450 ;
        RECT 265.290 92.510 265.750 92.515 ;
        RECT 267.200 92.510 267.700 97.450 ;
        RECT 267.930 92.350 269.430 93.400 ;
        RECT 269.660 92.510 270.160 96.450 ;
        RECT 271.590 92.510 272.090 93.100 ;
        RECT 272.690 92.350 273.560 134.950 ;
        RECT 273.910 127.850 274.210 136.510 ;
        RECT 274.635 136.100 274.995 136.520 ;
        RECT 274.685 128.850 274.985 134.475 ;
        RECT 276.400 131.850 276.890 151.850 ;
        RECT 278.440 150.350 278.740 151.740 ;
        RECT 278.410 149.930 278.770 150.350 ;
        RECT 277.425 148.120 277.725 149.850 ;
        RECT 278.415 149.030 278.775 149.450 ;
        RECT 278.360 148.120 278.660 148.520 ;
        RECT 279.110 144.795 279.410 149.440 ;
        RECT 278.275 143.765 278.635 144.185 ;
        RECT 277.425 129.850 277.725 136.510 ;
        RECT 278.295 136.100 278.655 136.520 ;
        RECT 279.060 135.145 279.460 135.645 ;
        RECT 278.305 130.850 278.605 134.475 ;
        RECT 279.060 125.850 279.360 135.145 ;
        RECT 279.730 132.850 280.220 150.410 ;
        RECT 284.870 150.215 285.380 150.815 ;
        RECT 287.330 150.215 287.840 150.815 ;
        RECT 281.870 149.765 282.330 149.815 ;
        RECT 284.330 149.765 284.790 149.815 ;
        RECT 280.870 132.850 281.250 149.765 ;
        RECT 281.850 148.875 282.350 149.765 ;
        RECT 282.580 148.670 282.750 149.765 ;
        RECT 281.450 147.170 281.820 148.670 ;
        RECT 282.380 147.170 282.750 148.670 ;
        RECT 281.450 146.530 281.620 147.170 ;
        RECT 281.870 146.735 282.330 146.965 ;
        RECT 282.580 146.530 282.750 147.170 ;
        RECT 281.450 145.030 281.820 146.530 ;
        RECT 282.380 145.030 282.750 146.530 ;
        RECT 281.450 144.390 281.620 145.030 ;
        RECT 281.870 144.595 282.330 144.825 ;
        RECT 282.580 144.390 282.750 145.030 ;
        RECT 281.450 142.890 281.820 144.390 ;
        RECT 282.380 142.890 282.750 144.390 ;
        RECT 281.450 142.250 281.620 142.890 ;
        RECT 281.870 142.455 282.330 142.685 ;
        RECT 282.580 142.250 282.750 142.890 ;
        RECT 281.450 140.750 281.820 142.250 ;
        RECT 282.380 140.750 282.750 142.250 ;
        RECT 281.450 139.740 281.620 140.750 ;
        RECT 281.870 140.315 282.330 140.545 ;
        RECT 282.580 139.740 282.750 140.750 ;
        RECT 281.450 139.570 282.750 139.740 ;
        RECT 281.450 138.605 281.620 139.570 ;
        RECT 281.870 138.765 282.330 138.995 ;
        RECT 282.580 138.605 282.750 139.570 ;
        RECT 281.450 138.105 281.820 138.605 ;
        RECT 282.380 138.105 282.750 138.605 ;
        RECT 281.450 137.555 281.620 138.105 ;
        RECT 281.870 137.715 282.330 137.945 ;
        RECT 282.580 137.555 282.750 138.105 ;
        RECT 281.450 137.055 281.820 137.555 ;
        RECT 282.380 137.055 282.750 137.555 ;
        RECT 281.450 136.505 281.620 137.055 ;
        RECT 281.870 136.665 282.330 136.895 ;
        RECT 282.580 136.505 282.750 137.055 ;
        RECT 281.450 136.005 281.820 136.505 ;
        RECT 282.380 136.005 282.750 136.505 ;
        RECT 281.450 135.455 281.620 136.005 ;
        RECT 281.870 135.615 282.330 135.845 ;
        RECT 282.580 135.455 282.750 136.005 ;
        RECT 281.450 134.955 281.820 135.455 ;
        RECT 282.380 134.955 282.750 135.455 ;
        RECT 281.450 127.450 281.620 134.955 ;
        RECT 281.850 133.905 282.350 134.795 ;
        RECT 282.580 133.905 282.750 134.955 ;
        RECT 281.870 133.855 282.330 133.905 ;
        RECT 282.950 131.850 283.710 149.765 ;
        RECT 283.910 148.715 284.080 149.765 ;
        RECT 284.310 148.875 284.810 149.765 ;
        RECT 285.040 148.715 285.210 150.215 ;
        RECT 283.910 148.215 284.280 148.715 ;
        RECT 284.840 148.215 285.210 148.715 ;
        RECT 283.910 147.665 284.080 148.215 ;
        RECT 284.330 147.825 284.790 148.055 ;
        RECT 285.040 147.665 285.210 148.215 ;
        RECT 283.910 147.165 284.280 147.665 ;
        RECT 284.840 147.165 285.210 147.665 ;
        RECT 283.910 146.615 284.080 147.165 ;
        RECT 284.330 146.775 284.790 147.005 ;
        RECT 285.040 146.615 285.210 147.165 ;
        RECT 283.910 146.115 284.280 146.615 ;
        RECT 284.840 146.115 285.210 146.615 ;
        RECT 283.910 145.565 284.080 146.115 ;
        RECT 284.330 145.725 284.790 145.955 ;
        RECT 285.040 145.565 285.210 146.115 ;
        RECT 283.910 145.065 284.280 145.565 ;
        RECT 284.840 145.065 285.210 145.565 ;
        RECT 283.910 142.920 284.080 145.065 ;
        RECT 284.330 144.675 284.790 144.905 ;
        RECT 284.330 143.125 284.790 143.355 ;
        RECT 285.040 142.920 285.210 145.065 ;
        RECT 283.910 141.420 284.280 142.920 ;
        RECT 284.840 141.420 285.210 142.920 ;
        RECT 283.910 140.780 284.080 141.420 ;
        RECT 284.330 140.985 284.790 141.215 ;
        RECT 285.040 140.780 285.210 141.420 ;
        RECT 283.910 139.280 284.280 140.780 ;
        RECT 284.840 139.280 285.210 140.780 ;
        RECT 283.910 138.640 284.080 139.280 ;
        RECT 284.330 138.845 284.790 139.075 ;
        RECT 285.040 138.640 285.210 139.280 ;
        RECT 283.910 137.140 284.280 138.640 ;
        RECT 284.840 137.140 285.210 138.640 ;
        RECT 283.910 136.500 284.080 137.140 ;
        RECT 284.330 136.705 284.790 136.935 ;
        RECT 285.040 136.500 285.210 137.140 ;
        RECT 283.910 135.000 284.280 136.500 ;
        RECT 284.840 135.000 285.210 136.500 ;
        RECT 285.410 149.760 285.790 149.765 ;
        RECT 286.790 149.760 287.250 149.815 ;
        RECT 283.910 127.450 284.080 135.000 ;
        RECT 284.310 133.905 284.810 134.795 ;
        RECT 284.330 127.850 284.790 133.905 ;
        RECT 285.410 132.850 286.170 149.760 ;
        RECT 286.770 148.870 287.270 149.760 ;
        RECT 287.500 148.665 287.670 150.215 ;
        RECT 286.370 147.165 286.740 148.665 ;
        RECT 287.300 147.165 287.670 148.665 ;
        RECT 286.370 146.525 286.540 147.165 ;
        RECT 286.790 146.730 287.250 146.960 ;
        RECT 287.500 146.525 287.670 147.165 ;
        RECT 286.370 145.025 286.740 146.525 ;
        RECT 287.300 145.025 287.670 146.525 ;
        RECT 286.370 144.385 286.540 145.025 ;
        RECT 286.790 144.590 287.250 144.820 ;
        RECT 287.500 144.385 287.670 145.025 ;
        RECT 286.370 142.885 286.740 144.385 ;
        RECT 287.300 142.885 287.670 144.385 ;
        RECT 286.370 142.245 286.540 142.885 ;
        RECT 286.790 142.450 287.250 142.680 ;
        RECT 287.500 142.245 287.670 142.885 ;
        RECT 286.370 140.745 286.740 142.245 ;
        RECT 287.300 140.745 287.670 142.245 ;
        RECT 286.370 139.735 286.540 140.745 ;
        RECT 286.790 140.310 287.250 140.540 ;
        RECT 287.500 139.735 287.670 140.745 ;
        RECT 286.370 139.565 287.670 139.735 ;
        RECT 286.370 138.600 286.540 139.565 ;
        RECT 286.790 138.760 287.250 138.990 ;
        RECT 287.500 138.600 287.670 139.565 ;
        RECT 286.370 138.100 286.740 138.600 ;
        RECT 287.300 138.100 287.670 138.600 ;
        RECT 286.370 137.550 286.540 138.100 ;
        RECT 286.790 137.710 287.250 137.940 ;
        RECT 287.500 137.550 287.670 138.100 ;
        RECT 286.370 137.050 286.740 137.550 ;
        RECT 287.300 137.050 287.670 137.550 ;
        RECT 286.370 136.500 286.540 137.050 ;
        RECT 286.790 136.660 287.250 136.890 ;
        RECT 287.500 136.500 287.670 137.050 ;
        RECT 286.370 136.000 286.740 136.500 ;
        RECT 287.300 136.000 287.670 136.500 ;
        RECT 286.370 135.450 286.540 136.000 ;
        RECT 286.790 135.610 287.250 135.840 ;
        RECT 287.500 135.450 287.670 136.000 ;
        RECT 286.370 134.950 286.740 135.450 ;
        RECT 287.300 134.950 287.670 135.450 ;
        RECT 286.370 133.900 286.540 134.950 ;
        RECT 286.770 133.900 287.270 134.790 ;
        RECT 287.500 133.900 287.670 134.950 ;
        RECT 287.870 144.010 288.250 149.760 ;
        RECT 287.870 142.915 288.630 144.010 ;
        RECT 289.250 143.120 289.710 143.350 ;
        RECT 291.180 143.120 291.640 143.350 ;
        RECT 291.890 142.915 293.390 150.815 ;
        RECT 287.870 141.415 289.200 142.915 ;
        RECT 289.760 141.415 291.130 142.915 ;
        RECT 291.690 141.685 293.390 142.915 ;
        RECT 291.690 141.415 293.385 141.685 ;
        RECT 287.870 140.775 289.000 141.415 ;
        RECT 289.250 140.980 289.710 141.210 ;
        RECT 289.960 140.775 290.930 141.415 ;
        RECT 291.180 140.980 291.640 141.210 ;
        RECT 291.890 140.775 293.385 141.415 ;
        RECT 287.870 139.275 289.200 140.775 ;
        RECT 289.760 139.275 291.130 140.775 ;
        RECT 291.690 139.275 293.385 140.775 ;
        RECT 297.030 139.600 297.520 151.850 ;
        RECT 298.565 151.330 298.925 151.750 ;
        RECT 298.485 149.030 298.845 149.450 ;
        RECT 298.560 148.110 298.920 148.530 ;
        RECT 299.525 148.120 299.825 149.850 ;
        RECT 298.610 144.785 298.970 145.205 ;
        RECT 287.870 138.635 289.000 139.275 ;
        RECT 289.250 138.840 289.710 139.070 ;
        RECT 289.960 138.635 290.930 139.275 ;
        RECT 291.180 138.840 291.640 139.070 ;
        RECT 291.890 138.635 293.385 139.275 ;
        RECT 293.640 138.760 294.100 138.990 ;
        RECT 295.570 138.760 296.030 138.990 ;
        RECT 287.870 137.135 289.200 138.635 ;
        RECT 289.760 137.135 291.130 138.635 ;
        RECT 291.690 138.600 293.385 138.635 ;
        RECT 296.650 138.600 297.520 139.600 ;
        RECT 291.690 138.100 293.590 138.600 ;
        RECT 294.150 138.100 295.520 138.600 ;
        RECT 296.080 138.100 297.520 138.600 ;
        RECT 291.690 137.550 293.385 138.100 ;
        RECT 293.640 137.710 294.100 137.940 ;
        RECT 294.350 137.550 295.320 138.100 ;
        RECT 295.570 137.710 296.030 137.940 ;
        RECT 296.280 137.550 297.520 138.100 ;
        RECT 291.690 137.135 293.590 137.550 ;
        RECT 287.870 136.495 289.000 137.135 ;
        RECT 289.250 136.700 289.710 136.930 ;
        RECT 289.960 136.495 290.930 137.135 ;
        RECT 291.890 137.050 293.590 137.135 ;
        RECT 294.150 137.050 295.520 137.550 ;
        RECT 296.080 137.050 297.520 137.550 ;
        RECT 291.180 136.700 291.640 136.930 ;
        RECT 291.890 136.500 293.385 137.050 ;
        RECT 293.640 136.660 294.100 136.890 ;
        RECT 294.350 136.500 295.320 137.050 ;
        RECT 295.570 136.660 296.030 136.890 ;
        RECT 296.280 136.500 297.520 137.050 ;
        RECT 291.890 136.495 293.590 136.500 ;
        RECT 287.870 134.995 289.200 136.495 ;
        RECT 289.760 134.995 291.130 136.495 ;
        RECT 291.690 136.000 293.590 136.495 ;
        RECT 294.150 136.000 295.520 136.500 ;
        RECT 296.080 136.000 297.520 136.500 ;
        RECT 291.690 135.450 293.385 136.000 ;
        RECT 293.640 135.610 294.100 135.840 ;
        RECT 294.350 135.450 295.320 136.000 ;
        RECT 295.570 135.610 296.030 135.840 ;
        RECT 296.280 135.450 297.520 136.000 ;
        RECT 291.690 134.995 293.590 135.450 ;
        RECT 286.790 133.855 287.250 133.900 ;
        RECT 281.280 126.850 281.790 127.450 ;
        RECT 283.740 126.850 284.250 127.450 ;
        RECT 280.870 110.900 281.370 126.450 ;
        RECT 281.870 119.900 282.370 125.450 ;
        RECT 281.820 119.400 282.420 119.900 ;
        RECT 280.820 110.400 281.420 110.900 ;
        RECT 267.930 92.305 269.630 92.350 ;
        RECT 263.910 90.805 265.240 92.305 ;
        RECT 265.800 90.805 267.170 92.305 ;
        RECT 267.730 91.850 269.630 92.305 ;
        RECT 270.190 91.850 271.560 92.350 ;
        RECT 272.120 91.850 273.560 92.350 ;
        RECT 267.730 91.300 269.430 91.850 ;
        RECT 269.680 91.460 270.140 91.690 ;
        RECT 270.390 91.300 271.360 91.850 ;
        RECT 271.610 91.460 272.070 91.690 ;
        RECT 272.320 91.300 273.560 91.850 ;
        RECT 267.730 90.805 269.630 91.300 ;
        RECT 263.910 90.165 265.040 90.805 ;
        RECT 265.290 90.370 265.750 90.600 ;
        RECT 266.000 90.165 266.970 90.805 ;
        RECT 267.930 90.800 269.630 90.805 ;
        RECT 270.190 90.800 271.560 91.300 ;
        RECT 272.120 90.800 273.560 91.300 ;
        RECT 267.220 90.370 267.680 90.600 ;
        RECT 267.930 90.250 269.430 90.800 ;
        RECT 269.680 90.410 270.140 90.640 ;
        RECT 270.390 90.250 271.360 90.800 ;
        RECT 271.610 90.410 272.070 90.640 ;
        RECT 272.320 90.250 273.560 90.800 ;
        RECT 273.910 90.790 274.210 99.450 ;
        RECT 274.685 92.825 274.985 98.450 ;
        RECT 274.635 90.780 274.995 91.200 ;
        RECT 267.930 90.165 269.630 90.250 ;
        RECT 263.910 88.665 265.240 90.165 ;
        RECT 265.800 88.665 267.170 90.165 ;
        RECT 267.730 89.750 269.630 90.165 ;
        RECT 270.190 89.750 271.560 90.250 ;
        RECT 272.120 89.750 273.560 90.250 ;
        RECT 267.730 89.200 269.430 89.750 ;
        RECT 269.680 89.360 270.140 89.590 ;
        RECT 270.390 89.200 271.360 89.750 ;
        RECT 271.610 89.360 272.070 89.590 ;
        RECT 272.320 89.200 273.560 89.750 ;
        RECT 267.730 88.700 269.630 89.200 ;
        RECT 270.190 88.700 271.560 89.200 ;
        RECT 272.120 88.700 273.560 89.200 ;
        RECT 267.730 88.665 269.430 88.700 ;
        RECT 263.910 88.025 265.040 88.665 ;
        RECT 265.290 88.230 265.750 88.460 ;
        RECT 266.000 88.025 266.970 88.665 ;
        RECT 267.220 88.230 267.680 88.460 ;
        RECT 267.930 88.025 269.430 88.665 ;
        RECT 269.680 88.310 270.140 88.540 ;
        RECT 271.610 88.310 272.070 88.540 ;
        RECT 263.910 86.525 265.240 88.025 ;
        RECT 265.800 86.525 267.170 88.025 ;
        RECT 267.730 86.525 269.430 88.025 ;
        RECT 272.690 87.700 273.560 88.700 ;
        RECT 263.910 85.885 265.040 86.525 ;
        RECT 265.290 86.090 265.750 86.320 ;
        RECT 266.000 85.885 266.970 86.525 ;
        RECT 267.220 86.090 267.680 86.320 ;
        RECT 267.930 85.885 269.430 86.525 ;
        RECT 263.910 84.385 265.240 85.885 ;
        RECT 265.800 84.385 267.170 85.885 ;
        RECT 267.730 84.385 269.430 85.885 ;
        RECT 263.910 83.290 264.670 84.385 ;
        RECT 265.290 83.950 265.750 84.180 ;
        RECT 267.220 83.950 267.680 84.180 ;
        RECT 263.910 77.540 264.290 83.290 ;
        RECT 260.910 76.485 261.420 77.085 ;
        RECT 263.370 76.485 263.880 77.085 ;
        RECT 267.930 76.485 269.430 84.385 ;
        RECT 273.070 75.450 273.560 87.700 ;
        RECT 274.650 82.095 275.010 82.515 ;
        RECT 274.600 78.770 274.960 79.190 ;
        RECT 274.525 77.850 274.885 78.270 ;
        RECT 275.565 77.450 275.865 79.180 ;
        RECT 274.605 75.550 274.965 75.970 ;
        RECT 276.400 75.450 276.890 95.450 ;
        RECT 277.425 90.790 277.725 97.450 ;
        RECT 278.305 92.825 278.605 96.450 ;
        RECT 279.060 92.155 279.360 101.450 ;
        RECT 280.870 100.850 281.370 110.400 ;
        RECT 281.870 101.850 282.370 103.100 ;
        RECT 281.280 99.850 281.790 100.450 ;
        RECT 283.740 99.850 284.250 100.450 ;
        RECT 279.060 91.655 279.460 92.155 ;
        RECT 278.295 90.780 278.655 91.200 ;
        RECT 278.275 83.115 278.635 83.535 ;
        RECT 277.425 77.450 277.725 79.180 ;
        RECT 278.360 78.780 278.660 79.180 ;
        RECT 278.415 77.850 278.775 78.270 ;
        RECT 279.110 77.860 279.410 82.505 ;
        RECT 278.410 76.950 278.770 77.370 ;
        RECT 278.440 75.560 278.740 76.950 ;
        RECT 279.730 76.890 280.220 94.450 ;
        RECT 280.870 77.535 281.250 94.450 ;
        RECT 281.450 92.345 281.620 99.850 ;
        RECT 281.870 93.395 282.330 93.445 ;
        RECT 281.850 92.505 282.350 93.395 ;
        RECT 282.580 92.345 282.750 93.395 ;
        RECT 281.450 91.845 281.820 92.345 ;
        RECT 282.380 91.845 282.750 92.345 ;
        RECT 281.450 91.295 281.620 91.845 ;
        RECT 281.870 91.455 282.330 91.685 ;
        RECT 282.580 91.295 282.750 91.845 ;
        RECT 281.450 90.795 281.820 91.295 ;
        RECT 282.380 90.795 282.750 91.295 ;
        RECT 281.450 90.245 281.620 90.795 ;
        RECT 281.870 90.405 282.330 90.635 ;
        RECT 282.580 90.245 282.750 90.795 ;
        RECT 281.450 89.745 281.820 90.245 ;
        RECT 282.380 89.745 282.750 90.245 ;
        RECT 281.450 89.195 281.620 89.745 ;
        RECT 281.870 89.355 282.330 89.585 ;
        RECT 282.580 89.195 282.750 89.745 ;
        RECT 281.450 88.695 281.820 89.195 ;
        RECT 282.380 88.695 282.750 89.195 ;
        RECT 281.450 87.730 281.620 88.695 ;
        RECT 281.870 88.305 282.330 88.535 ;
        RECT 282.580 87.730 282.750 88.695 ;
        RECT 281.450 87.560 282.750 87.730 ;
        RECT 281.450 86.550 281.620 87.560 ;
        RECT 281.870 86.755 282.330 86.985 ;
        RECT 282.580 86.550 282.750 87.560 ;
        RECT 281.450 85.050 281.820 86.550 ;
        RECT 282.380 85.050 282.750 86.550 ;
        RECT 281.450 84.410 281.620 85.050 ;
        RECT 281.870 84.615 282.330 84.845 ;
        RECT 282.580 84.410 282.750 85.050 ;
        RECT 281.450 82.910 281.820 84.410 ;
        RECT 282.380 82.910 282.750 84.410 ;
        RECT 281.450 82.270 281.620 82.910 ;
        RECT 281.870 82.475 282.330 82.705 ;
        RECT 282.580 82.270 282.750 82.910 ;
        RECT 281.450 80.770 281.820 82.270 ;
        RECT 282.380 80.770 282.750 82.270 ;
        RECT 281.450 80.130 281.620 80.770 ;
        RECT 281.870 80.335 282.330 80.565 ;
        RECT 282.580 80.130 282.750 80.770 ;
        RECT 281.450 78.630 281.820 80.130 ;
        RECT 282.380 78.630 282.750 80.130 ;
        RECT 281.850 77.535 282.350 78.425 ;
        RECT 282.580 77.535 282.750 78.630 ;
        RECT 282.950 77.535 283.710 95.450 ;
        RECT 283.910 92.300 284.080 99.850 ;
        RECT 284.330 93.395 284.790 99.450 ;
        RECT 284.310 92.505 284.810 93.395 ;
        RECT 283.910 90.800 284.280 92.300 ;
        RECT 284.840 90.800 285.210 92.300 ;
        RECT 283.910 90.160 284.080 90.800 ;
        RECT 284.330 90.365 284.790 90.595 ;
        RECT 285.040 90.160 285.210 90.800 ;
        RECT 283.910 88.660 284.280 90.160 ;
        RECT 284.840 88.660 285.210 90.160 ;
        RECT 283.910 88.020 284.080 88.660 ;
        RECT 284.330 88.225 284.790 88.455 ;
        RECT 285.040 88.020 285.210 88.660 ;
        RECT 283.910 86.520 284.280 88.020 ;
        RECT 284.840 86.520 285.210 88.020 ;
        RECT 283.910 85.880 284.080 86.520 ;
        RECT 284.330 86.085 284.790 86.315 ;
        RECT 285.040 85.880 285.210 86.520 ;
        RECT 283.910 84.380 284.280 85.880 ;
        RECT 284.840 84.380 285.210 85.880 ;
        RECT 283.910 82.235 284.080 84.380 ;
        RECT 284.330 83.945 284.790 84.175 ;
        RECT 284.330 82.395 284.790 82.625 ;
        RECT 285.040 82.235 285.210 84.380 ;
        RECT 283.910 81.735 284.280 82.235 ;
        RECT 284.840 81.735 285.210 82.235 ;
        RECT 283.910 81.185 284.080 81.735 ;
        RECT 284.330 81.345 284.790 81.575 ;
        RECT 285.040 81.185 285.210 81.735 ;
        RECT 283.910 80.685 284.280 81.185 ;
        RECT 284.840 80.685 285.210 81.185 ;
        RECT 283.910 80.135 284.080 80.685 ;
        RECT 284.330 80.295 284.790 80.525 ;
        RECT 285.040 80.135 285.210 80.685 ;
        RECT 283.910 79.635 284.280 80.135 ;
        RECT 284.840 79.635 285.210 80.135 ;
        RECT 283.910 79.085 284.080 79.635 ;
        RECT 284.330 79.245 284.790 79.475 ;
        RECT 285.040 79.085 285.210 79.635 ;
        RECT 283.910 78.585 284.280 79.085 ;
        RECT 284.840 78.585 285.210 79.085 ;
        RECT 283.910 77.535 284.080 78.585 ;
        RECT 284.310 77.535 284.810 78.425 ;
        RECT 281.870 77.485 282.330 77.535 ;
        RECT 284.330 77.485 284.790 77.535 ;
        RECT 285.040 77.085 285.210 78.585 ;
        RECT 285.410 77.540 286.170 94.450 ;
        RECT 286.790 93.400 287.250 93.445 ;
        RECT 286.370 92.350 286.540 93.400 ;
        RECT 286.770 92.510 287.270 93.400 ;
        RECT 287.500 92.350 287.670 93.400 ;
        RECT 286.370 91.850 286.740 92.350 ;
        RECT 287.300 91.850 287.670 92.350 ;
        RECT 286.370 91.300 286.540 91.850 ;
        RECT 286.790 91.460 287.250 91.690 ;
        RECT 287.500 91.300 287.670 91.850 ;
        RECT 286.370 90.800 286.740 91.300 ;
        RECT 287.300 90.800 287.670 91.300 ;
        RECT 286.370 90.250 286.540 90.800 ;
        RECT 286.790 90.410 287.250 90.640 ;
        RECT 287.500 90.250 287.670 90.800 ;
        RECT 286.370 89.750 286.740 90.250 ;
        RECT 287.300 89.750 287.670 90.250 ;
        RECT 286.370 89.200 286.540 89.750 ;
        RECT 286.790 89.360 287.250 89.590 ;
        RECT 287.500 89.200 287.670 89.750 ;
        RECT 286.370 88.700 286.740 89.200 ;
        RECT 287.300 88.700 287.670 89.200 ;
        RECT 286.370 87.735 286.540 88.700 ;
        RECT 286.790 88.310 287.250 88.540 ;
        RECT 287.500 87.735 287.670 88.700 ;
        RECT 286.370 87.565 287.670 87.735 ;
        RECT 286.370 86.555 286.540 87.565 ;
        RECT 286.790 86.760 287.250 86.990 ;
        RECT 287.500 86.555 287.670 87.565 ;
        RECT 286.370 85.055 286.740 86.555 ;
        RECT 287.300 85.055 287.670 86.555 ;
        RECT 286.370 84.415 286.540 85.055 ;
        RECT 286.790 84.620 287.250 84.850 ;
        RECT 287.500 84.415 287.670 85.055 ;
        RECT 286.370 82.915 286.740 84.415 ;
        RECT 287.300 82.915 287.670 84.415 ;
        RECT 286.370 82.275 286.540 82.915 ;
        RECT 286.790 82.480 287.250 82.710 ;
        RECT 287.500 82.275 287.670 82.915 ;
        RECT 286.370 80.775 286.740 82.275 ;
        RECT 287.300 80.775 287.670 82.275 ;
        RECT 286.370 80.135 286.540 80.775 ;
        RECT 286.790 80.340 287.250 80.570 ;
        RECT 287.500 80.135 287.670 80.775 ;
        RECT 286.370 78.635 286.740 80.135 ;
        RECT 287.300 78.635 287.670 80.135 ;
        RECT 286.770 77.540 287.270 78.430 ;
        RECT 285.410 77.535 285.790 77.540 ;
        RECT 286.790 77.485 287.250 77.540 ;
        RECT 287.500 77.085 287.670 78.635 ;
        RECT 287.870 92.305 288.630 134.995 ;
        RECT 291.890 134.950 293.590 134.995 ;
        RECT 294.150 134.950 295.520 135.450 ;
        RECT 296.080 134.950 297.520 135.450 ;
        RECT 289.250 134.785 289.710 134.790 ;
        RECT 289.230 124.850 289.730 134.785 ;
        RECT 291.160 129.850 291.660 134.790 ;
        RECT 291.890 133.900 293.385 134.950 ;
        RECT 293.620 130.850 294.120 134.790 ;
        RECT 295.550 134.200 296.050 134.790 ;
        RECT 289.230 92.515 289.730 102.450 ;
        RECT 289.250 92.510 289.710 92.515 ;
        RECT 291.160 92.510 291.660 97.450 ;
        RECT 291.890 92.350 293.385 93.400 ;
        RECT 293.620 92.510 294.120 96.450 ;
        RECT 295.550 92.510 296.050 93.100 ;
        RECT 296.650 92.350 297.520 134.950 ;
        RECT 297.870 127.850 298.170 136.510 ;
        RECT 298.595 136.100 298.955 136.520 ;
        RECT 298.645 128.850 298.945 134.475 ;
        RECT 300.360 131.850 300.850 151.850 ;
        RECT 302.400 150.350 302.700 151.740 ;
        RECT 302.370 149.930 302.730 150.350 ;
        RECT 301.385 148.120 301.685 149.850 ;
        RECT 302.375 149.030 302.735 149.450 ;
        RECT 302.320 148.120 302.620 148.520 ;
        RECT 303.070 144.795 303.370 149.440 ;
        RECT 302.235 143.765 302.595 144.185 ;
        RECT 301.385 129.850 301.685 136.510 ;
        RECT 302.255 136.100 302.615 136.520 ;
        RECT 303.020 135.145 303.420 135.645 ;
        RECT 302.265 130.850 302.565 134.475 ;
        RECT 303.020 125.850 303.320 135.145 ;
        RECT 303.690 132.850 304.180 150.410 ;
        RECT 308.880 150.215 309.390 150.815 ;
        RECT 311.340 150.215 311.850 150.815 ;
        RECT 305.880 149.765 306.340 149.815 ;
        RECT 308.340 149.765 308.800 149.815 ;
        RECT 304.880 132.850 305.260 149.765 ;
        RECT 305.860 148.875 306.360 149.765 ;
        RECT 306.590 148.670 306.760 149.765 ;
        RECT 305.460 147.170 305.830 148.670 ;
        RECT 306.390 147.170 306.760 148.670 ;
        RECT 305.460 146.530 305.630 147.170 ;
        RECT 305.880 146.735 306.340 146.965 ;
        RECT 306.590 146.530 306.760 147.170 ;
        RECT 305.460 145.030 305.830 146.530 ;
        RECT 306.390 145.030 306.760 146.530 ;
        RECT 305.460 144.390 305.630 145.030 ;
        RECT 305.880 144.595 306.340 144.825 ;
        RECT 306.590 144.390 306.760 145.030 ;
        RECT 305.460 142.890 305.830 144.390 ;
        RECT 306.390 142.890 306.760 144.390 ;
        RECT 305.460 142.250 305.630 142.890 ;
        RECT 305.880 142.455 306.340 142.685 ;
        RECT 306.590 142.250 306.760 142.890 ;
        RECT 305.460 140.750 305.830 142.250 ;
        RECT 306.390 140.750 306.760 142.250 ;
        RECT 305.460 139.740 305.630 140.750 ;
        RECT 305.880 140.315 306.340 140.545 ;
        RECT 306.590 139.740 306.760 140.750 ;
        RECT 305.460 139.570 306.760 139.740 ;
        RECT 305.460 138.605 305.630 139.570 ;
        RECT 305.880 138.765 306.340 138.995 ;
        RECT 306.590 138.605 306.760 139.570 ;
        RECT 305.460 138.105 305.830 138.605 ;
        RECT 306.390 138.105 306.760 138.605 ;
        RECT 305.460 137.555 305.630 138.105 ;
        RECT 305.880 137.715 306.340 137.945 ;
        RECT 306.590 137.555 306.760 138.105 ;
        RECT 305.460 137.055 305.830 137.555 ;
        RECT 306.390 137.055 306.760 137.555 ;
        RECT 305.460 136.505 305.630 137.055 ;
        RECT 305.880 136.665 306.340 136.895 ;
        RECT 306.590 136.505 306.760 137.055 ;
        RECT 305.460 136.005 305.830 136.505 ;
        RECT 306.390 136.005 306.760 136.505 ;
        RECT 305.460 135.455 305.630 136.005 ;
        RECT 305.880 135.615 306.340 135.845 ;
        RECT 306.590 135.455 306.760 136.005 ;
        RECT 305.460 134.955 305.830 135.455 ;
        RECT 306.390 134.955 306.760 135.455 ;
        RECT 305.460 127.450 305.630 134.955 ;
        RECT 305.860 133.905 306.360 134.795 ;
        RECT 306.590 133.905 306.760 134.955 ;
        RECT 305.880 133.855 306.340 133.905 ;
        RECT 306.960 131.850 307.720 149.765 ;
        RECT 307.920 148.715 308.090 149.765 ;
        RECT 308.320 148.875 308.820 149.765 ;
        RECT 309.050 148.715 309.220 150.215 ;
        RECT 307.920 148.215 308.290 148.715 ;
        RECT 308.850 148.215 309.220 148.715 ;
        RECT 307.920 147.665 308.090 148.215 ;
        RECT 308.340 147.825 308.800 148.055 ;
        RECT 309.050 147.665 309.220 148.215 ;
        RECT 307.920 147.165 308.290 147.665 ;
        RECT 308.850 147.165 309.220 147.665 ;
        RECT 307.920 146.615 308.090 147.165 ;
        RECT 308.340 146.775 308.800 147.005 ;
        RECT 309.050 146.615 309.220 147.165 ;
        RECT 307.920 146.115 308.290 146.615 ;
        RECT 308.850 146.115 309.220 146.615 ;
        RECT 307.920 145.565 308.090 146.115 ;
        RECT 308.340 145.725 308.800 145.955 ;
        RECT 309.050 145.565 309.220 146.115 ;
        RECT 307.920 145.065 308.290 145.565 ;
        RECT 308.850 145.065 309.220 145.565 ;
        RECT 307.920 142.920 308.090 145.065 ;
        RECT 308.340 144.675 308.800 144.905 ;
        RECT 308.340 143.125 308.800 143.355 ;
        RECT 309.050 142.920 309.220 145.065 ;
        RECT 307.920 141.420 308.290 142.920 ;
        RECT 308.850 141.420 309.220 142.920 ;
        RECT 307.920 140.780 308.090 141.420 ;
        RECT 308.340 140.985 308.800 141.215 ;
        RECT 309.050 140.780 309.220 141.420 ;
        RECT 307.920 139.280 308.290 140.780 ;
        RECT 308.850 139.280 309.220 140.780 ;
        RECT 307.920 138.640 308.090 139.280 ;
        RECT 308.340 138.845 308.800 139.075 ;
        RECT 309.050 138.640 309.220 139.280 ;
        RECT 307.920 137.140 308.290 138.640 ;
        RECT 308.850 137.140 309.220 138.640 ;
        RECT 307.920 136.500 308.090 137.140 ;
        RECT 308.340 136.705 308.800 136.935 ;
        RECT 309.050 136.500 309.220 137.140 ;
        RECT 307.920 135.000 308.290 136.500 ;
        RECT 308.850 135.000 309.220 136.500 ;
        RECT 309.420 149.760 309.800 149.765 ;
        RECT 310.800 149.760 311.260 149.815 ;
        RECT 307.920 127.450 308.090 135.000 ;
        RECT 308.320 133.905 308.820 134.795 ;
        RECT 308.340 127.850 308.800 133.905 ;
        RECT 309.420 132.850 310.180 149.760 ;
        RECT 310.780 148.870 311.280 149.760 ;
        RECT 311.510 148.665 311.680 150.215 ;
        RECT 310.380 147.165 310.750 148.665 ;
        RECT 311.310 147.165 311.680 148.665 ;
        RECT 310.380 146.525 310.550 147.165 ;
        RECT 310.800 146.730 311.260 146.960 ;
        RECT 311.510 146.525 311.680 147.165 ;
        RECT 310.380 145.025 310.750 146.525 ;
        RECT 311.310 145.025 311.680 146.525 ;
        RECT 310.380 144.385 310.550 145.025 ;
        RECT 310.800 144.590 311.260 144.820 ;
        RECT 311.510 144.385 311.680 145.025 ;
        RECT 310.380 142.885 310.750 144.385 ;
        RECT 311.310 142.885 311.680 144.385 ;
        RECT 310.380 142.245 310.550 142.885 ;
        RECT 310.800 142.450 311.260 142.680 ;
        RECT 311.510 142.245 311.680 142.885 ;
        RECT 310.380 140.745 310.750 142.245 ;
        RECT 311.310 140.745 311.680 142.245 ;
        RECT 310.380 139.735 310.550 140.745 ;
        RECT 310.800 140.310 311.260 140.540 ;
        RECT 311.510 139.735 311.680 140.745 ;
        RECT 310.380 139.565 311.680 139.735 ;
        RECT 310.380 138.600 310.550 139.565 ;
        RECT 310.800 138.760 311.260 138.990 ;
        RECT 311.510 138.600 311.680 139.565 ;
        RECT 310.380 138.100 310.750 138.600 ;
        RECT 311.310 138.100 311.680 138.600 ;
        RECT 310.380 137.550 310.550 138.100 ;
        RECT 310.800 137.710 311.260 137.940 ;
        RECT 311.510 137.550 311.680 138.100 ;
        RECT 310.380 137.050 310.750 137.550 ;
        RECT 311.310 137.050 311.680 137.550 ;
        RECT 310.380 136.500 310.550 137.050 ;
        RECT 310.800 136.660 311.260 136.890 ;
        RECT 311.510 136.500 311.680 137.050 ;
        RECT 310.380 136.000 310.750 136.500 ;
        RECT 311.310 136.000 311.680 136.500 ;
        RECT 310.380 135.450 310.550 136.000 ;
        RECT 310.800 135.610 311.260 135.840 ;
        RECT 311.510 135.450 311.680 136.000 ;
        RECT 310.380 134.950 310.750 135.450 ;
        RECT 311.310 134.950 311.680 135.450 ;
        RECT 310.380 133.900 310.550 134.950 ;
        RECT 310.780 133.900 311.280 134.790 ;
        RECT 311.510 133.900 311.680 134.950 ;
        RECT 311.880 144.010 312.260 149.760 ;
        RECT 311.880 142.915 312.640 144.010 ;
        RECT 313.260 143.120 313.720 143.350 ;
        RECT 315.190 143.120 315.650 143.350 ;
        RECT 315.900 142.915 317.400 150.815 ;
        RECT 311.880 141.415 313.210 142.915 ;
        RECT 313.770 141.415 315.140 142.915 ;
        RECT 315.700 141.855 317.400 142.915 ;
        RECT 315.700 141.415 317.450 141.855 ;
        RECT 311.880 140.775 313.010 141.415 ;
        RECT 313.260 140.980 313.720 141.210 ;
        RECT 313.970 140.775 314.940 141.415 ;
        RECT 315.190 140.980 315.650 141.210 ;
        RECT 315.900 140.775 317.450 141.415 ;
        RECT 311.880 139.275 313.210 140.775 ;
        RECT 313.770 139.275 315.140 140.775 ;
        RECT 315.700 139.275 317.450 140.775 ;
        RECT 321.040 139.600 321.530 151.850 ;
        RECT 322.575 151.330 322.935 151.750 ;
        RECT 322.495 149.030 322.855 149.450 ;
        RECT 322.570 148.110 322.930 148.530 ;
        RECT 323.535 148.120 323.835 149.850 ;
        RECT 322.620 144.785 322.980 145.205 ;
        RECT 311.880 138.635 313.010 139.275 ;
        RECT 313.260 138.840 313.720 139.070 ;
        RECT 313.970 138.635 314.940 139.275 ;
        RECT 315.190 138.840 315.650 139.070 ;
        RECT 315.900 138.635 317.450 139.275 ;
        RECT 317.650 138.760 318.110 138.990 ;
        RECT 319.580 138.760 320.040 138.990 ;
        RECT 311.880 137.135 313.210 138.635 ;
        RECT 313.770 137.135 315.140 138.635 ;
        RECT 315.700 138.600 317.450 138.635 ;
        RECT 320.660 138.600 321.530 139.600 ;
        RECT 315.700 138.100 317.600 138.600 ;
        RECT 318.160 138.100 319.530 138.600 ;
        RECT 320.090 138.100 321.530 138.600 ;
        RECT 315.700 137.550 317.450 138.100 ;
        RECT 317.650 137.710 318.110 137.940 ;
        RECT 318.360 137.550 319.330 138.100 ;
        RECT 319.580 137.710 320.040 137.940 ;
        RECT 320.290 137.550 321.530 138.100 ;
        RECT 315.700 137.135 317.600 137.550 ;
        RECT 311.880 136.495 313.010 137.135 ;
        RECT 313.260 136.700 313.720 136.930 ;
        RECT 313.970 136.495 314.940 137.135 ;
        RECT 315.900 137.050 317.600 137.135 ;
        RECT 318.160 137.050 319.530 137.550 ;
        RECT 320.090 137.050 321.530 137.550 ;
        RECT 315.190 136.700 315.650 136.930 ;
        RECT 315.900 136.500 317.450 137.050 ;
        RECT 317.650 136.660 318.110 136.890 ;
        RECT 318.360 136.500 319.330 137.050 ;
        RECT 319.580 136.660 320.040 136.890 ;
        RECT 320.290 136.500 321.530 137.050 ;
        RECT 315.900 136.495 317.600 136.500 ;
        RECT 311.880 134.995 313.210 136.495 ;
        RECT 313.770 134.995 315.140 136.495 ;
        RECT 315.700 136.000 317.600 136.495 ;
        RECT 318.160 136.000 319.530 136.500 ;
        RECT 320.090 136.000 321.530 136.500 ;
        RECT 315.700 135.450 317.450 136.000 ;
        RECT 317.650 135.610 318.110 135.840 ;
        RECT 318.360 135.450 319.330 136.000 ;
        RECT 319.580 135.610 320.040 135.840 ;
        RECT 320.290 135.450 321.530 136.000 ;
        RECT 315.700 134.995 317.600 135.450 ;
        RECT 310.800 133.855 311.260 133.900 ;
        RECT 305.290 126.850 305.800 127.450 ;
        RECT 307.750 126.850 308.260 127.450 ;
        RECT 304.880 109.900 305.380 126.450 ;
        RECT 305.880 118.900 306.380 125.450 ;
        RECT 305.830 118.400 306.430 118.900 ;
        RECT 304.830 109.400 305.430 109.900 ;
        RECT 291.890 92.305 293.590 92.350 ;
        RECT 287.870 90.805 289.200 92.305 ;
        RECT 289.760 90.805 291.130 92.305 ;
        RECT 291.690 91.850 293.590 92.305 ;
        RECT 294.150 91.850 295.520 92.350 ;
        RECT 296.080 91.850 297.520 92.350 ;
        RECT 291.690 91.300 293.385 91.850 ;
        RECT 293.640 91.460 294.100 91.690 ;
        RECT 294.350 91.300 295.320 91.850 ;
        RECT 295.570 91.460 296.030 91.690 ;
        RECT 296.280 91.300 297.520 91.850 ;
        RECT 291.690 90.805 293.590 91.300 ;
        RECT 287.870 90.165 289.000 90.805 ;
        RECT 289.250 90.370 289.710 90.600 ;
        RECT 289.960 90.165 290.930 90.805 ;
        RECT 291.890 90.800 293.590 90.805 ;
        RECT 294.150 90.800 295.520 91.300 ;
        RECT 296.080 90.800 297.520 91.300 ;
        RECT 291.180 90.370 291.640 90.600 ;
        RECT 291.890 90.250 293.385 90.800 ;
        RECT 293.640 90.410 294.100 90.640 ;
        RECT 294.350 90.250 295.320 90.800 ;
        RECT 295.570 90.410 296.030 90.640 ;
        RECT 296.280 90.250 297.520 90.800 ;
        RECT 297.870 90.790 298.170 99.450 ;
        RECT 298.645 92.825 298.945 98.450 ;
        RECT 298.595 90.780 298.955 91.200 ;
        RECT 291.890 90.165 293.590 90.250 ;
        RECT 287.870 88.665 289.200 90.165 ;
        RECT 289.760 88.665 291.130 90.165 ;
        RECT 291.690 89.750 293.590 90.165 ;
        RECT 294.150 89.750 295.520 90.250 ;
        RECT 296.080 89.750 297.520 90.250 ;
        RECT 291.690 89.200 293.385 89.750 ;
        RECT 293.640 89.360 294.100 89.590 ;
        RECT 294.350 89.200 295.320 89.750 ;
        RECT 295.570 89.360 296.030 89.590 ;
        RECT 296.280 89.200 297.520 89.750 ;
        RECT 291.690 88.700 293.590 89.200 ;
        RECT 294.150 88.700 295.520 89.200 ;
        RECT 296.080 88.700 297.520 89.200 ;
        RECT 291.690 88.665 293.385 88.700 ;
        RECT 287.870 88.025 289.000 88.665 ;
        RECT 289.250 88.230 289.710 88.460 ;
        RECT 289.960 88.025 290.930 88.665 ;
        RECT 291.180 88.230 291.640 88.460 ;
        RECT 291.890 88.025 293.385 88.665 ;
        RECT 293.640 88.310 294.100 88.540 ;
        RECT 295.570 88.310 296.030 88.540 ;
        RECT 287.870 86.525 289.200 88.025 ;
        RECT 289.760 86.525 291.130 88.025 ;
        RECT 291.690 86.525 293.385 88.025 ;
        RECT 296.650 87.700 297.520 88.700 ;
        RECT 287.870 85.885 289.000 86.525 ;
        RECT 289.250 86.090 289.710 86.320 ;
        RECT 289.960 85.885 290.930 86.525 ;
        RECT 291.180 86.090 291.640 86.320 ;
        RECT 291.890 85.885 293.385 86.525 ;
        RECT 287.870 84.385 289.200 85.885 ;
        RECT 289.760 84.385 291.130 85.885 ;
        RECT 291.690 85.615 293.385 85.885 ;
        RECT 291.690 84.385 293.390 85.615 ;
        RECT 287.870 83.290 288.630 84.385 ;
        RECT 289.250 83.950 289.710 84.180 ;
        RECT 291.180 83.950 291.640 84.180 ;
        RECT 287.870 77.540 288.250 83.290 ;
        RECT 284.870 76.485 285.380 77.085 ;
        RECT 287.330 76.485 287.840 77.085 ;
        RECT 291.890 76.485 293.390 84.385 ;
        RECT 297.030 75.450 297.520 87.700 ;
        RECT 298.610 82.095 298.970 82.515 ;
        RECT 298.560 78.770 298.920 79.190 ;
        RECT 298.485 77.850 298.845 78.270 ;
        RECT 299.525 77.450 299.825 79.180 ;
        RECT 298.565 75.550 298.925 75.970 ;
        RECT 300.360 75.450 300.850 95.450 ;
        RECT 301.385 90.790 301.685 97.450 ;
        RECT 302.265 92.825 302.565 96.450 ;
        RECT 303.020 92.155 303.320 101.450 ;
        RECT 304.880 100.850 305.380 109.400 ;
        RECT 305.880 101.850 306.380 103.100 ;
        RECT 305.290 99.850 305.800 100.450 ;
        RECT 307.750 99.850 308.260 100.450 ;
        RECT 303.020 91.655 303.420 92.155 ;
        RECT 302.255 90.780 302.615 91.200 ;
        RECT 302.235 83.115 302.595 83.535 ;
        RECT 301.385 77.450 301.685 79.180 ;
        RECT 302.320 78.780 302.620 79.180 ;
        RECT 302.375 77.850 302.735 78.270 ;
        RECT 303.070 77.860 303.370 82.505 ;
        RECT 302.370 76.950 302.730 77.370 ;
        RECT 302.400 75.560 302.700 76.950 ;
        RECT 303.690 76.890 304.180 94.450 ;
        RECT 304.880 77.535 305.260 94.450 ;
        RECT 305.460 92.345 305.630 99.850 ;
        RECT 305.880 93.395 306.340 93.445 ;
        RECT 305.860 92.505 306.360 93.395 ;
        RECT 306.590 92.345 306.760 93.395 ;
        RECT 305.460 91.845 305.830 92.345 ;
        RECT 306.390 91.845 306.760 92.345 ;
        RECT 305.460 91.295 305.630 91.845 ;
        RECT 305.880 91.455 306.340 91.685 ;
        RECT 306.590 91.295 306.760 91.845 ;
        RECT 305.460 90.795 305.830 91.295 ;
        RECT 306.390 90.795 306.760 91.295 ;
        RECT 305.460 90.245 305.630 90.795 ;
        RECT 305.880 90.405 306.340 90.635 ;
        RECT 306.590 90.245 306.760 90.795 ;
        RECT 305.460 89.745 305.830 90.245 ;
        RECT 306.390 89.745 306.760 90.245 ;
        RECT 305.460 89.195 305.630 89.745 ;
        RECT 305.880 89.355 306.340 89.585 ;
        RECT 306.590 89.195 306.760 89.745 ;
        RECT 305.460 88.695 305.830 89.195 ;
        RECT 306.390 88.695 306.760 89.195 ;
        RECT 305.460 87.730 305.630 88.695 ;
        RECT 305.880 88.305 306.340 88.535 ;
        RECT 306.590 87.730 306.760 88.695 ;
        RECT 305.460 87.560 306.760 87.730 ;
        RECT 305.460 86.550 305.630 87.560 ;
        RECT 305.880 86.755 306.340 86.985 ;
        RECT 306.590 86.550 306.760 87.560 ;
        RECT 305.460 85.050 305.830 86.550 ;
        RECT 306.390 85.050 306.760 86.550 ;
        RECT 305.460 84.410 305.630 85.050 ;
        RECT 305.880 84.615 306.340 84.845 ;
        RECT 306.590 84.410 306.760 85.050 ;
        RECT 305.460 82.910 305.830 84.410 ;
        RECT 306.390 82.910 306.760 84.410 ;
        RECT 305.460 82.270 305.630 82.910 ;
        RECT 305.880 82.475 306.340 82.705 ;
        RECT 306.590 82.270 306.760 82.910 ;
        RECT 305.460 80.770 305.830 82.270 ;
        RECT 306.390 80.770 306.760 82.270 ;
        RECT 305.460 80.130 305.630 80.770 ;
        RECT 305.880 80.335 306.340 80.565 ;
        RECT 306.590 80.130 306.760 80.770 ;
        RECT 305.460 78.630 305.830 80.130 ;
        RECT 306.390 78.630 306.760 80.130 ;
        RECT 305.860 77.535 306.360 78.425 ;
        RECT 306.590 77.535 306.760 78.630 ;
        RECT 306.960 77.535 307.720 95.450 ;
        RECT 307.920 92.300 308.090 99.850 ;
        RECT 308.340 93.395 308.800 99.450 ;
        RECT 308.320 92.505 308.820 93.395 ;
        RECT 307.920 90.800 308.290 92.300 ;
        RECT 308.850 90.800 309.220 92.300 ;
        RECT 307.920 90.160 308.090 90.800 ;
        RECT 308.340 90.365 308.800 90.595 ;
        RECT 309.050 90.160 309.220 90.800 ;
        RECT 307.920 88.660 308.290 90.160 ;
        RECT 308.850 88.660 309.220 90.160 ;
        RECT 307.920 88.020 308.090 88.660 ;
        RECT 308.340 88.225 308.800 88.455 ;
        RECT 309.050 88.020 309.220 88.660 ;
        RECT 307.920 86.520 308.290 88.020 ;
        RECT 308.850 86.520 309.220 88.020 ;
        RECT 307.920 85.880 308.090 86.520 ;
        RECT 308.340 86.085 308.800 86.315 ;
        RECT 309.050 85.880 309.220 86.520 ;
        RECT 307.920 84.380 308.290 85.880 ;
        RECT 308.850 84.380 309.220 85.880 ;
        RECT 307.920 82.235 308.090 84.380 ;
        RECT 308.340 83.945 308.800 84.175 ;
        RECT 308.340 82.395 308.800 82.625 ;
        RECT 309.050 82.235 309.220 84.380 ;
        RECT 307.920 81.735 308.290 82.235 ;
        RECT 308.850 81.735 309.220 82.235 ;
        RECT 307.920 81.185 308.090 81.735 ;
        RECT 308.340 81.345 308.800 81.575 ;
        RECT 309.050 81.185 309.220 81.735 ;
        RECT 307.920 80.685 308.290 81.185 ;
        RECT 308.850 80.685 309.220 81.185 ;
        RECT 307.920 80.135 308.090 80.685 ;
        RECT 308.340 80.295 308.800 80.525 ;
        RECT 309.050 80.135 309.220 80.685 ;
        RECT 307.920 79.635 308.290 80.135 ;
        RECT 308.850 79.635 309.220 80.135 ;
        RECT 307.920 79.085 308.090 79.635 ;
        RECT 308.340 79.245 308.800 79.475 ;
        RECT 309.050 79.085 309.220 79.635 ;
        RECT 307.920 78.585 308.290 79.085 ;
        RECT 308.850 78.585 309.220 79.085 ;
        RECT 307.920 77.535 308.090 78.585 ;
        RECT 308.320 77.535 308.820 78.425 ;
        RECT 305.880 77.485 306.340 77.535 ;
        RECT 308.340 77.485 308.800 77.535 ;
        RECT 309.050 77.085 309.220 78.585 ;
        RECT 309.420 77.540 310.180 94.450 ;
        RECT 310.800 93.400 311.260 93.445 ;
        RECT 310.380 92.350 310.550 93.400 ;
        RECT 310.780 92.510 311.280 93.400 ;
        RECT 311.510 92.350 311.680 93.400 ;
        RECT 310.380 91.850 310.750 92.350 ;
        RECT 311.310 91.850 311.680 92.350 ;
        RECT 310.380 91.300 310.550 91.850 ;
        RECT 310.800 91.460 311.260 91.690 ;
        RECT 311.510 91.300 311.680 91.850 ;
        RECT 310.380 90.800 310.750 91.300 ;
        RECT 311.310 90.800 311.680 91.300 ;
        RECT 310.380 90.250 310.550 90.800 ;
        RECT 310.800 90.410 311.260 90.640 ;
        RECT 311.510 90.250 311.680 90.800 ;
        RECT 310.380 89.750 310.750 90.250 ;
        RECT 311.310 89.750 311.680 90.250 ;
        RECT 310.380 89.200 310.550 89.750 ;
        RECT 310.800 89.360 311.260 89.590 ;
        RECT 311.510 89.200 311.680 89.750 ;
        RECT 310.380 88.700 310.750 89.200 ;
        RECT 311.310 88.700 311.680 89.200 ;
        RECT 310.380 87.735 310.550 88.700 ;
        RECT 310.800 88.310 311.260 88.540 ;
        RECT 311.510 87.735 311.680 88.700 ;
        RECT 310.380 87.565 311.680 87.735 ;
        RECT 310.380 86.555 310.550 87.565 ;
        RECT 310.800 86.760 311.260 86.990 ;
        RECT 311.510 86.555 311.680 87.565 ;
        RECT 310.380 85.055 310.750 86.555 ;
        RECT 311.310 85.055 311.680 86.555 ;
        RECT 310.380 84.415 310.550 85.055 ;
        RECT 310.800 84.620 311.260 84.850 ;
        RECT 311.510 84.415 311.680 85.055 ;
        RECT 310.380 82.915 310.750 84.415 ;
        RECT 311.310 82.915 311.680 84.415 ;
        RECT 310.380 82.275 310.550 82.915 ;
        RECT 310.800 82.480 311.260 82.710 ;
        RECT 311.510 82.275 311.680 82.915 ;
        RECT 310.380 80.775 310.750 82.275 ;
        RECT 311.310 80.775 311.680 82.275 ;
        RECT 310.380 80.135 310.550 80.775 ;
        RECT 310.800 80.340 311.260 80.570 ;
        RECT 311.510 80.135 311.680 80.775 ;
        RECT 310.380 78.635 310.750 80.135 ;
        RECT 311.310 78.635 311.680 80.135 ;
        RECT 310.780 77.540 311.280 78.430 ;
        RECT 309.420 77.535 309.800 77.540 ;
        RECT 310.800 77.485 311.260 77.540 ;
        RECT 311.510 77.085 311.680 78.635 ;
        RECT 311.880 92.305 312.640 134.995 ;
        RECT 315.900 134.950 317.600 134.995 ;
        RECT 318.160 134.950 319.530 135.450 ;
        RECT 320.090 134.950 321.530 135.450 ;
        RECT 313.260 134.785 313.720 134.790 ;
        RECT 313.240 124.850 313.740 134.785 ;
        RECT 315.170 129.850 315.670 134.790 ;
        RECT 315.900 133.900 317.450 134.950 ;
        RECT 317.630 130.850 318.130 134.790 ;
        RECT 319.560 134.200 320.060 134.790 ;
        RECT 313.240 92.515 313.740 102.450 ;
        RECT 313.260 92.510 313.720 92.515 ;
        RECT 315.170 92.510 315.670 97.450 ;
        RECT 315.900 92.350 317.450 93.400 ;
        RECT 317.630 92.510 318.130 96.450 ;
        RECT 319.560 92.510 320.060 93.100 ;
        RECT 320.660 92.350 321.530 134.950 ;
        RECT 321.880 127.850 322.180 136.510 ;
        RECT 322.605 136.100 322.965 136.520 ;
        RECT 322.655 128.850 322.955 134.475 ;
        RECT 324.370 131.850 324.860 151.850 ;
        RECT 326.410 150.350 326.710 151.740 ;
        RECT 326.380 149.930 326.740 150.350 ;
        RECT 325.395 148.120 325.695 149.850 ;
        RECT 326.385 149.030 326.745 149.450 ;
        RECT 326.330 148.120 326.630 148.520 ;
        RECT 327.080 144.795 327.380 149.440 ;
        RECT 326.245 143.765 326.605 144.185 ;
        RECT 325.395 129.850 325.695 136.510 ;
        RECT 326.265 136.100 326.625 136.520 ;
        RECT 327.030 135.145 327.430 135.645 ;
        RECT 326.275 130.850 326.575 134.475 ;
        RECT 327.030 125.850 327.330 135.145 ;
        RECT 327.700 132.850 328.190 150.410 ;
        RECT 315.900 92.305 317.600 92.350 ;
        RECT 311.880 90.805 313.210 92.305 ;
        RECT 313.770 90.805 315.140 92.305 ;
        RECT 315.700 91.850 317.600 92.305 ;
        RECT 318.160 91.850 319.530 92.350 ;
        RECT 320.090 91.850 321.530 92.350 ;
        RECT 315.700 91.300 317.450 91.850 ;
        RECT 317.650 91.460 318.110 91.690 ;
        RECT 318.360 91.300 319.330 91.850 ;
        RECT 319.580 91.460 320.040 91.690 ;
        RECT 320.290 91.300 321.530 91.850 ;
        RECT 315.700 90.805 317.600 91.300 ;
        RECT 311.880 90.165 313.010 90.805 ;
        RECT 313.260 90.370 313.720 90.600 ;
        RECT 313.970 90.165 314.940 90.805 ;
        RECT 315.900 90.800 317.600 90.805 ;
        RECT 318.160 90.800 319.530 91.300 ;
        RECT 320.090 90.800 321.530 91.300 ;
        RECT 315.190 90.370 315.650 90.600 ;
        RECT 315.900 90.250 317.450 90.800 ;
        RECT 317.650 90.410 318.110 90.640 ;
        RECT 318.360 90.250 319.330 90.800 ;
        RECT 319.580 90.410 320.040 90.640 ;
        RECT 320.290 90.250 321.530 90.800 ;
        RECT 321.880 90.790 322.180 99.450 ;
        RECT 322.655 92.825 322.955 98.450 ;
        RECT 322.605 90.780 322.965 91.200 ;
        RECT 315.900 90.165 317.600 90.250 ;
        RECT 311.880 88.665 313.210 90.165 ;
        RECT 313.770 88.665 315.140 90.165 ;
        RECT 315.700 89.750 317.600 90.165 ;
        RECT 318.160 89.750 319.530 90.250 ;
        RECT 320.090 89.750 321.530 90.250 ;
        RECT 315.700 89.200 317.450 89.750 ;
        RECT 317.650 89.360 318.110 89.590 ;
        RECT 318.360 89.200 319.330 89.750 ;
        RECT 319.580 89.360 320.040 89.590 ;
        RECT 320.290 89.200 321.530 89.750 ;
        RECT 315.700 88.700 317.600 89.200 ;
        RECT 318.160 88.700 319.530 89.200 ;
        RECT 320.090 88.700 321.530 89.200 ;
        RECT 315.700 88.665 317.450 88.700 ;
        RECT 311.880 88.025 313.010 88.665 ;
        RECT 313.260 88.230 313.720 88.460 ;
        RECT 313.970 88.025 314.940 88.665 ;
        RECT 315.190 88.230 315.650 88.460 ;
        RECT 315.900 88.025 317.450 88.665 ;
        RECT 317.650 88.310 318.110 88.540 ;
        RECT 319.580 88.310 320.040 88.540 ;
        RECT 311.880 86.525 313.210 88.025 ;
        RECT 313.770 86.525 315.140 88.025 ;
        RECT 315.700 86.525 317.450 88.025 ;
        RECT 320.660 87.700 321.530 88.700 ;
        RECT 311.880 85.885 313.010 86.525 ;
        RECT 313.260 86.090 313.720 86.320 ;
        RECT 313.970 85.885 314.940 86.525 ;
        RECT 315.190 86.090 315.650 86.320 ;
        RECT 315.900 85.885 317.450 86.525 ;
        RECT 311.880 84.385 313.210 85.885 ;
        RECT 313.770 84.385 315.140 85.885 ;
        RECT 315.700 85.445 317.450 85.885 ;
        RECT 315.700 84.385 317.400 85.445 ;
        RECT 311.880 83.290 312.640 84.385 ;
        RECT 313.260 83.950 313.720 84.180 ;
        RECT 315.190 83.950 315.650 84.180 ;
        RECT 311.880 77.540 312.260 83.290 ;
        RECT 308.880 76.485 309.390 77.085 ;
        RECT 311.340 76.485 311.850 77.085 ;
        RECT 315.900 76.485 317.400 84.385 ;
        RECT 321.040 75.450 321.530 87.700 ;
        RECT 322.620 82.095 322.980 82.515 ;
        RECT 322.570 78.770 322.930 79.190 ;
        RECT 322.495 77.850 322.855 78.270 ;
        RECT 323.535 77.450 323.835 79.180 ;
        RECT 322.575 75.550 322.935 75.970 ;
        RECT 324.370 75.450 324.860 95.450 ;
        RECT 325.395 90.790 325.695 97.450 ;
        RECT 326.275 92.825 326.575 96.450 ;
        RECT 327.030 92.155 327.330 101.450 ;
        RECT 327.030 91.655 327.430 92.155 ;
        RECT 326.265 90.780 326.625 91.200 ;
        RECT 326.245 83.115 326.605 83.535 ;
        RECT 325.395 77.450 325.695 79.180 ;
        RECT 326.330 78.780 326.630 79.180 ;
        RECT 326.385 77.850 326.745 78.270 ;
        RECT 327.080 77.860 327.380 82.505 ;
        RECT 326.380 76.950 326.740 77.370 ;
        RECT 326.410 75.560 326.710 76.950 ;
        RECT 327.700 76.890 328.190 94.450 ;
        RECT 111.750 73.460 330.185 73.980 ;
        RECT 112.800 72.420 330.185 72.940 ;
        RECT 83.115 71.100 83.615 71.500 ;
        RECT 112.800 71.380 330.185 71.900 ;
        RECT 53.930 70.705 54.310 70.760 ;
        RECT 26.090 70.360 26.470 70.640 ;
        RECT 53.930 70.505 83.075 70.705 ;
        RECT 53.930 70.450 54.310 70.505 ;
        RECT 26.170 70.005 26.370 70.360 ;
        RECT 26.170 69.805 82.015 70.005 ;
        RECT 71.475 41.155 71.955 69.395 ;
        RECT 72.435 42.115 72.915 68.435 ;
        RECT 80.315 67.235 80.795 69.395 ;
        RECT 73.395 52.965 73.875 54.345 ;
        RECT 74.460 53.755 74.950 59.555 ;
        RECT 76.230 58.260 76.490 59.605 ;
        RECT 76.755 58.260 77.015 59.085 ;
        RECT 76.160 57.930 76.490 58.260 ;
        RECT 76.685 57.930 77.015 58.260 ;
        RECT 75.260 57.490 76.260 57.720 ;
        RECT 77.000 57.490 80.000 57.720 ;
        RECT 75.260 57.050 76.260 57.280 ;
        RECT 77.000 57.050 80.000 57.280 ;
        RECT 75.260 56.610 76.260 56.840 ;
        RECT 77.000 56.610 80.000 56.840 ;
        RECT 77.000 56.170 80.000 56.400 ;
        RECT 75.940 55.180 76.270 55.510 ;
        RECT 76.685 55.180 77.015 55.510 ;
        RECT 76.010 54.275 76.270 55.180 ;
        RECT 76.755 53.340 77.015 55.180 ;
        RECT 80.310 53.805 80.800 67.235 ;
        RECT 81.815 67.070 82.015 69.805 ;
        RECT 81.785 66.750 82.045 67.070 ;
        RECT 81.085 58.725 81.385 64.220 ;
        RECT 81.685 59.245 81.985 65.030 ;
        RECT 82.160 64.620 82.520 65.040 ;
        RECT 82.240 63.810 82.600 64.230 ;
        RECT 82.370 62.720 82.630 62.780 ;
        RECT 82.875 62.720 83.075 70.505 ;
        RECT 83.270 62.750 83.470 71.100 ;
        RECT 93.635 69.900 103.495 70.400 ;
        RECT 112.800 70.340 330.185 70.860 ;
        RECT 82.370 62.520 83.075 62.720 ;
        RECT 82.370 62.460 82.630 62.520 ;
        RECT 82.305 61.550 82.665 61.970 ;
        RECT 82.305 60.980 82.665 61.400 ;
        RECT 82.875 61.310 83.075 62.520 ;
        RECT 83.240 62.430 83.500 62.750 ;
        RECT 82.845 60.990 83.105 61.310 ;
        RECT 82.370 60.430 82.630 60.490 ;
        RECT 83.270 60.430 83.470 62.430 ;
        RECT 82.370 60.230 83.470 60.430 ;
        RECT 82.370 60.170 82.630 60.230 ;
        RECT 83.640 60.035 84.130 67.235 ;
        RECT 83.650 59.985 84.130 60.035 ;
        RECT 84.165 58.260 84.425 59.605 ;
        RECT 84.690 58.260 84.950 59.085 ;
        RECT 84.095 57.930 84.425 58.260 ;
        RECT 84.620 57.930 84.950 58.260 ;
        RECT 81.110 57.490 84.110 57.720 ;
        RECT 84.850 57.490 85.850 57.720 ;
        RECT 81.110 57.050 84.110 57.280 ;
        RECT 84.850 57.050 85.850 57.280 ;
        RECT 81.110 56.610 84.110 56.840 ;
        RECT 84.850 56.610 85.850 56.840 ;
        RECT 81.110 56.170 84.110 56.400 ;
        RECT 84.095 55.180 84.425 55.510 ;
        RECT 84.840 55.180 85.170 55.510 ;
        RECT 73.395 52.805 75.630 52.965 ;
        RECT 73.395 44.755 73.875 52.805 ;
        RECT 75.140 50.565 75.630 52.805 ;
        RECT 76.755 52.820 77.070 53.340 ;
        RECT 80.315 52.965 80.795 53.805 ;
        RECT 84.165 53.340 84.425 55.180 ;
        RECT 84.910 53.755 85.170 55.180 ;
        RECT 86.160 53.755 86.650 60.565 ;
        RECT 76.755 52.750 77.015 52.820 ;
        RECT 78.470 52.810 82.640 52.965 ;
        RECT 84.040 52.820 84.425 53.340 ;
        RECT 87.235 52.965 87.715 54.345 ;
        RECT 76.735 51.590 77.065 52.020 ;
        RECT 78.470 50.565 78.960 52.810 ;
        RECT 74.485 49.385 75.485 49.615 ;
        RECT 76.325 49.385 79.325 49.615 ;
        RECT 75.890 48.585 76.120 49.125 ;
        RECT 74.485 48.095 75.485 48.325 ;
        RECT 76.325 48.095 79.325 48.325 ;
        RECT 74.095 47.295 74.325 47.835 ;
        RECT 79.530 47.295 80.100 47.835 ;
        RECT 74.125 44.475 74.295 47.295 ;
        RECT 74.485 46.805 75.485 47.035 ;
        RECT 76.325 46.805 79.325 47.035 ;
        RECT 79.515 45.955 79.775 46.595 ;
        RECT 74.485 45.515 75.485 45.745 ;
        RECT 76.325 45.515 79.325 45.745 ;
        RECT 74.080 44.115 74.340 44.475 ;
        RECT 79.560 43.435 79.730 45.955 ;
        RECT 79.930 43.955 80.100 47.295 ;
        RECT 79.885 43.595 80.145 43.955 ;
        RECT 79.515 43.075 79.775 43.435 ;
        RECT 79.560 41.205 79.730 43.075 ;
        RECT 63.505 39.920 64.125 40.440 ;
        RECT 44.610 39.070 56.190 39.560 ;
        RECT 48.395 37.905 55.075 38.135 ;
        RECT 42.325 37.585 42.705 37.650 ;
        RECT 45.525 37.585 45.815 37.615 ;
        RECT 16.805 37.415 45.815 37.585 ;
        RECT 48.000 37.535 54.665 37.765 ;
        RECT 42.325 37.350 42.705 37.415 ;
        RECT 45.525 37.385 45.815 37.415 ;
        RECT 54.835 37.320 55.940 37.580 ;
        RECT 55.580 36.705 55.940 36.965 ;
        RECT 44.610 36.225 55.650 36.230 ;
        RECT 63.555 36.225 64.075 39.920 ;
        RECT 79.930 36.225 80.100 43.595 ;
        RECT 80.315 41.155 80.795 52.810 ;
        RECT 82.150 50.565 82.640 52.810 ;
        RECT 84.165 52.750 84.425 52.820 ;
        RECT 85.480 52.805 87.715 52.965 ;
        RECT 84.045 51.590 84.375 52.020 ;
        RECT 85.480 50.565 85.970 52.805 ;
        RECT 81.785 49.385 84.785 49.615 ;
        RECT 85.625 49.385 86.625 49.615 ;
        RECT 84.990 48.585 85.220 49.125 ;
        RECT 81.785 48.095 84.785 48.325 ;
        RECT 85.625 48.095 86.625 48.325 ;
        RECT 81.010 47.295 81.580 47.835 ;
        RECT 86.785 47.295 87.015 47.835 ;
        RECT 81.010 44.475 81.180 47.295 ;
        RECT 81.785 46.805 84.785 47.035 ;
        RECT 85.625 46.805 86.625 47.035 ;
        RECT 81.335 45.955 81.595 46.595 ;
        RECT 80.965 44.115 81.225 44.475 ;
        RECT 3.955 35.745 58.580 36.225 ;
        RECT 44.610 35.740 55.650 35.745 ;
        RECT 51.590 34.070 52.380 35.740 ;
        RECT 51.480 33.810 53.420 34.070 ;
        RECT 51.050 33.500 51.340 33.530 ;
        RECT 52.630 33.500 52.920 33.530 ;
        RECT 57.260 33.500 57.620 33.545 ;
        RECT 51.050 33.330 57.620 33.500 ;
        RECT 51.050 33.300 51.340 33.330 ;
        RECT 52.630 33.300 52.920 33.330 ;
        RECT 57.260 33.285 57.620 33.330 ;
        RECT 50.550 31.140 51.090 33.140 ;
        RECT 51.300 31.140 51.840 33.140 ;
        RECT 52.130 25.640 52.670 33.140 ;
        RECT 52.880 25.640 53.420 33.140 ;
        RECT 53.710 25.950 54.250 29.950 ;
        RECT 54.460 28.080 54.690 29.950 ;
        RECT 58.050 28.555 58.530 35.745 ;
        RECT 62.200 34.945 80.100 36.225 ;
        RECT 81.010 36.225 81.180 44.115 ;
        RECT 81.380 43.435 81.550 45.955 ;
        RECT 81.785 45.515 84.785 45.745 ;
        RECT 85.625 45.515 86.625 45.745 ;
        RECT 86.815 43.955 86.985 47.295 ;
        RECT 87.235 44.755 87.715 52.805 ;
        RECT 86.770 43.595 87.030 43.955 ;
        RECT 81.335 43.075 81.595 43.435 ;
        RECT 88.195 42.115 88.675 68.435 ;
        RECT 89.155 41.155 89.635 69.395 ;
        RECT 102.995 44.000 103.495 69.900 ;
        RECT 112.800 69.300 330.185 69.820 ;
        RECT 112.800 68.260 330.185 68.780 ;
        RECT 112.800 67.220 330.185 67.740 ;
        RECT 112.800 66.180 330.185 66.700 ;
        RECT 112.800 65.140 330.185 65.660 ;
        RECT 112.800 64.100 330.185 64.620 ;
        RECT 241.475 55.620 249.115 56.100 ;
        RECT 241.475 44.820 249.115 45.300 ;
        RECT 102.995 43.500 119.440 44.000 ;
        RECT 97.145 41.250 97.765 41.770 ;
        RECT 97.195 36.225 97.715 41.250 ;
        RECT 104.930 39.070 116.510 39.560 ;
        RECT 106.045 37.905 112.725 38.135 ;
        RECT 106.455 37.535 113.120 37.765 ;
        RECT 115.305 37.585 115.595 37.615 ;
        RECT 118.940 37.585 119.440 43.500 ;
        RECT 241.475 37.620 249.115 38.100 ;
        RECT 104.160 37.225 106.285 37.485 ;
        RECT 115.305 37.415 144.315 37.585 ;
        RECT 115.305 37.385 115.595 37.415 ;
        RECT 248.535 36.360 252.535 36.840 ;
        RECT 105.470 36.225 116.510 36.230 ;
        RECT 81.010 34.945 98.920 36.225 ;
        RECT 102.540 35.745 144.315 36.225 ;
        RECT 62.200 34.045 63.480 34.945 ;
        RECT 64.760 34.045 66.040 34.945 ;
        RECT 67.320 34.045 68.600 34.945 ;
        RECT 69.880 34.045 71.160 34.945 ;
        RECT 72.440 34.045 73.720 34.945 ;
        RECT 75.000 34.045 76.280 34.945 ;
        RECT 84.840 34.045 86.120 34.945 ;
        RECT 87.400 34.045 88.680 34.945 ;
        RECT 89.960 34.045 91.240 34.945 ;
        RECT 92.520 34.045 93.800 34.945 ;
        RECT 95.080 34.045 96.360 34.945 ;
        RECT 97.640 34.045 98.920 34.945 ;
        RECT 59.640 33.105 79.520 34.045 ;
        RECT 58.730 29.430 58.990 32.950 ;
        RECT 59.160 32.590 59.420 32.950 ;
        RECT 59.580 32.875 79.580 33.105 ;
        RECT 59.640 32.665 79.520 32.875 ;
        RECT 59.580 32.435 79.580 32.665 ;
        RECT 59.640 31.525 79.520 32.435 ;
        RECT 59.160 31.010 59.420 31.370 ;
        RECT 59.580 31.295 79.580 31.525 ;
        RECT 59.580 30.855 79.580 31.085 ;
        RECT 59.640 29.945 79.520 30.855 ;
        RECT 59.160 29.430 59.420 29.790 ;
        RECT 59.580 29.715 79.580 29.945 ;
        RECT 59.640 29.505 79.520 29.715 ;
        RECT 59.580 29.275 79.580 29.505 ;
        RECT 59.640 28.335 79.520 29.275 ;
        RECT 80.320 28.555 80.800 33.825 ;
        RECT 81.600 33.105 101.480 34.045 ;
        RECT 81.540 32.875 101.540 33.105 ;
        RECT 81.600 32.665 101.480 32.875 ;
        RECT 81.540 32.435 101.540 32.665 ;
        RECT 101.700 32.590 101.960 32.950 ;
        RECT 81.600 31.525 101.480 32.435 ;
        RECT 81.540 31.295 101.540 31.525 ;
        RECT 81.540 30.855 101.540 31.085 ;
        RECT 101.700 31.010 101.960 31.370 ;
        RECT 81.600 29.945 101.480 30.855 ;
        RECT 81.540 29.715 101.540 29.945 ;
        RECT 81.600 29.505 101.480 29.715 ;
        RECT 81.540 29.275 101.540 29.505 ;
        RECT 101.700 29.430 101.960 29.790 ;
        RECT 102.130 29.430 102.390 32.950 ;
        RECT 81.600 28.335 101.480 29.275 ;
        RECT 102.590 28.555 103.070 35.745 ;
        RECT 105.470 35.740 116.510 35.745 ;
        RECT 108.740 34.070 109.530 35.740 ;
        RECT 241.475 34.560 253.335 35.040 ;
        RECT 107.700 33.810 109.640 34.070 ;
        RECT 103.500 33.500 103.860 33.545 ;
        RECT 108.200 33.500 108.490 33.530 ;
        RECT 109.780 33.500 110.070 33.530 ;
        RECT 103.500 33.330 110.070 33.500 ;
        RECT 103.500 33.285 103.860 33.330 ;
        RECT 108.200 33.300 108.490 33.330 ;
        RECT 109.780 33.300 110.070 33.330 ;
        RECT 67.320 28.080 68.600 28.335 ;
        RECT 54.460 27.820 68.600 28.080 ;
        RECT 69.880 27.820 71.160 28.335 ;
        RECT 72.440 27.820 73.720 28.335 ;
        RECT 75.000 27.820 76.280 28.335 ;
        RECT 84.840 27.820 86.120 28.335 ;
        RECT 87.400 27.820 88.680 28.335 ;
        RECT 89.960 27.820 91.240 28.335 ;
        RECT 92.520 28.080 93.800 28.335 ;
        RECT 106.430 28.080 106.660 29.950 ;
        RECT 92.520 27.820 106.660 28.080 ;
        RECT 54.460 25.950 54.690 27.820 ;
        RECT 67.270 26.540 76.330 27.820 ;
        RECT 84.790 26.540 93.850 27.820 ;
        RECT 106.430 25.950 106.660 27.820 ;
        RECT 106.870 25.950 107.410 29.950 ;
        RECT 54.175 25.530 54.535 25.790 ;
        RECT 106.585 25.530 106.945 25.790 ;
        RECT 107.700 25.640 108.240 33.140 ;
        RECT 108.450 25.640 108.990 33.140 ;
        RECT 109.280 31.140 109.820 33.140 ;
        RECT 110.030 31.140 110.570 33.140 ;
        RECT 241.475 32.760 252.535 33.240 ;
        RECT 248.535 30.960 254.135 31.440 ;
        RECT 241.475 26.820 249.115 27.300 ;
        RECT 50.550 25.080 54.070 25.340 ;
        RECT 107.050 25.080 110.570 25.340 ;
        RECT 53.060 24.690 57.620 24.800 ;
        RECT 50.550 17.190 51.090 17.690 ;
        RECT 51.300 17.190 51.840 17.690 ;
        RECT 52.130 17.190 52.670 24.690 ;
        RECT 52.880 24.540 57.620 24.690 ;
        RECT 103.500 24.690 108.060 24.800 ;
        RECT 103.500 24.540 108.240 24.690 ;
        RECT 52.880 17.450 53.420 24.540 ;
        RECT 53.710 20.380 54.250 24.380 ;
        RECT 54.460 20.380 55.000 24.380 ;
        RECT 106.120 20.380 106.660 24.380 ;
        RECT 106.870 20.380 107.410 24.380 ;
        RECT 107.700 17.450 108.240 24.540 ;
        RECT 52.880 17.190 70.530 17.450 ;
        RECT 90.590 17.190 108.240 17.450 ;
        RECT 108.450 17.190 108.990 24.690 ;
        RECT 241.475 23.220 249.115 23.700 ;
        RECT 109.280 17.190 109.820 17.690 ;
        RECT 110.030 17.190 110.570 17.690 ;
        RECT 51.015 16.770 51.375 17.030 ;
        RECT 52.595 16.770 52.955 17.030 ;
        RECT 108.165 16.770 108.525 17.030 ;
        RECT 109.745 16.770 110.105 17.030 ;
        RECT 49.000 16.050 49.620 16.570 ;
        RECT 51.480 16.310 70.065 16.570 ;
        RECT 91.055 16.310 109.640 16.570 ;
        RECT 111.500 16.050 112.120 16.570 ;
        RECT 49.000 15.790 69.275 16.050 ;
        RECT 91.845 15.790 112.120 16.050 ;
        RECT 49.000 15.270 49.620 15.790 ;
        RECT 51.015 15.250 51.375 15.510 ;
        RECT 51.050 15.245 51.340 15.250 ;
        RECT 51.480 15.040 51.840 15.045 ;
        RECT 50.860 13.930 51.090 15.040 ;
        RECT 51.300 14.295 51.840 15.040 ;
        RECT 51.300 14.290 51.530 14.295 ;
        RECT 50.740 13.700 51.650 13.930 ;
        RECT 50.800 13.290 51.590 13.700 ;
        RECT 50.800 13.030 52.955 13.290 ;
        RECT 50.800 10.660 51.590 13.030 ;
        RECT 67.660 11.400 68.200 15.400 ;
        RECT 68.410 15.040 68.640 15.400 ;
        RECT 69.705 15.245 70.065 15.505 ;
        RECT 91.055 15.245 91.415 15.505 ;
        RECT 92.480 15.040 92.710 15.400 ;
        RECT 68.410 13.040 69.780 15.040 ;
        RECT 69.990 13.040 70.530 15.040 ;
        RECT 90.590 13.040 91.130 15.040 ;
        RECT 91.340 13.040 92.710 15.040 ;
        RECT 68.410 11.400 68.640 13.040 ;
        RECT 92.480 11.400 92.710 13.040 ;
        RECT 92.920 11.400 93.460 15.400 ;
        RECT 109.745 15.250 110.105 15.510 ;
        RECT 111.500 15.270 112.120 15.790 ;
        RECT 109.780 15.245 110.070 15.250 ;
        RECT 109.280 15.040 109.640 15.045 ;
        RECT 109.280 14.295 109.820 15.040 ;
        RECT 109.590 14.290 109.820 14.295 ;
        RECT 110.030 13.930 110.260 15.040 ;
        RECT 109.470 13.700 110.380 13.930 ;
        RECT 109.530 13.290 110.320 13.700 ;
        RECT 108.165 13.030 110.320 13.290 ;
        RECT 67.660 10.660 68.020 11.400 ;
        RECT 68.160 10.935 70.530 11.195 ;
        RECT 90.590 10.935 92.960 11.195 ;
        RECT 50.800 10.300 68.020 10.660 ;
        RECT 93.100 10.660 93.460 11.400 ;
        RECT 109.530 10.660 110.320 13.030 ;
        RECT 241.475 12.420 249.115 12.900 ;
        RECT 93.100 10.300 110.320 10.660 ;
        RECT 50.800 6.155 51.590 10.300 ;
        RECT 109.530 6.155 110.320 10.300 ;
        RECT 0.950 5.675 144.315 6.155 ;
        RECT 134.530 -5.650 135.110 -5.170 ;
      LAYER met2 ;
        RECT 134.580 232.420 135.060 233.000 ;
        RECT 241.525 214.350 242.005 214.930 ;
        RECT 95.655 211.005 96.155 211.150 ;
        RECT 138.100 211.005 138.800 211.250 ;
        RECT 95.655 210.705 138.800 211.005 ;
        RECT 95.655 210.550 96.155 210.705 ;
        RECT 138.100 210.450 138.800 210.705 ;
        RECT 241.525 203.550 242.005 204.130 ;
        RECT 241.525 199.950 242.005 200.530 ;
        RECT 241.525 194.010 242.005 194.590 ;
        RECT 241.525 192.210 242.005 192.790 ;
        RECT 241.525 189.150 242.005 189.730 ;
        RECT 241.525 181.950 242.005 182.530 ;
        RECT 241.525 171.150 242.005 171.730 ;
        RECT 85.100 165.800 87.100 165.850 ;
        RECT 85.100 163.800 107.100 165.800 ;
        RECT 85.100 163.750 87.100 163.800 ;
        RECT 85.100 161.800 87.100 161.850 ;
        RECT 85.100 159.800 102.700 161.800 ;
        RECT 85.100 159.750 87.100 159.800 ;
        RECT 8.200 152.850 8.800 157.050 ;
        RECT 14.000 152.850 14.600 157.050 ;
        RECT 19.700 153.680 20.300 157.050 ;
        RECT 19.700 153.540 21.550 153.680 ;
        RECT 19.700 152.850 20.300 153.540 ;
        RECT 8.450 135.455 8.590 152.850 ;
        RECT 13.670 142.165 13.930 142.485 ;
        RECT 13.190 141.425 13.450 141.745 ;
        RECT 13.250 136.565 13.390 141.425 ;
        RECT 13.190 136.245 13.450 136.565 ;
        RECT 8.390 135.135 8.650 135.455 ;
        RECT 13.730 133.235 13.870 142.165 ;
        RECT 14.210 141.375 14.350 152.850 ;
        RECT 20.870 142.165 21.130 142.485 ;
        RECT 14.150 141.055 14.410 141.375 ;
        RECT 14.260 140.105 16.140 140.475 ;
        RECT 20.930 139.895 21.070 142.165 ;
        RECT 21.410 141.745 21.550 153.540 ;
        RECT 25.500 152.850 26.100 157.050 ;
        RECT 31.200 153.680 31.800 157.050 ;
        RECT 31.200 153.540 33.070 153.680 ;
        RECT 31.200 152.850 31.800 153.540 ;
        RECT 21.350 141.425 21.610 141.745 ;
        RECT 24.230 141.425 24.490 141.745 ;
        RECT 24.710 141.425 24.970 141.745 ;
        RECT 20.870 139.575 21.130 139.895 ;
        RECT 22.310 138.465 22.570 138.785 ;
        RECT 22.370 135.455 22.510 138.465 ;
        RECT 24.290 138.415 24.430 141.425 ;
        RECT 24.770 139.155 24.910 141.425 ;
        RECT 25.730 139.895 25.870 152.850 ;
        RECT 29.260 143.435 31.140 143.805 ;
        RECT 32.930 142.115 33.070 153.540 ;
        RECT 37.000 152.850 37.600 157.050 ;
        RECT 42.800 153.680 43.400 157.050 ;
        RECT 42.800 153.540 44.590 153.680 ;
        RECT 42.800 152.850 43.400 153.540 ;
        RECT 35.270 142.165 35.530 142.485 ;
        RECT 32.390 141.795 32.650 142.115 ;
        RECT 32.870 141.795 33.130 142.115 ;
        RECT 25.670 139.575 25.930 139.895 ;
        RECT 32.450 139.525 32.590 141.795 ;
        RECT 32.870 140.685 33.130 141.005 ;
        RECT 32.390 139.205 32.650 139.525 ;
        RECT 32.930 139.155 33.070 140.685 ;
        RECT 24.710 138.835 24.970 139.155 ;
        RECT 32.870 138.880 33.130 139.155 ;
        RECT 32.450 138.835 33.130 138.880 ;
        RECT 24.230 138.095 24.490 138.415 ;
        RECT 22.310 135.135 22.570 135.455 ;
        RECT 14.260 133.445 16.140 133.815 ;
        RECT 13.670 132.915 13.930 133.235 ;
        RECT 22.370 132.125 22.510 135.135 ;
        RECT 24.770 134.715 24.910 138.835 ;
        RECT 25.670 138.465 25.930 138.785 ;
        RECT 31.910 138.465 32.170 138.785 ;
        RECT 32.450 138.740 33.070 138.835 ;
        RECT 24.710 134.395 24.970 134.715 ;
        RECT 22.310 131.805 22.570 132.125 ;
        RECT 17.510 128.475 17.770 128.795 ;
        RECT 18.470 128.475 18.730 128.795 ;
        RECT 13.190 128.105 13.450 128.425 ;
        RECT 13.250 112.145 13.390 128.105 ;
        RECT 14.260 126.785 16.140 127.155 ;
        RECT 17.570 126.575 17.710 128.475 ;
        RECT 17.990 127.365 18.250 127.685 ;
        RECT 17.510 126.255 17.770 126.575 ;
        RECT 18.050 125.465 18.190 127.365 ;
        RECT 17.990 125.145 18.250 125.465 ;
        RECT 16.550 121.445 16.810 121.765 ;
        RECT 14.260 120.125 16.140 120.495 ;
        RECT 13.670 114.045 13.930 114.365 ;
        RECT 13.730 113.255 13.870 114.045 ;
        RECT 14.260 113.465 16.140 113.835 ;
        RECT 13.670 112.935 13.930 113.255 ;
        RECT 16.610 112.980 16.750 121.445 ;
        RECT 18.050 116.215 18.190 125.145 ;
        RECT 18.530 122.135 18.670 128.475 ;
        RECT 21.350 125.145 21.610 125.465 ;
        RECT 18.470 121.815 18.730 122.135 ;
        RECT 18.530 119.175 18.670 121.815 ;
        RECT 21.410 121.025 21.550 125.145 ;
        RECT 22.310 124.035 22.570 124.355 ;
        RECT 23.750 124.035 24.010 124.355 ;
        RECT 21.350 120.705 21.610 121.025 ;
        RECT 18.470 118.855 18.730 119.175 ;
        RECT 17.990 115.895 18.250 116.215 ;
        RECT 16.130 112.840 16.750 112.980 ;
        RECT 13.190 111.825 13.450 112.145 ;
        RECT 12.710 110.715 12.970 111.035 ;
        RECT 14.150 110.715 14.410 111.035 ;
        RECT 12.770 109.925 12.910 110.715 ;
        RECT 14.210 109.925 14.350 110.715 ;
        RECT 16.130 109.925 16.270 112.840 ;
        RECT 18.530 112.145 18.670 118.855 ;
        RECT 19.430 115.155 19.690 115.475 ;
        RECT 16.550 111.825 16.810 112.145 ;
        RECT 18.470 111.825 18.730 112.145 ;
        RECT 12.710 109.605 12.970 109.925 ;
        RECT 14.150 109.605 14.410 109.925 ;
        RECT 16.070 109.605 16.330 109.925 ;
        RECT 14.260 106.805 16.140 107.175 ;
        RECT 16.610 105.855 16.750 111.825 ;
        RECT 17.030 111.455 17.290 111.775 ;
        RECT 17.090 109.925 17.230 111.455 ;
        RECT 17.030 109.605 17.290 109.925 ;
        RECT 19.490 108.445 19.630 115.155 ;
        RECT 21.410 114.735 21.550 120.705 ;
        RECT 22.370 118.805 22.510 124.035 ;
        RECT 23.810 122.135 23.950 124.035 ;
        RECT 24.770 123.245 24.910 134.395 ;
        RECT 25.730 132.495 25.870 138.465 ;
        RECT 26.630 138.095 26.890 138.415 ;
        RECT 26.690 136.565 26.830 138.095 ;
        RECT 29.260 136.775 31.140 137.145 ;
        RECT 26.630 136.245 26.890 136.565 ;
        RECT 31.970 135.825 32.110 138.465 ;
        RECT 31.910 135.505 32.170 135.825 ;
        RECT 26.630 135.135 26.890 135.455 ;
        RECT 32.450 135.230 32.590 138.740 ;
        RECT 33.350 138.095 33.610 138.415 ;
        RECT 25.670 132.175 25.930 132.495 ;
        RECT 25.190 125.515 25.450 125.835 ;
        RECT 24.710 122.925 24.970 123.245 ;
        RECT 23.270 121.815 23.530 122.135 ;
        RECT 23.750 121.815 24.010 122.135 ;
        RECT 23.330 119.915 23.470 121.815 ;
        RECT 23.270 119.595 23.530 119.915 ;
        RECT 21.830 118.485 22.090 118.805 ;
        RECT 22.310 118.485 22.570 118.805 ;
        RECT 21.890 115.105 22.030 118.485 ;
        RECT 25.250 118.435 25.390 125.515 ;
        RECT 25.190 118.115 25.450 118.435 ;
        RECT 21.830 114.785 22.090 115.105 ;
        RECT 21.350 114.415 21.610 114.735 ;
        RECT 19.430 108.125 19.690 108.445 ;
        RECT 16.550 105.535 16.810 105.855 ;
        RECT 16.610 102.155 16.750 105.535 ;
        RECT 21.890 105.485 22.030 114.785 ;
        RECT 26.150 114.045 26.410 114.365 ;
        RECT 25.670 111.455 25.930 111.775 ;
        RECT 22.790 110.715 23.050 111.035 ;
        RECT 22.850 109.925 22.990 110.715 ;
        RECT 25.730 109.925 25.870 111.455 ;
        RECT 22.790 109.605 23.050 109.925 ;
        RECT 25.670 109.605 25.930 109.925 ;
        RECT 23.750 108.125 24.010 108.445 ;
        RECT 21.830 105.165 22.090 105.485 ;
        RECT 23.810 105.115 23.950 108.125 ;
        RECT 26.210 106.225 26.350 114.045 ;
        RECT 26.690 111.035 26.830 135.135 ;
        RECT 31.490 135.090 32.590 135.230 ;
        RECT 33.410 135.230 33.550 138.095 ;
        RECT 35.330 136.565 35.470 142.165 ;
        RECT 37.250 141.375 37.390 152.850 ;
        RECT 43.910 142.165 44.170 142.485 ;
        RECT 37.190 141.055 37.450 141.375 ;
        RECT 43.970 139.895 44.110 142.165 ;
        RECT 44.450 141.745 44.590 153.540 ;
        RECT 48.500 152.850 49.100 157.050 ;
        RECT 54.300 152.850 54.900 157.050 ;
        RECT 60.100 153.680 60.700 157.050 ;
        RECT 60.100 153.540 61.870 153.680 ;
        RECT 60.100 152.850 60.700 153.540 ;
        RECT 47.740 152.200 48.020 152.315 ;
        RECT 47.330 152.060 48.020 152.200 ;
        RECT 44.390 141.425 44.650 141.745 ;
        RECT 44.260 140.105 46.140 140.475 ;
        RECT 47.330 139.895 47.470 152.060 ;
        RECT 47.740 151.945 48.020 152.060 ;
        RECT 47.740 146.025 48.020 146.395 ;
        RECT 47.810 141.375 47.950 146.025 ;
        RECT 48.770 141.375 48.910 152.850 ;
        RECT 53.980 148.985 54.260 149.355 ;
        RECT 50.150 142.165 50.410 142.485 ;
        RECT 51.110 142.165 51.370 142.485 ;
        RECT 47.750 141.055 48.010 141.375 ;
        RECT 48.710 141.055 48.970 141.375 ;
        RECT 43.910 139.575 44.170 139.895 ;
        RECT 47.270 139.575 47.530 139.895 ;
        RECT 43.430 138.095 43.690 138.415 ;
        RECT 49.190 138.095 49.450 138.415 ;
        RECT 35.270 136.245 35.530 136.565 ;
        RECT 33.410 135.090 34.030 135.230 ;
        RECT 29.260 130.115 31.140 130.485 ;
        RECT 27.590 128.105 27.850 128.425 ;
        RECT 27.650 126.575 27.790 128.105 ;
        RECT 27.590 126.255 27.850 126.575 ;
        RECT 28.550 125.145 28.810 125.465 ;
        RECT 28.610 123.245 28.750 125.145 ;
        RECT 29.260 123.455 31.140 123.825 ;
        RECT 28.550 122.925 28.810 123.245 ;
        RECT 27.110 118.485 27.370 118.805 ;
        RECT 26.630 110.715 26.890 111.035 ;
        RECT 26.150 105.905 26.410 106.225 ;
        RECT 26.630 105.165 26.890 105.485 ;
        RECT 23.750 104.795 24.010 105.115 ;
        RECT 24.230 104.795 24.490 105.115 ;
        RECT 24.290 103.265 24.430 104.795 ;
        RECT 26.150 104.425 26.410 104.745 ;
        RECT 26.210 103.265 26.350 104.425 ;
        RECT 24.230 102.945 24.490 103.265 ;
        RECT 26.150 102.945 26.410 103.265 ;
        RECT 26.150 102.205 26.410 102.525 ;
        RECT 16.550 101.835 16.810 102.155 ;
        RECT 16.550 101.095 16.810 101.415 ;
        RECT 14.260 100.145 16.140 100.515 ;
        RECT 16.610 99.935 16.750 101.095 ;
        RECT 21.350 100.725 21.610 101.045 ;
        RECT 16.550 99.615 16.810 99.935 ;
        RECT 21.410 98.825 21.550 100.725 ;
        RECT 26.210 99.935 26.350 102.205 ;
        RECT 26.150 99.615 26.410 99.935 ;
        RECT 21.350 98.505 21.610 98.825 ;
        RECT 20.870 97.395 21.130 97.715 ;
        RECT 20.930 96.605 21.070 97.395 ;
        RECT 20.870 96.285 21.130 96.605 ;
        RECT 14.260 93.485 16.140 93.855 ;
        RECT 14.260 86.825 16.140 87.195 ;
        RECT 21.410 85.135 21.550 98.505 ;
        RECT 26.690 98.085 26.830 105.165 ;
        RECT 26.630 97.765 26.890 98.085 ;
        RECT 25.190 97.395 25.450 97.715 ;
        RECT 25.250 89.205 25.390 97.395 ;
        RECT 27.170 95.125 27.310 118.485 ;
        RECT 31.490 118.160 31.630 135.090 ;
        RECT 31.910 125.145 32.170 125.465 ;
        RECT 28.610 118.020 31.630 118.160 ;
        RECT 27.590 116.265 27.850 116.585 ;
        RECT 27.650 108.815 27.790 116.265 ;
        RECT 28.610 109.555 28.750 118.020 ;
        RECT 29.260 116.795 31.140 117.165 ;
        RECT 30.460 115.685 30.740 116.055 ;
        RECT 30.530 115.475 30.670 115.685 ;
        RECT 31.430 115.525 31.690 115.845 ;
        RECT 30.470 115.155 30.730 115.475 ;
        RECT 30.950 115.155 31.210 115.475 ;
        RECT 31.010 111.500 31.150 115.155 ;
        RECT 31.490 113.255 31.630 115.525 ;
        RECT 31.430 112.935 31.690 113.255 ;
        RECT 31.010 111.405 31.630 111.500 ;
        RECT 30.950 111.360 31.630 111.405 ;
        RECT 30.950 111.085 31.210 111.360 ;
        RECT 29.260 110.135 31.140 110.505 ;
        RECT 31.490 109.555 31.630 111.360 ;
        RECT 28.550 109.235 28.810 109.555 ;
        RECT 31.430 109.235 31.690 109.555 ;
        RECT 27.590 108.495 27.850 108.815 ;
        RECT 29.510 108.495 29.770 108.815 ;
        RECT 27.650 104.840 27.790 108.495 ;
        RECT 29.570 105.115 29.710 108.495 ;
        RECT 27.650 104.700 28.270 104.840 ;
        RECT 29.510 104.795 29.770 105.115 ;
        RECT 27.590 104.055 27.850 104.375 ;
        RECT 27.650 99.195 27.790 104.055 ;
        RECT 27.590 98.875 27.850 99.195 ;
        RECT 28.130 98.825 28.270 104.700 ;
        RECT 28.550 104.055 28.810 104.375 ;
        RECT 28.610 103.265 28.750 104.055 ;
        RECT 29.260 103.475 31.140 103.845 ;
        RECT 28.550 102.945 28.810 103.265 ;
        RECT 28.070 98.505 28.330 98.825 ;
        RECT 28.130 96.605 28.270 98.505 ;
        RECT 29.260 96.815 31.140 97.185 ;
        RECT 28.070 96.285 28.330 96.605 ;
        RECT 30.950 96.285 31.210 96.605 ;
        RECT 28.070 95.545 28.330 95.865 ;
        RECT 27.110 94.805 27.370 95.125 ;
        RECT 27.170 91.795 27.310 94.805 ;
        RECT 27.110 91.475 27.370 91.795 ;
        RECT 25.670 90.735 25.930 91.055 ;
        RECT 26.630 90.735 26.890 91.055 ;
        RECT 25.190 88.885 25.450 89.205 ;
        RECT 25.730 88.835 25.870 90.735 ;
        RECT 25.670 88.515 25.930 88.835 ;
        RECT 26.690 86.245 26.830 90.735 ;
        RECT 28.130 86.615 28.270 95.545 ;
        RECT 31.010 95.495 31.150 96.285 ;
        RECT 31.970 95.865 32.110 125.145 ;
        RECT 33.350 124.775 33.610 125.095 ;
        RECT 33.410 123.245 33.550 124.775 ;
        RECT 33.350 122.925 33.610 123.245 ;
        RECT 32.870 121.075 33.130 121.395 ;
        RECT 32.390 114.415 32.650 114.735 ;
        RECT 32.450 105.485 32.590 114.415 ;
        RECT 32.390 105.165 32.650 105.485 ;
        RECT 32.390 100.725 32.650 101.045 ;
        RECT 31.910 95.545 32.170 95.865 ;
        RECT 32.450 95.495 32.590 100.725 ;
        RECT 32.930 96.605 33.070 121.075 ;
        RECT 33.350 118.115 33.610 118.435 ;
        RECT 33.410 115.845 33.550 118.115 ;
        RECT 33.350 115.525 33.610 115.845 ;
        RECT 33.350 114.045 33.610 114.365 ;
        RECT 33.410 108.815 33.550 114.045 ;
        RECT 33.350 108.495 33.610 108.815 ;
        RECT 33.890 107.800 34.030 135.090 ;
        RECT 43.490 132.125 43.630 138.095 ;
        RECT 47.750 137.725 48.010 138.045 ;
        RECT 47.810 136.195 47.950 137.725 ;
        RECT 46.790 135.875 47.050 136.195 ;
        RECT 47.750 135.875 48.010 136.195 ;
        RECT 46.850 135.230 46.990 135.875 ;
        RECT 46.370 135.090 46.990 135.230 ;
        RECT 44.260 133.445 46.140 133.815 ;
        RECT 40.550 131.805 40.810 132.125 ;
        RECT 43.430 131.805 43.690 132.125 ;
        RECT 37.190 131.435 37.450 131.755 ;
        RECT 33.410 107.660 34.030 107.800 ;
        RECT 33.410 97.715 33.550 107.660 ;
        RECT 33.350 97.395 33.610 97.715 ;
        RECT 32.870 96.285 33.130 96.605 ;
        RECT 30.950 95.175 31.210 95.495 ;
        RECT 32.390 95.175 32.650 95.495 ;
        RECT 29.260 90.155 31.140 90.525 ;
        RECT 35.750 88.515 36.010 88.835 ;
        RECT 35.810 86.615 35.950 88.515 ;
        RECT 37.250 87.725 37.390 131.435 ;
        RECT 40.610 126.575 40.750 131.805 ;
        RECT 44.260 126.785 46.140 127.155 ;
        RECT 40.550 126.255 40.810 126.575 ;
        RECT 40.550 125.515 40.810 125.835 ;
        RECT 40.070 122.555 40.330 122.875 ;
        RECT 40.130 121.025 40.270 122.555 ;
        RECT 40.610 121.765 40.750 125.515 ;
        RECT 41.990 124.035 42.250 124.355 ;
        RECT 40.550 121.445 40.810 121.765 ;
        RECT 40.070 120.705 40.330 121.025 ;
        RECT 40.610 119.545 40.750 121.445 ;
        RECT 41.030 120.705 41.290 121.025 ;
        RECT 40.550 119.225 40.810 119.545 ;
        RECT 37.670 118.115 37.930 118.435 ;
        RECT 37.730 112.885 37.870 118.115 ;
        RECT 40.070 114.785 40.330 115.105 ;
        RECT 40.130 114.460 40.270 114.785 ;
        RECT 41.090 114.460 41.230 120.705 ;
        RECT 42.050 118.805 42.190 124.035 ;
        RECT 44.260 120.125 46.140 120.495 ;
        RECT 41.990 118.485 42.250 118.805 ;
        RECT 41.510 117.375 41.770 117.695 ;
        RECT 41.570 116.215 41.710 117.375 ;
        RECT 41.510 115.895 41.770 116.215 ;
        RECT 40.130 114.320 41.230 114.460 ;
        RECT 37.670 112.565 37.930 112.885 ;
        RECT 37.730 106.595 37.870 112.565 ;
        RECT 38.150 112.195 38.410 112.515 ;
        RECT 38.210 109.185 38.350 112.195 ;
        RECT 38.150 108.865 38.410 109.185 ;
        RECT 37.670 106.275 37.930 106.595 ;
        RECT 37.730 98.085 37.870 106.275 ;
        RECT 38.210 105.855 38.350 108.865 ;
        RECT 40.070 108.495 40.330 108.815 ;
        RECT 38.150 105.535 38.410 105.855 ;
        RECT 38.210 99.195 38.350 105.535 ;
        RECT 40.130 105.115 40.270 108.495 ;
        RECT 40.070 104.795 40.330 105.115 ;
        RECT 38.150 98.875 38.410 99.195 ;
        RECT 37.670 97.765 37.930 98.085 ;
        RECT 40.130 96.605 40.270 104.795 ;
        RECT 41.090 98.825 41.230 114.320 ;
        RECT 42.050 108.815 42.190 118.485 ;
        RECT 44.260 113.465 46.140 113.835 ;
        RECT 43.430 111.825 43.690 112.145 ;
        RECT 42.950 111.455 43.210 111.775 ;
        RECT 41.990 108.495 42.250 108.815 ;
        RECT 43.010 102.525 43.150 111.455 ;
        RECT 43.490 105.855 43.630 111.825 ;
        RECT 43.910 108.125 44.170 108.445 ;
        RECT 43.430 105.535 43.690 105.855 ;
        RECT 43.970 104.375 44.110 108.125 ;
        RECT 44.260 106.805 46.140 107.175 ;
        RECT 43.910 104.055 44.170 104.375 ;
        RECT 42.950 102.205 43.210 102.525 ;
        RECT 41.030 98.505 41.290 98.825 ;
        RECT 40.070 96.285 40.330 96.605 ;
        RECT 40.070 95.175 40.330 95.495 ;
        RECT 40.550 95.175 40.810 95.495 ;
        RECT 38.150 94.805 38.410 95.125 ;
        RECT 38.210 91.425 38.350 94.805 ;
        RECT 40.130 91.795 40.270 95.175 ;
        RECT 40.610 92.535 40.750 95.175 ;
        RECT 40.550 92.215 40.810 92.535 ;
        RECT 40.070 91.475 40.330 91.795 ;
        RECT 38.150 91.105 38.410 91.425 ;
        RECT 37.670 90.735 37.930 91.055 ;
        RECT 37.190 87.405 37.450 87.725 ;
        RECT 37.250 86.615 37.390 87.405 ;
        RECT 37.730 86.615 37.870 90.735 ;
        RECT 38.210 89.945 38.350 91.105 ;
        RECT 39.590 90.735 39.850 91.055 ;
        RECT 38.150 89.625 38.410 89.945 ;
        RECT 39.650 89.205 39.790 90.735 ;
        RECT 40.130 89.945 40.270 91.475 ;
        RECT 40.070 89.625 40.330 89.945 ;
        RECT 39.590 88.885 39.850 89.205 ;
        RECT 40.070 88.885 40.330 89.205 ;
        RECT 40.130 87.725 40.270 88.885 ;
        RECT 40.610 88.465 40.750 92.215 ;
        RECT 43.010 89.945 43.150 102.205 ;
        RECT 43.970 102.155 44.110 104.055 ;
        RECT 43.910 101.835 44.170 102.155 ;
        RECT 44.260 100.145 46.140 100.515 ;
        RECT 46.370 96.605 46.510 135.090 ;
        RECT 48.230 134.765 48.490 135.085 ;
        RECT 48.290 132.865 48.430 134.765 ;
        RECT 48.230 132.545 48.490 132.865 ;
        RECT 49.250 132.220 49.390 138.095 ;
        RECT 50.210 133.235 50.350 142.165 ;
        RECT 50.630 138.835 50.890 139.155 ;
        RECT 50.690 134.715 50.830 138.835 ;
        RECT 51.170 136.565 51.310 142.165 ;
        RECT 52.550 140.685 52.810 141.005 ;
        RECT 51.590 137.355 51.850 137.675 ;
        RECT 51.110 136.245 51.370 136.565 ;
        RECT 50.630 134.395 50.890 134.715 ;
        RECT 50.150 132.915 50.410 133.235 ;
        RECT 49.250 132.080 50.350 132.220 ;
        RECT 49.190 131.435 49.450 131.755 ;
        RECT 46.790 127.365 47.050 127.685 ;
        RECT 46.850 125.835 46.990 127.365 ;
        RECT 46.790 125.515 47.050 125.835 ;
        RECT 46.850 125.095 46.990 125.515 ;
        RECT 47.750 125.145 48.010 125.465 ;
        RECT 46.790 124.775 47.050 125.095 ;
        RECT 46.850 119.175 46.990 124.775 ;
        RECT 47.810 119.175 47.950 125.145 ;
        RECT 46.790 118.855 47.050 119.175 ;
        RECT 47.750 118.855 48.010 119.175 ;
        RECT 49.250 119.085 49.390 131.435 ;
        RECT 49.670 124.775 49.930 125.095 ;
        RECT 49.730 122.135 49.870 124.775 ;
        RECT 50.210 122.875 50.350 132.080 ;
        RECT 51.650 129.905 51.790 137.355 ;
        RECT 51.590 129.585 51.850 129.905 ;
        RECT 50.150 122.555 50.410 122.875 ;
        RECT 49.670 121.815 49.930 122.135 ;
        RECT 49.730 119.915 49.870 121.815 ;
        RECT 50.210 121.395 50.350 122.555 ;
        RECT 52.070 121.445 52.330 121.765 ;
        RECT 50.150 121.075 50.410 121.395 ;
        RECT 49.670 119.595 49.930 119.915 ;
        RECT 52.130 119.175 52.270 121.445 ;
        RECT 49.250 118.945 49.870 119.085 ;
        RECT 47.270 118.485 47.530 118.805 ;
        RECT 47.330 115.105 47.470 118.485 ;
        RECT 48.230 118.115 48.490 118.435 ;
        RECT 47.270 114.785 47.530 115.105 ;
        RECT 46.850 105.485 47.470 105.580 ;
        RECT 46.850 105.440 47.530 105.485 ;
        RECT 46.310 96.285 46.570 96.605 ;
        RECT 44.260 93.485 46.140 93.855 ;
        RECT 43.910 91.475 44.170 91.795 ;
        RECT 42.950 89.625 43.210 89.945 ;
        RECT 40.550 88.145 40.810 88.465 ;
        RECT 40.070 87.405 40.330 87.725 ;
        RECT 28.070 86.295 28.330 86.615 ;
        RECT 35.750 86.295 36.010 86.615 ;
        RECT 37.190 86.295 37.450 86.615 ;
        RECT 37.670 86.295 37.930 86.615 ;
        RECT 26.630 85.925 26.890 86.245 ;
        RECT 40.610 85.875 40.750 88.145 ;
        RECT 40.550 85.555 40.810 85.875 ;
        RECT 43.010 85.505 43.150 89.625 ;
        RECT 43.970 85.505 44.110 91.475 ;
        RECT 46.370 89.205 46.510 96.285 ;
        RECT 46.850 92.260 46.990 105.440 ;
        RECT 47.270 105.165 47.530 105.440 ;
        RECT 47.270 104.425 47.530 104.745 ;
        RECT 47.330 102.155 47.470 104.425 ;
        RECT 47.270 101.835 47.530 102.155 ;
        RECT 47.270 101.095 47.530 101.415 ;
        RECT 47.330 92.905 47.470 101.095 ;
        RECT 47.750 94.805 48.010 95.125 ;
        RECT 47.810 93.275 47.950 94.805 ;
        RECT 47.750 92.955 48.010 93.275 ;
        RECT 47.270 92.585 47.530 92.905 ;
        RECT 46.850 92.165 47.950 92.260 ;
        RECT 46.790 92.120 47.950 92.165 ;
        RECT 46.790 91.845 47.050 92.120 ;
        RECT 47.810 89.575 47.950 92.120 ;
        RECT 48.290 91.055 48.430 118.115 ;
        RECT 49.730 114.365 49.870 118.945 ;
        RECT 52.070 118.855 52.330 119.175 ;
        RECT 49.670 114.045 49.930 114.365 ;
        RECT 48.230 90.735 48.490 91.055 ;
        RECT 47.750 89.255 48.010 89.575 ;
        RECT 49.730 89.205 49.870 114.045 ;
        RECT 51.590 108.125 51.850 108.445 ;
        RECT 51.650 106.225 51.790 108.125 ;
        RECT 51.590 105.905 51.850 106.225 ;
        RECT 51.650 101.785 51.790 105.905 ;
        RECT 52.610 103.265 52.750 140.685 ;
        RECT 53.510 137.355 53.770 137.675 ;
        RECT 53.570 135.825 53.710 137.355 ;
        RECT 53.510 135.505 53.770 135.825 ;
        RECT 54.050 133.235 54.190 148.985 ;
        RECT 54.530 141.375 54.670 152.850 ;
        RECT 59.260 143.435 61.140 143.805 ;
        RECT 57.820 142.325 58.100 142.695 ;
        RECT 54.470 141.055 54.730 141.375 ;
        RECT 57.890 136.565 58.030 142.325 ;
        RECT 59.750 141.795 60.010 142.115 ;
        RECT 59.810 139.895 59.950 141.795 ;
        RECT 61.730 141.375 61.870 153.540 ;
        RECT 65.800 152.850 66.400 157.050 ;
        RECT 71.600 155.225 72.200 157.050 ;
        RECT 91.700 155.225 92.100 155.275 ;
        RECT 71.600 154.825 92.100 155.225 ;
        RECT 71.600 153.680 72.200 154.825 ;
        RECT 91.700 154.775 92.100 154.825 ;
        RECT 70.370 153.540 72.200 153.680 ;
        RECT 62.150 142.905 62.410 143.225 ;
        RECT 61.670 141.055 61.930 141.375 ;
        RECT 59.750 139.575 60.010 139.895 ;
        RECT 59.260 136.775 61.140 137.145 ;
        RECT 57.830 136.245 58.090 136.565 ;
        RECT 54.470 135.875 54.730 136.195 ;
        RECT 53.990 132.915 54.250 133.235 ;
        RECT 53.510 115.155 53.770 115.475 ;
        RECT 53.570 112.145 53.710 115.155 ;
        RECT 53.510 111.825 53.770 112.145 ;
        RECT 53.570 109.555 53.710 111.825 ;
        RECT 53.510 109.235 53.770 109.555 ;
        RECT 52.550 102.945 52.810 103.265 ;
        RECT 51.590 101.465 51.850 101.785 ;
        RECT 51.650 98.455 51.790 101.465 ;
        RECT 51.590 98.135 51.850 98.455 ;
        RECT 51.650 91.795 51.790 98.135 ;
        RECT 52.070 97.395 52.330 97.715 ;
        RECT 52.130 95.125 52.270 97.395 ;
        RECT 52.070 94.805 52.330 95.125 ;
        RECT 51.590 91.475 51.850 91.795 ;
        RECT 52.130 90.780 52.270 94.805 ;
        RECT 52.610 91.795 52.750 102.945 ;
        RECT 54.530 98.455 54.670 135.875 ;
        RECT 57.830 135.505 58.090 135.825 ;
        RECT 58.310 135.505 58.570 135.825 ;
        RECT 61.670 135.505 61.930 135.825 ;
        RECT 55.430 135.135 55.690 135.455 ;
        RECT 54.950 122.185 55.210 122.505 ;
        RECT 55.010 118.160 55.150 122.185 ;
        RECT 55.490 121.025 55.630 135.135 ;
        RECT 57.890 132.495 58.030 135.505 ;
        RECT 57.830 132.175 58.090 132.495 ;
        RECT 56.870 131.435 57.130 131.755 ;
        RECT 56.930 129.165 57.070 131.435 ;
        RECT 56.870 128.845 57.130 129.165 ;
        RECT 55.910 121.075 56.170 121.395 ;
        RECT 55.430 120.705 55.690 121.025 ;
        RECT 55.010 118.020 55.630 118.160 ;
        RECT 54.950 117.375 55.210 117.695 ;
        RECT 55.010 115.845 55.150 117.375 ;
        RECT 54.950 115.525 55.210 115.845 ;
        RECT 54.470 98.135 54.730 98.455 ;
        RECT 52.550 91.475 52.810 91.795 ;
        RECT 52.130 90.640 52.750 90.780 ;
        RECT 46.310 88.885 46.570 89.205 ;
        RECT 49.670 88.885 49.930 89.205 ;
        RECT 52.610 88.465 52.750 90.640 ;
        RECT 54.530 88.560 54.670 98.135 ;
        RECT 55.490 88.835 55.630 118.020 ;
        RECT 55.970 102.525 56.110 121.075 ;
        RECT 56.930 118.435 57.070 128.845 ;
        RECT 57.890 128.055 58.030 132.175 ;
        RECT 57.830 127.735 58.090 128.055 ;
        RECT 57.350 120.705 57.610 121.025 ;
        RECT 56.870 118.115 57.130 118.435 ;
        RECT 56.870 111.455 57.130 111.775 ;
        RECT 56.390 108.865 56.650 109.185 ;
        RECT 56.450 105.115 56.590 108.865 ;
        RECT 56.390 104.795 56.650 105.115 ;
        RECT 55.910 102.205 56.170 102.525 ;
        RECT 55.910 97.395 56.170 97.715 ;
        RECT 46.310 88.145 46.570 88.465 ;
        RECT 52.550 88.145 52.810 88.465 ;
        RECT 54.050 88.420 54.670 88.560 ;
        RECT 55.430 88.515 55.690 88.835 ;
        RECT 46.370 87.820 46.510 88.145 ;
        RECT 46.370 87.680 46.990 87.820 ;
        RECT 44.260 86.825 46.140 87.195 ;
        RECT 46.850 86.615 46.990 87.680 ;
        RECT 46.790 86.295 47.050 86.615 ;
        RECT 46.850 85.505 46.990 86.295 ;
        RECT 52.610 85.875 52.750 88.145 ;
        RECT 53.510 87.405 53.770 87.725 ;
        RECT 52.550 85.555 52.810 85.875 ;
        RECT 26.630 85.185 26.890 85.505 ;
        RECT 40.070 85.185 40.330 85.505 ;
        RECT 42.950 85.185 43.210 85.505 ;
        RECT 43.910 85.185 44.170 85.505 ;
        RECT 46.790 85.185 47.050 85.505 ;
        RECT 21.350 84.815 21.610 85.135 ;
        RECT 13.190 84.075 13.450 84.395 ;
        RECT 12.220 73.760 12.500 74.360 ;
        RECT 13.250 73.760 13.390 84.075 ;
        RECT 12.220 73.620 13.390 73.760 ;
        RECT 26.140 73.760 26.420 74.360 ;
        RECT 26.690 73.760 26.830 85.185 ;
        RECT 29.260 83.495 31.140 83.865 ;
        RECT 40.130 74.360 40.270 85.185 ;
        RECT 53.570 75.355 53.710 87.405 ;
        RECT 54.050 86.615 54.190 88.420 ;
        RECT 54.470 87.775 54.730 88.095 ;
        RECT 55.430 87.775 55.690 88.095 ;
        RECT 53.990 86.295 54.250 86.615 ;
        RECT 53.990 84.815 54.250 85.135 ;
        RECT 53.500 74.985 53.780 75.355 ;
        RECT 54.050 74.360 54.190 84.815 ;
        RECT 54.530 81.275 54.670 87.775 ;
        RECT 55.490 86.615 55.630 87.775 ;
        RECT 55.430 86.295 55.690 86.615 ;
        RECT 54.460 80.905 54.740 81.275 ;
        RECT 55.970 78.315 56.110 97.395 ;
        RECT 56.450 95.495 56.590 104.795 ;
        RECT 56.930 99.195 57.070 111.455 ;
        RECT 56.870 98.875 57.130 99.195 ;
        RECT 56.390 95.175 56.650 95.495 ;
        RECT 56.450 92.165 56.590 95.175 ;
        RECT 56.930 92.535 57.070 98.875 ;
        RECT 57.410 95.865 57.550 120.705 ;
        RECT 57.830 118.855 58.090 119.175 ;
        RECT 57.890 115.105 58.030 118.855 ;
        RECT 57.830 114.785 58.090 115.105 ;
        RECT 57.890 112.515 58.030 114.785 ;
        RECT 58.370 113.255 58.510 135.505 ;
        RECT 58.790 131.805 59.050 132.125 ;
        RECT 58.850 125.095 58.990 131.805 ;
        RECT 59.260 130.115 61.140 130.485 ;
        RECT 59.270 128.475 59.530 128.795 ;
        RECT 59.330 126.205 59.470 128.475 ;
        RECT 59.270 125.885 59.530 126.205 ;
        RECT 58.790 124.775 59.050 125.095 ;
        RECT 59.260 123.455 61.140 123.825 ;
        RECT 59.270 122.185 59.530 122.505 ;
        RECT 59.330 118.805 59.470 122.185 ;
        RECT 59.270 118.485 59.530 118.805 ;
        RECT 59.330 118.160 59.470 118.485 ;
        RECT 58.850 118.020 59.470 118.160 ;
        RECT 58.850 116.585 58.990 118.020 ;
        RECT 59.260 116.795 61.140 117.165 ;
        RECT 61.730 116.680 61.870 135.505 ;
        RECT 62.210 119.915 62.350 142.905 ;
        RECT 66.050 142.485 66.190 152.850 ;
        RECT 65.990 142.165 66.250 142.485 ;
        RECT 64.550 141.795 64.810 142.115 ;
        RECT 63.590 137.515 63.850 137.675 ;
        RECT 63.580 137.145 63.860 137.515 ;
        RECT 64.610 136.565 64.750 141.795 ;
        RECT 65.980 140.105 66.260 140.475 ;
        RECT 66.050 136.565 66.190 140.105 ;
        RECT 66.470 138.140 66.730 138.415 ;
        RECT 66.470 138.095 67.630 138.140 ;
        RECT 68.390 138.095 68.650 138.415 ;
        RECT 66.530 138.000 67.630 138.095 ;
        RECT 66.470 137.355 66.730 137.675 ;
        RECT 64.550 136.245 64.810 136.565 ;
        RECT 65.990 136.245 66.250 136.565 ;
        RECT 65.510 135.505 65.770 135.825 ;
        RECT 65.570 135.230 65.710 135.505 ;
        RECT 65.090 135.090 65.710 135.230 ;
        RECT 63.110 124.775 63.370 125.095 ;
        RECT 62.150 119.595 62.410 119.915 ;
        RECT 61.250 116.585 61.870 116.680 ;
        RECT 58.790 116.265 59.050 116.585 ;
        RECT 61.190 116.540 61.870 116.585 ;
        RECT 61.190 116.265 61.450 116.540 ;
        RECT 59.270 115.525 59.530 115.845 ;
        RECT 58.310 112.935 58.570 113.255 ;
        RECT 57.830 112.195 58.090 112.515 ;
        RECT 59.330 112.145 59.470 115.525 ;
        RECT 59.270 111.825 59.530 112.145 ;
        RECT 57.830 110.715 58.090 111.035 ;
        RECT 57.350 95.545 57.610 95.865 ;
        RECT 57.350 94.065 57.610 94.385 ;
        RECT 56.870 92.215 57.130 92.535 ;
        RECT 56.390 91.845 56.650 92.165 ;
        RECT 56.450 89.945 56.590 91.845 ;
        RECT 56.390 89.625 56.650 89.945 ;
        RECT 57.410 89.575 57.550 94.065 ;
        RECT 57.890 91.520 58.030 110.715 ;
        RECT 59.260 110.135 61.140 110.505 ;
        RECT 62.630 104.795 62.890 105.115 ;
        RECT 58.790 104.055 59.050 104.375 ;
        RECT 58.310 100.725 58.570 101.045 ;
        RECT 58.370 99.195 58.510 100.725 ;
        RECT 58.310 98.875 58.570 99.195 ;
        RECT 58.370 92.535 58.510 98.875 ;
        RECT 58.850 98.825 58.990 104.055 ;
        RECT 59.260 103.475 61.140 103.845 ;
        RECT 61.190 100.725 61.450 101.045 ;
        RECT 61.250 99.035 61.390 100.725 ;
        RECT 58.790 98.505 59.050 98.825 ;
        RECT 61.180 98.665 61.460 99.035 ;
        RECT 59.260 96.815 61.140 97.185 ;
        RECT 58.310 92.215 58.570 92.535 ;
        RECT 57.890 91.380 58.510 91.520 ;
        RECT 57.350 89.255 57.610 89.575 ;
        RECT 57.410 86.615 57.550 89.255 ;
        RECT 58.370 89.205 58.510 91.380 ;
        RECT 61.670 90.735 61.930 91.055 ;
        RECT 59.260 90.155 61.140 90.525 ;
        RECT 58.310 88.885 58.570 89.205 ;
        RECT 60.710 88.515 60.970 88.835 ;
        RECT 57.350 86.295 57.610 86.615 ;
        RECT 58.310 86.295 58.570 86.615 ;
        RECT 58.370 85.505 58.510 86.295 ;
        RECT 60.770 86.245 60.910 88.515 ;
        RECT 60.710 85.925 60.970 86.245 ;
        RECT 58.310 85.185 58.570 85.505 ;
        RECT 61.730 84.235 61.870 90.735 ;
        RECT 62.690 86.615 62.830 104.795 ;
        RECT 63.170 96.235 63.310 124.775 ;
        RECT 64.070 124.035 64.330 124.355 ;
        RECT 64.130 122.715 64.270 124.035 ;
        RECT 64.060 122.345 64.340 122.715 ;
        RECT 64.060 104.585 64.340 104.955 ;
        RECT 64.070 104.425 64.330 104.585 ;
        RECT 63.110 95.915 63.370 96.235 ;
        RECT 65.090 88.095 65.230 135.090 ;
        RECT 66.530 134.555 66.670 137.355 ;
        RECT 66.460 134.185 66.740 134.555 ;
        RECT 66.950 134.025 67.210 134.345 ;
        RECT 67.010 131.595 67.150 134.025 ;
        RECT 66.940 131.225 67.220 131.595 ;
        RECT 66.950 128.105 67.210 128.425 ;
        RECT 67.010 125.675 67.150 128.105 ;
        RECT 66.940 125.305 67.220 125.675 ;
        RECT 66.950 120.705 67.210 121.025 ;
        RECT 67.010 119.755 67.150 120.705 ;
        RECT 66.940 119.385 67.220 119.755 ;
        RECT 66.940 116.425 67.220 116.795 ;
        RECT 66.950 116.265 67.210 116.425 ;
        RECT 66.940 110.505 67.220 110.875 ;
        RECT 65.990 108.125 66.250 108.445 ;
        RECT 66.050 107.915 66.190 108.125 ;
        RECT 65.980 107.545 66.260 107.915 ;
        RECT 67.010 105.855 67.150 110.505 ;
        RECT 66.950 105.535 67.210 105.855 ;
        RECT 66.940 101.625 67.220 101.995 ;
        RECT 66.950 101.465 67.210 101.625 ;
        RECT 67.490 99.195 67.630 138.000 ;
        RECT 67.430 98.875 67.690 99.195 ;
        RECT 65.510 97.395 65.770 97.715 ;
        RECT 65.030 87.775 65.290 88.095 ;
        RECT 62.630 86.295 62.890 86.615 ;
        RECT 65.570 85.135 65.710 97.395 ;
        RECT 66.950 96.285 67.210 96.605 ;
        RECT 67.010 96.075 67.150 96.285 ;
        RECT 66.940 95.705 67.220 96.075 ;
        RECT 68.450 91.795 68.590 138.095 ;
        RECT 69.340 128.265 69.620 128.635 ;
        RECT 69.410 126.575 69.550 128.265 ;
        RECT 69.350 126.255 69.610 126.575 ;
        RECT 70.370 116.055 70.510 153.540 ;
        RECT 71.600 152.850 72.200 153.540 ;
        RECT 70.300 115.685 70.580 116.055 ;
        RECT 68.860 113.465 69.140 113.835 ;
        RECT 68.930 109.925 69.070 113.465 ;
        RECT 68.870 109.605 69.130 109.925 ;
        RECT 100.700 94.400 102.700 159.800 ;
        RECT 105.100 132.400 107.100 163.800 ;
        RECT 200.885 162.630 201.405 163.250 ;
        RECT 221.125 161.590 221.645 162.210 ;
        RECT 231.245 160.550 231.765 161.170 ;
        RECT 236.305 159.510 236.825 160.130 ;
        RECT 123.460 150.765 123.960 154.920 ;
        RECT 130.475 151.390 135.350 151.690 ;
        RECT 147.470 150.765 147.970 155.960 ;
        RECT 154.485 151.390 159.360 151.690 ;
        RECT 167.665 150.765 168.165 157.000 ;
        RECT 178.495 151.390 183.370 151.690 ;
        RECT 195.490 150.765 195.990 158.040 ;
        RECT 202.505 151.390 207.380 151.690 ;
        RECT 219.500 150.765 220.000 159.080 ;
        RECT 226.515 151.390 231.390 151.690 ;
        RECT 243.515 150.765 244.015 160.120 ;
        RECT 245.025 158.470 245.425 214.910 ;
        RECT 248.585 214.350 249.065 214.930 ;
        RECT 245.825 157.430 246.225 204.110 ;
        RECT 248.585 203.550 249.065 204.130 ;
        RECT 246.625 156.390 247.025 200.510 ;
        RECT 248.585 199.950 249.065 200.530 ;
        RECT 248.585 195.810 249.065 196.390 ;
        RECT 248.585 190.410 249.065 190.990 ;
        RECT 248.585 189.150 249.065 189.730 ;
        RECT 248.585 181.950 249.065 182.530 ;
        RECT 248.585 171.150 249.065 171.730 ;
        RECT 252.085 155.350 252.485 194.570 ;
        RECT 252.885 154.310 253.285 192.770 ;
        RECT 253.685 153.270 254.085 196.370 ;
        RECT 290.905 162.630 291.425 163.250 ;
        RECT 270.665 161.590 271.185 162.210 ;
        RECT 260.545 160.550 261.065 161.170 ;
        RECT 255.485 159.510 256.005 160.130 ;
        RECT 250.530 151.390 255.405 151.690 ;
        RECT 267.555 150.765 268.055 161.160 ;
        RECT 274.585 151.390 279.460 151.690 ;
        RECT 291.530 150.765 292.030 162.200 ;
        RECT 298.545 151.390 303.420 151.690 ;
        RECT 315.540 150.765 316.040 163.240 ;
        RECT 322.555 151.390 327.430 151.690 ;
        RECT 116.750 150.265 125.370 150.765 ;
        RECT 140.760 150.265 149.380 150.765 ;
        RECT 164.770 150.265 173.390 150.765 ;
        RECT 188.780 150.265 197.400 150.765 ;
        RECT 212.790 150.265 221.410 150.765 ;
        RECT 236.805 150.265 245.425 150.765 ;
        RECT 260.860 150.265 269.480 150.765 ;
        RECT 284.820 150.265 293.440 150.765 ;
        RECT 308.830 150.265 317.450 150.765 ;
        RECT 113.750 149.265 119.230 149.765 ;
        RECT 129.780 149.090 130.795 149.390 ;
        RECT 134.285 149.090 135.350 149.390 ;
        RECT 137.760 149.265 143.240 149.765 ;
        RECT 153.790 149.090 154.805 149.390 ;
        RECT 158.295 149.090 159.360 149.390 ;
        RECT 161.770 149.265 167.250 149.765 ;
        RECT 177.800 149.090 178.815 149.390 ;
        RECT 182.305 149.090 183.370 149.390 ;
        RECT 185.780 149.265 191.260 149.765 ;
        RECT 201.810 149.090 202.825 149.390 ;
        RECT 206.315 149.090 207.380 149.390 ;
        RECT 209.790 149.265 215.270 149.765 ;
        RECT 225.820 149.090 226.835 149.390 ;
        RECT 230.325 149.090 231.390 149.390 ;
        RECT 233.805 149.265 239.285 149.765 ;
        RECT 249.835 149.090 250.850 149.390 ;
        RECT 254.340 149.090 255.405 149.390 ;
        RECT 257.860 149.265 263.340 149.765 ;
        RECT 273.890 149.090 274.905 149.390 ;
        RECT 278.395 149.090 279.460 149.390 ;
        RECT 281.820 149.265 287.300 149.765 ;
        RECT 297.850 149.090 298.865 149.390 ;
        RECT 302.355 149.090 303.420 149.390 ;
        RECT 305.830 149.265 311.310 149.765 ;
        RECT 321.860 149.090 322.875 149.390 ;
        RECT 326.365 149.090 327.430 149.390 ;
        RECT 129.780 144.125 130.080 149.090 ;
        RECT 130.470 148.170 131.805 148.470 ;
        RECT 133.265 148.170 134.600 148.470 ;
        RECT 130.520 144.845 135.350 145.145 ;
        RECT 153.790 144.125 154.090 149.090 ;
        RECT 154.480 148.170 155.815 148.470 ;
        RECT 157.275 148.170 158.610 148.470 ;
        RECT 154.530 144.845 159.360 145.145 ;
        RECT 177.800 144.125 178.100 149.090 ;
        RECT 178.490 148.170 179.825 148.470 ;
        RECT 181.285 148.170 182.620 148.470 ;
        RECT 178.540 144.845 183.370 145.145 ;
        RECT 201.810 144.125 202.110 149.090 ;
        RECT 202.500 148.170 203.835 148.470 ;
        RECT 205.295 148.170 206.630 148.470 ;
        RECT 202.550 144.845 207.380 145.145 ;
        RECT 225.820 144.125 226.120 149.090 ;
        RECT 226.510 148.170 227.845 148.470 ;
        RECT 229.305 148.170 230.640 148.470 ;
        RECT 226.560 144.845 231.390 145.145 ;
        RECT 249.835 144.125 250.135 149.090 ;
        RECT 250.525 148.170 251.860 148.470 ;
        RECT 253.320 148.170 254.655 148.470 ;
        RECT 250.575 144.845 255.405 145.145 ;
        RECT 273.890 144.125 274.190 149.090 ;
        RECT 274.580 148.170 275.915 148.470 ;
        RECT 277.375 148.170 278.710 148.470 ;
        RECT 274.630 144.845 279.460 145.145 ;
        RECT 297.850 144.125 298.150 149.090 ;
        RECT 298.540 148.170 299.875 148.470 ;
        RECT 301.335 148.170 302.670 148.470 ;
        RECT 298.590 144.845 303.420 145.145 ;
        RECT 321.860 144.125 322.160 149.090 ;
        RECT 322.550 148.170 323.885 148.470 ;
        RECT 325.345 148.170 326.680 148.470 ;
        RECT 322.600 144.845 327.430 145.145 ;
        RECT 129.780 143.825 134.545 144.125 ;
        RECT 153.790 143.825 158.555 144.125 ;
        RECT 177.800 143.825 182.565 144.125 ;
        RECT 201.810 143.825 206.575 144.125 ;
        RECT 225.820 143.825 230.585 144.125 ;
        RECT 249.835 143.825 254.600 144.125 ;
        RECT 273.890 143.825 278.655 144.125 ;
        RECT 297.850 143.825 302.615 144.125 ;
        RECT 321.860 143.825 326.625 144.125 ;
        RECT 129.005 142.885 136.070 143.185 ;
        RECT 153.015 142.885 160.080 143.185 ;
        RECT 177.025 142.885 184.090 143.185 ;
        RECT 201.035 142.885 208.100 143.185 ;
        RECT 225.045 142.885 232.110 143.185 ;
        RECT 249.060 142.885 256.125 143.185 ;
        RECT 273.115 142.885 280.180 143.185 ;
        RECT 297.075 142.885 304.140 143.185 ;
        RECT 321.085 142.885 328.150 143.185 ;
        RECT 118.870 134.830 119.370 141.120 ;
        RECT 129.750 136.160 130.905 136.460 ;
        RECT 133.265 136.160 134.565 136.460 ;
        RECT 153.760 136.160 154.915 136.460 ;
        RECT 157.275 136.160 158.575 136.460 ;
        RECT 177.770 136.160 178.925 136.460 ;
        RECT 181.285 136.160 182.585 136.460 ;
        RECT 201.780 136.160 202.935 136.460 ;
        RECT 205.295 136.160 206.595 136.460 ;
        RECT 225.790 136.160 226.945 136.460 ;
        RECT 229.305 136.160 230.605 136.460 ;
        RECT 249.805 136.160 250.960 136.460 ;
        RECT 253.320 136.160 254.620 136.460 ;
        RECT 273.860 136.160 275.015 136.460 ;
        RECT 277.375 136.160 278.675 136.460 ;
        RECT 297.820 136.160 298.975 136.460 ;
        RECT 301.335 136.160 302.635 136.460 ;
        RECT 321.830 136.160 322.985 136.460 ;
        RECT 325.345 136.160 326.645 136.460 ;
        RECT 134.900 135.195 135.400 135.595 ;
        RECT 158.910 135.195 159.410 135.595 ;
        RECT 182.920 135.195 183.420 135.595 ;
        RECT 206.930 135.195 207.430 135.595 ;
        RECT 230.940 135.195 231.440 135.595 ;
        RECT 254.955 135.195 255.455 135.595 ;
        RECT 279.010 135.195 279.510 135.595 ;
        RECT 302.970 135.195 303.470 135.595 ;
        RECT 326.980 135.195 327.480 135.595 ;
        RECT 113.750 133.905 119.230 134.405 ;
        RECT 121.110 134.250 128.030 134.510 ;
        RECT 137.760 133.905 143.240 134.405 ;
        RECT 145.120 134.250 152.040 134.510 ;
        RECT 161.770 133.905 167.250 134.405 ;
        RECT 169.130 134.250 176.050 134.510 ;
        RECT 185.780 133.905 191.260 134.405 ;
        RECT 193.140 134.250 200.060 134.510 ;
        RECT 209.790 133.905 215.270 134.405 ;
        RECT 217.150 134.250 224.070 134.510 ;
        RECT 233.805 133.905 239.285 134.405 ;
        RECT 241.165 134.250 248.085 134.510 ;
        RECT 257.860 133.905 263.340 134.405 ;
        RECT 265.220 134.250 272.140 134.510 ;
        RECT 281.820 133.905 287.300 134.405 ;
        RECT 289.180 134.250 296.100 134.510 ;
        RECT 305.830 133.905 311.310 134.405 ;
        RECT 313.190 134.250 320.110 134.510 ;
        RECT 112.750 132.900 328.240 133.400 ;
        RECT 105.100 131.900 328.220 132.400 ;
        RECT 112.750 130.900 136.110 131.400 ;
        RECT 136.760 130.900 160.120 131.400 ;
        RECT 160.770 130.900 184.130 131.400 ;
        RECT 184.780 130.900 208.140 131.400 ;
        RECT 208.790 130.900 232.150 131.400 ;
        RECT 232.805 130.900 256.165 131.400 ;
        RECT 256.860 130.900 280.220 131.400 ;
        RECT 280.820 130.900 304.180 131.400 ;
        RECT 304.830 130.900 328.190 131.400 ;
        RECT 112.750 129.900 136.110 130.400 ;
        RECT 136.760 129.900 160.120 130.400 ;
        RECT 160.770 129.900 184.130 130.400 ;
        RECT 184.780 129.900 208.140 130.400 ;
        RECT 208.790 129.900 232.150 130.400 ;
        RECT 232.805 129.900 256.165 130.400 ;
        RECT 256.860 129.900 280.220 130.400 ;
        RECT 280.820 129.900 304.180 130.400 ;
        RECT 304.830 129.900 328.190 130.400 ;
        RECT 112.750 128.900 136.110 129.400 ;
        RECT 136.760 128.900 160.120 129.400 ;
        RECT 160.770 128.900 184.130 129.400 ;
        RECT 184.780 128.900 208.140 129.400 ;
        RECT 208.790 128.900 232.150 129.400 ;
        RECT 232.805 128.900 256.165 129.400 ;
        RECT 256.860 128.900 280.220 129.400 ;
        RECT 280.820 128.900 304.180 129.400 ;
        RECT 304.830 128.900 328.190 129.400 ;
        RECT 112.750 127.900 136.110 128.400 ;
        RECT 136.760 127.900 160.120 128.400 ;
        RECT 160.770 127.900 184.130 128.400 ;
        RECT 184.780 127.900 208.140 128.400 ;
        RECT 208.790 127.900 232.150 128.400 ;
        RECT 232.805 127.900 256.165 128.400 ;
        RECT 256.860 127.900 280.220 128.400 ;
        RECT 280.820 127.900 304.180 128.400 ;
        RECT 304.830 127.900 328.190 128.400 ;
        RECT 111.750 127.400 112.250 127.450 ;
        RECT 111.750 126.900 329.450 127.400 ;
        RECT 111.750 126.850 112.250 126.900 ;
        RECT 112.750 125.900 136.110 126.400 ;
        RECT 136.760 125.900 160.120 126.400 ;
        RECT 160.770 125.900 184.130 126.400 ;
        RECT 184.780 125.900 208.140 126.400 ;
        RECT 208.790 125.900 232.150 126.400 ;
        RECT 232.805 125.900 256.165 126.400 ;
        RECT 256.810 125.900 280.220 126.400 ;
        RECT 280.820 125.900 304.180 126.400 ;
        RECT 304.830 125.900 328.190 126.400 ;
        RECT 113.800 125.400 114.300 125.450 ;
        RECT 137.810 125.400 138.310 125.450 ;
        RECT 161.820 125.400 162.320 125.450 ;
        RECT 112.750 124.900 136.110 125.400 ;
        RECT 136.760 124.900 160.120 125.400 ;
        RECT 160.770 124.900 184.130 125.400 ;
        RECT 184.780 124.900 208.140 125.400 ;
        RECT 208.790 124.900 232.150 125.400 ;
        RECT 232.805 124.900 256.165 125.400 ;
        RECT 256.860 124.900 280.220 125.400 ;
        RECT 280.820 124.900 304.180 125.400 ;
        RECT 304.830 124.900 328.190 125.400 ;
        RECT 113.800 124.850 114.300 124.900 ;
        RECT 137.810 124.850 138.310 124.900 ;
        RECT 161.820 124.850 162.320 124.900 ;
        RECT 257.810 124.880 258.410 124.900 ;
        RECT 185.830 123.350 186.330 123.950 ;
        RECT 209.840 122.350 210.340 122.950 ;
        RECT 233.850 121.350 234.350 121.950 ;
        RECT 257.860 120.350 258.360 120.950 ;
        RECT 281.870 119.350 282.370 119.950 ;
        RECT 305.880 118.350 306.380 118.950 ;
        RECT 112.800 117.350 113.300 117.950 ;
        RECT 136.810 116.350 137.310 116.950 ;
        RECT 160.820 115.350 161.320 115.950 ;
        RECT 184.830 114.350 185.330 114.950 ;
        RECT 208.840 113.350 209.340 113.950 ;
        RECT 232.850 112.350 233.350 112.950 ;
        RECT 256.860 111.350 257.360 111.950 ;
        RECT 280.870 110.350 281.370 110.950 ;
        RECT 304.880 109.350 305.380 109.950 ;
        RECT 113.800 108.350 114.300 108.950 ;
        RECT 137.810 107.350 138.310 107.950 ;
        RECT 161.820 106.350 162.320 106.950 ;
        RECT 185.830 105.350 186.330 105.950 ;
        RECT 209.840 104.350 210.340 104.950 ;
        RECT 233.850 103.350 234.350 103.950 ;
        RECT 257.860 102.420 258.360 102.950 ;
        RECT 257.810 102.400 258.410 102.420 ;
        RECT 281.870 102.400 282.370 102.450 ;
        RECT 305.880 102.400 306.380 102.450 ;
        RECT 112.750 101.900 136.110 102.400 ;
        RECT 136.760 101.900 160.120 102.400 ;
        RECT 160.770 101.900 184.130 102.400 ;
        RECT 184.780 101.900 208.140 102.400 ;
        RECT 208.790 101.900 232.150 102.400 ;
        RECT 232.805 101.900 256.165 102.400 ;
        RECT 256.860 101.900 280.220 102.400 ;
        RECT 280.820 101.900 304.180 102.400 ;
        RECT 304.830 101.900 328.190 102.400 ;
        RECT 281.870 101.850 282.370 101.900 ;
        RECT 305.880 101.850 306.380 101.900 ;
        RECT 112.750 100.900 136.110 101.400 ;
        RECT 136.760 100.900 160.120 101.400 ;
        RECT 160.770 100.900 184.130 101.400 ;
        RECT 184.780 100.900 208.140 101.400 ;
        RECT 208.790 100.900 232.150 101.400 ;
        RECT 232.805 100.900 256.165 101.400 ;
        RECT 256.810 100.900 280.220 101.400 ;
        RECT 280.820 100.900 304.180 101.400 ;
        RECT 304.830 100.900 328.190 101.400 ;
        RECT 111.750 100.400 112.250 100.450 ;
        RECT 328.950 100.400 329.450 126.900 ;
        RECT 111.750 99.900 329.450 100.400 ;
        RECT 111.750 99.850 112.250 99.900 ;
        RECT 112.750 98.900 136.110 99.400 ;
        RECT 136.760 98.900 160.120 99.400 ;
        RECT 160.770 98.900 184.130 99.400 ;
        RECT 184.780 98.900 208.140 99.400 ;
        RECT 208.790 98.900 232.150 99.400 ;
        RECT 232.805 98.900 256.165 99.400 ;
        RECT 256.860 98.900 280.220 99.400 ;
        RECT 280.820 98.900 304.180 99.400 ;
        RECT 304.830 98.900 328.190 99.400 ;
        RECT 112.750 97.900 136.110 98.400 ;
        RECT 136.760 97.900 160.120 98.400 ;
        RECT 160.770 97.900 184.130 98.400 ;
        RECT 184.780 97.900 208.140 98.400 ;
        RECT 208.790 97.900 232.150 98.400 ;
        RECT 232.805 97.900 256.165 98.400 ;
        RECT 256.860 97.900 280.220 98.400 ;
        RECT 280.820 97.900 304.180 98.400 ;
        RECT 304.830 97.900 328.190 98.400 ;
        RECT 109.450 96.800 110.350 97.800 ;
        RECT 112.750 96.900 136.110 97.400 ;
        RECT 136.760 96.900 160.120 97.400 ;
        RECT 160.770 96.900 184.130 97.400 ;
        RECT 184.780 96.900 208.140 97.400 ;
        RECT 208.790 96.900 232.150 97.400 ;
        RECT 232.805 96.900 256.165 97.400 ;
        RECT 256.860 96.900 280.220 97.400 ;
        RECT 280.820 96.900 304.180 97.400 ;
        RECT 304.830 96.900 328.190 97.400 ;
        RECT 112.750 95.900 136.110 96.400 ;
        RECT 136.760 95.900 160.120 96.400 ;
        RECT 160.770 95.900 184.130 96.400 ;
        RECT 184.780 95.900 208.140 96.400 ;
        RECT 208.790 95.900 232.150 96.400 ;
        RECT 232.805 95.900 256.165 96.400 ;
        RECT 256.860 95.900 280.220 96.400 ;
        RECT 280.820 95.900 304.180 96.400 ;
        RECT 304.830 95.900 328.190 96.400 ;
        RECT 112.750 94.900 328.220 95.400 ;
        RECT 100.700 93.900 328.240 94.400 ;
        RECT 68.860 92.745 69.140 93.115 ;
        RECT 113.750 92.895 119.230 93.395 ;
        RECT 121.110 92.790 128.030 93.050 ;
        RECT 137.760 92.895 143.240 93.395 ;
        RECT 145.120 92.790 152.040 93.050 ;
        RECT 161.770 92.895 167.250 93.395 ;
        RECT 169.130 92.790 176.050 93.050 ;
        RECT 185.780 92.895 191.260 93.395 ;
        RECT 193.140 92.790 200.060 93.050 ;
        RECT 209.790 92.895 215.270 93.395 ;
        RECT 217.150 92.790 224.070 93.050 ;
        RECT 233.805 92.895 239.285 93.395 ;
        RECT 241.165 92.790 248.085 93.050 ;
        RECT 257.860 92.895 263.340 93.395 ;
        RECT 265.220 92.790 272.140 93.050 ;
        RECT 281.820 92.895 287.300 93.395 ;
        RECT 289.180 92.790 296.100 93.050 ;
        RECT 305.830 92.895 311.310 93.395 ;
        RECT 313.190 92.790 320.110 93.050 ;
        RECT 68.390 91.475 68.650 91.795 ;
        RECT 67.910 91.105 68.170 91.425 ;
        RECT 66.940 89.785 67.220 90.155 ;
        RECT 65.990 88.145 66.250 88.465 ;
        RECT 66.050 87.195 66.190 88.145 ;
        RECT 65.980 86.825 66.260 87.195 ;
        RECT 67.010 86.615 67.150 89.785 ;
        RECT 66.950 86.295 67.210 86.615 ;
        RECT 65.510 84.815 65.770 85.135 ;
        RECT 61.660 83.865 61.940 84.235 ;
        RECT 59.260 83.495 61.140 83.865 ;
        RECT 55.900 77.945 56.180 78.315 ;
        RECT 67.970 74.360 68.110 91.105 ;
        RECT 68.930 89.945 69.070 92.745 ;
        RECT 68.870 89.625 69.130 89.945 ;
        RECT 118.870 86.180 119.370 92.470 ;
        RECT 134.900 91.705 135.400 92.105 ;
        RECT 158.910 91.705 159.410 92.105 ;
        RECT 182.920 91.705 183.420 92.105 ;
        RECT 206.930 91.705 207.430 92.105 ;
        RECT 230.940 91.705 231.440 92.105 ;
        RECT 254.955 91.705 255.455 92.105 ;
        RECT 279.010 91.705 279.510 92.105 ;
        RECT 302.970 91.705 303.470 92.105 ;
        RECT 326.980 91.705 327.480 92.105 ;
        RECT 129.750 90.840 130.905 91.140 ;
        RECT 133.265 90.840 134.565 91.140 ;
        RECT 153.760 90.840 154.915 91.140 ;
        RECT 157.275 90.840 158.575 91.140 ;
        RECT 177.770 90.840 178.925 91.140 ;
        RECT 181.285 90.840 182.585 91.140 ;
        RECT 201.780 90.840 202.935 91.140 ;
        RECT 205.295 90.840 206.595 91.140 ;
        RECT 225.790 90.840 226.945 91.140 ;
        RECT 229.305 90.840 230.605 91.140 ;
        RECT 249.805 90.840 250.960 91.140 ;
        RECT 253.320 90.840 254.620 91.140 ;
        RECT 273.860 90.840 275.015 91.140 ;
        RECT 277.375 90.840 278.675 91.140 ;
        RECT 297.820 90.840 298.975 91.140 ;
        RECT 301.335 90.840 302.635 91.140 ;
        RECT 321.830 90.840 322.985 91.140 ;
        RECT 325.345 90.840 326.645 91.140 ;
        RECT 129.005 84.115 136.070 84.415 ;
        RECT 153.015 84.115 160.080 84.415 ;
        RECT 177.025 84.115 184.090 84.415 ;
        RECT 201.035 84.115 208.100 84.415 ;
        RECT 225.045 84.115 232.110 84.415 ;
        RECT 249.060 84.115 256.125 84.415 ;
        RECT 273.115 84.115 280.180 84.415 ;
        RECT 297.075 84.115 304.140 84.415 ;
        RECT 321.085 84.115 328.150 84.415 ;
        RECT 129.780 83.175 134.545 83.475 ;
        RECT 153.790 83.175 158.555 83.475 ;
        RECT 177.800 83.175 182.565 83.475 ;
        RECT 201.810 83.175 206.575 83.475 ;
        RECT 225.820 83.175 230.585 83.475 ;
        RECT 249.835 83.175 254.600 83.475 ;
        RECT 273.890 83.175 278.655 83.475 ;
        RECT 297.850 83.175 302.615 83.475 ;
        RECT 321.860 83.175 326.625 83.475 ;
        RECT 129.780 78.210 130.080 83.175 ;
        RECT 130.520 82.155 135.350 82.455 ;
        RECT 130.470 78.830 131.805 79.130 ;
        RECT 133.265 78.830 134.600 79.130 ;
        RECT 153.790 78.210 154.090 83.175 ;
        RECT 154.530 82.155 159.360 82.455 ;
        RECT 154.480 78.830 155.815 79.130 ;
        RECT 157.275 78.830 158.610 79.130 ;
        RECT 177.800 78.210 178.100 83.175 ;
        RECT 178.540 82.155 183.370 82.455 ;
        RECT 178.490 78.830 179.825 79.130 ;
        RECT 181.285 78.830 182.620 79.130 ;
        RECT 201.810 78.210 202.110 83.175 ;
        RECT 202.550 82.155 207.380 82.455 ;
        RECT 202.500 78.830 203.835 79.130 ;
        RECT 205.295 78.830 206.630 79.130 ;
        RECT 225.820 78.210 226.120 83.175 ;
        RECT 226.560 82.155 231.390 82.455 ;
        RECT 226.510 78.830 227.845 79.130 ;
        RECT 229.305 78.830 230.640 79.130 ;
        RECT 249.835 78.210 250.135 83.175 ;
        RECT 250.575 82.155 255.405 82.455 ;
        RECT 250.525 78.830 251.860 79.130 ;
        RECT 253.320 78.830 254.655 79.130 ;
        RECT 273.890 78.210 274.190 83.175 ;
        RECT 274.630 82.155 279.460 82.455 ;
        RECT 274.580 78.830 275.915 79.130 ;
        RECT 277.375 78.830 278.710 79.130 ;
        RECT 297.850 78.210 298.150 83.175 ;
        RECT 298.590 82.155 303.420 82.455 ;
        RECT 298.540 78.830 299.875 79.130 ;
        RECT 301.335 78.830 302.670 79.130 ;
        RECT 321.860 78.210 322.160 83.175 ;
        RECT 322.600 82.155 327.430 82.455 ;
        RECT 322.550 78.830 323.885 79.130 ;
        RECT 325.345 78.830 326.680 79.130 ;
        RECT 113.750 77.535 119.230 78.035 ;
        RECT 129.780 77.910 130.795 78.210 ;
        RECT 134.285 77.910 135.350 78.210 ;
        RECT 137.760 77.535 143.240 78.035 ;
        RECT 153.790 77.910 154.805 78.210 ;
        RECT 158.295 77.910 159.360 78.210 ;
        RECT 161.770 77.535 167.250 78.035 ;
        RECT 177.800 77.910 178.815 78.210 ;
        RECT 182.305 77.910 183.370 78.210 ;
        RECT 185.780 77.535 191.260 78.035 ;
        RECT 201.810 77.910 202.825 78.210 ;
        RECT 206.315 77.910 207.380 78.210 ;
        RECT 209.790 77.535 215.270 78.035 ;
        RECT 225.820 77.910 226.835 78.210 ;
        RECT 230.325 77.910 231.390 78.210 ;
        RECT 233.805 77.535 239.285 78.035 ;
        RECT 249.835 77.910 250.850 78.210 ;
        RECT 254.340 77.910 255.405 78.210 ;
        RECT 257.860 77.535 263.340 78.035 ;
        RECT 273.890 77.910 274.905 78.210 ;
        RECT 278.395 77.910 279.460 78.210 ;
        RECT 281.820 77.535 287.300 78.035 ;
        RECT 297.850 77.910 298.865 78.210 ;
        RECT 302.355 77.910 303.420 78.210 ;
        RECT 305.830 77.535 311.310 78.035 ;
        RECT 321.860 77.910 322.875 78.210 ;
        RECT 326.365 77.910 327.430 78.210 ;
        RECT 116.750 76.535 125.370 77.035 ;
        RECT 140.760 76.535 149.380 77.035 ;
        RECT 164.770 76.535 173.390 77.035 ;
        RECT 188.780 76.535 197.400 77.035 ;
        RECT 212.790 76.535 221.410 77.035 ;
        RECT 236.805 76.535 245.425 77.035 ;
        RECT 260.860 76.535 269.480 77.035 ;
        RECT 284.820 76.535 293.440 77.035 ;
        RECT 308.830 76.535 317.450 77.035 ;
        RECT 26.140 73.620 26.830 73.760 ;
        RECT 12.220 70.450 12.500 73.620 ;
        RECT 12.100 69.850 12.600 70.450 ;
        RECT 26.140 70.310 26.420 73.620 ;
        RECT 40.060 71.550 40.340 74.360 ;
        RECT 40.000 71.050 40.400 71.550 ;
        RECT 40.060 70.360 40.340 71.050 ;
        RECT 53.980 70.360 54.260 74.360 ;
        RECT 67.900 43.240 68.180 74.360 ;
        RECT 91.700 72.550 92.100 73.050 ;
        RECT 83.165 71.050 83.565 71.550 ;
        RECT 71.425 68.865 89.685 69.345 ;
        RECT 72.300 68.385 73.100 68.550 ;
        RECT 72.300 67.905 88.725 68.385 ;
        RECT 72.300 67.650 73.100 67.905 ;
        RECT 81.635 64.680 82.540 64.980 ;
        RECT 81.035 63.870 82.620 64.170 ;
        RECT 81.035 61.610 82.685 61.910 ;
        RECT 81.635 61.040 82.685 61.340 ;
        RECT 83.600 60.035 88.725 60.515 ;
        RECT 76.180 59.295 84.475 59.555 ;
        RECT 76.705 58.775 85.000 59.035 ;
        RECT 74.410 58.255 86.700 58.515 ;
        RECT 74.410 54.845 86.700 55.105 ;
        RECT 75.960 54.325 84.475 54.585 ;
        RECT 72.385 53.805 75.000 54.295 ;
        RECT 76.705 53.805 85.220 54.065 ;
        RECT 86.110 53.805 88.725 54.295 ;
        RECT 76.685 51.640 79.860 51.970 ;
        RECT 81.250 51.640 84.425 51.970 ;
        RECT 79.455 46.005 79.835 46.545 ;
        RECT 81.275 46.005 81.655 46.545 ;
        RECT 74.030 44.165 81.275 44.425 ;
        RECT 79.835 43.645 87.080 43.905 ;
        RECT 91.770 43.385 92.030 72.550 ;
        RECT 123.460 72.380 123.960 76.535 ;
        RECT 130.475 75.610 135.350 75.910 ;
        RECT 147.470 71.340 147.970 76.535 ;
        RECT 154.485 75.610 159.360 75.910 ;
        RECT 93.685 69.850 94.185 70.450 ;
        RECT 167.665 70.300 168.165 76.535 ;
        RECT 178.495 75.610 183.370 75.910 ;
        RECT 195.490 69.260 195.990 76.535 ;
        RECT 202.505 75.610 207.380 75.910 ;
        RECT 219.500 68.220 220.000 76.535 ;
        RECT 226.515 75.610 231.390 75.910 ;
        RECT 236.305 67.170 236.825 67.790 ;
        RECT 243.515 67.180 244.015 76.535 ;
        RECT 250.530 75.610 255.405 75.910 ;
        RECT 231.245 66.130 231.765 66.750 ;
        RECT 221.125 65.090 221.645 65.710 ;
        RECT 200.885 64.050 201.405 64.670 ;
        RECT 241.525 55.570 242.005 56.150 ;
        RECT 241.525 44.770 242.005 45.350 ;
        RECT 42.375 42.960 68.180 43.240 ;
        RECT 79.465 43.125 92.030 43.385 ;
        RECT 42.375 37.300 42.655 42.960 ;
        RECT 72.385 42.165 88.725 42.645 ;
        RECT 71.300 41.685 72.100 41.850 ;
        RECT 71.300 41.205 89.685 41.685 ;
        RECT 71.300 40.950 72.100 41.205 ;
        RECT 97.195 41.200 97.715 41.820 ;
        RECT 63.555 39.870 64.075 40.490 ;
        RECT 55.650 39.020 56.140 39.610 ;
        RECT 104.980 39.020 105.470 39.610 ;
        RECT 55.630 36.965 55.890 37.630 ;
        RECT 241.525 37.570 242.005 38.150 ;
        RECT 56.650 37.485 56.930 37.545 ;
        RECT 57.260 37.485 57.540 37.545 ;
        RECT 103.580 37.485 103.860 37.545 ;
        RECT 104.190 37.485 104.470 37.545 ;
        RECT 56.650 37.225 104.470 37.485 ;
        RECT 56.650 37.165 56.930 37.225 ;
        RECT 57.260 37.165 57.540 37.225 ;
        RECT 103.580 37.165 103.860 37.225 ;
        RECT 104.190 37.165 104.470 37.225 ;
        RECT 55.630 36.705 103.810 36.965 ;
        RECT 55.630 36.655 55.890 36.705 ;
        RECT 4.005 35.695 6.000 36.275 ;
        RECT 50.600 29.460 50.860 33.190 ;
        RECT 51.530 31.090 51.790 34.120 ;
        RECT 50.580 28.280 50.860 29.460 ;
        RECT 50.600 17.140 50.860 28.280 ;
        RECT 49.050 16.000 49.570 16.620 ;
        RECT 51.065 16.330 51.325 17.080 ;
        RECT 51.045 15.950 51.325 16.330 ;
        RECT 49.050 15.220 49.570 15.840 ;
        RECT 51.065 15.200 51.325 15.950 ;
        RECT 51.530 14.245 51.790 17.740 ;
        RECT 52.180 17.140 52.440 33.190 ;
        RECT 53.110 25.590 53.370 34.120 ;
        RECT 57.310 32.900 57.570 36.705 ;
        RECT 58.050 35.695 58.530 36.275 ;
        RECT 102.590 35.695 103.070 36.275 ;
        RECT 103.550 32.900 103.810 36.705 ;
        RECT 241.525 34.510 242.005 35.090 ;
        RECT 57.310 32.640 59.470 32.900 ;
        RECT 101.650 32.640 103.810 32.900 ;
        RECT 57.310 31.060 59.470 31.320 ;
        RECT 101.650 31.060 103.810 31.320 ;
        RECT 53.110 17.140 53.370 24.850 ;
        RECT 53.760 20.330 54.020 30.000 ;
        RECT 54.225 24.490 54.485 25.840 ;
        RECT 57.310 24.490 57.570 31.060 ;
        RECT 58.680 29.480 59.470 29.740 ;
        RECT 101.650 29.480 102.440 29.740 ;
        RECT 67.320 26.490 76.280 27.870 ;
        RECT 84.840 26.490 93.800 27.870 ;
        RECT 103.550 24.490 103.810 31.060 ;
        RECT 106.635 24.490 106.895 25.840 ;
        RECT 52.645 12.980 52.905 17.080 ;
        RECT 54.690 16.260 54.950 24.430 ;
        RECT 68.965 13.160 69.225 16.100 ;
        RECT 69.755 15.195 70.015 16.620 ;
        RECT 70.220 10.885 70.480 17.500 ;
        RECT 90.640 10.885 90.900 17.500 ;
        RECT 91.105 15.195 91.365 16.620 ;
        RECT 106.170 16.260 106.430 24.430 ;
        RECT 107.100 20.330 107.360 30.000 ;
        RECT 107.750 25.590 108.010 34.120 ;
        RECT 107.750 17.140 108.010 24.850 ;
        RECT 108.680 17.140 108.940 33.190 ;
        RECT 109.330 31.090 109.590 34.120 ;
        RECT 110.260 29.460 110.520 33.190 ;
        RECT 241.525 32.710 242.005 33.290 ;
        RECT 110.260 28.280 110.540 29.460 ;
        RECT 91.895 13.160 92.155 16.100 ;
        RECT 108.215 12.980 108.475 17.080 ;
        RECT 109.330 14.245 109.590 17.740 ;
        RECT 110.260 17.140 110.520 28.280 ;
        RECT 241.525 26.770 242.005 27.350 ;
        RECT 241.525 23.170 242.005 23.750 ;
        RECT 109.795 16.330 110.055 17.080 ;
        RECT 109.795 15.950 110.075 16.330 ;
        RECT 111.550 16.000 112.070 16.620 ;
        RECT 109.795 15.200 110.055 15.950 ;
        RECT 111.550 15.220 112.070 15.840 ;
        RECT 241.525 12.370 242.005 12.950 ;
        RECT 245.025 12.390 245.425 68.830 ;
        RECT 245.825 23.190 246.225 69.870 ;
        RECT 246.625 26.790 247.025 70.910 ;
        RECT 248.585 55.570 249.065 56.150 ;
        RECT 248.585 44.770 249.065 45.350 ;
        RECT 248.585 37.570 249.065 38.150 ;
        RECT 248.585 36.310 249.065 36.890 ;
        RECT 252.085 32.730 252.485 71.950 ;
        RECT 252.885 34.530 253.285 72.990 ;
        RECT 248.585 30.910 249.065 31.490 ;
        RECT 253.685 30.930 254.085 74.030 ;
        RECT 255.485 67.170 256.005 67.790 ;
        RECT 260.545 66.130 261.065 66.750 ;
        RECT 267.555 66.140 268.055 76.535 ;
        RECT 274.585 75.610 279.460 75.910 ;
        RECT 270.665 65.090 271.185 65.710 ;
        RECT 291.530 65.100 292.030 76.535 ;
        RECT 298.545 75.610 303.420 75.910 ;
        RECT 290.905 64.050 291.425 64.670 ;
        RECT 315.540 64.060 316.040 76.535 ;
        RECT 322.555 75.610 327.430 75.910 ;
        RECT 248.585 26.770 249.065 27.350 ;
        RECT 248.585 23.170 249.065 23.750 ;
        RECT 248.585 12.370 249.065 12.950 ;
        RECT 1.000 5.625 3.000 6.205 ;
        RECT 67.320 5.620 76.280 7.000 ;
        RECT 80.320 5.625 80.800 6.205 ;
        RECT 84.840 5.620 93.800 7.000 ;
        RECT 134.580 -5.700 135.060 -5.120 ;
      LAYER met3 ;
        RECT 134.530 232.445 135.110 232.975 ;
        RECT 97.195 222.720 167.785 223.240 ;
        RECT 47.050 221.800 47.650 222.300 ;
        RECT 49.850 221.800 50.450 222.300 ;
        RECT 47.100 215.125 47.600 221.800 ;
        RECT 49.900 215.125 50.400 221.800 ;
        RECT 0.950 213.125 50.400 215.125 ;
        RECT 8.220 211.005 8.820 211.100 ;
        RECT 95.605 211.005 96.205 211.125 ;
        RECT 8.220 210.705 96.205 211.005 ;
        RECT 8.220 210.600 8.820 210.705 ;
        RECT 95.605 210.575 96.205 210.705 ;
        RECT 85.050 165.800 87.150 165.825 ;
        RECT 0.950 163.800 87.150 165.800 ;
        RECT 85.050 163.775 87.150 163.800 ;
        RECT 85.050 161.800 87.150 161.825 ;
        RECT 3.950 159.800 87.150 161.800 ;
        RECT 85.050 159.775 87.150 159.800 ;
        RECT 8.150 152.875 8.850 157.025 ;
        RECT 13.950 152.875 14.650 157.025 ;
        RECT 19.650 152.875 20.350 157.025 ;
        RECT 25.450 152.875 26.150 157.025 ;
        RECT 31.150 152.875 31.850 157.025 ;
        RECT 36.950 152.875 37.650 157.025 ;
        RECT 42.750 152.875 43.450 157.025 ;
        RECT 48.450 152.875 49.150 157.025 ;
        RECT 54.250 152.875 54.950 157.025 ;
        RECT 60.050 152.875 60.750 157.025 ;
        RECT 65.750 152.875 66.450 157.025 ;
        RECT 71.550 152.875 72.250 157.025 ;
        RECT 91.650 154.800 92.150 155.250 ;
        RECT 47.715 152.280 48.045 152.295 ;
        RECT 71.880 152.280 75.980 152.430 ;
        RECT 47.715 151.980 75.980 152.280 ;
        RECT 47.715 151.965 48.045 151.980 ;
        RECT 71.880 151.830 75.980 151.980 ;
        RECT 53.955 149.320 54.285 149.335 ;
        RECT 71.880 149.320 75.980 149.470 ;
        RECT 53.955 149.020 75.980 149.320 ;
        RECT 53.955 149.005 54.285 149.020 ;
        RECT 0.950 146.900 16.250 148.900 ;
        RECT 71.880 148.870 75.980 149.020 ;
        RECT 47.715 146.360 48.045 146.375 ;
        RECT 71.880 146.360 75.980 146.510 ;
        RECT 47.715 146.060 75.980 146.360 ;
        RECT 47.715 146.045 48.045 146.060 ;
        RECT 71.880 145.910 75.980 146.060 ;
        RECT 29.210 143.455 31.190 143.785 ;
        RECT 59.210 143.455 61.190 143.785 ;
        RECT 71.880 143.400 75.980 143.550 ;
        RECT 62.370 143.100 75.980 143.400 ;
        RECT 57.795 142.660 58.125 142.675 ;
        RECT 62.370 142.660 62.670 143.100 ;
        RECT 71.880 142.950 75.980 143.100 ;
        RECT 57.795 142.360 62.670 142.660 ;
        RECT 57.795 142.345 58.125 142.360 ;
        RECT 14.210 140.125 16.190 140.455 ;
        RECT 44.210 140.125 46.190 140.455 ;
        RECT 65.955 140.440 66.285 140.455 ;
        RECT 71.880 140.440 75.980 140.590 ;
        RECT 65.955 140.140 75.980 140.440 ;
        RECT 65.955 140.125 66.285 140.140 ;
        RECT 71.880 139.990 75.980 140.140 ;
        RECT 63.555 137.480 63.885 137.495 ;
        RECT 71.880 137.480 75.980 137.630 ;
        RECT 63.555 137.180 75.980 137.480 ;
        RECT 63.555 137.165 63.885 137.180 ;
        RECT 29.210 136.795 31.190 137.125 ;
        RECT 59.210 136.795 61.190 137.125 ;
        RECT 71.880 137.030 75.980 137.180 ;
        RECT 66.435 134.520 66.765 134.535 ;
        RECT 71.880 134.520 75.980 134.670 ;
        RECT 66.435 134.220 75.980 134.520 ;
        RECT 66.435 134.205 66.765 134.220 ;
        RECT 71.880 134.070 75.980 134.220 ;
        RECT 14.210 133.465 16.190 133.795 ;
        RECT 44.210 133.465 46.190 133.795 ;
        RECT 66.915 131.560 67.245 131.575 ;
        RECT 71.880 131.560 75.980 131.710 ;
        RECT 66.915 131.260 75.980 131.560 ;
        RECT 66.915 131.245 67.245 131.260 ;
        RECT 71.880 131.110 75.980 131.260 ;
        RECT 29.210 130.135 31.190 130.465 ;
        RECT 59.210 130.135 61.190 130.465 ;
        RECT 69.315 128.600 69.645 128.615 ;
        RECT 71.880 128.600 75.980 128.750 ;
        RECT 69.315 128.300 75.980 128.600 ;
        RECT 69.315 128.285 69.645 128.300 ;
        RECT 71.880 128.150 75.980 128.300 ;
        RECT 14.210 126.805 16.190 127.135 ;
        RECT 44.210 126.805 46.190 127.135 ;
        RECT 66.915 125.640 67.245 125.655 ;
        RECT 71.880 125.640 75.980 125.790 ;
        RECT 66.915 125.340 75.980 125.640 ;
        RECT 66.915 125.325 67.245 125.340 ;
        RECT 71.880 125.190 75.980 125.340 ;
        RECT 29.210 123.475 31.190 123.805 ;
        RECT 59.210 123.475 61.190 123.805 ;
        RECT 64.035 122.680 64.365 122.695 ;
        RECT 71.880 122.680 75.980 122.830 ;
        RECT 64.035 122.380 75.980 122.680 ;
        RECT 64.035 122.365 64.365 122.380 ;
        RECT 71.880 122.230 75.980 122.380 ;
        RECT 14.210 120.145 16.190 120.475 ;
        RECT 44.210 120.145 46.190 120.475 ;
        RECT 66.915 119.720 67.245 119.735 ;
        RECT 71.880 119.720 75.980 119.870 ;
        RECT 66.915 119.420 75.980 119.720 ;
        RECT 66.915 119.405 67.245 119.420 ;
        RECT 71.880 119.270 75.980 119.420 ;
        RECT 29.210 116.815 31.190 117.145 ;
        RECT 59.210 116.815 61.190 117.145 ;
        RECT 66.915 116.760 67.245 116.775 ;
        RECT 71.880 116.760 75.980 116.910 ;
        RECT 66.915 116.460 75.980 116.760 ;
        RECT 66.915 116.445 67.245 116.460 ;
        RECT 71.880 116.310 75.980 116.460 ;
        RECT 30.435 116.020 30.765 116.035 ;
        RECT 70.275 116.020 70.605 116.035 ;
        RECT 30.435 115.720 70.605 116.020 ;
        RECT 30.435 115.705 30.765 115.720 ;
        RECT 70.275 115.705 70.605 115.720 ;
        RECT 14.210 113.485 16.190 113.815 ;
        RECT 44.210 113.485 46.190 113.815 ;
        RECT 68.835 113.800 69.165 113.815 ;
        RECT 71.880 113.800 75.980 113.950 ;
        RECT 68.835 113.500 75.980 113.800 ;
        RECT 68.835 113.485 69.165 113.500 ;
        RECT 71.880 113.350 75.980 113.500 ;
        RECT 66.915 110.840 67.245 110.855 ;
        RECT 71.880 110.840 75.980 110.990 ;
        RECT 66.915 110.540 75.980 110.840 ;
        RECT 66.915 110.525 67.245 110.540 ;
        RECT 29.210 110.155 31.190 110.485 ;
        RECT 59.210 110.155 61.190 110.485 ;
        RECT 71.880 110.390 75.980 110.540 ;
        RECT 65.955 107.880 66.285 107.895 ;
        RECT 71.880 107.880 75.980 108.030 ;
        RECT 65.955 107.580 75.980 107.880 ;
        RECT 65.955 107.565 66.285 107.580 ;
        RECT 71.880 107.430 75.980 107.580 ;
        RECT 14.210 106.825 16.190 107.155 ;
        RECT 44.210 106.825 46.190 107.155 ;
        RECT 64.035 104.920 64.365 104.935 ;
        RECT 71.880 104.920 75.980 105.070 ;
        RECT 64.035 104.620 75.980 104.920 ;
        RECT 64.035 104.605 64.365 104.620 ;
        RECT 71.880 104.470 75.980 104.620 ;
        RECT 29.210 103.495 31.190 103.825 ;
        RECT 59.210 103.495 61.190 103.825 ;
        RECT 66.915 101.960 67.245 101.975 ;
        RECT 71.880 101.960 75.980 102.110 ;
        RECT 66.915 101.660 75.980 101.960 ;
        RECT 66.915 101.645 67.245 101.660 ;
        RECT 71.880 101.510 75.980 101.660 ;
        RECT 14.210 100.165 16.190 100.495 ;
        RECT 44.210 100.165 46.190 100.495 ;
        RECT 61.155 99.000 61.485 99.015 ;
        RECT 71.880 99.000 75.980 99.150 ;
        RECT 61.155 98.700 75.980 99.000 ;
        RECT 61.155 98.685 61.485 98.700 ;
        RECT 71.880 98.550 75.980 98.700 ;
        RECT 29.210 96.835 31.190 97.165 ;
        RECT 59.210 96.835 61.190 97.165 ;
        RECT 66.915 96.040 67.245 96.055 ;
        RECT 71.880 96.040 75.980 96.190 ;
        RECT 66.915 95.740 75.980 96.040 ;
        RECT 66.915 95.725 67.245 95.740 ;
        RECT 71.880 95.590 75.980 95.740 ;
        RECT 14.210 93.505 16.190 93.835 ;
        RECT 44.210 93.505 46.190 93.835 ;
        RECT 68.835 93.080 69.165 93.095 ;
        RECT 71.880 93.080 75.980 93.230 ;
        RECT 68.835 92.780 75.980 93.080 ;
        RECT 68.835 92.765 69.165 92.780 ;
        RECT 71.880 92.630 75.980 92.780 ;
        RECT 29.210 90.175 31.190 90.505 ;
        RECT 59.210 90.175 61.190 90.505 ;
        RECT 66.915 90.120 67.245 90.135 ;
        RECT 71.880 90.120 75.980 90.270 ;
        RECT 66.915 89.820 75.980 90.120 ;
        RECT 66.915 89.805 67.245 89.820 ;
        RECT 71.880 89.670 75.980 89.820 ;
        RECT 14.210 86.845 16.190 87.175 ;
        RECT 44.210 86.845 46.190 87.175 ;
        RECT 65.955 87.160 66.285 87.175 ;
        RECT 71.880 87.160 75.980 87.310 ;
        RECT 65.955 86.860 75.980 87.160 ;
        RECT 65.955 86.845 66.285 86.860 ;
        RECT 71.880 86.710 75.980 86.860 ;
        RECT 61.635 84.200 61.965 84.215 ;
        RECT 71.880 84.200 75.980 84.350 ;
        RECT 61.635 83.900 75.980 84.200 ;
        RECT 61.635 83.885 61.965 83.900 ;
        RECT 29.210 83.515 31.190 83.845 ;
        RECT 59.210 83.515 61.190 83.845 ;
        RECT 71.880 83.750 75.980 83.900 ;
        RECT 54.435 81.240 54.765 81.255 ;
        RECT 71.880 81.240 75.980 81.390 ;
        RECT 54.435 80.940 75.980 81.240 ;
        RECT 54.435 80.925 54.765 80.940 ;
        RECT 71.880 80.790 75.980 80.940 ;
        RECT 55.875 78.280 56.205 78.295 ;
        RECT 71.880 78.280 75.980 78.430 ;
        RECT 55.875 77.980 75.980 78.280 ;
        RECT 55.875 77.965 56.205 77.980 ;
        RECT 71.880 77.830 75.980 77.980 ;
        RECT 53.475 75.320 53.805 75.335 ;
        RECT 71.880 75.320 75.980 75.470 ;
        RECT 53.475 75.020 75.980 75.320 ;
        RECT 53.475 75.005 53.805 75.020 ;
        RECT 71.880 74.870 75.980 75.020 ;
        RECT 91.700 73.025 92.100 154.800 ;
        RECT 91.650 72.575 92.150 73.025 ;
        RECT 39.950 71.500 40.450 71.525 ;
        RECT 83.115 71.500 83.615 71.525 ;
        RECT 39.950 71.100 83.615 71.500 ;
        RECT 39.950 71.075 40.450 71.100 ;
        RECT 83.115 71.075 83.615 71.100 ;
        RECT 12.050 70.400 12.650 70.425 ;
        RECT 93.635 70.400 94.235 70.425 ;
        RECT 12.050 69.900 94.235 70.400 ;
        RECT 12.050 69.875 12.650 69.900 ;
        RECT 93.635 69.875 94.235 69.900 ;
        RECT 72.250 68.500 73.150 68.525 ;
        RECT 3.950 67.700 73.150 68.500 ;
        RECT 72.250 67.675 73.150 67.700 ;
        RECT 79.455 51.590 79.835 52.020 ;
        RECT 81.275 51.590 81.655 52.020 ;
        RECT 79.480 45.955 79.810 51.590 ;
        RECT 81.300 45.955 81.630 51.590 ;
        RECT 71.250 41.800 72.150 41.825 ;
        RECT 0.950 41.000 72.150 41.800 ;
        RECT 97.195 41.795 97.715 222.720 ;
        RECT 165.465 219.200 169.325 221.600 ;
        RECT 170.525 219.200 174.385 221.600 ;
        RECT 175.585 219.200 179.445 221.600 ;
        RECT 180.645 219.200 184.505 221.600 ;
        RECT 185.705 219.200 189.565 221.600 ;
        RECT 190.765 219.200 194.625 221.600 ;
        RECT 195.825 219.200 199.685 221.600 ;
        RECT 200.885 219.200 204.745 221.600 ;
        RECT 205.945 219.200 209.805 221.600 ;
        RECT 211.005 219.200 214.865 221.600 ;
        RECT 216.065 219.200 219.925 221.600 ;
        RECT 221.125 219.200 224.985 221.600 ;
        RECT 226.185 219.200 230.045 221.600 ;
        RECT 231.245 219.200 235.105 221.600 ;
        RECT 236.305 219.200 240.165 221.600 ;
        RECT 243.365 219.200 247.225 221.600 ;
        RECT 250.425 219.200 254.285 221.600 ;
        RECT 255.485 219.200 259.345 221.600 ;
        RECT 260.545 219.200 264.405 221.600 ;
        RECT 265.605 219.200 269.465 221.600 ;
        RECT 270.665 219.200 274.525 221.600 ;
        RECT 275.725 219.200 279.585 221.600 ;
        RECT 280.785 219.200 284.645 221.600 ;
        RECT 285.845 219.200 289.705 221.600 ;
        RECT 290.905 219.200 294.765 221.600 ;
        RECT 295.965 219.200 299.825 221.600 ;
        RECT 301.025 219.200 304.885 221.600 ;
        RECT 306.085 219.200 309.945 221.600 ;
        RECT 311.145 219.200 315.005 221.600 ;
        RECT 316.205 219.200 320.065 221.600 ;
        RECT 321.265 219.200 325.125 221.600 ;
        RECT 326.325 219.200 330.185 221.600 ;
        RECT 165.465 215.600 169.325 218.000 ;
        RECT 170.525 215.600 174.385 218.000 ;
        RECT 175.585 215.600 179.445 218.000 ;
        RECT 180.645 215.600 184.505 218.000 ;
        RECT 185.705 215.600 189.565 218.000 ;
        RECT 190.765 215.600 194.625 218.000 ;
        RECT 195.825 215.600 199.685 218.000 ;
        RECT 200.885 215.600 204.745 218.000 ;
        RECT 205.945 215.600 209.805 218.000 ;
        RECT 211.005 215.600 214.865 218.000 ;
        RECT 216.065 215.600 219.925 218.000 ;
        RECT 221.125 215.600 224.985 218.000 ;
        RECT 226.185 215.600 230.045 218.000 ;
        RECT 231.245 215.600 235.105 218.000 ;
        RECT 236.305 215.600 240.165 218.000 ;
        RECT 243.365 215.600 247.225 218.000 ;
        RECT 250.425 215.600 254.285 218.000 ;
        RECT 255.485 215.600 259.345 218.000 ;
        RECT 260.545 215.600 264.405 218.000 ;
        RECT 265.605 215.600 269.465 218.000 ;
        RECT 270.665 215.600 274.525 218.000 ;
        RECT 275.725 215.600 279.585 218.000 ;
        RECT 280.785 215.600 284.645 218.000 ;
        RECT 285.845 215.600 289.705 218.000 ;
        RECT 290.905 215.600 294.765 218.000 ;
        RECT 295.965 215.600 299.825 218.000 ;
        RECT 301.025 215.600 304.885 218.000 ;
        RECT 306.085 215.600 309.945 218.000 ;
        RECT 311.145 215.600 315.005 218.000 ;
        RECT 316.205 215.600 320.065 218.000 ;
        RECT 321.265 215.600 325.125 218.000 ;
        RECT 326.325 215.600 330.185 218.000 ;
        RECT 165.465 212.000 169.325 214.400 ;
        RECT 170.525 212.000 174.385 214.400 ;
        RECT 175.585 212.000 179.445 214.400 ;
        RECT 180.645 212.000 184.505 214.400 ;
        RECT 185.705 212.000 189.565 214.400 ;
        RECT 190.765 212.000 194.625 214.400 ;
        RECT 195.825 212.000 199.685 214.400 ;
        RECT 200.885 212.000 204.745 214.400 ;
        RECT 205.945 212.000 209.805 214.400 ;
        RECT 211.005 212.000 214.865 214.400 ;
        RECT 216.065 212.000 219.925 214.400 ;
        RECT 221.125 212.000 224.985 214.400 ;
        RECT 226.185 212.000 230.045 214.400 ;
        RECT 231.245 212.000 235.105 214.400 ;
        RECT 236.305 212.000 240.165 214.400 ;
        RECT 241.475 214.375 242.055 214.905 ;
        RECT 243.365 212.000 247.225 214.400 ;
        RECT 248.535 214.375 249.115 214.905 ;
        RECT 250.425 212.000 254.285 214.400 ;
        RECT 255.485 212.000 259.345 214.400 ;
        RECT 260.545 212.000 264.405 214.400 ;
        RECT 265.605 212.000 269.465 214.400 ;
        RECT 270.665 212.000 274.525 214.400 ;
        RECT 275.725 212.000 279.585 214.400 ;
        RECT 280.785 212.000 284.645 214.400 ;
        RECT 285.845 212.000 289.705 214.400 ;
        RECT 290.905 212.000 294.765 214.400 ;
        RECT 295.965 212.000 299.825 214.400 ;
        RECT 301.025 212.000 304.885 214.400 ;
        RECT 306.085 212.000 309.945 214.400 ;
        RECT 311.145 212.000 315.005 214.400 ;
        RECT 316.205 212.000 320.065 214.400 ;
        RECT 321.265 212.000 325.125 214.400 ;
        RECT 326.325 212.000 330.185 214.400 ;
        RECT 138.050 210.475 138.850 211.225 ;
        RECT 165.465 208.400 169.325 210.800 ;
        RECT 170.525 208.400 174.385 210.800 ;
        RECT 175.585 208.400 179.445 210.800 ;
        RECT 180.645 208.400 184.505 210.800 ;
        RECT 185.705 208.400 189.565 210.800 ;
        RECT 190.765 208.400 194.625 210.800 ;
        RECT 195.825 208.400 199.685 210.800 ;
        RECT 200.885 208.400 204.745 210.800 ;
        RECT 205.945 208.400 209.805 210.800 ;
        RECT 211.005 208.400 214.865 210.800 ;
        RECT 216.065 208.400 219.925 210.800 ;
        RECT 221.125 208.400 224.985 210.800 ;
        RECT 226.185 208.400 230.045 210.800 ;
        RECT 231.245 208.400 235.105 210.800 ;
        RECT 236.305 208.400 240.165 210.800 ;
        RECT 243.365 208.400 247.225 210.800 ;
        RECT 250.425 208.400 254.285 210.800 ;
        RECT 255.485 208.400 259.345 210.800 ;
        RECT 260.545 208.400 264.405 210.800 ;
        RECT 265.605 208.400 269.465 210.800 ;
        RECT 270.665 208.400 274.525 210.800 ;
        RECT 275.725 208.400 279.585 210.800 ;
        RECT 280.785 208.400 284.645 210.800 ;
        RECT 285.845 208.400 289.705 210.800 ;
        RECT 290.905 208.400 294.765 210.800 ;
        RECT 295.965 208.400 299.825 210.800 ;
        RECT 301.025 208.400 304.885 210.800 ;
        RECT 306.085 208.400 309.945 210.800 ;
        RECT 311.145 208.400 315.005 210.800 ;
        RECT 316.205 208.400 320.065 210.800 ;
        RECT 321.265 208.400 325.125 210.800 ;
        RECT 326.325 208.400 330.185 210.800 ;
        RECT 165.465 204.800 169.325 207.200 ;
        RECT 170.525 204.800 174.385 207.200 ;
        RECT 175.585 204.800 179.445 207.200 ;
        RECT 180.645 204.800 184.505 207.200 ;
        RECT 185.705 204.800 189.565 207.200 ;
        RECT 190.765 204.800 194.625 207.200 ;
        RECT 195.825 204.800 199.685 207.200 ;
        RECT 200.885 204.800 204.745 207.200 ;
        RECT 205.945 204.800 209.805 207.200 ;
        RECT 211.005 204.800 214.865 207.200 ;
        RECT 216.065 204.800 219.925 207.200 ;
        RECT 221.125 204.800 224.985 207.200 ;
        RECT 226.185 204.800 230.045 207.200 ;
        RECT 231.245 204.800 235.105 207.200 ;
        RECT 236.305 204.800 240.165 207.200 ;
        RECT 243.365 204.800 247.225 207.200 ;
        RECT 250.425 204.800 254.285 207.200 ;
        RECT 255.485 204.800 259.345 207.200 ;
        RECT 260.545 204.800 264.405 207.200 ;
        RECT 265.605 204.800 269.465 207.200 ;
        RECT 270.665 204.800 274.525 207.200 ;
        RECT 275.725 204.800 279.585 207.200 ;
        RECT 280.785 204.800 284.645 207.200 ;
        RECT 285.845 204.800 289.705 207.200 ;
        RECT 290.905 204.800 294.765 207.200 ;
        RECT 295.965 204.800 299.825 207.200 ;
        RECT 301.025 204.800 304.885 207.200 ;
        RECT 306.085 204.800 309.945 207.200 ;
        RECT 311.145 204.800 315.005 207.200 ;
        RECT 316.205 204.800 320.065 207.200 ;
        RECT 321.265 204.800 325.125 207.200 ;
        RECT 326.325 204.800 330.185 207.200 ;
        RECT 165.465 201.200 169.325 203.600 ;
        RECT 170.525 201.200 174.385 203.600 ;
        RECT 175.585 201.200 179.445 203.600 ;
        RECT 180.645 201.200 184.505 203.600 ;
        RECT 185.705 201.200 189.565 203.600 ;
        RECT 190.765 201.200 194.625 203.600 ;
        RECT 195.825 201.200 199.685 203.600 ;
        RECT 200.885 201.200 204.745 203.600 ;
        RECT 205.945 201.200 209.805 203.600 ;
        RECT 211.005 201.200 214.865 203.600 ;
        RECT 216.065 201.200 219.925 203.600 ;
        RECT 221.125 201.200 224.985 203.600 ;
        RECT 226.185 201.200 230.045 203.600 ;
        RECT 231.245 201.200 235.105 203.600 ;
        RECT 236.305 201.200 240.165 203.600 ;
        RECT 241.475 203.575 242.055 204.105 ;
        RECT 243.365 201.200 247.225 203.600 ;
        RECT 248.535 203.575 249.115 204.105 ;
        RECT 250.425 201.200 254.285 203.600 ;
        RECT 255.485 201.200 259.345 203.600 ;
        RECT 260.545 201.200 264.405 203.600 ;
        RECT 265.605 201.200 269.465 203.600 ;
        RECT 270.665 201.200 274.525 203.600 ;
        RECT 275.725 201.200 279.585 203.600 ;
        RECT 280.785 201.200 284.645 203.600 ;
        RECT 285.845 201.200 289.705 203.600 ;
        RECT 290.905 201.200 294.765 203.600 ;
        RECT 295.965 201.200 299.825 203.600 ;
        RECT 301.025 201.200 304.885 203.600 ;
        RECT 306.085 201.200 309.945 203.600 ;
        RECT 311.145 201.200 315.005 203.600 ;
        RECT 316.205 201.200 320.065 203.600 ;
        RECT 321.265 201.200 325.125 203.600 ;
        RECT 326.325 201.200 330.185 203.600 ;
        RECT 165.465 197.600 169.325 200.000 ;
        RECT 170.525 197.600 174.385 200.000 ;
        RECT 175.585 197.600 179.445 200.000 ;
        RECT 180.645 197.600 184.505 200.000 ;
        RECT 185.705 197.600 189.565 200.000 ;
        RECT 190.765 197.600 194.625 200.000 ;
        RECT 195.825 197.600 199.685 200.000 ;
        RECT 200.885 197.600 204.745 200.000 ;
        RECT 205.945 197.600 209.805 200.000 ;
        RECT 211.005 197.600 214.865 200.000 ;
        RECT 216.065 197.600 219.925 200.000 ;
        RECT 221.125 197.600 224.985 200.000 ;
        RECT 226.185 197.600 230.045 200.000 ;
        RECT 231.245 197.600 235.105 200.000 ;
        RECT 236.305 197.600 240.165 200.000 ;
        RECT 241.475 199.975 242.055 200.505 ;
        RECT 243.365 197.600 247.225 200.000 ;
        RECT 248.535 199.975 249.115 200.505 ;
        RECT 250.425 197.600 254.285 200.000 ;
        RECT 255.485 197.600 259.345 200.000 ;
        RECT 260.545 197.600 264.405 200.000 ;
        RECT 265.605 197.600 269.465 200.000 ;
        RECT 270.665 197.600 274.525 200.000 ;
        RECT 275.725 197.600 279.585 200.000 ;
        RECT 280.785 197.600 284.645 200.000 ;
        RECT 285.845 197.600 289.705 200.000 ;
        RECT 290.905 197.600 294.765 200.000 ;
        RECT 295.965 197.600 299.825 200.000 ;
        RECT 301.025 197.600 304.885 200.000 ;
        RECT 306.085 197.600 309.945 200.000 ;
        RECT 311.145 197.600 315.005 200.000 ;
        RECT 316.205 197.600 320.065 200.000 ;
        RECT 321.265 197.600 325.125 200.000 ;
        RECT 326.325 197.600 330.185 200.000 ;
        RECT 165.465 194.000 169.325 196.400 ;
        RECT 170.525 194.000 174.385 196.400 ;
        RECT 175.585 194.000 179.445 196.400 ;
        RECT 180.645 194.000 184.505 196.400 ;
        RECT 185.705 194.000 189.565 196.400 ;
        RECT 190.765 194.000 194.625 196.400 ;
        RECT 195.825 194.000 199.685 196.400 ;
        RECT 200.885 194.000 204.745 196.400 ;
        RECT 205.945 194.000 209.805 196.400 ;
        RECT 211.005 194.000 214.865 196.400 ;
        RECT 216.065 194.000 219.925 196.400 ;
        RECT 221.125 194.000 224.985 196.400 ;
        RECT 226.185 194.000 230.045 196.400 ;
        RECT 231.245 194.000 235.105 196.400 ;
        RECT 236.305 194.000 240.165 196.400 ;
        RECT 241.475 194.035 242.055 194.565 ;
        RECT 243.365 194.000 247.225 196.400 ;
        RECT 248.535 195.835 249.115 196.365 ;
        RECT 250.425 194.000 254.285 196.400 ;
        RECT 255.485 194.000 259.345 196.400 ;
        RECT 260.545 194.000 264.405 196.400 ;
        RECT 265.605 194.000 269.465 196.400 ;
        RECT 270.665 194.000 274.525 196.400 ;
        RECT 275.725 194.000 279.585 196.400 ;
        RECT 280.785 194.000 284.645 196.400 ;
        RECT 285.845 194.000 289.705 196.400 ;
        RECT 290.905 194.000 294.765 196.400 ;
        RECT 295.965 194.000 299.825 196.400 ;
        RECT 301.025 194.000 304.885 196.400 ;
        RECT 306.085 194.000 309.945 196.400 ;
        RECT 311.145 194.000 315.005 196.400 ;
        RECT 316.205 194.000 320.065 196.400 ;
        RECT 321.265 194.000 325.125 196.400 ;
        RECT 326.325 194.000 330.185 196.400 ;
        RECT 165.465 190.400 169.325 192.800 ;
        RECT 170.525 190.400 174.385 192.800 ;
        RECT 175.585 190.400 179.445 192.800 ;
        RECT 180.645 190.400 184.505 192.800 ;
        RECT 185.705 190.400 189.565 192.800 ;
        RECT 190.765 190.400 194.625 192.800 ;
        RECT 195.825 190.400 199.685 192.800 ;
        RECT 200.885 190.400 204.745 192.800 ;
        RECT 205.945 190.400 209.805 192.800 ;
        RECT 211.005 190.400 214.865 192.800 ;
        RECT 216.065 190.400 219.925 192.800 ;
        RECT 221.125 190.400 224.985 192.800 ;
        RECT 226.185 190.400 230.045 192.800 ;
        RECT 231.245 190.400 235.105 192.800 ;
        RECT 236.305 190.400 240.165 192.800 ;
        RECT 241.475 192.235 242.055 192.765 ;
        RECT 243.365 190.400 247.225 192.800 ;
        RECT 248.535 190.435 249.115 190.965 ;
        RECT 250.425 190.400 254.285 192.800 ;
        RECT 255.485 190.400 259.345 192.800 ;
        RECT 260.545 190.400 264.405 192.800 ;
        RECT 265.605 190.400 269.465 192.800 ;
        RECT 270.665 190.400 274.525 192.800 ;
        RECT 275.725 190.400 279.585 192.800 ;
        RECT 280.785 190.400 284.645 192.800 ;
        RECT 285.845 190.400 289.705 192.800 ;
        RECT 290.905 190.400 294.765 192.800 ;
        RECT 295.965 190.400 299.825 192.800 ;
        RECT 301.025 190.400 304.885 192.800 ;
        RECT 306.085 190.400 309.945 192.800 ;
        RECT 311.145 190.400 315.005 192.800 ;
        RECT 316.205 190.400 320.065 192.800 ;
        RECT 321.265 190.400 325.125 192.800 ;
        RECT 326.325 190.400 330.185 192.800 ;
        RECT 165.465 186.800 169.325 189.200 ;
        RECT 170.525 186.800 174.385 189.200 ;
        RECT 175.585 186.800 179.445 189.200 ;
        RECT 180.645 186.800 184.505 189.200 ;
        RECT 185.705 186.800 189.565 189.200 ;
        RECT 190.765 186.800 194.625 189.200 ;
        RECT 195.825 186.800 199.685 189.200 ;
        RECT 200.885 186.800 204.745 189.200 ;
        RECT 205.945 186.800 209.805 189.200 ;
        RECT 211.005 186.800 214.865 189.200 ;
        RECT 216.065 186.800 219.925 189.200 ;
        RECT 221.125 186.800 224.985 189.200 ;
        RECT 226.185 186.800 230.045 189.200 ;
        RECT 231.245 186.800 235.105 189.200 ;
        RECT 236.305 186.800 240.165 189.200 ;
        RECT 241.475 189.175 242.055 189.705 ;
        RECT 243.365 186.800 247.225 189.200 ;
        RECT 248.535 189.175 249.115 189.705 ;
        RECT 250.425 186.800 254.285 189.200 ;
        RECT 255.485 186.800 259.345 189.200 ;
        RECT 260.545 186.800 264.405 189.200 ;
        RECT 265.605 186.800 269.465 189.200 ;
        RECT 270.665 186.800 274.525 189.200 ;
        RECT 275.725 186.800 279.585 189.200 ;
        RECT 280.785 186.800 284.645 189.200 ;
        RECT 285.845 186.800 289.705 189.200 ;
        RECT 290.905 186.800 294.765 189.200 ;
        RECT 295.965 186.800 299.825 189.200 ;
        RECT 301.025 186.800 304.885 189.200 ;
        RECT 306.085 186.800 309.945 189.200 ;
        RECT 311.145 186.800 315.005 189.200 ;
        RECT 316.205 186.800 320.065 189.200 ;
        RECT 321.265 186.800 325.125 189.200 ;
        RECT 326.325 186.800 330.185 189.200 ;
        RECT 165.465 183.200 169.325 185.600 ;
        RECT 170.525 183.200 174.385 185.600 ;
        RECT 175.585 183.200 179.445 185.600 ;
        RECT 180.645 183.200 184.505 185.600 ;
        RECT 185.705 183.200 189.565 185.600 ;
        RECT 190.765 183.200 194.625 185.600 ;
        RECT 195.825 183.200 199.685 185.600 ;
        RECT 200.885 183.200 204.745 185.600 ;
        RECT 205.945 183.200 209.805 185.600 ;
        RECT 211.005 183.200 214.865 185.600 ;
        RECT 216.065 183.200 219.925 185.600 ;
        RECT 221.125 183.200 224.985 185.600 ;
        RECT 226.185 183.200 230.045 185.600 ;
        RECT 231.245 183.200 235.105 185.600 ;
        RECT 236.305 183.200 240.165 185.600 ;
        RECT 243.365 183.200 247.225 185.600 ;
        RECT 250.425 183.200 254.285 185.600 ;
        RECT 255.485 183.200 259.345 185.600 ;
        RECT 260.545 183.200 264.405 185.600 ;
        RECT 265.605 183.200 269.465 185.600 ;
        RECT 270.665 183.200 274.525 185.600 ;
        RECT 275.725 183.200 279.585 185.600 ;
        RECT 280.785 183.200 284.645 185.600 ;
        RECT 285.845 183.200 289.705 185.600 ;
        RECT 290.905 183.200 294.765 185.600 ;
        RECT 295.965 183.200 299.825 185.600 ;
        RECT 301.025 183.200 304.885 185.600 ;
        RECT 306.085 183.200 309.945 185.600 ;
        RECT 311.145 183.200 315.005 185.600 ;
        RECT 316.205 183.200 320.065 185.600 ;
        RECT 321.265 183.200 325.125 185.600 ;
        RECT 326.325 183.200 330.185 185.600 ;
        RECT 165.465 179.600 169.325 182.000 ;
        RECT 170.525 179.600 174.385 182.000 ;
        RECT 175.585 179.600 179.445 182.000 ;
        RECT 180.645 179.600 184.505 182.000 ;
        RECT 185.705 179.600 189.565 182.000 ;
        RECT 190.765 179.600 194.625 182.000 ;
        RECT 195.825 179.600 199.685 182.000 ;
        RECT 200.885 179.600 204.745 182.000 ;
        RECT 205.945 179.600 209.805 182.000 ;
        RECT 211.005 179.600 214.865 182.000 ;
        RECT 216.065 179.600 219.925 182.000 ;
        RECT 221.125 179.600 224.985 182.000 ;
        RECT 226.185 179.600 230.045 182.000 ;
        RECT 231.245 179.600 235.105 182.000 ;
        RECT 236.305 179.600 240.165 182.000 ;
        RECT 241.475 181.975 242.055 182.505 ;
        RECT 243.365 179.600 247.225 182.000 ;
        RECT 248.535 181.975 249.115 182.505 ;
        RECT 250.425 179.600 254.285 182.000 ;
        RECT 255.485 179.600 259.345 182.000 ;
        RECT 260.545 179.600 264.405 182.000 ;
        RECT 265.605 179.600 269.465 182.000 ;
        RECT 270.665 179.600 274.525 182.000 ;
        RECT 275.725 179.600 279.585 182.000 ;
        RECT 280.785 179.600 284.645 182.000 ;
        RECT 285.845 179.600 289.705 182.000 ;
        RECT 290.905 179.600 294.765 182.000 ;
        RECT 295.965 179.600 299.825 182.000 ;
        RECT 301.025 179.600 304.885 182.000 ;
        RECT 306.085 179.600 309.945 182.000 ;
        RECT 311.145 179.600 315.005 182.000 ;
        RECT 316.205 179.600 320.065 182.000 ;
        RECT 321.265 179.600 325.125 182.000 ;
        RECT 326.325 179.600 330.185 182.000 ;
        RECT 165.465 176.000 169.325 178.400 ;
        RECT 170.525 176.000 174.385 178.400 ;
        RECT 175.585 176.000 179.445 178.400 ;
        RECT 180.645 176.000 184.505 178.400 ;
        RECT 185.705 176.000 189.565 178.400 ;
        RECT 190.765 176.000 194.625 178.400 ;
        RECT 195.825 176.000 199.685 178.400 ;
        RECT 200.885 176.000 204.745 178.400 ;
        RECT 205.945 176.000 209.805 178.400 ;
        RECT 211.005 176.000 214.865 178.400 ;
        RECT 216.065 176.000 219.925 178.400 ;
        RECT 221.125 176.000 224.985 178.400 ;
        RECT 226.185 176.000 230.045 178.400 ;
        RECT 231.245 176.000 235.105 178.400 ;
        RECT 236.305 176.000 240.165 178.400 ;
        RECT 243.365 176.000 247.225 178.400 ;
        RECT 250.425 176.000 254.285 178.400 ;
        RECT 255.485 176.000 259.345 178.400 ;
        RECT 260.545 176.000 264.405 178.400 ;
        RECT 265.605 176.000 269.465 178.400 ;
        RECT 270.665 176.000 274.525 178.400 ;
        RECT 275.725 176.000 279.585 178.400 ;
        RECT 280.785 176.000 284.645 178.400 ;
        RECT 285.845 176.000 289.705 178.400 ;
        RECT 290.905 176.000 294.765 178.400 ;
        RECT 295.965 176.000 299.825 178.400 ;
        RECT 301.025 176.000 304.885 178.400 ;
        RECT 306.085 176.000 309.945 178.400 ;
        RECT 311.145 176.000 315.005 178.400 ;
        RECT 316.205 176.000 320.065 178.400 ;
        RECT 321.265 176.000 325.125 178.400 ;
        RECT 326.325 176.000 330.185 178.400 ;
        RECT 165.465 172.400 169.325 174.800 ;
        RECT 170.525 172.400 174.385 174.800 ;
        RECT 175.585 172.400 179.445 174.800 ;
        RECT 180.645 172.400 184.505 174.800 ;
        RECT 185.705 172.400 189.565 174.800 ;
        RECT 190.765 172.400 194.625 174.800 ;
        RECT 195.825 172.400 199.685 174.800 ;
        RECT 200.885 172.400 204.745 174.800 ;
        RECT 205.945 172.400 209.805 174.800 ;
        RECT 211.005 172.400 214.865 174.800 ;
        RECT 216.065 172.400 219.925 174.800 ;
        RECT 221.125 172.400 224.985 174.800 ;
        RECT 226.185 172.400 230.045 174.800 ;
        RECT 231.245 172.400 235.105 174.800 ;
        RECT 236.305 172.400 240.165 174.800 ;
        RECT 243.365 172.400 247.225 174.800 ;
        RECT 250.425 172.400 254.285 174.800 ;
        RECT 255.485 172.400 259.345 174.800 ;
        RECT 260.545 172.400 264.405 174.800 ;
        RECT 265.605 172.400 269.465 174.800 ;
        RECT 270.665 172.400 274.525 174.800 ;
        RECT 275.725 172.400 279.585 174.800 ;
        RECT 280.785 172.400 284.645 174.800 ;
        RECT 285.845 172.400 289.705 174.800 ;
        RECT 290.905 172.400 294.765 174.800 ;
        RECT 295.965 172.400 299.825 174.800 ;
        RECT 301.025 172.400 304.885 174.800 ;
        RECT 306.085 172.400 309.945 174.800 ;
        RECT 311.145 172.400 315.005 174.800 ;
        RECT 316.205 172.400 320.065 174.800 ;
        RECT 321.265 172.400 325.125 174.800 ;
        RECT 326.325 172.400 330.185 174.800 ;
        RECT 165.465 168.800 169.325 171.200 ;
        RECT 170.525 168.800 174.385 171.200 ;
        RECT 175.585 168.800 179.445 171.200 ;
        RECT 180.645 168.800 184.505 171.200 ;
        RECT 185.705 168.800 189.565 171.200 ;
        RECT 190.765 168.800 194.625 171.200 ;
        RECT 195.825 168.800 199.685 171.200 ;
        RECT 200.885 168.800 204.745 171.200 ;
        RECT 205.945 168.800 209.805 171.200 ;
        RECT 211.005 168.800 214.865 171.200 ;
        RECT 216.065 168.800 219.925 171.200 ;
        RECT 221.125 168.800 224.985 171.200 ;
        RECT 226.185 168.800 230.045 171.200 ;
        RECT 231.245 168.800 235.105 171.200 ;
        RECT 236.305 168.800 240.165 171.200 ;
        RECT 241.475 171.175 242.055 171.705 ;
        RECT 243.365 168.800 247.225 171.200 ;
        RECT 248.535 171.175 249.115 171.705 ;
        RECT 250.425 168.800 254.285 171.200 ;
        RECT 255.485 168.800 259.345 171.200 ;
        RECT 260.545 168.800 264.405 171.200 ;
        RECT 265.605 168.800 269.465 171.200 ;
        RECT 270.665 168.800 274.525 171.200 ;
        RECT 275.725 168.800 279.585 171.200 ;
        RECT 280.785 168.800 284.645 171.200 ;
        RECT 285.845 168.800 289.705 171.200 ;
        RECT 290.905 168.800 294.765 171.200 ;
        RECT 295.965 168.800 299.825 171.200 ;
        RECT 301.025 168.800 304.885 171.200 ;
        RECT 306.085 168.800 309.945 171.200 ;
        RECT 311.145 168.800 315.005 171.200 ;
        RECT 316.205 168.800 320.065 171.200 ;
        RECT 321.265 168.800 325.125 171.200 ;
        RECT 326.325 168.800 330.185 171.200 ;
        RECT 165.465 165.200 169.325 167.600 ;
        RECT 170.525 165.200 174.385 167.600 ;
        RECT 175.585 165.200 179.445 167.600 ;
        RECT 180.645 165.200 184.505 167.600 ;
        RECT 185.705 165.200 189.565 167.600 ;
        RECT 190.765 165.200 194.625 167.600 ;
        RECT 195.825 165.200 199.685 167.600 ;
        RECT 200.885 165.200 204.745 167.600 ;
        RECT 205.945 165.200 209.805 167.600 ;
        RECT 211.005 165.200 214.865 167.600 ;
        RECT 216.065 165.200 219.925 167.600 ;
        RECT 221.125 165.200 224.985 167.600 ;
        RECT 226.185 165.200 230.045 167.600 ;
        RECT 231.245 165.200 235.105 167.600 ;
        RECT 236.305 165.200 240.165 167.600 ;
        RECT 243.365 165.200 247.225 167.600 ;
        RECT 250.425 165.200 254.285 167.600 ;
        RECT 255.485 165.200 259.345 167.600 ;
        RECT 260.545 165.200 264.405 167.600 ;
        RECT 265.605 165.200 269.465 167.600 ;
        RECT 270.665 165.200 274.525 167.600 ;
        RECT 275.725 165.200 279.585 167.600 ;
        RECT 280.785 165.200 284.645 167.600 ;
        RECT 285.845 165.200 289.705 167.600 ;
        RECT 290.905 165.200 294.765 167.600 ;
        RECT 295.965 165.200 299.825 167.600 ;
        RECT 301.025 165.200 304.885 167.600 ;
        RECT 306.085 165.200 309.945 167.600 ;
        RECT 311.145 165.200 315.005 167.600 ;
        RECT 316.205 165.200 320.065 167.600 ;
        RECT 321.265 165.200 325.125 167.600 ;
        RECT 326.325 165.200 330.185 167.600 ;
        RECT 200.835 162.655 201.455 163.225 ;
        RECT 290.855 162.655 291.475 163.225 ;
        RECT 221.075 161.615 221.695 162.185 ;
        RECT 270.615 161.615 271.235 162.185 ;
        RECT 231.195 160.575 231.815 161.145 ;
        RECT 260.495 160.575 261.115 161.145 ;
        RECT 236.255 159.535 236.875 160.105 ;
        RECT 255.435 159.535 256.055 160.105 ;
        RECT 118.695 149.215 119.205 149.815 ;
        RECT 118.720 129.450 119.180 149.215 ;
        RECT 134.950 135.645 135.350 151.740 ;
        RECT 142.705 149.215 143.215 149.815 ;
        RECT 134.925 135.145 135.375 135.645 ;
        RECT 142.730 129.450 143.190 149.215 ;
        RECT 158.960 135.645 159.360 151.740 ;
        RECT 166.715 149.215 167.225 149.815 ;
        RECT 158.935 135.145 159.385 135.645 ;
        RECT 166.740 129.450 167.200 149.215 ;
        RECT 182.970 135.645 183.370 151.740 ;
        RECT 190.725 149.215 191.235 149.815 ;
        RECT 182.945 135.145 183.395 135.645 ;
        RECT 190.750 129.450 191.210 149.215 ;
        RECT 206.980 135.645 207.380 151.740 ;
        RECT 214.735 149.215 215.245 149.815 ;
        RECT 206.955 135.145 207.405 135.645 ;
        RECT 214.760 129.450 215.220 149.215 ;
        RECT 230.990 135.645 231.390 151.740 ;
        RECT 238.750 149.215 239.260 149.815 ;
        RECT 230.965 135.145 231.415 135.645 ;
        RECT 238.775 129.450 239.235 149.215 ;
        RECT 255.005 135.645 255.405 151.740 ;
        RECT 262.805 149.215 263.315 149.815 ;
        RECT 254.980 135.145 255.430 135.645 ;
        RECT 262.830 129.450 263.290 149.215 ;
        RECT 279.060 135.645 279.460 151.740 ;
        RECT 286.765 149.215 287.275 149.815 ;
        RECT 279.035 135.145 279.485 135.645 ;
        RECT 286.790 129.450 287.250 149.215 ;
        RECT 303.020 135.645 303.420 151.740 ;
        RECT 310.775 149.215 311.285 149.815 ;
        RECT 302.995 135.145 303.445 135.645 ;
        RECT 310.800 129.450 311.260 149.215 ;
        RECT 327.030 135.645 327.430 151.740 ;
        RECT 327.005 135.145 327.455 135.645 ;
        RECT 118.695 128.850 119.205 129.450 ;
        RECT 142.705 128.850 143.215 129.450 ;
        RECT 166.715 128.850 167.225 129.450 ;
        RECT 190.725 128.850 191.235 129.450 ;
        RECT 214.735 128.850 215.245 129.450 ;
        RECT 238.750 128.850 239.260 129.450 ;
        RECT 262.805 128.850 263.315 129.450 ;
        RECT 286.765 128.850 287.275 129.450 ;
        RECT 310.775 128.850 311.285 129.450 ;
        RECT 113.750 126.400 114.350 126.900 ;
        RECT 113.800 125.425 114.300 126.400 ;
        RECT 113.750 124.875 114.350 125.425 ;
        RECT 137.760 124.875 138.360 125.900 ;
        RECT 161.770 124.875 162.370 125.425 ;
        RECT 185.780 123.375 186.380 123.925 ;
        RECT 209.790 122.375 210.390 122.925 ;
        RECT 233.800 121.375 234.400 121.925 ;
        RECT 257.810 120.375 258.410 120.925 ;
        RECT 281.820 119.375 282.420 119.925 ;
        RECT 305.830 118.375 306.430 118.925 ;
        RECT 112.750 117.375 113.350 117.925 ;
        RECT 136.760 116.375 137.360 116.925 ;
        RECT 160.770 115.375 161.370 115.925 ;
        RECT 184.780 114.375 185.380 114.925 ;
        RECT 208.790 113.375 209.390 113.925 ;
        RECT 232.800 112.375 233.400 112.925 ;
        RECT 256.810 111.375 257.410 111.925 ;
        RECT 280.820 110.375 281.420 110.925 ;
        RECT 304.830 109.375 305.430 109.925 ;
        RECT 113.750 108.375 114.350 108.925 ;
        RECT 137.760 107.375 138.360 107.925 ;
        RECT 161.770 106.375 162.370 106.925 ;
        RECT 185.780 105.375 186.380 105.925 ;
        RECT 209.790 104.375 210.390 104.925 ;
        RECT 233.800 103.375 234.400 103.925 ;
        RECT 257.810 102.375 258.410 102.925 ;
        RECT 281.820 101.875 282.420 102.425 ;
        RECT 305.830 101.875 306.430 102.425 ;
        RECT 118.695 97.850 119.205 98.450 ;
        RECT 142.705 97.850 143.215 98.450 ;
        RECT 166.715 97.850 167.225 98.450 ;
        RECT 190.725 97.850 191.235 98.450 ;
        RECT 214.735 97.850 215.245 98.450 ;
        RECT 238.750 97.850 239.260 98.450 ;
        RECT 262.805 97.850 263.315 98.450 ;
        RECT 286.765 97.850 287.275 98.450 ;
        RECT 310.775 97.850 311.285 98.450 ;
        RECT 109.400 96.825 110.400 97.775 ;
        RECT 118.720 78.085 119.180 97.850 ;
        RECT 134.925 91.655 135.375 92.155 ;
        RECT 118.695 77.485 119.205 78.085 ;
        RECT 134.950 75.560 135.350 91.655 ;
        RECT 142.730 78.085 143.190 97.850 ;
        RECT 158.935 91.655 159.385 92.155 ;
        RECT 142.705 77.485 143.215 78.085 ;
        RECT 158.960 75.560 159.360 91.655 ;
        RECT 166.740 78.085 167.200 97.850 ;
        RECT 182.945 91.655 183.395 92.155 ;
        RECT 166.715 77.485 167.225 78.085 ;
        RECT 182.970 75.560 183.370 91.655 ;
        RECT 190.750 78.085 191.210 97.850 ;
        RECT 206.955 91.655 207.405 92.155 ;
        RECT 190.725 77.485 191.235 78.085 ;
        RECT 206.980 75.560 207.380 91.655 ;
        RECT 214.760 78.085 215.220 97.850 ;
        RECT 230.965 91.655 231.415 92.155 ;
        RECT 214.735 77.485 215.245 78.085 ;
        RECT 230.990 75.560 231.390 91.655 ;
        RECT 238.775 78.085 239.235 97.850 ;
        RECT 254.980 91.655 255.430 92.155 ;
        RECT 238.750 77.485 239.260 78.085 ;
        RECT 255.005 75.560 255.405 91.655 ;
        RECT 262.830 78.085 263.290 97.850 ;
        RECT 279.035 91.655 279.485 92.155 ;
        RECT 262.805 77.485 263.315 78.085 ;
        RECT 279.060 75.560 279.460 91.655 ;
        RECT 286.790 78.085 287.250 97.850 ;
        RECT 302.995 91.655 303.445 92.155 ;
        RECT 286.765 77.485 287.275 78.085 ;
        RECT 303.020 75.560 303.420 91.655 ;
        RECT 310.800 78.085 311.260 97.850 ;
        RECT 327.005 91.655 327.455 92.155 ;
        RECT 310.775 77.485 311.285 78.085 ;
        RECT 327.030 75.560 327.430 91.655 ;
        RECT 236.255 67.195 236.875 67.765 ;
        RECT 255.435 67.195 256.055 67.765 ;
        RECT 231.195 66.155 231.815 66.725 ;
        RECT 260.495 66.155 261.115 66.725 ;
        RECT 221.075 65.115 221.695 65.685 ;
        RECT 270.615 65.115 271.235 65.685 ;
        RECT 200.835 64.075 201.455 64.645 ;
        RECT 290.855 64.075 291.475 64.645 ;
        RECT 165.465 59.700 169.325 62.100 ;
        RECT 170.525 59.700 174.385 62.100 ;
        RECT 175.585 59.700 179.445 62.100 ;
        RECT 180.645 59.700 184.505 62.100 ;
        RECT 185.705 59.700 189.565 62.100 ;
        RECT 190.765 59.700 194.625 62.100 ;
        RECT 195.825 59.700 199.685 62.100 ;
        RECT 200.885 59.700 204.745 62.100 ;
        RECT 205.945 59.700 209.805 62.100 ;
        RECT 211.005 59.700 214.865 62.100 ;
        RECT 216.065 59.700 219.925 62.100 ;
        RECT 221.125 59.700 224.985 62.100 ;
        RECT 226.185 59.700 230.045 62.100 ;
        RECT 231.245 59.700 235.105 62.100 ;
        RECT 236.305 59.700 240.165 62.100 ;
        RECT 243.365 59.700 247.225 62.100 ;
        RECT 250.425 59.700 254.285 62.100 ;
        RECT 255.485 59.700 259.345 62.100 ;
        RECT 260.545 59.700 264.405 62.100 ;
        RECT 265.605 59.700 269.465 62.100 ;
        RECT 270.665 59.700 274.525 62.100 ;
        RECT 275.725 59.700 279.585 62.100 ;
        RECT 280.785 59.700 284.645 62.100 ;
        RECT 285.845 59.700 289.705 62.100 ;
        RECT 290.905 59.700 294.765 62.100 ;
        RECT 295.965 59.700 299.825 62.100 ;
        RECT 301.025 59.700 304.885 62.100 ;
        RECT 306.085 59.700 309.945 62.100 ;
        RECT 311.145 59.700 315.005 62.100 ;
        RECT 316.205 59.700 320.065 62.100 ;
        RECT 321.265 59.700 325.125 62.100 ;
        RECT 326.325 59.700 330.185 62.100 ;
        RECT 165.465 56.100 169.325 58.500 ;
        RECT 170.525 56.100 174.385 58.500 ;
        RECT 175.585 56.100 179.445 58.500 ;
        RECT 180.645 56.100 184.505 58.500 ;
        RECT 185.705 56.100 189.565 58.500 ;
        RECT 190.765 56.100 194.625 58.500 ;
        RECT 195.825 56.100 199.685 58.500 ;
        RECT 200.885 56.100 204.745 58.500 ;
        RECT 205.945 56.100 209.805 58.500 ;
        RECT 211.005 56.100 214.865 58.500 ;
        RECT 216.065 56.100 219.925 58.500 ;
        RECT 221.125 56.100 224.985 58.500 ;
        RECT 226.185 56.100 230.045 58.500 ;
        RECT 231.245 56.100 235.105 58.500 ;
        RECT 236.305 56.100 240.165 58.500 ;
        RECT 241.475 55.595 242.055 56.125 ;
        RECT 243.365 56.100 247.225 58.500 ;
        RECT 248.535 55.595 249.115 56.125 ;
        RECT 250.425 56.100 254.285 58.500 ;
        RECT 255.485 56.100 259.345 58.500 ;
        RECT 260.545 56.100 264.405 58.500 ;
        RECT 265.605 56.100 269.465 58.500 ;
        RECT 270.665 56.100 274.525 58.500 ;
        RECT 275.725 56.100 279.585 58.500 ;
        RECT 280.785 56.100 284.645 58.500 ;
        RECT 285.845 56.100 289.705 58.500 ;
        RECT 290.905 56.100 294.765 58.500 ;
        RECT 295.965 56.100 299.825 58.500 ;
        RECT 301.025 56.100 304.885 58.500 ;
        RECT 306.085 56.100 309.945 58.500 ;
        RECT 311.145 56.100 315.005 58.500 ;
        RECT 316.205 56.100 320.065 58.500 ;
        RECT 321.265 56.100 325.125 58.500 ;
        RECT 326.325 56.100 330.185 58.500 ;
        RECT 165.465 52.500 169.325 54.900 ;
        RECT 170.525 52.500 174.385 54.900 ;
        RECT 175.585 52.500 179.445 54.900 ;
        RECT 180.645 52.500 184.505 54.900 ;
        RECT 185.705 52.500 189.565 54.900 ;
        RECT 190.765 52.500 194.625 54.900 ;
        RECT 195.825 52.500 199.685 54.900 ;
        RECT 200.885 52.500 204.745 54.900 ;
        RECT 205.945 52.500 209.805 54.900 ;
        RECT 211.005 52.500 214.865 54.900 ;
        RECT 216.065 52.500 219.925 54.900 ;
        RECT 221.125 52.500 224.985 54.900 ;
        RECT 226.185 52.500 230.045 54.900 ;
        RECT 231.245 52.500 235.105 54.900 ;
        RECT 236.305 52.500 240.165 54.900 ;
        RECT 243.365 52.500 247.225 54.900 ;
        RECT 250.425 52.500 254.285 54.900 ;
        RECT 255.485 52.500 259.345 54.900 ;
        RECT 260.545 52.500 264.405 54.900 ;
        RECT 265.605 52.500 269.465 54.900 ;
        RECT 270.665 52.500 274.525 54.900 ;
        RECT 275.725 52.500 279.585 54.900 ;
        RECT 280.785 52.500 284.645 54.900 ;
        RECT 285.845 52.500 289.705 54.900 ;
        RECT 290.905 52.500 294.765 54.900 ;
        RECT 295.965 52.500 299.825 54.900 ;
        RECT 301.025 52.500 304.885 54.900 ;
        RECT 306.085 52.500 309.945 54.900 ;
        RECT 311.145 52.500 315.005 54.900 ;
        RECT 316.205 52.500 320.065 54.900 ;
        RECT 321.265 52.500 325.125 54.900 ;
        RECT 326.325 52.500 330.185 54.900 ;
        RECT 165.465 48.900 169.325 51.300 ;
        RECT 170.525 48.900 174.385 51.300 ;
        RECT 175.585 48.900 179.445 51.300 ;
        RECT 180.645 48.900 184.505 51.300 ;
        RECT 185.705 48.900 189.565 51.300 ;
        RECT 190.765 48.900 194.625 51.300 ;
        RECT 195.825 48.900 199.685 51.300 ;
        RECT 200.885 48.900 204.745 51.300 ;
        RECT 205.945 48.900 209.805 51.300 ;
        RECT 211.005 48.900 214.865 51.300 ;
        RECT 216.065 48.900 219.925 51.300 ;
        RECT 221.125 48.900 224.985 51.300 ;
        RECT 226.185 48.900 230.045 51.300 ;
        RECT 231.245 48.900 235.105 51.300 ;
        RECT 236.305 48.900 240.165 51.300 ;
        RECT 243.365 48.900 247.225 51.300 ;
        RECT 250.425 48.900 254.285 51.300 ;
        RECT 255.485 48.900 259.345 51.300 ;
        RECT 260.545 48.900 264.405 51.300 ;
        RECT 265.605 48.900 269.465 51.300 ;
        RECT 270.665 48.900 274.525 51.300 ;
        RECT 275.725 48.900 279.585 51.300 ;
        RECT 280.785 48.900 284.645 51.300 ;
        RECT 285.845 48.900 289.705 51.300 ;
        RECT 290.905 48.900 294.765 51.300 ;
        RECT 295.965 48.900 299.825 51.300 ;
        RECT 301.025 48.900 304.885 51.300 ;
        RECT 306.085 48.900 309.945 51.300 ;
        RECT 311.145 48.900 315.005 51.300 ;
        RECT 316.205 48.900 320.065 51.300 ;
        RECT 321.265 48.900 325.125 51.300 ;
        RECT 326.325 48.900 330.185 51.300 ;
        RECT 165.465 45.300 169.325 47.700 ;
        RECT 170.525 45.300 174.385 47.700 ;
        RECT 175.585 45.300 179.445 47.700 ;
        RECT 180.645 45.300 184.505 47.700 ;
        RECT 185.705 45.300 189.565 47.700 ;
        RECT 190.765 45.300 194.625 47.700 ;
        RECT 195.825 45.300 199.685 47.700 ;
        RECT 200.885 45.300 204.745 47.700 ;
        RECT 205.945 45.300 209.805 47.700 ;
        RECT 211.005 45.300 214.865 47.700 ;
        RECT 216.065 45.300 219.925 47.700 ;
        RECT 221.125 45.300 224.985 47.700 ;
        RECT 226.185 45.300 230.045 47.700 ;
        RECT 231.245 45.300 235.105 47.700 ;
        RECT 236.305 45.300 240.165 47.700 ;
        RECT 241.475 44.795 242.055 45.325 ;
        RECT 243.365 45.300 247.225 47.700 ;
        RECT 248.535 44.795 249.115 45.325 ;
        RECT 250.425 45.300 254.285 47.700 ;
        RECT 255.485 45.300 259.345 47.700 ;
        RECT 260.545 45.300 264.405 47.700 ;
        RECT 265.605 45.300 269.465 47.700 ;
        RECT 270.665 45.300 274.525 47.700 ;
        RECT 275.725 45.300 279.585 47.700 ;
        RECT 280.785 45.300 284.645 47.700 ;
        RECT 285.845 45.300 289.705 47.700 ;
        RECT 290.905 45.300 294.765 47.700 ;
        RECT 295.965 45.300 299.825 47.700 ;
        RECT 301.025 45.300 304.885 47.700 ;
        RECT 306.085 45.300 309.945 47.700 ;
        RECT 311.145 45.300 315.005 47.700 ;
        RECT 316.205 45.300 320.065 47.700 ;
        RECT 321.265 45.300 325.125 47.700 ;
        RECT 326.325 45.300 330.185 47.700 ;
        RECT 97.145 41.225 97.765 41.795 ;
        RECT 165.465 41.700 169.325 44.100 ;
        RECT 170.525 41.700 174.385 44.100 ;
        RECT 175.585 41.700 179.445 44.100 ;
        RECT 180.645 41.700 184.505 44.100 ;
        RECT 185.705 41.700 189.565 44.100 ;
        RECT 190.765 41.700 194.625 44.100 ;
        RECT 195.825 41.700 199.685 44.100 ;
        RECT 200.885 41.700 204.745 44.100 ;
        RECT 205.945 41.700 209.805 44.100 ;
        RECT 211.005 41.700 214.865 44.100 ;
        RECT 216.065 41.700 219.925 44.100 ;
        RECT 221.125 41.700 224.985 44.100 ;
        RECT 226.185 41.700 230.045 44.100 ;
        RECT 231.245 41.700 235.105 44.100 ;
        RECT 236.305 41.700 240.165 44.100 ;
        RECT 243.365 41.700 247.225 44.100 ;
        RECT 250.425 41.700 254.285 44.100 ;
        RECT 255.485 41.700 259.345 44.100 ;
        RECT 260.545 41.700 264.405 44.100 ;
        RECT 265.605 41.700 269.465 44.100 ;
        RECT 270.665 41.700 274.525 44.100 ;
        RECT 275.725 41.700 279.585 44.100 ;
        RECT 280.785 41.700 284.645 44.100 ;
        RECT 285.845 41.700 289.705 44.100 ;
        RECT 290.905 41.700 294.765 44.100 ;
        RECT 295.965 41.700 299.825 44.100 ;
        RECT 301.025 41.700 304.885 44.100 ;
        RECT 306.085 41.700 309.945 44.100 ;
        RECT 311.145 41.700 315.005 44.100 ;
        RECT 316.205 41.700 320.065 44.100 ;
        RECT 321.265 41.700 325.125 44.100 ;
        RECT 326.325 41.700 330.185 44.100 ;
        RECT 71.250 40.975 72.150 41.000 ;
        RECT 63.505 40.440 64.125 40.465 ;
        RECT 63.505 39.920 162.930 40.440 ;
        RECT 63.505 39.895 64.125 39.920 ;
        RECT 55.600 39.560 56.190 39.585 ;
        RECT 104.930 39.560 105.520 39.585 ;
        RECT 55.600 39.070 105.520 39.560 ;
        RECT 55.600 39.045 56.190 39.070 ;
        RECT 104.930 39.045 105.520 39.070 ;
        RECT 56.600 37.190 57.590 37.520 ;
        RECT 103.530 37.190 104.520 37.520 ;
        RECT 3.955 35.720 6.050 36.250 ;
        RECT 18.635 28.605 21.035 32.465 ;
        RECT 22.235 28.605 24.635 32.465 ;
        RECT 25.835 28.605 28.235 32.465 ;
        RECT 29.435 28.605 31.835 32.465 ;
        RECT 33.035 28.605 35.435 32.465 ;
        RECT 36.635 28.605 39.035 32.465 ;
        RECT 40.235 28.605 42.635 32.465 ;
        RECT 43.835 28.605 46.235 32.465 ;
        RECT 50.530 29.130 50.910 29.435 ;
        RECT 47.880 28.610 50.910 29.130 ;
        RECT 50.530 28.305 50.910 28.610 ;
        RECT 18.635 23.545 21.035 27.405 ;
        RECT 22.235 23.545 24.635 27.405 ;
        RECT 25.835 23.545 28.235 27.405 ;
        RECT 29.435 23.545 31.835 27.405 ;
        RECT 33.035 23.545 35.435 27.405 ;
        RECT 36.635 23.545 39.035 27.405 ;
        RECT 40.235 23.545 42.635 27.405 ;
        RECT 43.835 23.545 46.235 27.405 ;
        RECT 18.635 18.485 21.035 22.345 ;
        RECT 22.235 18.485 24.635 22.345 ;
        RECT 25.835 18.485 28.235 22.345 ;
        RECT 29.435 18.485 31.835 22.345 ;
        RECT 33.035 18.485 35.435 22.345 ;
        RECT 36.635 18.485 39.035 22.345 ;
        RECT 40.235 18.485 42.635 22.345 ;
        RECT 43.835 18.485 46.235 22.345 ;
        RECT 18.635 13.425 21.035 17.285 ;
        RECT 22.235 13.425 24.635 17.285 ;
        RECT 25.835 13.425 28.235 17.285 ;
        RECT 29.435 13.425 31.835 17.285 ;
        RECT 33.035 13.425 35.435 17.285 ;
        RECT 36.635 13.425 39.035 17.285 ;
        RECT 40.235 13.425 42.635 17.285 ;
        RECT 43.835 13.425 46.235 17.285 ;
        RECT 49.000 15.245 49.620 16.595 ;
        RECT 56.930 16.305 57.260 37.190 ;
        RECT 58.000 36.225 58.580 36.250 ;
        RECT 102.540 36.225 103.120 36.250 ;
        RECT 58.000 35.745 103.120 36.225 ;
        RECT 58.000 35.720 58.580 35.745 ;
        RECT 102.540 35.720 103.120 35.745 ;
        RECT 80.270 33.825 80.850 34.305 ;
        RECT 67.270 26.515 76.330 27.845 ;
        RECT 50.995 15.975 57.570 16.305 ;
        RECT 67.320 6.975 68.600 26.515 ;
        RECT 69.880 6.975 71.160 26.515 ;
        RECT 72.440 6.975 73.720 26.515 ;
        RECT 75.000 6.975 76.280 26.515 ;
        RECT 0.950 5.650 3.050 6.180 ;
        RECT 67.270 5.645 76.330 6.975 ;
        RECT 80.320 6.180 80.800 33.825 ;
        RECT 84.790 26.515 93.850 27.845 ;
        RECT 84.840 6.975 86.120 26.515 ;
        RECT 87.400 6.975 88.680 26.515 ;
        RECT 89.960 6.975 91.240 26.515 ;
        RECT 92.520 6.975 93.800 26.515 ;
        RECT 103.860 16.305 104.190 37.190 ;
        RECT 110.210 29.130 110.590 29.435 ;
        RECT 110.210 28.610 113.240 29.130 ;
        RECT 110.210 28.305 110.590 28.610 ;
        RECT 114.885 28.605 117.285 32.465 ;
        RECT 118.485 28.605 120.885 32.465 ;
        RECT 122.085 28.605 124.485 32.465 ;
        RECT 125.685 28.605 128.085 32.465 ;
        RECT 129.285 28.605 131.685 32.465 ;
        RECT 132.885 28.605 135.285 32.465 ;
        RECT 136.485 28.605 138.885 32.465 ;
        RECT 140.085 28.605 142.485 32.465 ;
        RECT 114.885 23.545 117.285 27.405 ;
        RECT 118.485 23.545 120.885 27.405 ;
        RECT 122.085 23.545 124.485 27.405 ;
        RECT 125.685 23.545 128.085 27.405 ;
        RECT 129.285 23.545 131.685 27.405 ;
        RECT 132.885 23.545 135.285 27.405 ;
        RECT 136.485 23.545 138.885 27.405 ;
        RECT 140.085 23.545 142.485 27.405 ;
        RECT 114.885 18.485 117.285 22.345 ;
        RECT 118.485 18.485 120.885 22.345 ;
        RECT 122.085 18.485 124.485 22.345 ;
        RECT 125.685 18.485 128.085 22.345 ;
        RECT 129.285 18.485 131.685 22.345 ;
        RECT 132.885 18.485 135.285 22.345 ;
        RECT 136.485 18.485 138.885 22.345 ;
        RECT 140.085 18.485 142.485 22.345 ;
        RECT 103.550 15.975 110.125 16.305 ;
        RECT 111.500 15.245 112.120 16.595 ;
        RECT 114.885 13.425 117.285 17.285 ;
        RECT 118.485 13.425 120.885 17.285 ;
        RECT 122.085 13.425 124.485 17.285 ;
        RECT 125.685 13.425 128.085 17.285 ;
        RECT 129.285 13.425 131.685 17.285 ;
        RECT 132.885 13.425 135.285 17.285 ;
        RECT 136.485 13.425 138.885 17.285 ;
        RECT 140.085 13.425 142.485 17.285 ;
        RECT 80.270 5.650 80.850 6.180 ;
        RECT 84.790 5.645 93.850 6.975 ;
        RECT 162.410 4.580 162.930 39.920 ;
        RECT 165.465 38.100 169.325 40.500 ;
        RECT 170.525 38.100 174.385 40.500 ;
        RECT 175.585 38.100 179.445 40.500 ;
        RECT 180.645 38.100 184.505 40.500 ;
        RECT 185.705 38.100 189.565 40.500 ;
        RECT 190.765 38.100 194.625 40.500 ;
        RECT 195.825 38.100 199.685 40.500 ;
        RECT 200.885 38.100 204.745 40.500 ;
        RECT 205.945 38.100 209.805 40.500 ;
        RECT 211.005 38.100 214.865 40.500 ;
        RECT 216.065 38.100 219.925 40.500 ;
        RECT 221.125 38.100 224.985 40.500 ;
        RECT 226.185 38.100 230.045 40.500 ;
        RECT 231.245 38.100 235.105 40.500 ;
        RECT 236.305 38.100 240.165 40.500 ;
        RECT 241.475 37.595 242.055 38.125 ;
        RECT 243.365 38.100 247.225 40.500 ;
        RECT 248.535 37.595 249.115 38.125 ;
        RECT 250.425 38.100 254.285 40.500 ;
        RECT 255.485 38.100 259.345 40.500 ;
        RECT 260.545 38.100 264.405 40.500 ;
        RECT 265.605 38.100 269.465 40.500 ;
        RECT 270.665 38.100 274.525 40.500 ;
        RECT 275.725 38.100 279.585 40.500 ;
        RECT 280.785 38.100 284.645 40.500 ;
        RECT 285.845 38.100 289.705 40.500 ;
        RECT 290.905 38.100 294.765 40.500 ;
        RECT 295.965 38.100 299.825 40.500 ;
        RECT 301.025 38.100 304.885 40.500 ;
        RECT 306.085 38.100 309.945 40.500 ;
        RECT 311.145 38.100 315.005 40.500 ;
        RECT 316.205 38.100 320.065 40.500 ;
        RECT 321.265 38.100 325.125 40.500 ;
        RECT 326.325 38.100 330.185 40.500 ;
        RECT 165.465 34.500 169.325 36.900 ;
        RECT 170.525 34.500 174.385 36.900 ;
        RECT 175.585 34.500 179.445 36.900 ;
        RECT 180.645 34.500 184.505 36.900 ;
        RECT 185.705 34.500 189.565 36.900 ;
        RECT 190.765 34.500 194.625 36.900 ;
        RECT 195.825 34.500 199.685 36.900 ;
        RECT 200.885 34.500 204.745 36.900 ;
        RECT 205.945 34.500 209.805 36.900 ;
        RECT 211.005 34.500 214.865 36.900 ;
        RECT 216.065 34.500 219.925 36.900 ;
        RECT 221.125 34.500 224.985 36.900 ;
        RECT 226.185 34.500 230.045 36.900 ;
        RECT 231.245 34.500 235.105 36.900 ;
        RECT 236.305 34.500 240.165 36.900 ;
        RECT 241.475 34.535 242.055 35.065 ;
        RECT 243.365 34.500 247.225 36.900 ;
        RECT 248.535 36.335 249.115 36.865 ;
        RECT 250.425 34.500 254.285 36.900 ;
        RECT 255.485 34.500 259.345 36.900 ;
        RECT 260.545 34.500 264.405 36.900 ;
        RECT 265.605 34.500 269.465 36.900 ;
        RECT 270.665 34.500 274.525 36.900 ;
        RECT 275.725 34.500 279.585 36.900 ;
        RECT 280.785 34.500 284.645 36.900 ;
        RECT 285.845 34.500 289.705 36.900 ;
        RECT 290.905 34.500 294.765 36.900 ;
        RECT 295.965 34.500 299.825 36.900 ;
        RECT 301.025 34.500 304.885 36.900 ;
        RECT 306.085 34.500 309.945 36.900 ;
        RECT 311.145 34.500 315.005 36.900 ;
        RECT 316.205 34.500 320.065 36.900 ;
        RECT 321.265 34.500 325.125 36.900 ;
        RECT 326.325 34.500 330.185 36.900 ;
        RECT 165.465 30.900 169.325 33.300 ;
        RECT 170.525 30.900 174.385 33.300 ;
        RECT 175.585 30.900 179.445 33.300 ;
        RECT 180.645 30.900 184.505 33.300 ;
        RECT 185.705 30.900 189.565 33.300 ;
        RECT 190.765 30.900 194.625 33.300 ;
        RECT 195.825 30.900 199.685 33.300 ;
        RECT 200.885 30.900 204.745 33.300 ;
        RECT 205.945 30.900 209.805 33.300 ;
        RECT 211.005 30.900 214.865 33.300 ;
        RECT 216.065 30.900 219.925 33.300 ;
        RECT 221.125 30.900 224.985 33.300 ;
        RECT 226.185 30.900 230.045 33.300 ;
        RECT 231.245 30.900 235.105 33.300 ;
        RECT 236.305 30.900 240.165 33.300 ;
        RECT 241.475 32.735 242.055 33.265 ;
        RECT 243.365 30.900 247.225 33.300 ;
        RECT 248.535 30.935 249.115 31.465 ;
        RECT 250.425 30.900 254.285 33.300 ;
        RECT 255.485 30.900 259.345 33.300 ;
        RECT 260.545 30.900 264.405 33.300 ;
        RECT 265.605 30.900 269.465 33.300 ;
        RECT 270.665 30.900 274.525 33.300 ;
        RECT 275.725 30.900 279.585 33.300 ;
        RECT 280.785 30.900 284.645 33.300 ;
        RECT 285.845 30.900 289.705 33.300 ;
        RECT 290.905 30.900 294.765 33.300 ;
        RECT 295.965 30.900 299.825 33.300 ;
        RECT 301.025 30.900 304.885 33.300 ;
        RECT 306.085 30.900 309.945 33.300 ;
        RECT 311.145 30.900 315.005 33.300 ;
        RECT 316.205 30.900 320.065 33.300 ;
        RECT 321.265 30.900 325.125 33.300 ;
        RECT 326.325 30.900 330.185 33.300 ;
        RECT 165.465 27.300 169.325 29.700 ;
        RECT 170.525 27.300 174.385 29.700 ;
        RECT 175.585 27.300 179.445 29.700 ;
        RECT 180.645 27.300 184.505 29.700 ;
        RECT 185.705 27.300 189.565 29.700 ;
        RECT 190.765 27.300 194.625 29.700 ;
        RECT 195.825 27.300 199.685 29.700 ;
        RECT 200.885 27.300 204.745 29.700 ;
        RECT 205.945 27.300 209.805 29.700 ;
        RECT 211.005 27.300 214.865 29.700 ;
        RECT 216.065 27.300 219.925 29.700 ;
        RECT 221.125 27.300 224.985 29.700 ;
        RECT 226.185 27.300 230.045 29.700 ;
        RECT 231.245 27.300 235.105 29.700 ;
        RECT 236.305 27.300 240.165 29.700 ;
        RECT 241.475 26.795 242.055 27.325 ;
        RECT 243.365 27.300 247.225 29.700 ;
        RECT 248.535 26.795 249.115 27.325 ;
        RECT 250.425 27.300 254.285 29.700 ;
        RECT 255.485 27.300 259.345 29.700 ;
        RECT 260.545 27.300 264.405 29.700 ;
        RECT 265.605 27.300 269.465 29.700 ;
        RECT 270.665 27.300 274.525 29.700 ;
        RECT 275.725 27.300 279.585 29.700 ;
        RECT 280.785 27.300 284.645 29.700 ;
        RECT 285.845 27.300 289.705 29.700 ;
        RECT 290.905 27.300 294.765 29.700 ;
        RECT 295.965 27.300 299.825 29.700 ;
        RECT 301.025 27.300 304.885 29.700 ;
        RECT 306.085 27.300 309.945 29.700 ;
        RECT 311.145 27.300 315.005 29.700 ;
        RECT 316.205 27.300 320.065 29.700 ;
        RECT 321.265 27.300 325.125 29.700 ;
        RECT 326.325 27.300 330.185 29.700 ;
        RECT 165.465 23.700 169.325 26.100 ;
        RECT 170.525 23.700 174.385 26.100 ;
        RECT 175.585 23.700 179.445 26.100 ;
        RECT 180.645 23.700 184.505 26.100 ;
        RECT 185.705 23.700 189.565 26.100 ;
        RECT 190.765 23.700 194.625 26.100 ;
        RECT 195.825 23.700 199.685 26.100 ;
        RECT 200.885 23.700 204.745 26.100 ;
        RECT 205.945 23.700 209.805 26.100 ;
        RECT 211.005 23.700 214.865 26.100 ;
        RECT 216.065 23.700 219.925 26.100 ;
        RECT 221.125 23.700 224.985 26.100 ;
        RECT 226.185 23.700 230.045 26.100 ;
        RECT 231.245 23.700 235.105 26.100 ;
        RECT 236.305 23.700 240.165 26.100 ;
        RECT 241.475 23.195 242.055 23.725 ;
        RECT 243.365 23.700 247.225 26.100 ;
        RECT 248.535 23.195 249.115 23.725 ;
        RECT 250.425 23.700 254.285 26.100 ;
        RECT 255.485 23.700 259.345 26.100 ;
        RECT 260.545 23.700 264.405 26.100 ;
        RECT 265.605 23.700 269.465 26.100 ;
        RECT 270.665 23.700 274.525 26.100 ;
        RECT 275.725 23.700 279.585 26.100 ;
        RECT 280.785 23.700 284.645 26.100 ;
        RECT 285.845 23.700 289.705 26.100 ;
        RECT 290.905 23.700 294.765 26.100 ;
        RECT 295.965 23.700 299.825 26.100 ;
        RECT 301.025 23.700 304.885 26.100 ;
        RECT 306.085 23.700 309.945 26.100 ;
        RECT 311.145 23.700 315.005 26.100 ;
        RECT 316.205 23.700 320.065 26.100 ;
        RECT 321.265 23.700 325.125 26.100 ;
        RECT 326.325 23.700 330.185 26.100 ;
        RECT 165.465 20.100 169.325 22.500 ;
        RECT 170.525 20.100 174.385 22.500 ;
        RECT 175.585 20.100 179.445 22.500 ;
        RECT 180.645 20.100 184.505 22.500 ;
        RECT 185.705 20.100 189.565 22.500 ;
        RECT 190.765 20.100 194.625 22.500 ;
        RECT 195.825 20.100 199.685 22.500 ;
        RECT 200.885 20.100 204.745 22.500 ;
        RECT 205.945 20.100 209.805 22.500 ;
        RECT 211.005 20.100 214.865 22.500 ;
        RECT 216.065 20.100 219.925 22.500 ;
        RECT 221.125 20.100 224.985 22.500 ;
        RECT 226.185 20.100 230.045 22.500 ;
        RECT 231.245 20.100 235.105 22.500 ;
        RECT 236.305 20.100 240.165 22.500 ;
        RECT 243.365 20.100 247.225 22.500 ;
        RECT 250.425 20.100 254.285 22.500 ;
        RECT 255.485 20.100 259.345 22.500 ;
        RECT 260.545 20.100 264.405 22.500 ;
        RECT 265.605 20.100 269.465 22.500 ;
        RECT 270.665 20.100 274.525 22.500 ;
        RECT 275.725 20.100 279.585 22.500 ;
        RECT 280.785 20.100 284.645 22.500 ;
        RECT 285.845 20.100 289.705 22.500 ;
        RECT 290.905 20.100 294.765 22.500 ;
        RECT 295.965 20.100 299.825 22.500 ;
        RECT 301.025 20.100 304.885 22.500 ;
        RECT 306.085 20.100 309.945 22.500 ;
        RECT 311.145 20.100 315.005 22.500 ;
        RECT 316.205 20.100 320.065 22.500 ;
        RECT 321.265 20.100 325.125 22.500 ;
        RECT 326.325 20.100 330.185 22.500 ;
        RECT 165.465 16.500 169.325 18.900 ;
        RECT 170.525 16.500 174.385 18.900 ;
        RECT 175.585 16.500 179.445 18.900 ;
        RECT 180.645 16.500 184.505 18.900 ;
        RECT 185.705 16.500 189.565 18.900 ;
        RECT 190.765 16.500 194.625 18.900 ;
        RECT 195.825 16.500 199.685 18.900 ;
        RECT 200.885 16.500 204.745 18.900 ;
        RECT 205.945 16.500 209.805 18.900 ;
        RECT 211.005 16.500 214.865 18.900 ;
        RECT 216.065 16.500 219.925 18.900 ;
        RECT 221.125 16.500 224.985 18.900 ;
        RECT 226.185 16.500 230.045 18.900 ;
        RECT 231.245 16.500 235.105 18.900 ;
        RECT 236.305 16.500 240.165 18.900 ;
        RECT 243.365 16.500 247.225 18.900 ;
        RECT 250.425 16.500 254.285 18.900 ;
        RECT 255.485 16.500 259.345 18.900 ;
        RECT 260.545 16.500 264.405 18.900 ;
        RECT 265.605 16.500 269.465 18.900 ;
        RECT 270.665 16.500 274.525 18.900 ;
        RECT 275.725 16.500 279.585 18.900 ;
        RECT 280.785 16.500 284.645 18.900 ;
        RECT 285.845 16.500 289.705 18.900 ;
        RECT 290.905 16.500 294.765 18.900 ;
        RECT 295.965 16.500 299.825 18.900 ;
        RECT 301.025 16.500 304.885 18.900 ;
        RECT 306.085 16.500 309.945 18.900 ;
        RECT 311.145 16.500 315.005 18.900 ;
        RECT 316.205 16.500 320.065 18.900 ;
        RECT 321.265 16.500 325.125 18.900 ;
        RECT 326.325 16.500 330.185 18.900 ;
        RECT 165.465 12.900 169.325 15.300 ;
        RECT 170.525 12.900 174.385 15.300 ;
        RECT 175.585 12.900 179.445 15.300 ;
        RECT 180.645 12.900 184.505 15.300 ;
        RECT 185.705 12.900 189.565 15.300 ;
        RECT 190.765 12.900 194.625 15.300 ;
        RECT 195.825 12.900 199.685 15.300 ;
        RECT 200.885 12.900 204.745 15.300 ;
        RECT 205.945 12.900 209.805 15.300 ;
        RECT 211.005 12.900 214.865 15.300 ;
        RECT 216.065 12.900 219.925 15.300 ;
        RECT 221.125 12.900 224.985 15.300 ;
        RECT 226.185 12.900 230.045 15.300 ;
        RECT 231.245 12.900 235.105 15.300 ;
        RECT 236.305 12.900 240.165 15.300 ;
        RECT 241.475 12.395 242.055 12.925 ;
        RECT 243.365 12.900 247.225 15.300 ;
        RECT 248.535 12.395 249.115 12.925 ;
        RECT 250.425 12.900 254.285 15.300 ;
        RECT 255.485 12.900 259.345 15.300 ;
        RECT 260.545 12.900 264.405 15.300 ;
        RECT 265.605 12.900 269.465 15.300 ;
        RECT 270.665 12.900 274.525 15.300 ;
        RECT 275.725 12.900 279.585 15.300 ;
        RECT 280.785 12.900 284.645 15.300 ;
        RECT 285.845 12.900 289.705 15.300 ;
        RECT 290.905 12.900 294.765 15.300 ;
        RECT 295.965 12.900 299.825 15.300 ;
        RECT 301.025 12.900 304.885 15.300 ;
        RECT 306.085 12.900 309.945 15.300 ;
        RECT 311.145 12.900 315.005 15.300 ;
        RECT 316.205 12.900 320.065 15.300 ;
        RECT 321.265 12.900 325.125 15.300 ;
        RECT 326.325 12.900 330.185 15.300 ;
        RECT 165.465 9.300 169.325 11.700 ;
        RECT 170.525 9.300 174.385 11.700 ;
        RECT 175.585 9.300 179.445 11.700 ;
        RECT 180.645 9.300 184.505 11.700 ;
        RECT 185.705 9.300 189.565 11.700 ;
        RECT 190.765 9.300 194.625 11.700 ;
        RECT 195.825 9.300 199.685 11.700 ;
        RECT 200.885 9.300 204.745 11.700 ;
        RECT 205.945 9.300 209.805 11.700 ;
        RECT 211.005 9.300 214.865 11.700 ;
        RECT 216.065 9.300 219.925 11.700 ;
        RECT 221.125 9.300 224.985 11.700 ;
        RECT 226.185 9.300 230.045 11.700 ;
        RECT 231.245 9.300 235.105 11.700 ;
        RECT 236.305 9.300 240.165 11.700 ;
        RECT 243.365 9.300 247.225 11.700 ;
        RECT 250.425 9.300 254.285 11.700 ;
        RECT 255.485 9.300 259.345 11.700 ;
        RECT 260.545 9.300 264.405 11.700 ;
        RECT 265.605 9.300 269.465 11.700 ;
        RECT 270.665 9.300 274.525 11.700 ;
        RECT 275.725 9.300 279.585 11.700 ;
        RECT 280.785 9.300 284.645 11.700 ;
        RECT 285.845 9.300 289.705 11.700 ;
        RECT 290.905 9.300 294.765 11.700 ;
        RECT 295.965 9.300 299.825 11.700 ;
        RECT 301.025 9.300 304.885 11.700 ;
        RECT 306.085 9.300 309.945 11.700 ;
        RECT 311.145 9.300 315.005 11.700 ;
        RECT 316.205 9.300 320.065 11.700 ;
        RECT 321.265 9.300 325.125 11.700 ;
        RECT 326.325 9.300 330.185 11.700 ;
        RECT 165.465 5.700 169.325 8.100 ;
        RECT 170.525 5.700 174.385 8.100 ;
        RECT 175.585 5.700 179.445 8.100 ;
        RECT 180.645 5.700 184.505 8.100 ;
        RECT 185.705 5.700 189.565 8.100 ;
        RECT 190.765 5.700 194.625 8.100 ;
        RECT 195.825 5.700 199.685 8.100 ;
        RECT 200.885 5.700 204.745 8.100 ;
        RECT 205.945 5.700 209.805 8.100 ;
        RECT 211.005 5.700 214.865 8.100 ;
        RECT 216.065 5.700 219.925 8.100 ;
        RECT 221.125 5.700 224.985 8.100 ;
        RECT 226.185 5.700 230.045 8.100 ;
        RECT 231.245 5.700 235.105 8.100 ;
        RECT 236.305 5.700 240.165 8.100 ;
        RECT 243.365 5.700 247.225 8.100 ;
        RECT 250.425 5.700 254.285 8.100 ;
        RECT 255.485 5.700 259.345 8.100 ;
        RECT 260.545 5.700 264.405 8.100 ;
        RECT 265.605 5.700 269.465 8.100 ;
        RECT 270.665 5.700 274.525 8.100 ;
        RECT 275.725 5.700 279.585 8.100 ;
        RECT 280.785 5.700 284.645 8.100 ;
        RECT 285.845 5.700 289.705 8.100 ;
        RECT 290.905 5.700 294.765 8.100 ;
        RECT 295.965 5.700 299.825 8.100 ;
        RECT 301.025 5.700 304.885 8.100 ;
        RECT 306.085 5.700 309.945 8.100 ;
        RECT 311.145 5.700 315.005 8.100 ;
        RECT 316.205 5.700 320.065 8.100 ;
        RECT 321.265 5.700 325.125 8.100 ;
        RECT 326.325 5.700 330.185 8.100 ;
        RECT 162.410 4.060 167.785 4.580 ;
        RECT 134.530 -5.675 135.110 -5.145 ;
      LAYER met4 ;
        RECT 134.575 232.950 135.065 232.955 ;
        RECT 134.575 232.470 136.440 232.950 ;
        RECT 134.575 232.465 135.065 232.470 ;
        RECT 30.670 219.215 30.970 224.760 ;
        RECT 33.430 219.215 33.730 224.760 ;
        RECT 36.190 219.215 36.490 224.760 ;
        RECT 38.950 219.215 39.250 224.760 ;
        RECT 41.710 219.215 42.010 224.760 ;
        RECT 44.470 219.215 44.770 224.760 ;
        RECT 47.230 222.305 47.530 224.760 ;
        RECT 49.990 222.305 50.290 224.760 ;
        RECT 47.095 221.795 47.605 222.305 ;
        RECT 49.895 221.795 50.405 222.305 ;
        RECT 52.750 219.215 53.050 224.760 ;
        RECT 55.510 219.215 55.810 224.760 ;
        RECT 58.270 219.215 58.570 224.760 ;
        RECT 61.030 219.215 61.330 224.760 ;
        RECT 63.790 219.215 64.090 224.760 ;
        RECT 66.550 219.215 66.850 224.760 ;
        RECT 6.000 217.215 66.850 219.215 ;
        RECT 0.995 213.120 1.000 215.130 ;
        RECT 3.000 213.120 3.005 215.130 ;
        RECT 8.265 210.595 8.775 211.105 ;
        RECT 0.995 163.795 1.000 165.805 ;
        RECT 3.000 163.795 3.005 165.805 ;
        RECT 3.995 159.795 4.000 161.805 ;
        RECT 6.000 159.795 6.005 161.805 ;
        RECT 8.370 157.005 8.670 210.595 ;
        RECT 69.310 205.900 69.610 224.760 ;
        RECT 14.125 205.600 69.610 205.900 ;
        RECT 14.125 157.005 14.425 205.600 ;
        RECT 72.070 202.455 72.370 224.760 ;
        RECT 19.890 202.155 72.370 202.455 ;
        RECT 19.890 157.005 20.190 202.155 ;
        RECT 74.830 199.160 75.130 224.760 ;
        RECT 25.650 198.860 75.130 199.160 ;
        RECT 25.650 157.005 25.950 198.860 ;
        RECT 77.590 196.200 77.890 224.760 ;
        RECT 31.410 195.900 77.890 196.200 ;
        RECT 31.410 157.005 31.710 195.900 ;
        RECT 80.350 193.165 80.650 224.760 ;
        RECT 37.170 192.865 80.650 193.165 ;
        RECT 37.170 157.005 37.470 192.865 ;
        RECT 83.110 190.300 83.410 224.760 ;
        RECT 42.930 190.000 83.410 190.300 ;
        RECT 42.930 157.005 43.230 190.000 ;
        RECT 85.870 187.780 86.170 224.760 ;
        RECT 48.690 187.480 86.170 187.780 ;
        RECT 48.690 157.005 48.990 187.480 ;
        RECT 88.630 185.855 88.930 224.760 ;
        RECT 54.450 185.555 88.930 185.855 ;
        RECT 54.450 157.005 54.750 185.555 ;
        RECT 91.390 183.790 91.690 224.760 ;
        RECT 60.210 183.490 91.690 183.790 ;
        RECT 60.210 157.005 60.510 183.490 ;
        RECT 94.150 182.200 94.450 224.760 ;
        RECT 138.310 211.205 138.610 224.760 ;
        RECT 138.095 210.495 138.805 211.205 ;
        RECT 65.970 181.900 94.450 182.200 ;
        RECT 65.970 157.005 66.270 181.900 ;
        RECT 143.830 169.835 144.130 224.760 ;
        RECT 167.210 223.240 167.740 223.245 ;
        RECT 317.525 223.240 318.045 223.390 ;
        RECT 165.215 222.720 330.185 223.240 ;
        RECT 167.210 222.715 167.740 222.720 ;
        RECT 71.730 169.535 144.130 169.835 ;
        RECT 71.730 157.005 72.030 169.535 ;
        RECT 165.465 164.080 165.985 222.200 ;
        RECT 167.865 221.205 168.385 222.720 ;
        RECT 167.320 219.595 168.930 221.205 ;
        RECT 167.865 217.605 168.385 219.595 ;
        RECT 167.320 215.995 168.930 217.605 ;
        RECT 167.865 214.005 168.385 215.995 ;
        RECT 167.320 212.395 168.930 214.005 ;
        RECT 167.865 210.405 168.385 212.395 ;
        RECT 167.320 208.795 168.930 210.405 ;
        RECT 167.865 206.805 168.385 208.795 ;
        RECT 167.320 205.195 168.930 206.805 ;
        RECT 167.865 203.205 168.385 205.195 ;
        RECT 167.320 201.595 168.930 203.205 ;
        RECT 167.865 199.605 168.385 201.595 ;
        RECT 167.320 197.995 168.930 199.605 ;
        RECT 167.865 196.005 168.385 197.995 ;
        RECT 167.320 194.395 168.930 196.005 ;
        RECT 167.865 192.405 168.385 194.395 ;
        RECT 167.320 190.795 168.930 192.405 ;
        RECT 167.865 188.805 168.385 190.795 ;
        RECT 167.320 187.195 168.930 188.805 ;
        RECT 167.865 185.205 168.385 187.195 ;
        RECT 167.320 183.595 168.930 185.205 ;
        RECT 167.865 181.605 168.385 183.595 ;
        RECT 167.320 179.995 168.930 181.605 ;
        RECT 167.865 178.005 168.385 179.995 ;
        RECT 167.320 176.395 168.930 178.005 ;
        RECT 167.865 174.405 168.385 176.395 ;
        RECT 167.320 172.795 168.930 174.405 ;
        RECT 167.865 170.805 168.385 172.795 ;
        RECT 167.320 169.195 168.930 170.805 ;
        RECT 167.865 167.205 168.385 169.195 ;
        RECT 167.320 165.595 168.930 167.205 ;
        RECT 167.865 164.600 168.385 165.595 ;
        RECT 170.525 164.080 171.045 222.200 ;
        RECT 172.925 221.205 173.445 222.720 ;
        RECT 172.380 219.595 173.990 221.205 ;
        RECT 172.925 217.605 173.445 219.595 ;
        RECT 172.380 215.995 173.990 217.605 ;
        RECT 172.925 214.005 173.445 215.995 ;
        RECT 172.380 212.395 173.990 214.005 ;
        RECT 172.925 210.405 173.445 212.395 ;
        RECT 172.380 208.795 173.990 210.405 ;
        RECT 172.925 206.805 173.445 208.795 ;
        RECT 172.380 205.195 173.990 206.805 ;
        RECT 172.925 203.205 173.445 205.195 ;
        RECT 172.380 201.595 173.990 203.205 ;
        RECT 172.925 199.605 173.445 201.595 ;
        RECT 172.380 197.995 173.990 199.605 ;
        RECT 172.925 196.005 173.445 197.995 ;
        RECT 172.380 194.395 173.990 196.005 ;
        RECT 172.925 192.405 173.445 194.395 ;
        RECT 172.380 190.795 173.990 192.405 ;
        RECT 172.925 188.805 173.445 190.795 ;
        RECT 172.380 187.195 173.990 188.805 ;
        RECT 172.925 185.205 173.445 187.195 ;
        RECT 172.380 183.595 173.990 185.205 ;
        RECT 172.925 181.605 173.445 183.595 ;
        RECT 172.380 179.995 173.990 181.605 ;
        RECT 172.925 178.005 173.445 179.995 ;
        RECT 172.380 176.395 173.990 178.005 ;
        RECT 172.925 174.405 173.445 176.395 ;
        RECT 172.380 172.795 173.990 174.405 ;
        RECT 172.925 170.805 173.445 172.795 ;
        RECT 172.380 169.195 173.990 170.805 ;
        RECT 172.925 167.205 173.445 169.195 ;
        RECT 172.380 165.595 173.990 167.205 ;
        RECT 172.925 164.600 173.445 165.595 ;
        RECT 175.585 164.080 176.105 222.200 ;
        RECT 177.985 221.205 178.505 222.720 ;
        RECT 177.440 219.595 179.050 221.205 ;
        RECT 177.985 217.605 178.505 219.595 ;
        RECT 177.440 215.995 179.050 217.605 ;
        RECT 177.985 214.005 178.505 215.995 ;
        RECT 177.440 212.395 179.050 214.005 ;
        RECT 177.985 210.405 178.505 212.395 ;
        RECT 177.440 208.795 179.050 210.405 ;
        RECT 177.985 206.805 178.505 208.795 ;
        RECT 177.440 205.195 179.050 206.805 ;
        RECT 177.985 203.205 178.505 205.195 ;
        RECT 177.440 201.595 179.050 203.205 ;
        RECT 177.985 199.605 178.505 201.595 ;
        RECT 177.440 197.995 179.050 199.605 ;
        RECT 177.985 196.005 178.505 197.995 ;
        RECT 177.440 194.395 179.050 196.005 ;
        RECT 177.985 192.405 178.505 194.395 ;
        RECT 177.440 190.795 179.050 192.405 ;
        RECT 177.985 188.805 178.505 190.795 ;
        RECT 177.440 187.195 179.050 188.805 ;
        RECT 177.985 185.205 178.505 187.195 ;
        RECT 177.440 183.595 179.050 185.205 ;
        RECT 177.985 181.605 178.505 183.595 ;
        RECT 177.440 179.995 179.050 181.605 ;
        RECT 177.985 178.005 178.505 179.995 ;
        RECT 177.440 176.395 179.050 178.005 ;
        RECT 177.985 174.405 178.505 176.395 ;
        RECT 177.440 172.795 179.050 174.405 ;
        RECT 177.985 170.805 178.505 172.795 ;
        RECT 177.440 169.195 179.050 170.805 ;
        RECT 177.985 167.205 178.505 169.195 ;
        RECT 177.440 165.595 179.050 167.205 ;
        RECT 177.985 164.600 178.505 165.595 ;
        RECT 180.645 164.080 181.165 222.200 ;
        RECT 183.045 221.205 183.565 222.720 ;
        RECT 182.500 219.595 184.110 221.205 ;
        RECT 183.045 217.605 183.565 219.595 ;
        RECT 182.500 215.995 184.110 217.605 ;
        RECT 183.045 214.005 183.565 215.995 ;
        RECT 182.500 212.395 184.110 214.005 ;
        RECT 183.045 210.405 183.565 212.395 ;
        RECT 182.500 208.795 184.110 210.405 ;
        RECT 183.045 206.805 183.565 208.795 ;
        RECT 182.500 205.195 184.110 206.805 ;
        RECT 183.045 203.205 183.565 205.195 ;
        RECT 182.500 201.595 184.110 203.205 ;
        RECT 183.045 199.605 183.565 201.595 ;
        RECT 182.500 197.995 184.110 199.605 ;
        RECT 183.045 196.005 183.565 197.995 ;
        RECT 182.500 194.395 184.110 196.005 ;
        RECT 183.045 192.405 183.565 194.395 ;
        RECT 182.500 190.795 184.110 192.405 ;
        RECT 183.045 188.805 183.565 190.795 ;
        RECT 182.500 187.195 184.110 188.805 ;
        RECT 183.045 185.205 183.565 187.195 ;
        RECT 182.500 183.595 184.110 185.205 ;
        RECT 183.045 181.605 183.565 183.595 ;
        RECT 182.500 179.995 184.110 181.605 ;
        RECT 183.045 178.005 183.565 179.995 ;
        RECT 182.500 176.395 184.110 178.005 ;
        RECT 183.045 174.405 183.565 176.395 ;
        RECT 182.500 172.795 184.110 174.405 ;
        RECT 183.045 170.805 183.565 172.795 ;
        RECT 182.500 169.195 184.110 170.805 ;
        RECT 183.045 167.205 183.565 169.195 ;
        RECT 182.500 165.595 184.110 167.205 ;
        RECT 183.045 164.600 183.565 165.595 ;
        RECT 185.705 164.080 186.225 222.200 ;
        RECT 188.105 221.205 188.625 222.720 ;
        RECT 187.560 219.595 189.170 221.205 ;
        RECT 188.105 217.605 188.625 219.595 ;
        RECT 187.560 215.995 189.170 217.605 ;
        RECT 188.105 214.005 188.625 215.995 ;
        RECT 187.560 212.395 189.170 214.005 ;
        RECT 188.105 210.405 188.625 212.395 ;
        RECT 187.560 208.795 189.170 210.405 ;
        RECT 188.105 206.805 188.625 208.795 ;
        RECT 187.560 205.195 189.170 206.805 ;
        RECT 188.105 203.205 188.625 205.195 ;
        RECT 187.560 201.595 189.170 203.205 ;
        RECT 188.105 199.605 188.625 201.595 ;
        RECT 187.560 197.995 189.170 199.605 ;
        RECT 188.105 196.005 188.625 197.995 ;
        RECT 187.560 194.395 189.170 196.005 ;
        RECT 188.105 192.405 188.625 194.395 ;
        RECT 187.560 190.795 189.170 192.405 ;
        RECT 188.105 188.805 188.625 190.795 ;
        RECT 187.560 187.195 189.170 188.805 ;
        RECT 188.105 185.205 188.625 187.195 ;
        RECT 187.560 183.595 189.170 185.205 ;
        RECT 188.105 181.605 188.625 183.595 ;
        RECT 187.560 179.995 189.170 181.605 ;
        RECT 188.105 178.005 188.625 179.995 ;
        RECT 187.560 176.395 189.170 178.005 ;
        RECT 188.105 174.405 188.625 176.395 ;
        RECT 187.560 172.795 189.170 174.405 ;
        RECT 188.105 170.805 188.625 172.795 ;
        RECT 187.560 169.195 189.170 170.805 ;
        RECT 188.105 167.205 188.625 169.195 ;
        RECT 187.560 165.595 189.170 167.205 ;
        RECT 188.105 164.600 188.625 165.595 ;
        RECT 190.765 164.080 191.285 222.200 ;
        RECT 193.165 221.205 193.685 222.720 ;
        RECT 192.620 219.595 194.230 221.205 ;
        RECT 193.165 217.605 193.685 219.595 ;
        RECT 192.620 215.995 194.230 217.605 ;
        RECT 193.165 214.005 193.685 215.995 ;
        RECT 192.620 212.395 194.230 214.005 ;
        RECT 193.165 210.405 193.685 212.395 ;
        RECT 192.620 208.795 194.230 210.405 ;
        RECT 193.165 206.805 193.685 208.795 ;
        RECT 192.620 205.195 194.230 206.805 ;
        RECT 193.165 203.205 193.685 205.195 ;
        RECT 192.620 201.595 194.230 203.205 ;
        RECT 193.165 199.605 193.685 201.595 ;
        RECT 192.620 197.995 194.230 199.605 ;
        RECT 193.165 196.005 193.685 197.995 ;
        RECT 192.620 194.395 194.230 196.005 ;
        RECT 193.165 192.405 193.685 194.395 ;
        RECT 192.620 190.795 194.230 192.405 ;
        RECT 193.165 188.805 193.685 190.795 ;
        RECT 192.620 187.195 194.230 188.805 ;
        RECT 193.165 185.205 193.685 187.195 ;
        RECT 192.620 183.595 194.230 185.205 ;
        RECT 193.165 181.605 193.685 183.595 ;
        RECT 192.620 179.995 194.230 181.605 ;
        RECT 193.165 178.005 193.685 179.995 ;
        RECT 192.620 176.395 194.230 178.005 ;
        RECT 193.165 174.405 193.685 176.395 ;
        RECT 192.620 172.795 194.230 174.405 ;
        RECT 193.165 170.805 193.685 172.795 ;
        RECT 192.620 169.195 194.230 170.805 ;
        RECT 193.165 167.205 193.685 169.195 ;
        RECT 192.620 165.595 194.230 167.205 ;
        RECT 193.165 164.600 193.685 165.595 ;
        RECT 195.825 164.080 196.345 222.200 ;
        RECT 198.225 221.205 198.745 222.720 ;
        RECT 197.680 219.595 199.290 221.205 ;
        RECT 198.225 217.605 198.745 219.595 ;
        RECT 197.680 215.995 199.290 217.605 ;
        RECT 198.225 214.005 198.745 215.995 ;
        RECT 197.680 212.395 199.290 214.005 ;
        RECT 198.225 210.405 198.745 212.395 ;
        RECT 197.680 208.795 199.290 210.405 ;
        RECT 198.225 206.805 198.745 208.795 ;
        RECT 197.680 205.195 199.290 206.805 ;
        RECT 198.225 203.205 198.745 205.195 ;
        RECT 197.680 201.595 199.290 203.205 ;
        RECT 198.225 199.605 198.745 201.595 ;
        RECT 197.680 197.995 199.290 199.605 ;
        RECT 198.225 196.005 198.745 197.995 ;
        RECT 197.680 194.395 199.290 196.005 ;
        RECT 198.225 192.405 198.745 194.395 ;
        RECT 197.680 190.795 199.290 192.405 ;
        RECT 198.225 188.805 198.745 190.795 ;
        RECT 197.680 187.195 199.290 188.805 ;
        RECT 198.225 185.205 198.745 187.195 ;
        RECT 197.680 183.595 199.290 185.205 ;
        RECT 198.225 181.605 198.745 183.595 ;
        RECT 197.680 179.995 199.290 181.605 ;
        RECT 198.225 178.005 198.745 179.995 ;
        RECT 197.680 176.395 199.290 178.005 ;
        RECT 198.225 174.405 198.745 176.395 ;
        RECT 197.680 172.795 199.290 174.405 ;
        RECT 198.225 170.805 198.745 172.795 ;
        RECT 197.680 169.195 199.290 170.805 ;
        RECT 198.225 167.205 198.745 169.195 ;
        RECT 197.680 165.595 199.290 167.205 ;
        RECT 198.225 164.600 198.745 165.595 ;
        RECT 200.885 164.080 201.405 222.200 ;
        RECT 203.285 221.205 203.805 222.720 ;
        RECT 202.740 219.595 204.350 221.205 ;
        RECT 203.285 217.605 203.805 219.595 ;
        RECT 202.740 215.995 204.350 217.605 ;
        RECT 203.285 214.005 203.805 215.995 ;
        RECT 202.740 212.395 204.350 214.005 ;
        RECT 203.285 210.405 203.805 212.395 ;
        RECT 202.740 208.795 204.350 210.405 ;
        RECT 203.285 206.805 203.805 208.795 ;
        RECT 202.740 205.195 204.350 206.805 ;
        RECT 203.285 203.205 203.805 205.195 ;
        RECT 202.740 201.595 204.350 203.205 ;
        RECT 203.285 199.605 203.805 201.595 ;
        RECT 202.740 197.995 204.350 199.605 ;
        RECT 203.285 196.005 203.805 197.995 ;
        RECT 202.740 194.395 204.350 196.005 ;
        RECT 203.285 192.405 203.805 194.395 ;
        RECT 202.740 190.795 204.350 192.405 ;
        RECT 203.285 188.805 203.805 190.795 ;
        RECT 202.740 187.195 204.350 188.805 ;
        RECT 203.285 185.205 203.805 187.195 ;
        RECT 202.740 183.595 204.350 185.205 ;
        RECT 203.285 181.605 203.805 183.595 ;
        RECT 202.740 179.995 204.350 181.605 ;
        RECT 203.285 178.005 203.805 179.995 ;
        RECT 202.740 176.395 204.350 178.005 ;
        RECT 203.285 174.405 203.805 176.395 ;
        RECT 202.740 172.795 204.350 174.405 ;
        RECT 203.285 170.805 203.805 172.795 ;
        RECT 202.740 169.195 204.350 170.805 ;
        RECT 203.285 167.205 203.805 169.195 ;
        RECT 202.740 165.595 204.350 167.205 ;
        RECT 203.285 164.600 203.805 165.595 ;
        RECT 165.465 163.560 201.405 164.080 ;
        RECT 205.945 164.080 206.465 222.200 ;
        RECT 208.345 221.205 208.865 222.720 ;
        RECT 207.800 219.595 209.410 221.205 ;
        RECT 208.345 217.605 208.865 219.595 ;
        RECT 207.800 215.995 209.410 217.605 ;
        RECT 208.345 214.005 208.865 215.995 ;
        RECT 207.800 212.395 209.410 214.005 ;
        RECT 208.345 210.405 208.865 212.395 ;
        RECT 207.800 208.795 209.410 210.405 ;
        RECT 208.345 206.805 208.865 208.795 ;
        RECT 207.800 205.195 209.410 206.805 ;
        RECT 208.345 203.205 208.865 205.195 ;
        RECT 207.800 201.595 209.410 203.205 ;
        RECT 208.345 199.605 208.865 201.595 ;
        RECT 207.800 197.995 209.410 199.605 ;
        RECT 208.345 196.005 208.865 197.995 ;
        RECT 207.800 194.395 209.410 196.005 ;
        RECT 208.345 192.405 208.865 194.395 ;
        RECT 207.800 190.795 209.410 192.405 ;
        RECT 208.345 188.805 208.865 190.795 ;
        RECT 207.800 187.195 209.410 188.805 ;
        RECT 208.345 185.205 208.865 187.195 ;
        RECT 207.800 183.595 209.410 185.205 ;
        RECT 208.345 181.605 208.865 183.595 ;
        RECT 207.800 179.995 209.410 181.605 ;
        RECT 208.345 178.005 208.865 179.995 ;
        RECT 207.800 176.395 209.410 178.005 ;
        RECT 208.345 174.405 208.865 176.395 ;
        RECT 207.800 172.795 209.410 174.405 ;
        RECT 208.345 170.805 208.865 172.795 ;
        RECT 207.800 169.195 209.410 170.805 ;
        RECT 208.345 167.205 208.865 169.195 ;
        RECT 207.800 165.595 209.410 167.205 ;
        RECT 208.345 164.600 208.865 165.595 ;
        RECT 211.005 164.080 211.525 222.200 ;
        RECT 213.405 221.205 213.925 222.720 ;
        RECT 212.860 219.595 214.470 221.205 ;
        RECT 213.405 217.605 213.925 219.595 ;
        RECT 212.860 215.995 214.470 217.605 ;
        RECT 213.405 214.005 213.925 215.995 ;
        RECT 212.860 212.395 214.470 214.005 ;
        RECT 213.405 210.405 213.925 212.395 ;
        RECT 212.860 208.795 214.470 210.405 ;
        RECT 213.405 206.805 213.925 208.795 ;
        RECT 212.860 205.195 214.470 206.805 ;
        RECT 213.405 203.205 213.925 205.195 ;
        RECT 212.860 201.595 214.470 203.205 ;
        RECT 213.405 199.605 213.925 201.595 ;
        RECT 212.860 197.995 214.470 199.605 ;
        RECT 213.405 196.005 213.925 197.995 ;
        RECT 212.860 194.395 214.470 196.005 ;
        RECT 213.405 192.405 213.925 194.395 ;
        RECT 212.860 190.795 214.470 192.405 ;
        RECT 213.405 188.805 213.925 190.795 ;
        RECT 212.860 187.195 214.470 188.805 ;
        RECT 213.405 185.205 213.925 187.195 ;
        RECT 212.860 183.595 214.470 185.205 ;
        RECT 213.405 181.605 213.925 183.595 ;
        RECT 212.860 179.995 214.470 181.605 ;
        RECT 213.405 178.005 213.925 179.995 ;
        RECT 212.860 176.395 214.470 178.005 ;
        RECT 213.405 174.405 213.925 176.395 ;
        RECT 212.860 172.795 214.470 174.405 ;
        RECT 213.405 170.805 213.925 172.795 ;
        RECT 212.860 169.195 214.470 170.805 ;
        RECT 213.405 167.205 213.925 169.195 ;
        RECT 212.860 165.595 214.470 167.205 ;
        RECT 213.405 164.600 213.925 165.595 ;
        RECT 216.065 164.080 216.585 222.200 ;
        RECT 218.465 221.205 218.985 222.720 ;
        RECT 217.920 219.595 219.530 221.205 ;
        RECT 218.465 217.605 218.985 219.595 ;
        RECT 217.920 215.995 219.530 217.605 ;
        RECT 218.465 214.005 218.985 215.995 ;
        RECT 217.920 212.395 219.530 214.005 ;
        RECT 218.465 210.405 218.985 212.395 ;
        RECT 217.920 208.795 219.530 210.405 ;
        RECT 218.465 206.805 218.985 208.795 ;
        RECT 217.920 205.195 219.530 206.805 ;
        RECT 218.465 203.205 218.985 205.195 ;
        RECT 217.920 201.595 219.530 203.205 ;
        RECT 218.465 199.605 218.985 201.595 ;
        RECT 217.920 197.995 219.530 199.605 ;
        RECT 218.465 196.005 218.985 197.995 ;
        RECT 217.920 194.395 219.530 196.005 ;
        RECT 218.465 192.405 218.985 194.395 ;
        RECT 217.920 190.795 219.530 192.405 ;
        RECT 218.465 188.805 218.985 190.795 ;
        RECT 217.920 187.195 219.530 188.805 ;
        RECT 218.465 185.205 218.985 187.195 ;
        RECT 217.920 183.595 219.530 185.205 ;
        RECT 218.465 181.605 218.985 183.595 ;
        RECT 217.920 179.995 219.530 181.605 ;
        RECT 218.465 178.005 218.985 179.995 ;
        RECT 217.920 176.395 219.530 178.005 ;
        RECT 218.465 174.405 218.985 176.395 ;
        RECT 217.920 172.795 219.530 174.405 ;
        RECT 218.465 170.805 218.985 172.795 ;
        RECT 217.920 169.195 219.530 170.805 ;
        RECT 218.465 167.205 218.985 169.195 ;
        RECT 217.920 165.595 219.530 167.205 ;
        RECT 218.465 164.600 218.985 165.595 ;
        RECT 221.125 164.080 221.645 222.200 ;
        RECT 223.525 221.205 224.045 222.720 ;
        RECT 222.980 219.595 224.590 221.205 ;
        RECT 223.525 217.605 224.045 219.595 ;
        RECT 222.980 215.995 224.590 217.605 ;
        RECT 223.525 214.005 224.045 215.995 ;
        RECT 222.980 212.395 224.590 214.005 ;
        RECT 223.525 210.405 224.045 212.395 ;
        RECT 222.980 208.795 224.590 210.405 ;
        RECT 223.525 206.805 224.045 208.795 ;
        RECT 222.980 205.195 224.590 206.805 ;
        RECT 223.525 203.205 224.045 205.195 ;
        RECT 222.980 201.595 224.590 203.205 ;
        RECT 223.525 199.605 224.045 201.595 ;
        RECT 222.980 197.995 224.590 199.605 ;
        RECT 223.525 196.005 224.045 197.995 ;
        RECT 222.980 194.395 224.590 196.005 ;
        RECT 223.525 192.405 224.045 194.395 ;
        RECT 222.980 190.795 224.590 192.405 ;
        RECT 223.525 188.805 224.045 190.795 ;
        RECT 222.980 187.195 224.590 188.805 ;
        RECT 223.525 185.205 224.045 187.195 ;
        RECT 222.980 183.595 224.590 185.205 ;
        RECT 223.525 181.605 224.045 183.595 ;
        RECT 222.980 179.995 224.590 181.605 ;
        RECT 223.525 178.005 224.045 179.995 ;
        RECT 222.980 176.395 224.590 178.005 ;
        RECT 223.525 174.405 224.045 176.395 ;
        RECT 222.980 172.795 224.590 174.405 ;
        RECT 223.525 170.805 224.045 172.795 ;
        RECT 222.980 169.195 224.590 170.805 ;
        RECT 223.525 167.205 224.045 169.195 ;
        RECT 222.980 165.595 224.590 167.205 ;
        RECT 223.525 164.600 224.045 165.595 ;
        RECT 205.945 163.560 221.645 164.080 ;
        RECT 226.185 164.080 226.705 222.200 ;
        RECT 228.585 221.205 229.105 222.720 ;
        RECT 228.040 219.595 229.650 221.205 ;
        RECT 228.585 217.605 229.105 219.595 ;
        RECT 228.040 215.995 229.650 217.605 ;
        RECT 228.585 214.005 229.105 215.995 ;
        RECT 228.040 212.395 229.650 214.005 ;
        RECT 228.585 210.405 229.105 212.395 ;
        RECT 228.040 208.795 229.650 210.405 ;
        RECT 228.585 206.805 229.105 208.795 ;
        RECT 228.040 205.195 229.650 206.805 ;
        RECT 228.585 203.205 229.105 205.195 ;
        RECT 228.040 201.595 229.650 203.205 ;
        RECT 228.585 199.605 229.105 201.595 ;
        RECT 228.040 197.995 229.650 199.605 ;
        RECT 228.585 196.005 229.105 197.995 ;
        RECT 228.040 194.395 229.650 196.005 ;
        RECT 228.585 192.405 229.105 194.395 ;
        RECT 228.040 190.795 229.650 192.405 ;
        RECT 228.585 188.805 229.105 190.795 ;
        RECT 228.040 187.195 229.650 188.805 ;
        RECT 228.585 185.205 229.105 187.195 ;
        RECT 228.040 183.595 229.650 185.205 ;
        RECT 228.585 181.605 229.105 183.595 ;
        RECT 228.040 179.995 229.650 181.605 ;
        RECT 228.585 178.005 229.105 179.995 ;
        RECT 228.040 176.395 229.650 178.005 ;
        RECT 228.585 174.405 229.105 176.395 ;
        RECT 228.040 172.795 229.650 174.405 ;
        RECT 228.585 170.805 229.105 172.795 ;
        RECT 228.040 169.195 229.650 170.805 ;
        RECT 228.585 167.205 229.105 169.195 ;
        RECT 228.040 165.595 229.650 167.205 ;
        RECT 228.585 164.600 229.105 165.595 ;
        RECT 231.245 164.080 231.765 222.200 ;
        RECT 233.645 221.205 234.165 222.720 ;
        RECT 233.100 219.595 234.710 221.205 ;
        RECT 233.645 217.605 234.165 219.595 ;
        RECT 233.100 215.995 234.710 217.605 ;
        RECT 233.645 214.005 234.165 215.995 ;
        RECT 233.100 212.395 234.710 214.005 ;
        RECT 233.645 210.405 234.165 212.395 ;
        RECT 233.100 208.795 234.710 210.405 ;
        RECT 233.645 206.805 234.165 208.795 ;
        RECT 233.100 205.195 234.710 206.805 ;
        RECT 233.645 203.205 234.165 205.195 ;
        RECT 233.100 201.595 234.710 203.205 ;
        RECT 233.645 199.605 234.165 201.595 ;
        RECT 233.100 197.995 234.710 199.605 ;
        RECT 233.645 196.005 234.165 197.995 ;
        RECT 233.100 194.395 234.710 196.005 ;
        RECT 233.645 192.405 234.165 194.395 ;
        RECT 233.100 190.795 234.710 192.405 ;
        RECT 233.645 188.805 234.165 190.795 ;
        RECT 233.100 187.195 234.710 188.805 ;
        RECT 233.645 185.205 234.165 187.195 ;
        RECT 233.100 183.595 234.710 185.205 ;
        RECT 233.645 181.605 234.165 183.595 ;
        RECT 233.100 179.995 234.710 181.605 ;
        RECT 233.645 178.005 234.165 179.995 ;
        RECT 233.100 176.395 234.710 178.005 ;
        RECT 233.645 174.405 234.165 176.395 ;
        RECT 233.100 172.795 234.710 174.405 ;
        RECT 233.645 170.805 234.165 172.795 ;
        RECT 233.100 169.195 234.710 170.805 ;
        RECT 233.645 167.205 234.165 169.195 ;
        RECT 233.100 165.595 234.710 167.205 ;
        RECT 233.645 164.600 234.165 165.595 ;
        RECT 226.185 163.560 231.765 164.080 ;
        RECT 200.885 163.205 201.405 163.560 ;
        RECT 200.880 162.675 201.410 163.205 ;
        RECT 221.125 162.165 221.645 163.560 ;
        RECT 221.120 161.635 221.650 162.165 ;
        RECT 231.245 161.125 231.765 163.560 ;
        RECT 231.240 160.595 231.770 161.125 ;
        RECT 236.305 160.085 236.825 222.200 ;
        RECT 238.705 221.205 239.225 222.720 ;
        RECT 238.160 219.595 239.770 221.205 ;
        RECT 238.705 217.605 239.225 219.595 ;
        RECT 238.160 215.995 239.770 217.605 ;
        RECT 238.705 214.005 239.225 215.995 ;
        RECT 241.520 214.880 242.010 214.885 ;
        RECT 243.385 214.880 243.865 221.540 ;
        RECT 245.765 221.205 246.285 222.720 ;
        RECT 245.220 219.595 246.830 221.205 ;
        RECT 245.765 217.605 246.285 219.595 ;
        RECT 245.220 215.995 246.830 217.605 ;
        RECT 241.520 214.400 243.865 214.880 ;
        RECT 241.520 214.395 242.010 214.400 ;
        RECT 238.160 212.395 239.770 214.005 ;
        RECT 238.705 210.405 239.225 212.395 ;
        RECT 238.160 208.795 239.770 210.405 ;
        RECT 238.705 206.805 239.225 208.795 ;
        RECT 243.385 208.460 243.865 214.400 ;
        RECT 245.765 214.005 246.285 215.995 ;
        RECT 248.580 214.880 249.070 214.885 ;
        RECT 250.445 214.880 250.925 221.540 ;
        RECT 252.825 221.205 253.345 222.720 ;
        RECT 252.280 219.595 253.890 221.205 ;
        RECT 252.825 217.605 253.345 219.595 ;
        RECT 252.280 215.995 253.890 217.605 ;
        RECT 248.580 214.400 250.925 214.880 ;
        RECT 248.580 214.395 249.070 214.400 ;
        RECT 245.220 212.395 246.830 214.005 ;
        RECT 245.765 210.405 246.285 212.395 ;
        RECT 245.220 208.795 246.830 210.405 ;
        RECT 238.160 205.195 239.770 206.805 ;
        RECT 238.705 203.205 239.225 205.195 ;
        RECT 241.520 204.080 242.010 204.085 ;
        RECT 243.385 204.080 243.865 207.140 ;
        RECT 245.765 206.805 246.285 208.795 ;
        RECT 250.445 208.460 250.925 214.400 ;
        RECT 252.825 214.005 253.345 215.995 ;
        RECT 252.280 212.395 253.890 214.005 ;
        RECT 252.825 210.405 253.345 212.395 ;
        RECT 252.280 208.795 253.890 210.405 ;
        RECT 245.220 205.195 246.830 206.805 ;
        RECT 241.520 203.600 243.865 204.080 ;
        RECT 241.520 203.595 242.010 203.600 ;
        RECT 238.160 201.595 239.770 203.205 ;
        RECT 238.705 199.605 239.225 201.595 ;
        RECT 243.385 201.260 243.865 203.600 ;
        RECT 245.765 203.205 246.285 205.195 ;
        RECT 248.580 204.080 249.070 204.085 ;
        RECT 250.445 204.080 250.925 207.140 ;
        RECT 252.825 206.805 253.345 208.795 ;
        RECT 252.280 205.195 253.890 206.805 ;
        RECT 248.580 203.600 250.925 204.080 ;
        RECT 248.580 203.595 249.070 203.600 ;
        RECT 245.220 201.595 246.830 203.205 ;
        RECT 241.520 200.480 242.010 200.485 ;
        RECT 241.520 200.000 243.865 200.480 ;
        RECT 241.520 199.995 242.010 200.000 ;
        RECT 238.160 197.995 239.770 199.605 ;
        RECT 238.705 196.005 239.225 197.995 ;
        RECT 243.385 197.660 243.865 200.000 ;
        RECT 245.765 199.605 246.285 201.595 ;
        RECT 250.445 201.260 250.925 203.600 ;
        RECT 252.825 203.205 253.345 205.195 ;
        RECT 252.280 201.595 253.890 203.205 ;
        RECT 248.580 200.480 249.070 200.485 ;
        RECT 248.580 200.000 250.925 200.480 ;
        RECT 248.580 199.995 249.070 200.000 ;
        RECT 245.220 197.995 246.830 199.605 ;
        RECT 238.160 194.395 239.770 196.005 ;
        RECT 241.520 194.540 242.010 194.545 ;
        RECT 243.385 194.540 243.865 196.340 ;
        RECT 245.765 196.005 246.285 197.995 ;
        RECT 250.445 197.660 250.925 200.000 ;
        RECT 252.825 199.605 253.345 201.595 ;
        RECT 252.280 197.995 253.890 199.605 ;
        RECT 248.580 196.340 249.070 196.345 ;
        RECT 238.705 192.405 239.225 194.395 ;
        RECT 241.520 194.060 243.865 194.540 ;
        RECT 245.220 194.395 246.830 196.005 ;
        RECT 248.580 195.860 250.925 196.340 ;
        RECT 252.825 196.005 253.345 197.995 ;
        RECT 248.580 195.855 249.070 195.860 ;
        RECT 241.520 194.055 242.010 194.060 ;
        RECT 241.520 192.740 242.010 192.745 ;
        RECT 238.160 190.795 239.770 192.405 ;
        RECT 241.520 192.260 243.865 192.740 ;
        RECT 245.765 192.405 246.285 194.395 ;
        RECT 250.445 194.060 250.925 195.860 ;
        RECT 252.280 194.395 253.890 196.005 ;
        RECT 241.520 192.255 242.010 192.260 ;
        RECT 238.705 188.805 239.225 190.795 ;
        RECT 243.385 190.460 243.865 192.260 ;
        RECT 245.220 190.795 246.830 192.405 ;
        RECT 248.580 190.940 249.070 190.945 ;
        RECT 250.445 190.940 250.925 192.740 ;
        RECT 252.825 192.405 253.345 194.395 ;
        RECT 241.520 189.680 242.010 189.685 ;
        RECT 241.520 189.200 243.865 189.680 ;
        RECT 241.520 189.195 242.010 189.200 ;
        RECT 238.160 187.195 239.770 188.805 ;
        RECT 238.705 185.205 239.225 187.195 ;
        RECT 243.385 186.860 243.865 189.200 ;
        RECT 245.765 188.805 246.285 190.795 ;
        RECT 248.580 190.460 250.925 190.940 ;
        RECT 252.280 190.795 253.890 192.405 ;
        RECT 248.580 190.455 249.070 190.460 ;
        RECT 248.580 189.680 249.070 189.685 ;
        RECT 248.580 189.200 250.925 189.680 ;
        RECT 248.580 189.195 249.070 189.200 ;
        RECT 245.220 187.195 246.830 188.805 ;
        RECT 238.160 183.595 239.770 185.205 ;
        RECT 238.705 181.605 239.225 183.595 ;
        RECT 241.520 182.480 242.010 182.485 ;
        RECT 243.385 182.480 243.865 185.540 ;
        RECT 245.765 185.205 246.285 187.195 ;
        RECT 250.445 186.860 250.925 189.200 ;
        RECT 252.825 188.805 253.345 190.795 ;
        RECT 252.280 187.195 253.890 188.805 ;
        RECT 245.220 183.595 246.830 185.205 ;
        RECT 241.520 182.000 243.865 182.480 ;
        RECT 241.520 181.995 242.010 182.000 ;
        RECT 238.160 179.995 239.770 181.605 ;
        RECT 238.705 178.005 239.225 179.995 ;
        RECT 243.385 179.660 243.865 182.000 ;
        RECT 245.765 181.605 246.285 183.595 ;
        RECT 248.580 182.480 249.070 182.485 ;
        RECT 250.445 182.480 250.925 185.540 ;
        RECT 252.825 185.205 253.345 187.195 ;
        RECT 252.280 183.595 253.890 185.205 ;
        RECT 248.580 182.000 250.925 182.480 ;
        RECT 248.580 181.995 249.070 182.000 ;
        RECT 245.220 179.995 246.830 181.605 ;
        RECT 238.160 176.395 239.770 178.005 ;
        RECT 238.705 174.405 239.225 176.395 ;
        RECT 238.160 172.795 239.770 174.405 ;
        RECT 238.705 170.805 239.225 172.795 ;
        RECT 241.520 171.680 242.010 171.685 ;
        RECT 243.385 171.680 243.865 178.340 ;
        RECT 245.765 178.005 246.285 179.995 ;
        RECT 250.445 179.660 250.925 182.000 ;
        RECT 252.825 181.605 253.345 183.595 ;
        RECT 252.280 179.995 253.890 181.605 ;
        RECT 245.220 176.395 246.830 178.005 ;
        RECT 245.765 174.405 246.285 176.395 ;
        RECT 245.220 172.795 246.830 174.405 ;
        RECT 241.520 171.200 243.865 171.680 ;
        RECT 241.520 171.195 242.010 171.200 ;
        RECT 238.160 169.195 239.770 170.805 ;
        RECT 238.705 167.205 239.225 169.195 ;
        RECT 238.160 165.595 239.770 167.205 ;
        RECT 238.705 164.600 239.225 165.595 ;
        RECT 243.385 165.260 243.865 171.200 ;
        RECT 245.765 170.805 246.285 172.795 ;
        RECT 248.580 171.680 249.070 171.685 ;
        RECT 250.445 171.680 250.925 178.340 ;
        RECT 252.825 178.005 253.345 179.995 ;
        RECT 252.280 176.395 253.890 178.005 ;
        RECT 252.825 174.405 253.345 176.395 ;
        RECT 252.280 172.795 253.890 174.405 ;
        RECT 248.580 171.200 250.925 171.680 ;
        RECT 248.580 171.195 249.070 171.200 ;
        RECT 245.220 169.195 246.830 170.805 ;
        RECT 245.765 167.205 246.285 169.195 ;
        RECT 245.220 165.595 246.830 167.205 ;
        RECT 245.765 164.600 246.285 165.595 ;
        RECT 250.445 165.260 250.925 171.200 ;
        RECT 252.825 170.805 253.345 172.795 ;
        RECT 252.280 169.195 253.890 170.805 ;
        RECT 252.825 167.205 253.345 169.195 ;
        RECT 252.280 165.595 253.890 167.205 ;
        RECT 252.825 164.600 253.345 165.595 ;
        RECT 255.485 160.085 256.005 222.200 ;
        RECT 257.885 221.205 258.405 222.720 ;
        RECT 257.340 219.595 258.950 221.205 ;
        RECT 257.885 217.605 258.405 219.595 ;
        RECT 257.340 215.995 258.950 217.605 ;
        RECT 257.885 214.005 258.405 215.995 ;
        RECT 257.340 212.395 258.950 214.005 ;
        RECT 257.885 210.405 258.405 212.395 ;
        RECT 257.340 208.795 258.950 210.405 ;
        RECT 257.885 206.805 258.405 208.795 ;
        RECT 257.340 205.195 258.950 206.805 ;
        RECT 257.885 203.205 258.405 205.195 ;
        RECT 257.340 201.595 258.950 203.205 ;
        RECT 257.885 199.605 258.405 201.595 ;
        RECT 257.340 197.995 258.950 199.605 ;
        RECT 257.885 196.005 258.405 197.995 ;
        RECT 257.340 194.395 258.950 196.005 ;
        RECT 257.885 192.405 258.405 194.395 ;
        RECT 257.340 190.795 258.950 192.405 ;
        RECT 257.885 188.805 258.405 190.795 ;
        RECT 257.340 187.195 258.950 188.805 ;
        RECT 257.885 185.205 258.405 187.195 ;
        RECT 257.340 183.595 258.950 185.205 ;
        RECT 257.885 181.605 258.405 183.595 ;
        RECT 257.340 179.995 258.950 181.605 ;
        RECT 257.885 178.005 258.405 179.995 ;
        RECT 257.340 176.395 258.950 178.005 ;
        RECT 257.885 174.405 258.405 176.395 ;
        RECT 257.340 172.795 258.950 174.405 ;
        RECT 257.885 170.805 258.405 172.795 ;
        RECT 257.340 169.195 258.950 170.805 ;
        RECT 257.885 167.205 258.405 169.195 ;
        RECT 257.340 165.595 258.950 167.205 ;
        RECT 257.885 164.600 258.405 165.595 ;
        RECT 260.545 164.080 261.065 222.200 ;
        RECT 262.945 221.205 263.465 222.720 ;
        RECT 262.400 219.595 264.010 221.205 ;
        RECT 262.945 217.605 263.465 219.595 ;
        RECT 262.400 215.995 264.010 217.605 ;
        RECT 262.945 214.005 263.465 215.995 ;
        RECT 262.400 212.395 264.010 214.005 ;
        RECT 262.945 210.405 263.465 212.395 ;
        RECT 262.400 208.795 264.010 210.405 ;
        RECT 262.945 206.805 263.465 208.795 ;
        RECT 262.400 205.195 264.010 206.805 ;
        RECT 262.945 203.205 263.465 205.195 ;
        RECT 262.400 201.595 264.010 203.205 ;
        RECT 262.945 199.605 263.465 201.595 ;
        RECT 262.400 197.995 264.010 199.605 ;
        RECT 262.945 196.005 263.465 197.995 ;
        RECT 262.400 194.395 264.010 196.005 ;
        RECT 262.945 192.405 263.465 194.395 ;
        RECT 262.400 190.795 264.010 192.405 ;
        RECT 262.945 188.805 263.465 190.795 ;
        RECT 262.400 187.195 264.010 188.805 ;
        RECT 262.945 185.205 263.465 187.195 ;
        RECT 262.400 183.595 264.010 185.205 ;
        RECT 262.945 181.605 263.465 183.595 ;
        RECT 262.400 179.995 264.010 181.605 ;
        RECT 262.945 178.005 263.465 179.995 ;
        RECT 262.400 176.395 264.010 178.005 ;
        RECT 262.945 174.405 263.465 176.395 ;
        RECT 262.400 172.795 264.010 174.405 ;
        RECT 262.945 170.805 263.465 172.795 ;
        RECT 262.400 169.195 264.010 170.805 ;
        RECT 262.945 167.205 263.465 169.195 ;
        RECT 262.400 165.595 264.010 167.205 ;
        RECT 262.945 164.600 263.465 165.595 ;
        RECT 265.605 164.080 266.125 222.200 ;
        RECT 268.005 221.205 268.525 222.720 ;
        RECT 267.460 219.595 269.070 221.205 ;
        RECT 268.005 217.605 268.525 219.595 ;
        RECT 267.460 215.995 269.070 217.605 ;
        RECT 268.005 214.005 268.525 215.995 ;
        RECT 267.460 212.395 269.070 214.005 ;
        RECT 268.005 210.405 268.525 212.395 ;
        RECT 267.460 208.795 269.070 210.405 ;
        RECT 268.005 206.805 268.525 208.795 ;
        RECT 267.460 205.195 269.070 206.805 ;
        RECT 268.005 203.205 268.525 205.195 ;
        RECT 267.460 201.595 269.070 203.205 ;
        RECT 268.005 199.605 268.525 201.595 ;
        RECT 267.460 197.995 269.070 199.605 ;
        RECT 268.005 196.005 268.525 197.995 ;
        RECT 267.460 194.395 269.070 196.005 ;
        RECT 268.005 192.405 268.525 194.395 ;
        RECT 267.460 190.795 269.070 192.405 ;
        RECT 268.005 188.805 268.525 190.795 ;
        RECT 267.460 187.195 269.070 188.805 ;
        RECT 268.005 185.205 268.525 187.195 ;
        RECT 267.460 183.595 269.070 185.205 ;
        RECT 268.005 181.605 268.525 183.595 ;
        RECT 267.460 179.995 269.070 181.605 ;
        RECT 268.005 178.005 268.525 179.995 ;
        RECT 267.460 176.395 269.070 178.005 ;
        RECT 268.005 174.405 268.525 176.395 ;
        RECT 267.460 172.795 269.070 174.405 ;
        RECT 268.005 170.805 268.525 172.795 ;
        RECT 267.460 169.195 269.070 170.805 ;
        RECT 268.005 167.205 268.525 169.195 ;
        RECT 267.460 165.595 269.070 167.205 ;
        RECT 268.005 164.600 268.525 165.595 ;
        RECT 260.545 163.560 266.125 164.080 ;
        RECT 270.665 164.080 271.185 222.200 ;
        RECT 273.065 221.205 273.585 222.720 ;
        RECT 272.520 219.595 274.130 221.205 ;
        RECT 273.065 217.605 273.585 219.595 ;
        RECT 272.520 215.995 274.130 217.605 ;
        RECT 273.065 214.005 273.585 215.995 ;
        RECT 272.520 212.395 274.130 214.005 ;
        RECT 273.065 210.405 273.585 212.395 ;
        RECT 272.520 208.795 274.130 210.405 ;
        RECT 273.065 206.805 273.585 208.795 ;
        RECT 272.520 205.195 274.130 206.805 ;
        RECT 273.065 203.205 273.585 205.195 ;
        RECT 272.520 201.595 274.130 203.205 ;
        RECT 273.065 199.605 273.585 201.595 ;
        RECT 272.520 197.995 274.130 199.605 ;
        RECT 273.065 196.005 273.585 197.995 ;
        RECT 272.520 194.395 274.130 196.005 ;
        RECT 273.065 192.405 273.585 194.395 ;
        RECT 272.520 190.795 274.130 192.405 ;
        RECT 273.065 188.805 273.585 190.795 ;
        RECT 272.520 187.195 274.130 188.805 ;
        RECT 273.065 185.205 273.585 187.195 ;
        RECT 272.520 183.595 274.130 185.205 ;
        RECT 273.065 181.605 273.585 183.595 ;
        RECT 272.520 179.995 274.130 181.605 ;
        RECT 273.065 178.005 273.585 179.995 ;
        RECT 272.520 176.395 274.130 178.005 ;
        RECT 273.065 174.405 273.585 176.395 ;
        RECT 272.520 172.795 274.130 174.405 ;
        RECT 273.065 170.805 273.585 172.795 ;
        RECT 272.520 169.195 274.130 170.805 ;
        RECT 273.065 167.205 273.585 169.195 ;
        RECT 272.520 165.595 274.130 167.205 ;
        RECT 273.065 164.600 273.585 165.595 ;
        RECT 275.725 164.080 276.245 222.200 ;
        RECT 278.125 221.205 278.645 222.720 ;
        RECT 277.580 219.595 279.190 221.205 ;
        RECT 278.125 217.605 278.645 219.595 ;
        RECT 277.580 215.995 279.190 217.605 ;
        RECT 278.125 214.005 278.645 215.995 ;
        RECT 277.580 212.395 279.190 214.005 ;
        RECT 278.125 210.405 278.645 212.395 ;
        RECT 277.580 208.795 279.190 210.405 ;
        RECT 278.125 206.805 278.645 208.795 ;
        RECT 277.580 205.195 279.190 206.805 ;
        RECT 278.125 203.205 278.645 205.195 ;
        RECT 277.580 201.595 279.190 203.205 ;
        RECT 278.125 199.605 278.645 201.595 ;
        RECT 277.580 197.995 279.190 199.605 ;
        RECT 278.125 196.005 278.645 197.995 ;
        RECT 277.580 194.395 279.190 196.005 ;
        RECT 278.125 192.405 278.645 194.395 ;
        RECT 277.580 190.795 279.190 192.405 ;
        RECT 278.125 188.805 278.645 190.795 ;
        RECT 277.580 187.195 279.190 188.805 ;
        RECT 278.125 185.205 278.645 187.195 ;
        RECT 277.580 183.595 279.190 185.205 ;
        RECT 278.125 181.605 278.645 183.595 ;
        RECT 277.580 179.995 279.190 181.605 ;
        RECT 278.125 178.005 278.645 179.995 ;
        RECT 277.580 176.395 279.190 178.005 ;
        RECT 278.125 174.405 278.645 176.395 ;
        RECT 277.580 172.795 279.190 174.405 ;
        RECT 278.125 170.805 278.645 172.795 ;
        RECT 277.580 169.195 279.190 170.805 ;
        RECT 278.125 167.205 278.645 169.195 ;
        RECT 277.580 165.595 279.190 167.205 ;
        RECT 278.125 164.600 278.645 165.595 ;
        RECT 280.785 164.080 281.305 222.200 ;
        RECT 283.185 221.205 283.705 222.720 ;
        RECT 282.640 219.595 284.250 221.205 ;
        RECT 283.185 217.605 283.705 219.595 ;
        RECT 282.640 215.995 284.250 217.605 ;
        RECT 283.185 214.005 283.705 215.995 ;
        RECT 282.640 212.395 284.250 214.005 ;
        RECT 283.185 210.405 283.705 212.395 ;
        RECT 282.640 208.795 284.250 210.405 ;
        RECT 283.185 206.805 283.705 208.795 ;
        RECT 282.640 205.195 284.250 206.805 ;
        RECT 283.185 203.205 283.705 205.195 ;
        RECT 282.640 201.595 284.250 203.205 ;
        RECT 283.185 199.605 283.705 201.595 ;
        RECT 282.640 197.995 284.250 199.605 ;
        RECT 283.185 196.005 283.705 197.995 ;
        RECT 282.640 194.395 284.250 196.005 ;
        RECT 283.185 192.405 283.705 194.395 ;
        RECT 282.640 190.795 284.250 192.405 ;
        RECT 283.185 188.805 283.705 190.795 ;
        RECT 282.640 187.195 284.250 188.805 ;
        RECT 283.185 185.205 283.705 187.195 ;
        RECT 282.640 183.595 284.250 185.205 ;
        RECT 283.185 181.605 283.705 183.595 ;
        RECT 282.640 179.995 284.250 181.605 ;
        RECT 283.185 178.005 283.705 179.995 ;
        RECT 282.640 176.395 284.250 178.005 ;
        RECT 283.185 174.405 283.705 176.395 ;
        RECT 282.640 172.795 284.250 174.405 ;
        RECT 283.185 170.805 283.705 172.795 ;
        RECT 282.640 169.195 284.250 170.805 ;
        RECT 283.185 167.205 283.705 169.195 ;
        RECT 282.640 165.595 284.250 167.205 ;
        RECT 283.185 164.600 283.705 165.595 ;
        RECT 285.845 164.080 286.365 222.200 ;
        RECT 288.245 221.205 288.765 222.720 ;
        RECT 287.700 219.595 289.310 221.205 ;
        RECT 288.245 217.605 288.765 219.595 ;
        RECT 287.700 215.995 289.310 217.605 ;
        RECT 288.245 214.005 288.765 215.995 ;
        RECT 287.700 212.395 289.310 214.005 ;
        RECT 288.245 210.405 288.765 212.395 ;
        RECT 287.700 208.795 289.310 210.405 ;
        RECT 288.245 206.805 288.765 208.795 ;
        RECT 287.700 205.195 289.310 206.805 ;
        RECT 288.245 203.205 288.765 205.195 ;
        RECT 287.700 201.595 289.310 203.205 ;
        RECT 288.245 199.605 288.765 201.595 ;
        RECT 287.700 197.995 289.310 199.605 ;
        RECT 288.245 196.005 288.765 197.995 ;
        RECT 287.700 194.395 289.310 196.005 ;
        RECT 288.245 192.405 288.765 194.395 ;
        RECT 287.700 190.795 289.310 192.405 ;
        RECT 288.245 188.805 288.765 190.795 ;
        RECT 287.700 187.195 289.310 188.805 ;
        RECT 288.245 185.205 288.765 187.195 ;
        RECT 287.700 183.595 289.310 185.205 ;
        RECT 288.245 181.605 288.765 183.595 ;
        RECT 287.700 179.995 289.310 181.605 ;
        RECT 288.245 178.005 288.765 179.995 ;
        RECT 287.700 176.395 289.310 178.005 ;
        RECT 288.245 174.405 288.765 176.395 ;
        RECT 287.700 172.795 289.310 174.405 ;
        RECT 288.245 170.805 288.765 172.795 ;
        RECT 287.700 169.195 289.310 170.805 ;
        RECT 288.245 167.205 288.765 169.195 ;
        RECT 287.700 165.595 289.310 167.205 ;
        RECT 288.245 164.600 288.765 165.595 ;
        RECT 270.665 163.560 286.365 164.080 ;
        RECT 290.905 164.080 291.425 222.200 ;
        RECT 293.305 221.205 293.825 222.720 ;
        RECT 292.760 219.595 294.370 221.205 ;
        RECT 293.305 217.605 293.825 219.595 ;
        RECT 292.760 215.995 294.370 217.605 ;
        RECT 293.305 214.005 293.825 215.995 ;
        RECT 292.760 212.395 294.370 214.005 ;
        RECT 293.305 210.405 293.825 212.395 ;
        RECT 292.760 208.795 294.370 210.405 ;
        RECT 293.305 206.805 293.825 208.795 ;
        RECT 292.760 205.195 294.370 206.805 ;
        RECT 293.305 203.205 293.825 205.195 ;
        RECT 292.760 201.595 294.370 203.205 ;
        RECT 293.305 199.605 293.825 201.595 ;
        RECT 292.760 197.995 294.370 199.605 ;
        RECT 293.305 196.005 293.825 197.995 ;
        RECT 292.760 194.395 294.370 196.005 ;
        RECT 293.305 192.405 293.825 194.395 ;
        RECT 292.760 190.795 294.370 192.405 ;
        RECT 293.305 188.805 293.825 190.795 ;
        RECT 292.760 187.195 294.370 188.805 ;
        RECT 293.305 185.205 293.825 187.195 ;
        RECT 292.760 183.595 294.370 185.205 ;
        RECT 293.305 181.605 293.825 183.595 ;
        RECT 292.760 179.995 294.370 181.605 ;
        RECT 293.305 178.005 293.825 179.995 ;
        RECT 292.760 176.395 294.370 178.005 ;
        RECT 293.305 174.405 293.825 176.395 ;
        RECT 292.760 172.795 294.370 174.405 ;
        RECT 293.305 170.805 293.825 172.795 ;
        RECT 292.760 169.195 294.370 170.805 ;
        RECT 293.305 167.205 293.825 169.195 ;
        RECT 292.760 165.595 294.370 167.205 ;
        RECT 293.305 164.600 293.825 165.595 ;
        RECT 295.965 164.080 296.485 222.200 ;
        RECT 298.365 221.205 298.885 222.720 ;
        RECT 297.820 219.595 299.430 221.205 ;
        RECT 298.365 217.605 298.885 219.595 ;
        RECT 297.820 215.995 299.430 217.605 ;
        RECT 298.365 214.005 298.885 215.995 ;
        RECT 297.820 212.395 299.430 214.005 ;
        RECT 298.365 210.405 298.885 212.395 ;
        RECT 297.820 208.795 299.430 210.405 ;
        RECT 298.365 206.805 298.885 208.795 ;
        RECT 297.820 205.195 299.430 206.805 ;
        RECT 298.365 203.205 298.885 205.195 ;
        RECT 297.820 201.595 299.430 203.205 ;
        RECT 298.365 199.605 298.885 201.595 ;
        RECT 297.820 197.995 299.430 199.605 ;
        RECT 298.365 196.005 298.885 197.995 ;
        RECT 297.820 194.395 299.430 196.005 ;
        RECT 298.365 192.405 298.885 194.395 ;
        RECT 297.820 190.795 299.430 192.405 ;
        RECT 298.365 188.805 298.885 190.795 ;
        RECT 297.820 187.195 299.430 188.805 ;
        RECT 298.365 185.205 298.885 187.195 ;
        RECT 297.820 183.595 299.430 185.205 ;
        RECT 298.365 181.605 298.885 183.595 ;
        RECT 297.820 179.995 299.430 181.605 ;
        RECT 298.365 178.005 298.885 179.995 ;
        RECT 297.820 176.395 299.430 178.005 ;
        RECT 298.365 174.405 298.885 176.395 ;
        RECT 297.820 172.795 299.430 174.405 ;
        RECT 298.365 170.805 298.885 172.795 ;
        RECT 297.820 169.195 299.430 170.805 ;
        RECT 298.365 167.205 298.885 169.195 ;
        RECT 297.820 165.595 299.430 167.205 ;
        RECT 298.365 164.600 298.885 165.595 ;
        RECT 301.025 164.080 301.545 222.200 ;
        RECT 303.425 221.205 303.945 222.720 ;
        RECT 302.880 219.595 304.490 221.205 ;
        RECT 303.425 217.605 303.945 219.595 ;
        RECT 302.880 215.995 304.490 217.605 ;
        RECT 303.425 214.005 303.945 215.995 ;
        RECT 302.880 212.395 304.490 214.005 ;
        RECT 303.425 210.405 303.945 212.395 ;
        RECT 302.880 208.795 304.490 210.405 ;
        RECT 303.425 206.805 303.945 208.795 ;
        RECT 302.880 205.195 304.490 206.805 ;
        RECT 303.425 203.205 303.945 205.195 ;
        RECT 302.880 201.595 304.490 203.205 ;
        RECT 303.425 199.605 303.945 201.595 ;
        RECT 302.880 197.995 304.490 199.605 ;
        RECT 303.425 196.005 303.945 197.995 ;
        RECT 302.880 194.395 304.490 196.005 ;
        RECT 303.425 192.405 303.945 194.395 ;
        RECT 302.880 190.795 304.490 192.405 ;
        RECT 303.425 188.805 303.945 190.795 ;
        RECT 302.880 187.195 304.490 188.805 ;
        RECT 303.425 185.205 303.945 187.195 ;
        RECT 302.880 183.595 304.490 185.205 ;
        RECT 303.425 181.605 303.945 183.595 ;
        RECT 302.880 179.995 304.490 181.605 ;
        RECT 303.425 178.005 303.945 179.995 ;
        RECT 302.880 176.395 304.490 178.005 ;
        RECT 303.425 174.405 303.945 176.395 ;
        RECT 302.880 172.795 304.490 174.405 ;
        RECT 303.425 170.805 303.945 172.795 ;
        RECT 302.880 169.195 304.490 170.805 ;
        RECT 303.425 167.205 303.945 169.195 ;
        RECT 302.880 165.595 304.490 167.205 ;
        RECT 303.425 164.600 303.945 165.595 ;
        RECT 306.085 164.080 306.605 222.200 ;
        RECT 308.485 221.205 309.005 222.720 ;
        RECT 307.940 219.595 309.550 221.205 ;
        RECT 308.485 217.605 309.005 219.595 ;
        RECT 307.940 215.995 309.550 217.605 ;
        RECT 308.485 214.005 309.005 215.995 ;
        RECT 307.940 212.395 309.550 214.005 ;
        RECT 308.485 210.405 309.005 212.395 ;
        RECT 307.940 208.795 309.550 210.405 ;
        RECT 308.485 206.805 309.005 208.795 ;
        RECT 307.940 205.195 309.550 206.805 ;
        RECT 308.485 203.205 309.005 205.195 ;
        RECT 307.940 201.595 309.550 203.205 ;
        RECT 308.485 199.605 309.005 201.595 ;
        RECT 307.940 197.995 309.550 199.605 ;
        RECT 308.485 196.005 309.005 197.995 ;
        RECT 307.940 194.395 309.550 196.005 ;
        RECT 308.485 192.405 309.005 194.395 ;
        RECT 307.940 190.795 309.550 192.405 ;
        RECT 308.485 188.805 309.005 190.795 ;
        RECT 307.940 187.195 309.550 188.805 ;
        RECT 308.485 185.205 309.005 187.195 ;
        RECT 307.940 183.595 309.550 185.205 ;
        RECT 308.485 181.605 309.005 183.595 ;
        RECT 307.940 179.995 309.550 181.605 ;
        RECT 308.485 178.005 309.005 179.995 ;
        RECT 307.940 176.395 309.550 178.005 ;
        RECT 308.485 174.405 309.005 176.395 ;
        RECT 307.940 172.795 309.550 174.405 ;
        RECT 308.485 170.805 309.005 172.795 ;
        RECT 307.940 169.195 309.550 170.805 ;
        RECT 308.485 167.205 309.005 169.195 ;
        RECT 307.940 165.595 309.550 167.205 ;
        RECT 308.485 164.600 309.005 165.595 ;
        RECT 311.145 164.080 311.665 222.200 ;
        RECT 313.545 221.205 314.065 222.720 ;
        RECT 313.000 219.595 314.610 221.205 ;
        RECT 313.545 217.605 314.065 219.595 ;
        RECT 313.000 215.995 314.610 217.605 ;
        RECT 313.545 214.005 314.065 215.995 ;
        RECT 313.000 212.395 314.610 214.005 ;
        RECT 313.545 210.405 314.065 212.395 ;
        RECT 313.000 208.795 314.610 210.405 ;
        RECT 313.545 206.805 314.065 208.795 ;
        RECT 313.000 205.195 314.610 206.805 ;
        RECT 313.545 203.205 314.065 205.195 ;
        RECT 313.000 201.595 314.610 203.205 ;
        RECT 313.545 199.605 314.065 201.595 ;
        RECT 313.000 197.995 314.610 199.605 ;
        RECT 313.545 196.005 314.065 197.995 ;
        RECT 313.000 194.395 314.610 196.005 ;
        RECT 313.545 192.405 314.065 194.395 ;
        RECT 313.000 190.795 314.610 192.405 ;
        RECT 313.545 188.805 314.065 190.795 ;
        RECT 313.000 187.195 314.610 188.805 ;
        RECT 313.545 185.205 314.065 187.195 ;
        RECT 313.000 183.595 314.610 185.205 ;
        RECT 313.545 181.605 314.065 183.595 ;
        RECT 313.000 179.995 314.610 181.605 ;
        RECT 313.545 178.005 314.065 179.995 ;
        RECT 313.000 176.395 314.610 178.005 ;
        RECT 313.545 174.405 314.065 176.395 ;
        RECT 313.000 172.795 314.610 174.405 ;
        RECT 313.545 170.805 314.065 172.795 ;
        RECT 313.000 169.195 314.610 170.805 ;
        RECT 313.545 167.205 314.065 169.195 ;
        RECT 313.000 165.595 314.610 167.205 ;
        RECT 313.545 164.600 314.065 165.595 ;
        RECT 316.205 164.080 316.725 222.200 ;
        RECT 318.605 221.205 319.125 222.720 ;
        RECT 318.060 219.595 319.670 221.205 ;
        RECT 318.605 217.605 319.125 219.595 ;
        RECT 318.060 215.995 319.670 217.605 ;
        RECT 318.605 214.005 319.125 215.995 ;
        RECT 318.060 212.395 319.670 214.005 ;
        RECT 318.605 210.405 319.125 212.395 ;
        RECT 318.060 208.795 319.670 210.405 ;
        RECT 318.605 206.805 319.125 208.795 ;
        RECT 318.060 205.195 319.670 206.805 ;
        RECT 318.605 203.205 319.125 205.195 ;
        RECT 318.060 201.595 319.670 203.205 ;
        RECT 318.605 199.605 319.125 201.595 ;
        RECT 318.060 197.995 319.670 199.605 ;
        RECT 318.605 196.005 319.125 197.995 ;
        RECT 318.060 194.395 319.670 196.005 ;
        RECT 318.605 192.405 319.125 194.395 ;
        RECT 318.060 190.795 319.670 192.405 ;
        RECT 318.605 188.805 319.125 190.795 ;
        RECT 318.060 187.195 319.670 188.805 ;
        RECT 318.605 185.205 319.125 187.195 ;
        RECT 318.060 183.595 319.670 185.205 ;
        RECT 318.605 181.605 319.125 183.595 ;
        RECT 318.060 179.995 319.670 181.605 ;
        RECT 318.605 178.005 319.125 179.995 ;
        RECT 318.060 176.395 319.670 178.005 ;
        RECT 318.605 174.405 319.125 176.395 ;
        RECT 318.060 172.795 319.670 174.405 ;
        RECT 318.605 170.805 319.125 172.795 ;
        RECT 318.060 169.195 319.670 170.805 ;
        RECT 318.605 167.205 319.125 169.195 ;
        RECT 318.060 165.595 319.670 167.205 ;
        RECT 318.605 164.600 319.125 165.595 ;
        RECT 321.265 164.080 321.785 222.200 ;
        RECT 323.665 221.205 324.185 222.720 ;
        RECT 323.120 219.595 324.730 221.205 ;
        RECT 323.665 217.605 324.185 219.595 ;
        RECT 323.120 215.995 324.730 217.605 ;
        RECT 323.665 214.005 324.185 215.995 ;
        RECT 323.120 212.395 324.730 214.005 ;
        RECT 323.665 210.405 324.185 212.395 ;
        RECT 323.120 208.795 324.730 210.405 ;
        RECT 323.665 206.805 324.185 208.795 ;
        RECT 323.120 205.195 324.730 206.805 ;
        RECT 323.665 203.205 324.185 205.195 ;
        RECT 323.120 201.595 324.730 203.205 ;
        RECT 323.665 199.605 324.185 201.595 ;
        RECT 323.120 197.995 324.730 199.605 ;
        RECT 323.665 196.005 324.185 197.995 ;
        RECT 323.120 194.395 324.730 196.005 ;
        RECT 323.665 192.405 324.185 194.395 ;
        RECT 323.120 190.795 324.730 192.405 ;
        RECT 323.665 188.805 324.185 190.795 ;
        RECT 323.120 187.195 324.730 188.805 ;
        RECT 323.665 185.205 324.185 187.195 ;
        RECT 323.120 183.595 324.730 185.205 ;
        RECT 323.665 181.605 324.185 183.595 ;
        RECT 323.120 179.995 324.730 181.605 ;
        RECT 323.665 178.005 324.185 179.995 ;
        RECT 323.120 176.395 324.730 178.005 ;
        RECT 323.665 174.405 324.185 176.395 ;
        RECT 323.120 172.795 324.730 174.405 ;
        RECT 323.665 170.805 324.185 172.795 ;
        RECT 323.120 169.195 324.730 170.805 ;
        RECT 323.665 167.205 324.185 169.195 ;
        RECT 323.120 165.595 324.730 167.205 ;
        RECT 323.665 164.600 324.185 165.595 ;
        RECT 326.325 164.080 326.845 222.200 ;
        RECT 328.725 221.205 329.245 222.720 ;
        RECT 328.180 219.595 329.790 221.205 ;
        RECT 328.725 217.605 329.245 219.595 ;
        RECT 328.180 215.995 329.790 217.605 ;
        RECT 328.725 214.005 329.245 215.995 ;
        RECT 328.180 212.395 329.790 214.005 ;
        RECT 328.725 210.405 329.245 212.395 ;
        RECT 328.180 208.795 329.790 210.405 ;
        RECT 328.725 206.805 329.245 208.795 ;
        RECT 328.180 205.195 329.790 206.805 ;
        RECT 328.725 203.205 329.245 205.195 ;
        RECT 328.180 201.595 329.790 203.205 ;
        RECT 328.725 199.605 329.245 201.595 ;
        RECT 328.180 197.995 329.790 199.605 ;
        RECT 328.725 196.005 329.245 197.995 ;
        RECT 328.180 194.395 329.790 196.005 ;
        RECT 328.725 192.405 329.245 194.395 ;
        RECT 328.180 190.795 329.790 192.405 ;
        RECT 328.725 188.805 329.245 190.795 ;
        RECT 328.180 187.195 329.790 188.805 ;
        RECT 328.725 185.205 329.245 187.195 ;
        RECT 328.180 183.595 329.790 185.205 ;
        RECT 328.725 181.605 329.245 183.595 ;
        RECT 328.180 179.995 329.790 181.605 ;
        RECT 328.725 178.005 329.245 179.995 ;
        RECT 328.180 176.395 329.790 178.005 ;
        RECT 328.725 174.405 329.245 176.395 ;
        RECT 328.180 172.795 329.790 174.405 ;
        RECT 328.725 170.805 329.245 172.795 ;
        RECT 328.180 169.195 329.790 170.805 ;
        RECT 328.725 167.205 329.245 169.195 ;
        RECT 328.180 165.595 329.790 167.205 ;
        RECT 328.725 164.600 329.245 165.595 ;
        RECT 290.905 163.560 326.845 164.080 ;
        RECT 260.545 161.125 261.065 163.560 ;
        RECT 270.665 162.165 271.185 163.560 ;
        RECT 290.905 163.205 291.425 163.560 ;
        RECT 290.900 162.675 291.430 163.205 ;
        RECT 270.660 161.635 271.190 162.165 ;
        RECT 260.540 160.595 261.070 161.125 ;
        RECT 236.300 159.555 236.830 160.085 ;
        RECT 255.480 159.555 256.010 160.085 ;
        RECT 8.195 152.895 8.805 157.005 ;
        RECT 13.995 152.895 14.605 157.005 ;
        RECT 19.695 152.895 20.305 157.005 ;
        RECT 25.495 152.895 26.105 157.005 ;
        RECT 31.195 152.895 31.805 157.005 ;
        RECT 36.995 152.895 37.605 157.005 ;
        RECT 42.795 152.895 43.405 157.005 ;
        RECT 48.495 152.895 49.105 157.005 ;
        RECT 54.295 152.895 54.905 157.005 ;
        RECT 60.095 152.895 60.705 157.005 ;
        RECT 65.795 152.895 66.405 157.005 ;
        RECT 71.595 152.895 72.205 157.005 ;
        RECT 71.925 152.380 75.935 152.435 ;
        RECT 71.925 151.880 93.750 152.380 ;
        RECT 71.925 151.825 75.935 151.880 ;
        RECT 71.925 149.425 75.935 149.475 ;
        RECT 71.925 148.925 92.150 149.425 ;
        RECT 0.995 146.895 1.000 148.905 ;
        RECT 3.000 146.895 3.005 148.905 ;
        RECT 14.195 146.895 16.205 148.905 ;
        RECT 71.925 148.865 75.935 148.925 ;
        RECT 14.200 83.440 16.200 146.895 ;
        RECT 71.925 146.455 75.935 146.515 ;
        RECT 71.925 145.955 90.650 146.455 ;
        RECT 71.925 145.905 75.935 145.955 ;
        RECT 29.200 80.500 31.200 143.860 ;
        RECT 44.200 83.440 46.200 143.860 ;
        RECT 59.200 83.440 61.200 143.860 ;
        RECT 71.925 143.500 75.935 143.555 ;
        RECT 71.925 143.000 89.250 143.500 ;
        RECT 71.925 142.945 75.935 143.000 ;
        RECT 71.925 140.540 75.935 140.595 ;
        RECT 71.925 140.040 87.750 140.540 ;
        RECT 71.925 139.985 75.935 140.040 ;
        RECT 71.925 137.580 75.935 137.635 ;
        RECT 71.925 137.080 86.450 137.580 ;
        RECT 71.925 137.025 75.935 137.080 ;
        RECT 71.925 134.630 75.935 134.675 ;
        RECT 71.925 134.130 85.150 134.630 ;
        RECT 71.925 134.065 75.935 134.130 ;
        RECT 71.925 131.655 75.935 131.715 ;
        RECT 71.925 131.155 83.950 131.655 ;
        RECT 71.925 131.105 75.935 131.155 ;
        RECT 71.925 128.700 75.935 128.755 ;
        RECT 71.925 128.200 82.650 128.700 ;
        RECT 71.925 128.145 75.935 128.200 ;
        RECT 71.925 125.745 75.935 125.795 ;
        RECT 71.925 125.245 81.350 125.745 ;
        RECT 71.925 125.185 75.935 125.245 ;
        RECT 71.925 122.770 75.935 122.835 ;
        RECT 71.925 122.270 80.150 122.770 ;
        RECT 71.925 122.225 75.935 122.270 ;
        RECT 71.925 119.820 75.935 119.875 ;
        RECT 71.925 119.320 79.050 119.820 ;
        RECT 71.925 119.265 75.935 119.320 ;
        RECT 71.925 116.850 75.935 116.915 ;
        RECT 71.925 116.350 77.900 116.850 ;
        RECT 71.925 116.305 75.935 116.350 ;
        RECT 77.400 114.900 77.900 116.350 ;
        RECT 78.550 115.900 79.050 119.320 ;
        RECT 79.650 116.900 80.150 122.270 ;
        RECT 80.850 117.900 81.350 125.245 ;
        RECT 82.150 118.900 82.650 128.200 ;
        RECT 83.450 119.900 83.950 131.155 ;
        RECT 84.650 120.900 85.150 134.130 ;
        RECT 85.950 121.900 86.450 137.080 ;
        RECT 87.250 122.900 87.750 140.040 ;
        RECT 88.750 123.900 89.250 143.000 ;
        RECT 90.150 124.900 90.650 145.955 ;
        RECT 91.650 125.900 92.150 148.925 ;
        RECT 93.250 126.900 93.750 151.880 ;
        RECT 113.795 126.900 114.305 126.905 ;
        RECT 93.250 126.400 114.305 126.900 ;
        RECT 113.795 126.395 114.305 126.400 ;
        RECT 137.805 125.900 138.315 125.905 ;
        RECT 91.650 125.400 138.315 125.900 ;
        RECT 137.805 125.395 138.315 125.400 ;
        RECT 161.815 124.900 162.325 125.405 ;
        RECT 90.150 124.895 162.325 124.900 ;
        RECT 90.150 124.400 162.320 124.895 ;
        RECT 185.825 123.900 186.335 123.905 ;
        RECT 88.750 123.400 186.335 123.900 ;
        RECT 185.825 123.395 186.335 123.400 ;
        RECT 209.835 122.900 210.345 122.905 ;
        RECT 87.250 122.400 210.345 122.900 ;
        RECT 209.835 122.395 210.345 122.400 ;
        RECT 233.845 121.900 234.355 121.905 ;
        RECT 85.950 121.400 234.355 121.900 ;
        RECT 233.845 121.395 234.355 121.400 ;
        RECT 257.855 120.900 258.365 120.905 ;
        RECT 84.650 120.400 258.365 120.900 ;
        RECT 257.855 120.395 258.365 120.400 ;
        RECT 281.865 119.900 282.375 119.905 ;
        RECT 83.450 119.400 282.375 119.900 ;
        RECT 281.865 119.395 282.375 119.400 ;
        RECT 305.875 118.900 306.385 118.905 ;
        RECT 82.150 118.400 306.385 118.900 ;
        RECT 305.875 118.395 306.385 118.400 ;
        RECT 112.795 117.900 113.305 117.905 ;
        RECT 80.850 117.400 113.305 117.900 ;
        RECT 112.795 117.395 113.305 117.400 ;
        RECT 136.805 116.900 137.315 116.905 ;
        RECT 79.650 116.400 137.315 116.900 ;
        RECT 136.805 116.395 137.315 116.400 ;
        RECT 160.815 115.900 161.325 115.905 ;
        RECT 78.550 115.400 161.325 115.900 ;
        RECT 160.815 115.395 161.325 115.400 ;
        RECT 184.825 114.900 185.335 114.905 ;
        RECT 77.400 114.400 185.335 114.900 ;
        RECT 184.825 114.395 185.335 114.400 ;
        RECT 71.925 113.900 75.935 113.955 ;
        RECT 208.835 113.900 209.345 113.905 ;
        RECT 71.925 113.400 209.345 113.900 ;
        RECT 71.925 113.345 75.935 113.400 ;
        RECT 208.835 113.395 209.345 113.400 ;
        RECT 232.845 112.900 233.355 112.905 ;
        RECT 77.400 112.400 233.355 112.900 ;
        RECT 71.925 110.950 75.935 110.995 ;
        RECT 77.400 110.950 77.900 112.400 ;
        RECT 232.845 112.395 233.355 112.400 ;
        RECT 256.855 111.900 257.365 111.905 ;
        RECT 71.925 110.450 77.900 110.950 ;
        RECT 78.550 111.400 257.365 111.900 ;
        RECT 71.925 110.385 75.935 110.450 ;
        RECT 71.925 107.980 75.935 108.035 ;
        RECT 78.550 107.980 79.050 111.400 ;
        RECT 256.855 111.395 257.365 111.400 ;
        RECT 280.865 110.900 281.375 110.905 ;
        RECT 71.925 107.480 79.050 107.980 ;
        RECT 79.650 110.400 281.375 110.900 ;
        RECT 71.925 107.425 75.935 107.480 ;
        RECT 71.925 105.030 75.935 105.075 ;
        RECT 79.650 105.030 80.150 110.400 ;
        RECT 280.865 110.395 281.375 110.400 ;
        RECT 304.875 109.900 305.385 109.905 ;
        RECT 71.925 104.530 80.150 105.030 ;
        RECT 80.850 109.400 305.385 109.900 ;
        RECT 71.925 104.465 75.935 104.530 ;
        RECT 71.925 102.055 75.935 102.115 ;
        RECT 80.850 102.055 81.350 109.400 ;
        RECT 304.875 109.395 305.385 109.400 ;
        RECT 113.795 108.900 114.305 108.905 ;
        RECT 71.925 101.555 81.350 102.055 ;
        RECT 82.150 108.400 114.305 108.900 ;
        RECT 71.925 101.505 75.935 101.555 ;
        RECT 71.925 99.100 75.935 99.155 ;
        RECT 82.150 99.100 82.650 108.400 ;
        RECT 113.795 108.395 114.305 108.400 ;
        RECT 137.805 107.900 138.315 107.905 ;
        RECT 71.925 98.600 82.650 99.100 ;
        RECT 83.450 107.400 138.315 107.900 ;
        RECT 71.925 98.545 75.935 98.600 ;
        RECT 71.925 96.145 75.935 96.195 ;
        RECT 83.450 96.145 83.950 107.400 ;
        RECT 137.805 107.395 138.315 107.400 ;
        RECT 161.815 106.900 162.325 106.905 ;
        RECT 71.925 95.645 83.950 96.145 ;
        RECT 84.650 106.400 162.325 106.900 ;
        RECT 71.925 95.585 75.935 95.645 ;
        RECT 71.925 93.170 75.935 93.235 ;
        RECT 84.650 93.170 85.150 106.400 ;
        RECT 161.815 106.395 162.325 106.400 ;
        RECT 185.825 105.900 186.335 105.905 ;
        RECT 71.925 92.670 85.150 93.170 ;
        RECT 85.950 105.400 186.335 105.900 ;
        RECT 71.925 92.625 75.935 92.670 ;
        RECT 71.925 90.220 75.935 90.275 ;
        RECT 85.950 90.220 86.450 105.400 ;
        RECT 185.825 105.395 186.335 105.400 ;
        RECT 209.835 104.900 210.345 104.905 ;
        RECT 71.925 89.720 86.450 90.220 ;
        RECT 87.250 104.400 210.345 104.900 ;
        RECT 71.925 89.665 75.935 89.720 ;
        RECT 71.925 87.260 75.935 87.315 ;
        RECT 87.250 87.260 87.750 104.400 ;
        RECT 209.835 104.395 210.345 104.400 ;
        RECT 233.845 103.900 234.355 103.905 ;
        RECT 71.925 86.760 87.750 87.260 ;
        RECT 88.750 103.400 234.355 103.900 ;
        RECT 71.925 86.705 75.935 86.760 ;
        RECT 71.925 84.300 75.935 84.355 ;
        RECT 88.750 84.300 89.250 103.400 ;
        RECT 233.845 103.395 234.355 103.400 ;
        RECT 257.855 102.900 258.365 102.905 ;
        RECT 71.925 83.800 89.250 84.300 ;
        RECT 90.150 102.400 258.365 102.900 ;
        RECT 71.925 83.745 75.935 83.800 ;
        RECT 71.925 81.345 75.935 81.395 ;
        RECT 90.150 81.345 90.650 102.400 ;
        RECT 257.855 102.395 258.365 102.400 ;
        RECT 281.865 101.900 282.375 102.405 ;
        RECT 71.925 80.845 90.650 81.345 ;
        RECT 91.650 101.895 282.375 101.900 ;
        RECT 305.875 101.895 306.385 102.405 ;
        RECT 91.650 101.400 282.370 101.895 ;
        RECT 71.925 80.785 75.935 80.845 ;
        RECT 6.000 78.500 31.200 80.500 ;
        RECT 71.925 78.375 75.935 78.435 ;
        RECT 91.650 78.375 92.150 101.400 ;
        RECT 305.880 100.900 306.380 101.895 ;
        RECT 71.925 77.875 92.150 78.375 ;
        RECT 93.250 100.400 306.380 100.900 ;
        RECT 71.925 77.825 75.935 77.875 ;
        RECT 71.925 75.420 75.935 75.475 ;
        RECT 93.250 75.420 93.750 100.400 ;
        RECT 109.445 96.845 110.355 97.755 ;
        RECT 71.925 74.920 93.750 75.420 ;
        RECT 71.925 74.865 75.935 74.920 ;
        RECT 3.995 67.695 4.000 68.505 ;
        RECT 6.000 67.695 6.005 68.505 ;
        RECT 109.450 55.750 110.350 96.845 ;
        RECT 236.300 67.215 236.830 67.745 ;
        RECT 255.480 67.215 256.010 67.745 ;
        RECT 231.240 66.175 231.770 66.705 ;
        RECT 221.120 65.135 221.650 65.665 ;
        RECT 200.880 64.095 201.410 64.625 ;
        RECT 200.885 63.740 201.405 64.095 ;
        RECT 221.125 63.740 221.645 65.135 ;
        RECT 231.245 63.740 231.765 66.175 ;
        RECT 165.465 63.220 201.405 63.740 ;
        RECT 109.450 54.850 152.710 55.750 ;
        RECT 0.995 40.995 1.000 41.805 ;
        RECT 3.000 40.995 3.005 41.805 ;
        RECT 80.315 39.075 80.805 39.565 ;
        RECT 6.000 35.740 6.005 36.230 ;
        RECT 80.320 34.310 80.800 39.075 ;
        RECT 80.315 33.820 80.805 34.310 ;
        RECT 19.030 31.525 20.640 32.070 ;
        RECT 22.630 31.525 24.240 32.070 ;
        RECT 26.230 31.525 27.840 32.070 ;
        RECT 29.830 31.525 31.440 32.070 ;
        RECT 33.430 31.525 35.040 32.070 ;
        RECT 37.030 31.525 38.640 32.070 ;
        RECT 40.630 31.525 42.240 32.070 ;
        RECT 44.230 31.525 45.840 32.070 ;
        RECT 115.280 31.525 116.890 32.070 ;
        RECT 118.880 31.525 120.490 32.070 ;
        RECT 122.480 31.525 124.090 32.070 ;
        RECT 126.080 31.525 127.690 32.070 ;
        RECT 129.680 31.525 131.290 32.070 ;
        RECT 133.280 31.525 134.890 32.070 ;
        RECT 136.880 31.525 138.490 32.070 ;
        RECT 140.480 31.525 142.090 32.070 ;
        RECT 18.035 31.005 49.570 31.525 ;
        RECT 19.030 30.460 20.640 31.005 ;
        RECT 22.630 30.460 24.240 31.005 ;
        RECT 26.230 30.460 27.840 31.005 ;
        RECT 29.830 30.460 31.440 31.005 ;
        RECT 33.430 30.460 35.040 31.005 ;
        RECT 37.030 30.460 38.640 31.005 ;
        RECT 40.630 30.460 42.240 31.005 ;
        RECT 44.230 30.460 45.840 31.005 ;
        RECT 47.925 29.125 48.535 29.135 ;
        RECT 16.755 28.605 48.535 29.125 ;
        RECT 16.755 24.065 17.275 28.605 ;
        RECT 19.030 26.465 20.640 27.010 ;
        RECT 22.630 26.465 24.240 27.010 ;
        RECT 26.230 26.465 27.840 27.010 ;
        RECT 29.830 26.465 31.440 27.010 ;
        RECT 33.430 26.465 35.040 27.010 ;
        RECT 37.030 26.465 38.640 27.010 ;
        RECT 40.630 26.465 42.240 27.010 ;
        RECT 44.230 26.465 45.840 27.010 ;
        RECT 49.050 26.465 49.570 31.005 ;
        RECT 18.035 25.945 49.570 26.465 ;
        RECT 19.030 25.400 20.640 25.945 ;
        RECT 22.630 25.400 24.240 25.945 ;
        RECT 26.230 25.400 27.840 25.945 ;
        RECT 29.830 25.400 31.440 25.945 ;
        RECT 33.430 25.400 35.040 25.945 ;
        RECT 37.030 25.400 38.640 25.945 ;
        RECT 40.630 25.400 42.240 25.945 ;
        RECT 44.230 25.400 45.840 25.945 ;
        RECT 16.755 23.545 46.835 24.065 ;
        RECT 16.755 19.005 17.275 23.545 ;
        RECT 19.030 21.405 20.640 21.950 ;
        RECT 22.630 21.405 24.240 21.950 ;
        RECT 26.230 21.405 27.840 21.950 ;
        RECT 29.830 21.405 31.440 21.950 ;
        RECT 33.430 21.405 35.040 21.950 ;
        RECT 37.030 21.405 38.640 21.950 ;
        RECT 40.630 21.405 42.240 21.950 ;
        RECT 44.230 21.405 45.840 21.950 ;
        RECT 49.050 21.405 49.570 25.945 ;
        RECT 18.035 20.885 49.570 21.405 ;
        RECT 19.030 20.340 20.640 20.885 ;
        RECT 22.630 20.340 24.240 20.885 ;
        RECT 26.230 20.340 27.840 20.885 ;
        RECT 29.830 20.340 31.440 20.885 ;
        RECT 33.430 20.340 35.040 20.885 ;
        RECT 37.030 20.340 38.640 20.885 ;
        RECT 40.630 20.340 42.240 20.885 ;
        RECT 44.230 20.340 45.840 20.885 ;
        RECT 16.755 18.485 46.835 19.005 ;
        RECT 16.755 13.945 17.275 18.485 ;
        RECT 19.030 16.345 20.640 16.890 ;
        RECT 22.630 16.345 24.240 16.890 ;
        RECT 26.230 16.345 27.840 16.890 ;
        RECT 29.830 16.345 31.440 16.890 ;
        RECT 33.430 16.345 35.040 16.890 ;
        RECT 37.030 16.345 38.640 16.890 ;
        RECT 40.630 16.345 42.240 16.890 ;
        RECT 44.230 16.345 45.840 16.890 ;
        RECT 49.050 16.575 49.570 20.885 ;
        RECT 111.550 31.005 143.085 31.525 ;
        RECT 111.550 26.465 112.070 31.005 ;
        RECT 115.280 30.460 116.890 31.005 ;
        RECT 118.880 30.460 120.490 31.005 ;
        RECT 122.480 30.460 124.090 31.005 ;
        RECT 126.080 30.460 127.690 31.005 ;
        RECT 129.680 30.460 131.290 31.005 ;
        RECT 133.280 30.460 134.890 31.005 ;
        RECT 136.880 30.460 138.490 31.005 ;
        RECT 140.480 30.460 142.090 31.005 ;
        RECT 112.585 29.125 113.195 29.135 ;
        RECT 112.585 28.605 144.365 29.125 ;
        RECT 115.280 26.465 116.890 27.010 ;
        RECT 118.880 26.465 120.490 27.010 ;
        RECT 122.480 26.465 124.090 27.010 ;
        RECT 126.080 26.465 127.690 27.010 ;
        RECT 129.680 26.465 131.290 27.010 ;
        RECT 133.280 26.465 134.890 27.010 ;
        RECT 136.880 26.465 138.490 27.010 ;
        RECT 140.480 26.465 142.090 27.010 ;
        RECT 111.550 25.945 143.085 26.465 ;
        RECT 111.550 21.405 112.070 25.945 ;
        RECT 115.280 25.400 116.890 25.945 ;
        RECT 118.880 25.400 120.490 25.945 ;
        RECT 122.480 25.400 124.090 25.945 ;
        RECT 126.080 25.400 127.690 25.945 ;
        RECT 129.680 25.400 131.290 25.945 ;
        RECT 133.280 25.400 134.890 25.945 ;
        RECT 136.880 25.400 138.490 25.945 ;
        RECT 140.480 25.400 142.090 25.945 ;
        RECT 143.845 24.065 144.365 28.605 ;
        RECT 114.285 23.545 144.365 24.065 ;
        RECT 115.280 21.405 116.890 21.950 ;
        RECT 118.880 21.405 120.490 21.950 ;
        RECT 122.480 21.405 124.090 21.950 ;
        RECT 126.080 21.405 127.690 21.950 ;
        RECT 129.680 21.405 131.290 21.950 ;
        RECT 133.280 21.405 134.890 21.950 ;
        RECT 136.880 21.405 138.490 21.950 ;
        RECT 140.480 21.405 142.090 21.950 ;
        RECT 111.550 20.885 143.085 21.405 ;
        RECT 111.550 16.575 112.070 20.885 ;
        RECT 115.280 20.340 116.890 20.885 ;
        RECT 118.880 20.340 120.490 20.885 ;
        RECT 122.480 20.340 124.090 20.885 ;
        RECT 126.080 20.340 127.690 20.885 ;
        RECT 129.680 20.340 131.290 20.885 ;
        RECT 133.280 20.340 134.890 20.885 ;
        RECT 136.880 20.340 138.490 20.885 ;
        RECT 140.480 20.340 142.090 20.885 ;
        RECT 143.845 19.005 144.365 23.545 ;
        RECT 114.285 18.485 144.365 19.005 ;
        RECT 49.045 16.345 49.575 16.575 ;
        RECT 18.035 15.825 49.575 16.345 ;
        RECT 19.030 15.280 20.640 15.825 ;
        RECT 22.630 15.280 24.240 15.825 ;
        RECT 26.230 15.280 27.840 15.825 ;
        RECT 29.830 15.280 31.440 15.825 ;
        RECT 33.430 15.280 35.040 15.825 ;
        RECT 37.030 15.280 38.640 15.825 ;
        RECT 40.630 15.280 42.240 15.825 ;
        RECT 44.230 15.280 45.840 15.825 ;
        RECT 49.045 15.265 49.575 15.825 ;
        RECT 111.545 16.345 112.075 16.575 ;
        RECT 115.280 16.345 116.890 16.890 ;
        RECT 118.880 16.345 120.490 16.890 ;
        RECT 122.480 16.345 124.090 16.890 ;
        RECT 126.080 16.345 127.690 16.890 ;
        RECT 129.680 16.345 131.290 16.890 ;
        RECT 133.280 16.345 134.890 16.890 ;
        RECT 136.880 16.345 138.490 16.890 ;
        RECT 140.480 16.345 142.090 16.890 ;
        RECT 111.545 15.825 143.085 16.345 ;
        RECT 111.545 15.265 112.075 15.825 ;
        RECT 115.280 15.280 116.890 15.825 ;
        RECT 118.880 15.280 120.490 15.825 ;
        RECT 122.480 15.280 124.090 15.825 ;
        RECT 126.080 15.280 127.690 15.825 ;
        RECT 129.680 15.280 131.290 15.825 ;
        RECT 133.280 15.280 134.890 15.825 ;
        RECT 136.880 15.280 138.490 15.825 ;
        RECT 140.480 15.280 142.090 15.825 ;
        RECT 143.845 13.945 144.365 18.485 ;
        RECT 16.755 13.425 46.835 13.945 ;
        RECT 114.285 13.425 144.365 13.945 ;
        RECT 0.995 5.670 1.000 6.160 ;
        RECT 3.000 5.670 3.005 6.160 ;
        RECT 67.455 5.765 76.145 6.855 ;
        RECT 84.975 5.765 93.665 6.855 ;
        RECT 71.250 2.655 72.150 5.765 ;
        RECT 88.950 4.200 89.850 5.765 ;
        RECT 88.950 3.300 133.390 4.200 ;
        RECT 113.170 2.655 114.070 2.660 ;
        RECT 71.250 1.755 114.070 2.655 ;
        RECT 113.170 1.000 114.070 1.755 ;
        RECT 132.490 1.000 133.390 3.300 ;
        RECT 151.810 1.000 152.710 54.850 ;
        RECT 165.465 5.100 165.985 63.220 ;
        RECT 167.865 61.705 168.385 62.700 ;
        RECT 167.320 60.095 168.930 61.705 ;
        RECT 167.865 58.105 168.385 60.095 ;
        RECT 167.320 56.495 168.930 58.105 ;
        RECT 167.865 54.505 168.385 56.495 ;
        RECT 167.320 52.895 168.930 54.505 ;
        RECT 167.865 50.905 168.385 52.895 ;
        RECT 167.320 49.295 168.930 50.905 ;
        RECT 167.865 47.305 168.385 49.295 ;
        RECT 167.320 45.695 168.930 47.305 ;
        RECT 167.865 43.705 168.385 45.695 ;
        RECT 167.320 42.095 168.930 43.705 ;
        RECT 167.865 40.105 168.385 42.095 ;
        RECT 167.320 38.495 168.930 40.105 ;
        RECT 167.865 36.505 168.385 38.495 ;
        RECT 167.320 34.895 168.930 36.505 ;
        RECT 167.865 32.905 168.385 34.895 ;
        RECT 167.320 31.295 168.930 32.905 ;
        RECT 167.865 29.305 168.385 31.295 ;
        RECT 167.320 27.695 168.930 29.305 ;
        RECT 167.865 25.705 168.385 27.695 ;
        RECT 167.320 24.095 168.930 25.705 ;
        RECT 167.865 22.105 168.385 24.095 ;
        RECT 167.320 20.495 168.930 22.105 ;
        RECT 167.865 18.505 168.385 20.495 ;
        RECT 167.320 16.895 168.930 18.505 ;
        RECT 167.865 14.905 168.385 16.895 ;
        RECT 167.320 13.295 168.930 14.905 ;
        RECT 167.865 11.305 168.385 13.295 ;
        RECT 167.320 9.695 168.930 11.305 ;
        RECT 167.865 7.705 168.385 9.695 ;
        RECT 167.320 6.095 168.930 7.705 ;
        RECT 167.210 4.580 167.740 4.585 ;
        RECT 167.865 4.580 168.385 6.095 ;
        RECT 170.525 5.100 171.045 63.220 ;
        RECT 172.925 61.705 173.445 62.700 ;
        RECT 172.380 60.095 173.990 61.705 ;
        RECT 172.925 58.105 173.445 60.095 ;
        RECT 172.380 56.495 173.990 58.105 ;
        RECT 172.925 54.505 173.445 56.495 ;
        RECT 172.380 52.895 173.990 54.505 ;
        RECT 172.925 50.905 173.445 52.895 ;
        RECT 172.380 49.295 173.990 50.905 ;
        RECT 172.925 47.305 173.445 49.295 ;
        RECT 172.380 45.695 173.990 47.305 ;
        RECT 172.925 43.705 173.445 45.695 ;
        RECT 172.380 42.095 173.990 43.705 ;
        RECT 172.925 40.105 173.445 42.095 ;
        RECT 172.380 38.495 173.990 40.105 ;
        RECT 172.925 36.505 173.445 38.495 ;
        RECT 172.380 34.895 173.990 36.505 ;
        RECT 172.925 32.905 173.445 34.895 ;
        RECT 172.380 31.295 173.990 32.905 ;
        RECT 172.925 29.305 173.445 31.295 ;
        RECT 172.380 27.695 173.990 29.305 ;
        RECT 172.925 25.705 173.445 27.695 ;
        RECT 172.380 24.095 173.990 25.705 ;
        RECT 172.925 22.105 173.445 24.095 ;
        RECT 172.380 20.495 173.990 22.105 ;
        RECT 172.925 18.505 173.445 20.495 ;
        RECT 172.380 16.895 173.990 18.505 ;
        RECT 172.925 14.905 173.445 16.895 ;
        RECT 172.380 13.295 173.990 14.905 ;
        RECT 172.925 11.305 173.445 13.295 ;
        RECT 172.380 9.695 173.990 11.305 ;
        RECT 172.925 7.705 173.445 9.695 ;
        RECT 172.380 6.095 173.990 7.705 ;
        RECT 172.925 4.580 173.445 6.095 ;
        RECT 175.585 5.100 176.105 63.220 ;
        RECT 177.985 61.705 178.505 62.700 ;
        RECT 177.440 60.095 179.050 61.705 ;
        RECT 177.985 58.105 178.505 60.095 ;
        RECT 177.440 56.495 179.050 58.105 ;
        RECT 177.985 54.505 178.505 56.495 ;
        RECT 177.440 52.895 179.050 54.505 ;
        RECT 177.985 50.905 178.505 52.895 ;
        RECT 177.440 49.295 179.050 50.905 ;
        RECT 177.985 47.305 178.505 49.295 ;
        RECT 177.440 45.695 179.050 47.305 ;
        RECT 177.985 43.705 178.505 45.695 ;
        RECT 177.440 42.095 179.050 43.705 ;
        RECT 177.985 40.105 178.505 42.095 ;
        RECT 177.440 38.495 179.050 40.105 ;
        RECT 177.985 36.505 178.505 38.495 ;
        RECT 177.440 34.895 179.050 36.505 ;
        RECT 177.985 32.905 178.505 34.895 ;
        RECT 177.440 31.295 179.050 32.905 ;
        RECT 177.985 29.305 178.505 31.295 ;
        RECT 177.440 27.695 179.050 29.305 ;
        RECT 177.985 25.705 178.505 27.695 ;
        RECT 177.440 24.095 179.050 25.705 ;
        RECT 177.985 22.105 178.505 24.095 ;
        RECT 177.440 20.495 179.050 22.105 ;
        RECT 177.985 18.505 178.505 20.495 ;
        RECT 177.440 16.895 179.050 18.505 ;
        RECT 177.985 14.905 178.505 16.895 ;
        RECT 177.440 13.295 179.050 14.905 ;
        RECT 177.985 11.305 178.505 13.295 ;
        RECT 177.440 9.695 179.050 11.305 ;
        RECT 177.985 7.705 178.505 9.695 ;
        RECT 177.440 6.095 179.050 7.705 ;
        RECT 177.985 4.580 178.505 6.095 ;
        RECT 180.645 5.100 181.165 63.220 ;
        RECT 183.045 61.705 183.565 62.700 ;
        RECT 182.500 60.095 184.110 61.705 ;
        RECT 183.045 58.105 183.565 60.095 ;
        RECT 182.500 56.495 184.110 58.105 ;
        RECT 183.045 54.505 183.565 56.495 ;
        RECT 182.500 52.895 184.110 54.505 ;
        RECT 183.045 50.905 183.565 52.895 ;
        RECT 182.500 49.295 184.110 50.905 ;
        RECT 183.045 47.305 183.565 49.295 ;
        RECT 182.500 45.695 184.110 47.305 ;
        RECT 183.045 43.705 183.565 45.695 ;
        RECT 182.500 42.095 184.110 43.705 ;
        RECT 183.045 40.105 183.565 42.095 ;
        RECT 182.500 38.495 184.110 40.105 ;
        RECT 183.045 36.505 183.565 38.495 ;
        RECT 182.500 34.895 184.110 36.505 ;
        RECT 183.045 32.905 183.565 34.895 ;
        RECT 182.500 31.295 184.110 32.905 ;
        RECT 183.045 29.305 183.565 31.295 ;
        RECT 182.500 27.695 184.110 29.305 ;
        RECT 183.045 25.705 183.565 27.695 ;
        RECT 182.500 24.095 184.110 25.705 ;
        RECT 183.045 22.105 183.565 24.095 ;
        RECT 182.500 20.495 184.110 22.105 ;
        RECT 183.045 18.505 183.565 20.495 ;
        RECT 182.500 16.895 184.110 18.505 ;
        RECT 183.045 14.905 183.565 16.895 ;
        RECT 182.500 13.295 184.110 14.905 ;
        RECT 183.045 11.305 183.565 13.295 ;
        RECT 182.500 9.695 184.110 11.305 ;
        RECT 183.045 7.705 183.565 9.695 ;
        RECT 182.500 6.095 184.110 7.705 ;
        RECT 183.045 4.580 183.565 6.095 ;
        RECT 185.705 5.100 186.225 63.220 ;
        RECT 188.105 61.705 188.625 62.700 ;
        RECT 187.560 60.095 189.170 61.705 ;
        RECT 188.105 58.105 188.625 60.095 ;
        RECT 187.560 56.495 189.170 58.105 ;
        RECT 188.105 54.505 188.625 56.495 ;
        RECT 187.560 52.895 189.170 54.505 ;
        RECT 188.105 50.905 188.625 52.895 ;
        RECT 187.560 49.295 189.170 50.905 ;
        RECT 188.105 47.305 188.625 49.295 ;
        RECT 187.560 45.695 189.170 47.305 ;
        RECT 188.105 43.705 188.625 45.695 ;
        RECT 187.560 42.095 189.170 43.705 ;
        RECT 188.105 40.105 188.625 42.095 ;
        RECT 187.560 38.495 189.170 40.105 ;
        RECT 188.105 36.505 188.625 38.495 ;
        RECT 187.560 34.895 189.170 36.505 ;
        RECT 188.105 32.905 188.625 34.895 ;
        RECT 187.560 31.295 189.170 32.905 ;
        RECT 188.105 29.305 188.625 31.295 ;
        RECT 187.560 27.695 189.170 29.305 ;
        RECT 188.105 25.705 188.625 27.695 ;
        RECT 187.560 24.095 189.170 25.705 ;
        RECT 188.105 22.105 188.625 24.095 ;
        RECT 187.560 20.495 189.170 22.105 ;
        RECT 188.105 18.505 188.625 20.495 ;
        RECT 187.560 16.895 189.170 18.505 ;
        RECT 188.105 14.905 188.625 16.895 ;
        RECT 187.560 13.295 189.170 14.905 ;
        RECT 188.105 11.305 188.625 13.295 ;
        RECT 187.560 9.695 189.170 11.305 ;
        RECT 188.105 7.705 188.625 9.695 ;
        RECT 187.560 6.095 189.170 7.705 ;
        RECT 188.105 4.580 188.625 6.095 ;
        RECT 190.765 5.100 191.285 63.220 ;
        RECT 193.165 61.705 193.685 62.700 ;
        RECT 192.620 60.095 194.230 61.705 ;
        RECT 193.165 58.105 193.685 60.095 ;
        RECT 192.620 56.495 194.230 58.105 ;
        RECT 193.165 54.505 193.685 56.495 ;
        RECT 192.620 52.895 194.230 54.505 ;
        RECT 193.165 50.905 193.685 52.895 ;
        RECT 192.620 49.295 194.230 50.905 ;
        RECT 193.165 47.305 193.685 49.295 ;
        RECT 192.620 45.695 194.230 47.305 ;
        RECT 193.165 43.705 193.685 45.695 ;
        RECT 192.620 42.095 194.230 43.705 ;
        RECT 193.165 40.105 193.685 42.095 ;
        RECT 192.620 38.495 194.230 40.105 ;
        RECT 193.165 36.505 193.685 38.495 ;
        RECT 192.620 34.895 194.230 36.505 ;
        RECT 193.165 32.905 193.685 34.895 ;
        RECT 192.620 31.295 194.230 32.905 ;
        RECT 193.165 29.305 193.685 31.295 ;
        RECT 192.620 27.695 194.230 29.305 ;
        RECT 193.165 25.705 193.685 27.695 ;
        RECT 192.620 24.095 194.230 25.705 ;
        RECT 193.165 22.105 193.685 24.095 ;
        RECT 192.620 20.495 194.230 22.105 ;
        RECT 193.165 18.505 193.685 20.495 ;
        RECT 192.620 16.895 194.230 18.505 ;
        RECT 193.165 14.905 193.685 16.895 ;
        RECT 192.620 13.295 194.230 14.905 ;
        RECT 193.165 11.305 193.685 13.295 ;
        RECT 192.620 9.695 194.230 11.305 ;
        RECT 193.165 7.705 193.685 9.695 ;
        RECT 192.620 6.095 194.230 7.705 ;
        RECT 193.165 4.580 193.685 6.095 ;
        RECT 195.825 5.100 196.345 63.220 ;
        RECT 198.225 61.705 198.745 62.700 ;
        RECT 197.680 60.095 199.290 61.705 ;
        RECT 198.225 58.105 198.745 60.095 ;
        RECT 197.680 56.495 199.290 58.105 ;
        RECT 198.225 54.505 198.745 56.495 ;
        RECT 197.680 52.895 199.290 54.505 ;
        RECT 198.225 50.905 198.745 52.895 ;
        RECT 197.680 49.295 199.290 50.905 ;
        RECT 198.225 47.305 198.745 49.295 ;
        RECT 197.680 45.695 199.290 47.305 ;
        RECT 198.225 43.705 198.745 45.695 ;
        RECT 197.680 42.095 199.290 43.705 ;
        RECT 198.225 40.105 198.745 42.095 ;
        RECT 197.680 38.495 199.290 40.105 ;
        RECT 198.225 36.505 198.745 38.495 ;
        RECT 197.680 34.895 199.290 36.505 ;
        RECT 198.225 32.905 198.745 34.895 ;
        RECT 197.680 31.295 199.290 32.905 ;
        RECT 198.225 29.305 198.745 31.295 ;
        RECT 197.680 27.695 199.290 29.305 ;
        RECT 198.225 25.705 198.745 27.695 ;
        RECT 197.680 24.095 199.290 25.705 ;
        RECT 198.225 22.105 198.745 24.095 ;
        RECT 197.680 20.495 199.290 22.105 ;
        RECT 198.225 18.505 198.745 20.495 ;
        RECT 197.680 16.895 199.290 18.505 ;
        RECT 198.225 14.905 198.745 16.895 ;
        RECT 197.680 13.295 199.290 14.905 ;
        RECT 198.225 11.305 198.745 13.295 ;
        RECT 197.680 9.695 199.290 11.305 ;
        RECT 198.225 7.705 198.745 9.695 ;
        RECT 197.680 6.095 199.290 7.705 ;
        RECT 198.225 4.580 198.745 6.095 ;
        RECT 200.885 5.100 201.405 63.220 ;
        RECT 205.945 63.220 221.645 63.740 ;
        RECT 203.285 61.705 203.805 62.700 ;
        RECT 202.740 60.095 204.350 61.705 ;
        RECT 203.285 58.105 203.805 60.095 ;
        RECT 202.740 56.495 204.350 58.105 ;
        RECT 203.285 54.505 203.805 56.495 ;
        RECT 202.740 52.895 204.350 54.505 ;
        RECT 203.285 50.905 203.805 52.895 ;
        RECT 202.740 49.295 204.350 50.905 ;
        RECT 203.285 47.305 203.805 49.295 ;
        RECT 202.740 45.695 204.350 47.305 ;
        RECT 203.285 43.705 203.805 45.695 ;
        RECT 202.740 42.095 204.350 43.705 ;
        RECT 203.285 40.105 203.805 42.095 ;
        RECT 202.740 38.495 204.350 40.105 ;
        RECT 203.285 36.505 203.805 38.495 ;
        RECT 202.740 34.895 204.350 36.505 ;
        RECT 203.285 32.905 203.805 34.895 ;
        RECT 202.740 31.295 204.350 32.905 ;
        RECT 203.285 29.305 203.805 31.295 ;
        RECT 202.740 27.695 204.350 29.305 ;
        RECT 203.285 25.705 203.805 27.695 ;
        RECT 202.740 24.095 204.350 25.705 ;
        RECT 203.285 22.105 203.805 24.095 ;
        RECT 202.740 20.495 204.350 22.105 ;
        RECT 203.285 18.505 203.805 20.495 ;
        RECT 202.740 16.895 204.350 18.505 ;
        RECT 203.285 14.905 203.805 16.895 ;
        RECT 202.740 13.295 204.350 14.905 ;
        RECT 203.285 11.305 203.805 13.295 ;
        RECT 202.740 9.695 204.350 11.305 ;
        RECT 203.285 7.705 203.805 9.695 ;
        RECT 202.740 6.095 204.350 7.705 ;
        RECT 203.285 4.580 203.805 6.095 ;
        RECT 205.945 5.100 206.465 63.220 ;
        RECT 208.345 61.705 208.865 62.700 ;
        RECT 207.800 60.095 209.410 61.705 ;
        RECT 208.345 58.105 208.865 60.095 ;
        RECT 207.800 56.495 209.410 58.105 ;
        RECT 208.345 54.505 208.865 56.495 ;
        RECT 207.800 52.895 209.410 54.505 ;
        RECT 208.345 50.905 208.865 52.895 ;
        RECT 207.800 49.295 209.410 50.905 ;
        RECT 208.345 47.305 208.865 49.295 ;
        RECT 207.800 45.695 209.410 47.305 ;
        RECT 208.345 43.705 208.865 45.695 ;
        RECT 207.800 42.095 209.410 43.705 ;
        RECT 208.345 40.105 208.865 42.095 ;
        RECT 207.800 38.495 209.410 40.105 ;
        RECT 208.345 36.505 208.865 38.495 ;
        RECT 207.800 34.895 209.410 36.505 ;
        RECT 208.345 32.905 208.865 34.895 ;
        RECT 207.800 31.295 209.410 32.905 ;
        RECT 208.345 29.305 208.865 31.295 ;
        RECT 207.800 27.695 209.410 29.305 ;
        RECT 208.345 25.705 208.865 27.695 ;
        RECT 207.800 24.095 209.410 25.705 ;
        RECT 208.345 22.105 208.865 24.095 ;
        RECT 207.800 20.495 209.410 22.105 ;
        RECT 208.345 18.505 208.865 20.495 ;
        RECT 207.800 16.895 209.410 18.505 ;
        RECT 208.345 14.905 208.865 16.895 ;
        RECT 207.800 13.295 209.410 14.905 ;
        RECT 208.345 11.305 208.865 13.295 ;
        RECT 207.800 9.695 209.410 11.305 ;
        RECT 208.345 7.705 208.865 9.695 ;
        RECT 207.800 6.095 209.410 7.705 ;
        RECT 208.345 4.580 208.865 6.095 ;
        RECT 211.005 5.100 211.525 63.220 ;
        RECT 213.405 61.705 213.925 62.700 ;
        RECT 212.860 60.095 214.470 61.705 ;
        RECT 213.405 58.105 213.925 60.095 ;
        RECT 212.860 56.495 214.470 58.105 ;
        RECT 213.405 54.505 213.925 56.495 ;
        RECT 212.860 52.895 214.470 54.505 ;
        RECT 213.405 50.905 213.925 52.895 ;
        RECT 212.860 49.295 214.470 50.905 ;
        RECT 213.405 47.305 213.925 49.295 ;
        RECT 212.860 45.695 214.470 47.305 ;
        RECT 213.405 43.705 213.925 45.695 ;
        RECT 212.860 42.095 214.470 43.705 ;
        RECT 213.405 40.105 213.925 42.095 ;
        RECT 212.860 38.495 214.470 40.105 ;
        RECT 213.405 36.505 213.925 38.495 ;
        RECT 212.860 34.895 214.470 36.505 ;
        RECT 213.405 32.905 213.925 34.895 ;
        RECT 212.860 31.295 214.470 32.905 ;
        RECT 213.405 29.305 213.925 31.295 ;
        RECT 212.860 27.695 214.470 29.305 ;
        RECT 213.405 25.705 213.925 27.695 ;
        RECT 212.860 24.095 214.470 25.705 ;
        RECT 213.405 22.105 213.925 24.095 ;
        RECT 212.860 20.495 214.470 22.105 ;
        RECT 213.405 18.505 213.925 20.495 ;
        RECT 212.860 16.895 214.470 18.505 ;
        RECT 213.405 14.905 213.925 16.895 ;
        RECT 212.860 13.295 214.470 14.905 ;
        RECT 213.405 11.305 213.925 13.295 ;
        RECT 212.860 9.695 214.470 11.305 ;
        RECT 213.405 7.705 213.925 9.695 ;
        RECT 212.860 6.095 214.470 7.705 ;
        RECT 213.405 4.580 213.925 6.095 ;
        RECT 216.065 5.100 216.585 63.220 ;
        RECT 218.465 61.705 218.985 62.700 ;
        RECT 217.920 60.095 219.530 61.705 ;
        RECT 218.465 58.105 218.985 60.095 ;
        RECT 217.920 56.495 219.530 58.105 ;
        RECT 218.465 54.505 218.985 56.495 ;
        RECT 217.920 52.895 219.530 54.505 ;
        RECT 218.465 50.905 218.985 52.895 ;
        RECT 217.920 49.295 219.530 50.905 ;
        RECT 218.465 47.305 218.985 49.295 ;
        RECT 217.920 45.695 219.530 47.305 ;
        RECT 218.465 43.705 218.985 45.695 ;
        RECT 217.920 42.095 219.530 43.705 ;
        RECT 218.465 40.105 218.985 42.095 ;
        RECT 217.920 38.495 219.530 40.105 ;
        RECT 218.465 36.505 218.985 38.495 ;
        RECT 217.920 34.895 219.530 36.505 ;
        RECT 218.465 32.905 218.985 34.895 ;
        RECT 217.920 31.295 219.530 32.905 ;
        RECT 218.465 29.305 218.985 31.295 ;
        RECT 217.920 27.695 219.530 29.305 ;
        RECT 218.465 25.705 218.985 27.695 ;
        RECT 217.920 24.095 219.530 25.705 ;
        RECT 218.465 22.105 218.985 24.095 ;
        RECT 217.920 20.495 219.530 22.105 ;
        RECT 218.465 18.505 218.985 20.495 ;
        RECT 217.920 16.895 219.530 18.505 ;
        RECT 218.465 14.905 218.985 16.895 ;
        RECT 217.920 13.295 219.530 14.905 ;
        RECT 218.465 11.305 218.985 13.295 ;
        RECT 217.920 9.695 219.530 11.305 ;
        RECT 218.465 7.705 218.985 9.695 ;
        RECT 217.920 6.095 219.530 7.705 ;
        RECT 218.465 4.580 218.985 6.095 ;
        RECT 221.125 5.100 221.645 63.220 ;
        RECT 226.185 63.220 231.765 63.740 ;
        RECT 223.525 61.705 224.045 62.700 ;
        RECT 222.980 60.095 224.590 61.705 ;
        RECT 223.525 58.105 224.045 60.095 ;
        RECT 222.980 56.495 224.590 58.105 ;
        RECT 223.525 54.505 224.045 56.495 ;
        RECT 222.980 52.895 224.590 54.505 ;
        RECT 223.525 50.905 224.045 52.895 ;
        RECT 222.980 49.295 224.590 50.905 ;
        RECT 223.525 47.305 224.045 49.295 ;
        RECT 222.980 45.695 224.590 47.305 ;
        RECT 223.525 43.705 224.045 45.695 ;
        RECT 222.980 42.095 224.590 43.705 ;
        RECT 223.525 40.105 224.045 42.095 ;
        RECT 222.980 38.495 224.590 40.105 ;
        RECT 223.525 36.505 224.045 38.495 ;
        RECT 222.980 34.895 224.590 36.505 ;
        RECT 223.525 32.905 224.045 34.895 ;
        RECT 222.980 31.295 224.590 32.905 ;
        RECT 223.525 29.305 224.045 31.295 ;
        RECT 222.980 27.695 224.590 29.305 ;
        RECT 223.525 25.705 224.045 27.695 ;
        RECT 222.980 24.095 224.590 25.705 ;
        RECT 223.525 22.105 224.045 24.095 ;
        RECT 222.980 20.495 224.590 22.105 ;
        RECT 223.525 18.505 224.045 20.495 ;
        RECT 222.980 16.895 224.590 18.505 ;
        RECT 223.525 14.905 224.045 16.895 ;
        RECT 222.980 13.295 224.590 14.905 ;
        RECT 223.525 11.305 224.045 13.295 ;
        RECT 222.980 9.695 224.590 11.305 ;
        RECT 223.525 7.705 224.045 9.695 ;
        RECT 222.980 6.095 224.590 7.705 ;
        RECT 223.525 4.580 224.045 6.095 ;
        RECT 226.185 5.100 226.705 63.220 ;
        RECT 228.585 61.705 229.105 62.700 ;
        RECT 228.040 60.095 229.650 61.705 ;
        RECT 228.585 58.105 229.105 60.095 ;
        RECT 228.040 56.495 229.650 58.105 ;
        RECT 228.585 54.505 229.105 56.495 ;
        RECT 228.040 52.895 229.650 54.505 ;
        RECT 228.585 50.905 229.105 52.895 ;
        RECT 228.040 49.295 229.650 50.905 ;
        RECT 228.585 47.305 229.105 49.295 ;
        RECT 228.040 45.695 229.650 47.305 ;
        RECT 228.585 43.705 229.105 45.695 ;
        RECT 228.040 42.095 229.650 43.705 ;
        RECT 228.585 40.105 229.105 42.095 ;
        RECT 228.040 38.495 229.650 40.105 ;
        RECT 228.585 36.505 229.105 38.495 ;
        RECT 228.040 34.895 229.650 36.505 ;
        RECT 228.585 32.905 229.105 34.895 ;
        RECT 228.040 31.295 229.650 32.905 ;
        RECT 228.585 29.305 229.105 31.295 ;
        RECT 228.040 27.695 229.650 29.305 ;
        RECT 228.585 25.705 229.105 27.695 ;
        RECT 228.040 24.095 229.650 25.705 ;
        RECT 228.585 22.105 229.105 24.095 ;
        RECT 228.040 20.495 229.650 22.105 ;
        RECT 228.585 18.505 229.105 20.495 ;
        RECT 228.040 16.895 229.650 18.505 ;
        RECT 228.585 14.905 229.105 16.895 ;
        RECT 228.040 13.295 229.650 14.905 ;
        RECT 228.585 11.305 229.105 13.295 ;
        RECT 228.040 9.695 229.650 11.305 ;
        RECT 228.585 7.705 229.105 9.695 ;
        RECT 228.040 6.095 229.650 7.705 ;
        RECT 228.585 4.580 229.105 6.095 ;
        RECT 231.245 5.100 231.765 63.220 ;
        RECT 233.645 61.705 234.165 62.700 ;
        RECT 233.100 60.095 234.710 61.705 ;
        RECT 233.645 58.105 234.165 60.095 ;
        RECT 233.100 56.495 234.710 58.105 ;
        RECT 233.645 54.505 234.165 56.495 ;
        RECT 233.100 52.895 234.710 54.505 ;
        RECT 233.645 50.905 234.165 52.895 ;
        RECT 233.100 49.295 234.710 50.905 ;
        RECT 233.645 47.305 234.165 49.295 ;
        RECT 233.100 45.695 234.710 47.305 ;
        RECT 233.645 43.705 234.165 45.695 ;
        RECT 233.100 42.095 234.710 43.705 ;
        RECT 233.645 40.105 234.165 42.095 ;
        RECT 233.100 38.495 234.710 40.105 ;
        RECT 233.645 36.505 234.165 38.495 ;
        RECT 233.100 34.895 234.710 36.505 ;
        RECT 233.645 32.905 234.165 34.895 ;
        RECT 233.100 31.295 234.710 32.905 ;
        RECT 233.645 29.305 234.165 31.295 ;
        RECT 233.100 27.695 234.710 29.305 ;
        RECT 233.645 25.705 234.165 27.695 ;
        RECT 233.100 24.095 234.710 25.705 ;
        RECT 233.645 22.105 234.165 24.095 ;
        RECT 233.100 20.495 234.710 22.105 ;
        RECT 233.645 18.505 234.165 20.495 ;
        RECT 233.100 16.895 234.710 18.505 ;
        RECT 233.645 14.905 234.165 16.895 ;
        RECT 233.100 13.295 234.710 14.905 ;
        RECT 233.645 11.305 234.165 13.295 ;
        RECT 233.100 9.695 234.710 11.305 ;
        RECT 233.645 7.705 234.165 9.695 ;
        RECT 233.100 6.095 234.710 7.705 ;
        RECT 233.645 4.580 234.165 6.095 ;
        RECT 236.305 5.100 236.825 67.215 ;
        RECT 238.705 61.705 239.225 62.700 ;
        RECT 238.160 60.095 239.770 61.705 ;
        RECT 238.705 58.105 239.225 60.095 ;
        RECT 238.160 56.495 239.770 58.105 ;
        RECT 238.705 54.505 239.225 56.495 ;
        RECT 241.520 56.100 242.010 56.105 ;
        RECT 243.385 56.100 243.865 62.040 ;
        RECT 245.765 61.705 246.285 62.700 ;
        RECT 245.220 60.095 246.830 61.705 ;
        RECT 245.765 58.105 246.285 60.095 ;
        RECT 245.220 56.495 246.830 58.105 ;
        RECT 241.520 55.620 243.865 56.100 ;
        RECT 241.520 55.615 242.010 55.620 ;
        RECT 238.160 52.895 239.770 54.505 ;
        RECT 238.705 50.905 239.225 52.895 ;
        RECT 238.160 49.295 239.770 50.905 ;
        RECT 238.705 47.305 239.225 49.295 ;
        RECT 243.385 48.960 243.865 55.620 ;
        RECT 245.765 54.505 246.285 56.495 ;
        RECT 248.580 56.100 249.070 56.105 ;
        RECT 250.445 56.100 250.925 62.040 ;
        RECT 252.825 61.705 253.345 62.700 ;
        RECT 252.280 60.095 253.890 61.705 ;
        RECT 252.825 58.105 253.345 60.095 ;
        RECT 252.280 56.495 253.890 58.105 ;
        RECT 248.580 55.620 250.925 56.100 ;
        RECT 248.580 55.615 249.070 55.620 ;
        RECT 245.220 52.895 246.830 54.505 ;
        RECT 245.765 50.905 246.285 52.895 ;
        RECT 245.220 49.295 246.830 50.905 ;
        RECT 238.160 45.695 239.770 47.305 ;
        RECT 238.705 43.705 239.225 45.695 ;
        RECT 241.520 45.300 242.010 45.305 ;
        RECT 243.385 45.300 243.865 47.640 ;
        RECT 245.765 47.305 246.285 49.295 ;
        RECT 250.445 48.960 250.925 55.620 ;
        RECT 252.825 54.505 253.345 56.495 ;
        RECT 252.280 52.895 253.890 54.505 ;
        RECT 252.825 50.905 253.345 52.895 ;
        RECT 252.280 49.295 253.890 50.905 ;
        RECT 245.220 45.695 246.830 47.305 ;
        RECT 241.520 44.820 243.865 45.300 ;
        RECT 241.520 44.815 242.010 44.820 ;
        RECT 238.160 42.095 239.770 43.705 ;
        RECT 238.705 40.105 239.225 42.095 ;
        RECT 243.385 41.760 243.865 44.820 ;
        RECT 245.765 43.705 246.285 45.695 ;
        RECT 248.580 45.300 249.070 45.305 ;
        RECT 250.445 45.300 250.925 47.640 ;
        RECT 252.825 47.305 253.345 49.295 ;
        RECT 252.280 45.695 253.890 47.305 ;
        RECT 248.580 44.820 250.925 45.300 ;
        RECT 248.580 44.815 249.070 44.820 ;
        RECT 245.220 42.095 246.830 43.705 ;
        RECT 238.160 38.495 239.770 40.105 ;
        RECT 238.705 36.505 239.225 38.495 ;
        RECT 241.520 38.100 242.010 38.105 ;
        RECT 243.385 38.100 243.865 40.440 ;
        RECT 245.765 40.105 246.285 42.095 ;
        RECT 250.445 41.760 250.925 44.820 ;
        RECT 252.825 43.705 253.345 45.695 ;
        RECT 252.280 42.095 253.890 43.705 ;
        RECT 245.220 38.495 246.830 40.105 ;
        RECT 241.520 37.620 243.865 38.100 ;
        RECT 241.520 37.615 242.010 37.620 ;
        RECT 238.160 34.895 239.770 36.505 ;
        RECT 241.520 35.040 242.010 35.045 ;
        RECT 243.385 35.040 243.865 36.840 ;
        RECT 245.765 36.505 246.285 38.495 ;
        RECT 248.580 38.100 249.070 38.105 ;
        RECT 250.445 38.100 250.925 40.440 ;
        RECT 252.825 40.105 253.345 42.095 ;
        RECT 252.280 38.495 253.890 40.105 ;
        RECT 248.580 37.620 250.925 38.100 ;
        RECT 248.580 37.615 249.070 37.620 ;
        RECT 248.580 36.840 249.070 36.845 ;
        RECT 238.705 32.905 239.225 34.895 ;
        RECT 241.520 34.560 243.865 35.040 ;
        RECT 245.220 34.895 246.830 36.505 ;
        RECT 248.580 36.360 250.925 36.840 ;
        RECT 252.825 36.505 253.345 38.495 ;
        RECT 248.580 36.355 249.070 36.360 ;
        RECT 241.520 34.555 242.010 34.560 ;
        RECT 241.520 33.240 242.010 33.245 ;
        RECT 238.160 31.295 239.770 32.905 ;
        RECT 241.520 32.760 243.865 33.240 ;
        RECT 245.765 32.905 246.285 34.895 ;
        RECT 250.445 34.560 250.925 36.360 ;
        RECT 252.280 34.895 253.890 36.505 ;
        RECT 241.520 32.755 242.010 32.760 ;
        RECT 238.705 29.305 239.225 31.295 ;
        RECT 243.385 30.960 243.865 32.760 ;
        RECT 245.220 31.295 246.830 32.905 ;
        RECT 248.580 31.440 249.070 31.445 ;
        RECT 250.445 31.440 250.925 33.240 ;
        RECT 252.825 32.905 253.345 34.895 ;
        RECT 238.160 27.695 239.770 29.305 ;
        RECT 238.705 25.705 239.225 27.695 ;
        RECT 241.520 27.300 242.010 27.305 ;
        RECT 243.385 27.300 243.865 29.640 ;
        RECT 245.765 29.305 246.285 31.295 ;
        RECT 248.580 30.960 250.925 31.440 ;
        RECT 252.280 31.295 253.890 32.905 ;
        RECT 248.580 30.955 249.070 30.960 ;
        RECT 245.220 27.695 246.830 29.305 ;
        RECT 241.520 26.820 243.865 27.300 ;
        RECT 241.520 26.815 242.010 26.820 ;
        RECT 238.160 24.095 239.770 25.705 ;
        RECT 238.705 22.105 239.225 24.095 ;
        RECT 241.520 23.700 242.010 23.705 ;
        RECT 243.385 23.700 243.865 26.040 ;
        RECT 245.765 25.705 246.285 27.695 ;
        RECT 248.580 27.300 249.070 27.305 ;
        RECT 250.445 27.300 250.925 29.640 ;
        RECT 252.825 29.305 253.345 31.295 ;
        RECT 252.280 27.695 253.890 29.305 ;
        RECT 248.580 26.820 250.925 27.300 ;
        RECT 248.580 26.815 249.070 26.820 ;
        RECT 245.220 24.095 246.830 25.705 ;
        RECT 241.520 23.220 243.865 23.700 ;
        RECT 241.520 23.215 242.010 23.220 ;
        RECT 238.160 20.495 239.770 22.105 ;
        RECT 238.705 18.505 239.225 20.495 ;
        RECT 243.385 20.160 243.865 23.220 ;
        RECT 245.765 22.105 246.285 24.095 ;
        RECT 248.580 23.700 249.070 23.705 ;
        RECT 250.445 23.700 250.925 26.040 ;
        RECT 252.825 25.705 253.345 27.695 ;
        RECT 252.280 24.095 253.890 25.705 ;
        RECT 248.580 23.220 250.925 23.700 ;
        RECT 248.580 23.215 249.070 23.220 ;
        RECT 245.220 20.495 246.830 22.105 ;
        RECT 238.160 16.895 239.770 18.505 ;
        RECT 238.705 14.905 239.225 16.895 ;
        RECT 238.160 13.295 239.770 14.905 ;
        RECT 238.705 11.305 239.225 13.295 ;
        RECT 241.520 12.900 242.010 12.905 ;
        RECT 243.385 12.900 243.865 18.840 ;
        RECT 245.765 18.505 246.285 20.495 ;
        RECT 250.445 20.160 250.925 23.220 ;
        RECT 252.825 22.105 253.345 24.095 ;
        RECT 252.280 20.495 253.890 22.105 ;
        RECT 245.220 16.895 246.830 18.505 ;
        RECT 245.765 14.905 246.285 16.895 ;
        RECT 245.220 13.295 246.830 14.905 ;
        RECT 241.520 12.420 243.865 12.900 ;
        RECT 241.520 12.415 242.010 12.420 ;
        RECT 238.160 9.695 239.770 11.305 ;
        RECT 238.705 7.705 239.225 9.695 ;
        RECT 238.160 6.095 239.770 7.705 ;
        RECT 238.705 4.580 239.225 6.095 ;
        RECT 243.385 5.760 243.865 12.420 ;
        RECT 245.765 11.305 246.285 13.295 ;
        RECT 248.580 12.900 249.070 12.905 ;
        RECT 250.445 12.900 250.925 18.840 ;
        RECT 252.825 18.505 253.345 20.495 ;
        RECT 252.280 16.895 253.890 18.505 ;
        RECT 252.825 14.905 253.345 16.895 ;
        RECT 252.280 13.295 253.890 14.905 ;
        RECT 248.580 12.420 250.925 12.900 ;
        RECT 248.580 12.415 249.070 12.420 ;
        RECT 245.220 9.695 246.830 11.305 ;
        RECT 245.765 7.705 246.285 9.695 ;
        RECT 245.220 6.095 246.830 7.705 ;
        RECT 245.765 4.580 246.285 6.095 ;
        RECT 250.445 5.760 250.925 12.420 ;
        RECT 252.825 11.305 253.345 13.295 ;
        RECT 252.280 9.695 253.890 11.305 ;
        RECT 252.825 7.705 253.345 9.695 ;
        RECT 252.280 6.095 253.890 7.705 ;
        RECT 252.825 4.580 253.345 6.095 ;
        RECT 255.485 5.100 256.005 67.215 ;
        RECT 260.540 66.175 261.070 66.705 ;
        RECT 260.545 63.740 261.065 66.175 ;
        RECT 270.660 65.135 271.190 65.665 ;
        RECT 270.665 63.740 271.185 65.135 ;
        RECT 290.900 64.095 291.430 64.625 ;
        RECT 290.905 63.740 291.425 64.095 ;
        RECT 260.545 63.220 266.125 63.740 ;
        RECT 257.885 61.705 258.405 62.700 ;
        RECT 257.340 60.095 258.950 61.705 ;
        RECT 257.885 58.105 258.405 60.095 ;
        RECT 257.340 56.495 258.950 58.105 ;
        RECT 257.885 54.505 258.405 56.495 ;
        RECT 257.340 52.895 258.950 54.505 ;
        RECT 257.885 50.905 258.405 52.895 ;
        RECT 257.340 49.295 258.950 50.905 ;
        RECT 257.885 47.305 258.405 49.295 ;
        RECT 257.340 45.695 258.950 47.305 ;
        RECT 257.885 43.705 258.405 45.695 ;
        RECT 257.340 42.095 258.950 43.705 ;
        RECT 257.885 40.105 258.405 42.095 ;
        RECT 257.340 38.495 258.950 40.105 ;
        RECT 257.885 36.505 258.405 38.495 ;
        RECT 257.340 34.895 258.950 36.505 ;
        RECT 257.885 32.905 258.405 34.895 ;
        RECT 257.340 31.295 258.950 32.905 ;
        RECT 257.885 29.305 258.405 31.295 ;
        RECT 257.340 27.695 258.950 29.305 ;
        RECT 257.885 25.705 258.405 27.695 ;
        RECT 257.340 24.095 258.950 25.705 ;
        RECT 257.885 22.105 258.405 24.095 ;
        RECT 257.340 20.495 258.950 22.105 ;
        RECT 257.885 18.505 258.405 20.495 ;
        RECT 257.340 16.895 258.950 18.505 ;
        RECT 257.885 14.905 258.405 16.895 ;
        RECT 257.340 13.295 258.950 14.905 ;
        RECT 257.885 11.305 258.405 13.295 ;
        RECT 257.340 9.695 258.950 11.305 ;
        RECT 257.885 7.705 258.405 9.695 ;
        RECT 257.340 6.095 258.950 7.705 ;
        RECT 257.885 4.580 258.405 6.095 ;
        RECT 260.545 5.100 261.065 63.220 ;
        RECT 262.945 61.705 263.465 62.700 ;
        RECT 262.400 60.095 264.010 61.705 ;
        RECT 262.945 58.105 263.465 60.095 ;
        RECT 262.400 56.495 264.010 58.105 ;
        RECT 262.945 54.505 263.465 56.495 ;
        RECT 262.400 52.895 264.010 54.505 ;
        RECT 262.945 50.905 263.465 52.895 ;
        RECT 262.400 49.295 264.010 50.905 ;
        RECT 262.945 47.305 263.465 49.295 ;
        RECT 262.400 45.695 264.010 47.305 ;
        RECT 262.945 43.705 263.465 45.695 ;
        RECT 262.400 42.095 264.010 43.705 ;
        RECT 262.945 40.105 263.465 42.095 ;
        RECT 262.400 38.495 264.010 40.105 ;
        RECT 262.945 36.505 263.465 38.495 ;
        RECT 262.400 34.895 264.010 36.505 ;
        RECT 262.945 32.905 263.465 34.895 ;
        RECT 262.400 31.295 264.010 32.905 ;
        RECT 262.945 29.305 263.465 31.295 ;
        RECT 262.400 27.695 264.010 29.305 ;
        RECT 262.945 25.705 263.465 27.695 ;
        RECT 262.400 24.095 264.010 25.705 ;
        RECT 262.945 22.105 263.465 24.095 ;
        RECT 262.400 20.495 264.010 22.105 ;
        RECT 262.945 18.505 263.465 20.495 ;
        RECT 262.400 16.895 264.010 18.505 ;
        RECT 262.945 14.905 263.465 16.895 ;
        RECT 262.400 13.295 264.010 14.905 ;
        RECT 262.945 11.305 263.465 13.295 ;
        RECT 262.400 9.695 264.010 11.305 ;
        RECT 262.945 7.705 263.465 9.695 ;
        RECT 262.400 6.095 264.010 7.705 ;
        RECT 262.945 4.580 263.465 6.095 ;
        RECT 265.605 5.100 266.125 63.220 ;
        RECT 270.665 63.220 286.365 63.740 ;
        RECT 268.005 61.705 268.525 62.700 ;
        RECT 267.460 60.095 269.070 61.705 ;
        RECT 268.005 58.105 268.525 60.095 ;
        RECT 267.460 56.495 269.070 58.105 ;
        RECT 268.005 54.505 268.525 56.495 ;
        RECT 267.460 52.895 269.070 54.505 ;
        RECT 268.005 50.905 268.525 52.895 ;
        RECT 267.460 49.295 269.070 50.905 ;
        RECT 268.005 47.305 268.525 49.295 ;
        RECT 267.460 45.695 269.070 47.305 ;
        RECT 268.005 43.705 268.525 45.695 ;
        RECT 267.460 42.095 269.070 43.705 ;
        RECT 268.005 40.105 268.525 42.095 ;
        RECT 267.460 38.495 269.070 40.105 ;
        RECT 268.005 36.505 268.525 38.495 ;
        RECT 267.460 34.895 269.070 36.505 ;
        RECT 268.005 32.905 268.525 34.895 ;
        RECT 267.460 31.295 269.070 32.905 ;
        RECT 268.005 29.305 268.525 31.295 ;
        RECT 267.460 27.695 269.070 29.305 ;
        RECT 268.005 25.705 268.525 27.695 ;
        RECT 267.460 24.095 269.070 25.705 ;
        RECT 268.005 22.105 268.525 24.095 ;
        RECT 267.460 20.495 269.070 22.105 ;
        RECT 268.005 18.505 268.525 20.495 ;
        RECT 267.460 16.895 269.070 18.505 ;
        RECT 268.005 14.905 268.525 16.895 ;
        RECT 267.460 13.295 269.070 14.905 ;
        RECT 268.005 11.305 268.525 13.295 ;
        RECT 267.460 9.695 269.070 11.305 ;
        RECT 268.005 7.705 268.525 9.695 ;
        RECT 267.460 6.095 269.070 7.705 ;
        RECT 268.005 4.580 268.525 6.095 ;
        RECT 270.665 5.100 271.185 63.220 ;
        RECT 273.065 61.705 273.585 62.700 ;
        RECT 272.520 60.095 274.130 61.705 ;
        RECT 273.065 58.105 273.585 60.095 ;
        RECT 272.520 56.495 274.130 58.105 ;
        RECT 273.065 54.505 273.585 56.495 ;
        RECT 272.520 52.895 274.130 54.505 ;
        RECT 273.065 50.905 273.585 52.895 ;
        RECT 272.520 49.295 274.130 50.905 ;
        RECT 273.065 47.305 273.585 49.295 ;
        RECT 272.520 45.695 274.130 47.305 ;
        RECT 273.065 43.705 273.585 45.695 ;
        RECT 272.520 42.095 274.130 43.705 ;
        RECT 273.065 40.105 273.585 42.095 ;
        RECT 272.520 38.495 274.130 40.105 ;
        RECT 273.065 36.505 273.585 38.495 ;
        RECT 272.520 34.895 274.130 36.505 ;
        RECT 273.065 32.905 273.585 34.895 ;
        RECT 272.520 31.295 274.130 32.905 ;
        RECT 273.065 29.305 273.585 31.295 ;
        RECT 272.520 27.695 274.130 29.305 ;
        RECT 273.065 25.705 273.585 27.695 ;
        RECT 272.520 24.095 274.130 25.705 ;
        RECT 273.065 22.105 273.585 24.095 ;
        RECT 272.520 20.495 274.130 22.105 ;
        RECT 273.065 18.505 273.585 20.495 ;
        RECT 272.520 16.895 274.130 18.505 ;
        RECT 273.065 14.905 273.585 16.895 ;
        RECT 272.520 13.295 274.130 14.905 ;
        RECT 273.065 11.305 273.585 13.295 ;
        RECT 272.520 9.695 274.130 11.305 ;
        RECT 273.065 7.705 273.585 9.695 ;
        RECT 272.520 6.095 274.130 7.705 ;
        RECT 273.065 4.580 273.585 6.095 ;
        RECT 275.725 5.100 276.245 63.220 ;
        RECT 278.125 61.705 278.645 62.700 ;
        RECT 277.580 60.095 279.190 61.705 ;
        RECT 278.125 58.105 278.645 60.095 ;
        RECT 277.580 56.495 279.190 58.105 ;
        RECT 278.125 54.505 278.645 56.495 ;
        RECT 277.580 52.895 279.190 54.505 ;
        RECT 278.125 50.905 278.645 52.895 ;
        RECT 277.580 49.295 279.190 50.905 ;
        RECT 278.125 47.305 278.645 49.295 ;
        RECT 277.580 45.695 279.190 47.305 ;
        RECT 278.125 43.705 278.645 45.695 ;
        RECT 277.580 42.095 279.190 43.705 ;
        RECT 278.125 40.105 278.645 42.095 ;
        RECT 277.580 38.495 279.190 40.105 ;
        RECT 278.125 36.505 278.645 38.495 ;
        RECT 277.580 34.895 279.190 36.505 ;
        RECT 278.125 32.905 278.645 34.895 ;
        RECT 277.580 31.295 279.190 32.905 ;
        RECT 278.125 29.305 278.645 31.295 ;
        RECT 277.580 27.695 279.190 29.305 ;
        RECT 278.125 25.705 278.645 27.695 ;
        RECT 277.580 24.095 279.190 25.705 ;
        RECT 278.125 22.105 278.645 24.095 ;
        RECT 277.580 20.495 279.190 22.105 ;
        RECT 278.125 18.505 278.645 20.495 ;
        RECT 277.580 16.895 279.190 18.505 ;
        RECT 278.125 14.905 278.645 16.895 ;
        RECT 277.580 13.295 279.190 14.905 ;
        RECT 278.125 11.305 278.645 13.295 ;
        RECT 277.580 9.695 279.190 11.305 ;
        RECT 278.125 7.705 278.645 9.695 ;
        RECT 277.580 6.095 279.190 7.705 ;
        RECT 278.125 4.580 278.645 6.095 ;
        RECT 280.785 5.100 281.305 63.220 ;
        RECT 283.185 61.705 283.705 62.700 ;
        RECT 282.640 60.095 284.250 61.705 ;
        RECT 283.185 58.105 283.705 60.095 ;
        RECT 282.640 56.495 284.250 58.105 ;
        RECT 283.185 54.505 283.705 56.495 ;
        RECT 282.640 52.895 284.250 54.505 ;
        RECT 283.185 50.905 283.705 52.895 ;
        RECT 282.640 49.295 284.250 50.905 ;
        RECT 283.185 47.305 283.705 49.295 ;
        RECT 282.640 45.695 284.250 47.305 ;
        RECT 283.185 43.705 283.705 45.695 ;
        RECT 282.640 42.095 284.250 43.705 ;
        RECT 283.185 40.105 283.705 42.095 ;
        RECT 282.640 38.495 284.250 40.105 ;
        RECT 283.185 36.505 283.705 38.495 ;
        RECT 282.640 34.895 284.250 36.505 ;
        RECT 283.185 32.905 283.705 34.895 ;
        RECT 282.640 31.295 284.250 32.905 ;
        RECT 283.185 29.305 283.705 31.295 ;
        RECT 282.640 27.695 284.250 29.305 ;
        RECT 283.185 25.705 283.705 27.695 ;
        RECT 282.640 24.095 284.250 25.705 ;
        RECT 283.185 22.105 283.705 24.095 ;
        RECT 282.640 20.495 284.250 22.105 ;
        RECT 283.185 18.505 283.705 20.495 ;
        RECT 282.640 16.895 284.250 18.505 ;
        RECT 283.185 14.905 283.705 16.895 ;
        RECT 282.640 13.295 284.250 14.905 ;
        RECT 283.185 11.305 283.705 13.295 ;
        RECT 282.640 9.695 284.250 11.305 ;
        RECT 283.185 7.705 283.705 9.695 ;
        RECT 282.640 6.095 284.250 7.705 ;
        RECT 283.185 4.580 283.705 6.095 ;
        RECT 285.845 5.100 286.365 63.220 ;
        RECT 290.905 63.220 326.845 63.740 ;
        RECT 288.245 61.705 288.765 62.700 ;
        RECT 287.700 60.095 289.310 61.705 ;
        RECT 288.245 58.105 288.765 60.095 ;
        RECT 287.700 56.495 289.310 58.105 ;
        RECT 288.245 54.505 288.765 56.495 ;
        RECT 287.700 52.895 289.310 54.505 ;
        RECT 288.245 50.905 288.765 52.895 ;
        RECT 287.700 49.295 289.310 50.905 ;
        RECT 288.245 47.305 288.765 49.295 ;
        RECT 287.700 45.695 289.310 47.305 ;
        RECT 288.245 43.705 288.765 45.695 ;
        RECT 287.700 42.095 289.310 43.705 ;
        RECT 288.245 40.105 288.765 42.095 ;
        RECT 287.700 38.495 289.310 40.105 ;
        RECT 288.245 36.505 288.765 38.495 ;
        RECT 287.700 34.895 289.310 36.505 ;
        RECT 288.245 32.905 288.765 34.895 ;
        RECT 287.700 31.295 289.310 32.905 ;
        RECT 288.245 29.305 288.765 31.295 ;
        RECT 287.700 27.695 289.310 29.305 ;
        RECT 288.245 25.705 288.765 27.695 ;
        RECT 287.700 24.095 289.310 25.705 ;
        RECT 288.245 22.105 288.765 24.095 ;
        RECT 287.700 20.495 289.310 22.105 ;
        RECT 288.245 18.505 288.765 20.495 ;
        RECT 287.700 16.895 289.310 18.505 ;
        RECT 288.245 14.905 288.765 16.895 ;
        RECT 287.700 13.295 289.310 14.905 ;
        RECT 288.245 11.305 288.765 13.295 ;
        RECT 287.700 9.695 289.310 11.305 ;
        RECT 288.245 7.705 288.765 9.695 ;
        RECT 287.700 6.095 289.310 7.705 ;
        RECT 288.245 4.580 288.765 6.095 ;
        RECT 290.905 5.100 291.425 63.220 ;
        RECT 293.305 61.705 293.825 62.700 ;
        RECT 292.760 60.095 294.370 61.705 ;
        RECT 293.305 58.105 293.825 60.095 ;
        RECT 292.760 56.495 294.370 58.105 ;
        RECT 293.305 54.505 293.825 56.495 ;
        RECT 292.760 52.895 294.370 54.505 ;
        RECT 293.305 50.905 293.825 52.895 ;
        RECT 292.760 49.295 294.370 50.905 ;
        RECT 293.305 47.305 293.825 49.295 ;
        RECT 292.760 45.695 294.370 47.305 ;
        RECT 293.305 43.705 293.825 45.695 ;
        RECT 292.760 42.095 294.370 43.705 ;
        RECT 293.305 40.105 293.825 42.095 ;
        RECT 292.760 38.495 294.370 40.105 ;
        RECT 293.305 36.505 293.825 38.495 ;
        RECT 292.760 34.895 294.370 36.505 ;
        RECT 293.305 32.905 293.825 34.895 ;
        RECT 292.760 31.295 294.370 32.905 ;
        RECT 293.305 29.305 293.825 31.295 ;
        RECT 292.760 27.695 294.370 29.305 ;
        RECT 293.305 25.705 293.825 27.695 ;
        RECT 292.760 24.095 294.370 25.705 ;
        RECT 293.305 22.105 293.825 24.095 ;
        RECT 292.760 20.495 294.370 22.105 ;
        RECT 293.305 18.505 293.825 20.495 ;
        RECT 292.760 16.895 294.370 18.505 ;
        RECT 293.305 14.905 293.825 16.895 ;
        RECT 292.760 13.295 294.370 14.905 ;
        RECT 293.305 11.305 293.825 13.295 ;
        RECT 292.760 9.695 294.370 11.305 ;
        RECT 293.305 7.705 293.825 9.695 ;
        RECT 292.760 6.095 294.370 7.705 ;
        RECT 293.305 4.580 293.825 6.095 ;
        RECT 295.965 5.100 296.485 63.220 ;
        RECT 298.365 61.705 298.885 62.700 ;
        RECT 297.820 60.095 299.430 61.705 ;
        RECT 298.365 58.105 298.885 60.095 ;
        RECT 297.820 56.495 299.430 58.105 ;
        RECT 298.365 54.505 298.885 56.495 ;
        RECT 297.820 52.895 299.430 54.505 ;
        RECT 298.365 50.905 298.885 52.895 ;
        RECT 297.820 49.295 299.430 50.905 ;
        RECT 298.365 47.305 298.885 49.295 ;
        RECT 297.820 45.695 299.430 47.305 ;
        RECT 298.365 43.705 298.885 45.695 ;
        RECT 297.820 42.095 299.430 43.705 ;
        RECT 298.365 40.105 298.885 42.095 ;
        RECT 297.820 38.495 299.430 40.105 ;
        RECT 298.365 36.505 298.885 38.495 ;
        RECT 297.820 34.895 299.430 36.505 ;
        RECT 298.365 32.905 298.885 34.895 ;
        RECT 297.820 31.295 299.430 32.905 ;
        RECT 298.365 29.305 298.885 31.295 ;
        RECT 297.820 27.695 299.430 29.305 ;
        RECT 298.365 25.705 298.885 27.695 ;
        RECT 297.820 24.095 299.430 25.705 ;
        RECT 298.365 22.105 298.885 24.095 ;
        RECT 297.820 20.495 299.430 22.105 ;
        RECT 298.365 18.505 298.885 20.495 ;
        RECT 297.820 16.895 299.430 18.505 ;
        RECT 298.365 14.905 298.885 16.895 ;
        RECT 297.820 13.295 299.430 14.905 ;
        RECT 298.365 11.305 298.885 13.295 ;
        RECT 297.820 9.695 299.430 11.305 ;
        RECT 298.365 7.705 298.885 9.695 ;
        RECT 297.820 6.095 299.430 7.705 ;
        RECT 298.365 4.580 298.885 6.095 ;
        RECT 301.025 5.100 301.545 63.220 ;
        RECT 303.425 61.705 303.945 62.700 ;
        RECT 302.880 60.095 304.490 61.705 ;
        RECT 303.425 58.105 303.945 60.095 ;
        RECT 302.880 56.495 304.490 58.105 ;
        RECT 303.425 54.505 303.945 56.495 ;
        RECT 302.880 52.895 304.490 54.505 ;
        RECT 303.425 50.905 303.945 52.895 ;
        RECT 302.880 49.295 304.490 50.905 ;
        RECT 303.425 47.305 303.945 49.295 ;
        RECT 302.880 45.695 304.490 47.305 ;
        RECT 303.425 43.705 303.945 45.695 ;
        RECT 302.880 42.095 304.490 43.705 ;
        RECT 303.425 40.105 303.945 42.095 ;
        RECT 302.880 38.495 304.490 40.105 ;
        RECT 303.425 36.505 303.945 38.495 ;
        RECT 302.880 34.895 304.490 36.505 ;
        RECT 303.425 32.905 303.945 34.895 ;
        RECT 302.880 31.295 304.490 32.905 ;
        RECT 303.425 29.305 303.945 31.295 ;
        RECT 302.880 27.695 304.490 29.305 ;
        RECT 303.425 25.705 303.945 27.695 ;
        RECT 302.880 24.095 304.490 25.705 ;
        RECT 303.425 22.105 303.945 24.095 ;
        RECT 302.880 20.495 304.490 22.105 ;
        RECT 303.425 18.505 303.945 20.495 ;
        RECT 302.880 16.895 304.490 18.505 ;
        RECT 303.425 14.905 303.945 16.895 ;
        RECT 302.880 13.295 304.490 14.905 ;
        RECT 303.425 11.305 303.945 13.295 ;
        RECT 302.880 9.695 304.490 11.305 ;
        RECT 303.425 7.705 303.945 9.695 ;
        RECT 302.880 6.095 304.490 7.705 ;
        RECT 303.425 4.580 303.945 6.095 ;
        RECT 306.085 5.100 306.605 63.220 ;
        RECT 308.485 61.705 309.005 62.700 ;
        RECT 307.940 60.095 309.550 61.705 ;
        RECT 308.485 58.105 309.005 60.095 ;
        RECT 307.940 56.495 309.550 58.105 ;
        RECT 308.485 54.505 309.005 56.495 ;
        RECT 307.940 52.895 309.550 54.505 ;
        RECT 308.485 50.905 309.005 52.895 ;
        RECT 307.940 49.295 309.550 50.905 ;
        RECT 308.485 47.305 309.005 49.295 ;
        RECT 307.940 45.695 309.550 47.305 ;
        RECT 308.485 43.705 309.005 45.695 ;
        RECT 307.940 42.095 309.550 43.705 ;
        RECT 308.485 40.105 309.005 42.095 ;
        RECT 307.940 38.495 309.550 40.105 ;
        RECT 308.485 36.505 309.005 38.495 ;
        RECT 307.940 34.895 309.550 36.505 ;
        RECT 308.485 32.905 309.005 34.895 ;
        RECT 307.940 31.295 309.550 32.905 ;
        RECT 308.485 29.305 309.005 31.295 ;
        RECT 307.940 27.695 309.550 29.305 ;
        RECT 308.485 25.705 309.005 27.695 ;
        RECT 307.940 24.095 309.550 25.705 ;
        RECT 308.485 22.105 309.005 24.095 ;
        RECT 307.940 20.495 309.550 22.105 ;
        RECT 308.485 18.505 309.005 20.495 ;
        RECT 307.940 16.895 309.550 18.505 ;
        RECT 308.485 14.905 309.005 16.895 ;
        RECT 307.940 13.295 309.550 14.905 ;
        RECT 308.485 11.305 309.005 13.295 ;
        RECT 307.940 9.695 309.550 11.305 ;
        RECT 308.485 7.705 309.005 9.695 ;
        RECT 307.940 6.095 309.550 7.705 ;
        RECT 308.485 4.580 309.005 6.095 ;
        RECT 311.145 5.100 311.665 63.220 ;
        RECT 313.545 61.705 314.065 62.700 ;
        RECT 313.000 60.095 314.610 61.705 ;
        RECT 313.545 58.105 314.065 60.095 ;
        RECT 313.000 56.495 314.610 58.105 ;
        RECT 313.545 54.505 314.065 56.495 ;
        RECT 313.000 52.895 314.610 54.505 ;
        RECT 313.545 50.905 314.065 52.895 ;
        RECT 313.000 49.295 314.610 50.905 ;
        RECT 313.545 47.305 314.065 49.295 ;
        RECT 313.000 45.695 314.610 47.305 ;
        RECT 313.545 43.705 314.065 45.695 ;
        RECT 313.000 42.095 314.610 43.705 ;
        RECT 313.545 40.105 314.065 42.095 ;
        RECT 313.000 38.495 314.610 40.105 ;
        RECT 313.545 36.505 314.065 38.495 ;
        RECT 313.000 34.895 314.610 36.505 ;
        RECT 313.545 32.905 314.065 34.895 ;
        RECT 313.000 31.295 314.610 32.905 ;
        RECT 313.545 29.305 314.065 31.295 ;
        RECT 313.000 27.695 314.610 29.305 ;
        RECT 313.545 25.705 314.065 27.695 ;
        RECT 313.000 24.095 314.610 25.705 ;
        RECT 313.545 22.105 314.065 24.095 ;
        RECT 313.000 20.495 314.610 22.105 ;
        RECT 313.545 18.505 314.065 20.495 ;
        RECT 313.000 16.895 314.610 18.505 ;
        RECT 313.545 14.905 314.065 16.895 ;
        RECT 313.000 13.295 314.610 14.905 ;
        RECT 313.545 11.305 314.065 13.295 ;
        RECT 313.000 9.695 314.610 11.305 ;
        RECT 313.545 7.705 314.065 9.695 ;
        RECT 313.000 6.095 314.610 7.705 ;
        RECT 313.545 4.580 314.065 6.095 ;
        RECT 316.205 5.100 316.725 63.220 ;
        RECT 318.605 61.705 319.125 62.700 ;
        RECT 318.060 60.095 319.670 61.705 ;
        RECT 318.605 58.105 319.125 60.095 ;
        RECT 318.060 56.495 319.670 58.105 ;
        RECT 318.605 54.505 319.125 56.495 ;
        RECT 318.060 52.895 319.670 54.505 ;
        RECT 318.605 50.905 319.125 52.895 ;
        RECT 318.060 49.295 319.670 50.905 ;
        RECT 318.605 47.305 319.125 49.295 ;
        RECT 318.060 45.695 319.670 47.305 ;
        RECT 318.605 43.705 319.125 45.695 ;
        RECT 318.060 42.095 319.670 43.705 ;
        RECT 318.605 40.105 319.125 42.095 ;
        RECT 318.060 38.495 319.670 40.105 ;
        RECT 318.605 36.505 319.125 38.495 ;
        RECT 318.060 34.895 319.670 36.505 ;
        RECT 318.605 32.905 319.125 34.895 ;
        RECT 318.060 31.295 319.670 32.905 ;
        RECT 318.605 29.305 319.125 31.295 ;
        RECT 318.060 27.695 319.670 29.305 ;
        RECT 318.605 25.705 319.125 27.695 ;
        RECT 318.060 24.095 319.670 25.705 ;
        RECT 318.605 22.105 319.125 24.095 ;
        RECT 318.060 20.495 319.670 22.105 ;
        RECT 318.605 18.505 319.125 20.495 ;
        RECT 318.060 16.895 319.670 18.505 ;
        RECT 318.605 14.905 319.125 16.895 ;
        RECT 318.060 13.295 319.670 14.905 ;
        RECT 318.605 11.305 319.125 13.295 ;
        RECT 318.060 9.695 319.670 11.305 ;
        RECT 318.605 7.705 319.125 9.695 ;
        RECT 318.060 6.095 319.670 7.705 ;
        RECT 318.605 4.580 319.125 6.095 ;
        RECT 321.265 5.100 321.785 63.220 ;
        RECT 323.665 61.705 324.185 62.700 ;
        RECT 323.120 60.095 324.730 61.705 ;
        RECT 323.665 58.105 324.185 60.095 ;
        RECT 323.120 56.495 324.730 58.105 ;
        RECT 323.665 54.505 324.185 56.495 ;
        RECT 323.120 52.895 324.730 54.505 ;
        RECT 323.665 50.905 324.185 52.895 ;
        RECT 323.120 49.295 324.730 50.905 ;
        RECT 323.665 47.305 324.185 49.295 ;
        RECT 323.120 45.695 324.730 47.305 ;
        RECT 323.665 43.705 324.185 45.695 ;
        RECT 323.120 42.095 324.730 43.705 ;
        RECT 323.665 40.105 324.185 42.095 ;
        RECT 323.120 38.495 324.730 40.105 ;
        RECT 323.665 36.505 324.185 38.495 ;
        RECT 323.120 34.895 324.730 36.505 ;
        RECT 323.665 32.905 324.185 34.895 ;
        RECT 323.120 31.295 324.730 32.905 ;
        RECT 323.665 29.305 324.185 31.295 ;
        RECT 323.120 27.695 324.730 29.305 ;
        RECT 323.665 25.705 324.185 27.695 ;
        RECT 323.120 24.095 324.730 25.705 ;
        RECT 323.665 22.105 324.185 24.095 ;
        RECT 323.120 20.495 324.730 22.105 ;
        RECT 323.665 18.505 324.185 20.495 ;
        RECT 323.120 16.895 324.730 18.505 ;
        RECT 323.665 14.905 324.185 16.895 ;
        RECT 323.120 13.295 324.730 14.905 ;
        RECT 323.665 11.305 324.185 13.295 ;
        RECT 323.120 9.695 324.730 11.305 ;
        RECT 323.665 7.705 324.185 9.695 ;
        RECT 323.120 6.095 324.730 7.705 ;
        RECT 323.665 4.580 324.185 6.095 ;
        RECT 326.325 5.100 326.845 63.220 ;
        RECT 328.725 61.705 329.245 62.700 ;
        RECT 328.180 60.095 329.790 61.705 ;
        RECT 328.725 58.105 329.245 60.095 ;
        RECT 328.180 56.495 329.790 58.105 ;
        RECT 328.725 54.505 329.245 56.495 ;
        RECT 328.180 52.895 329.790 54.505 ;
        RECT 328.725 50.905 329.245 52.895 ;
        RECT 328.180 49.295 329.790 50.905 ;
        RECT 328.725 47.305 329.245 49.295 ;
        RECT 328.180 45.695 329.790 47.305 ;
        RECT 328.725 43.705 329.245 45.695 ;
        RECT 328.180 42.095 329.790 43.705 ;
        RECT 328.725 40.105 329.245 42.095 ;
        RECT 328.180 38.495 329.790 40.105 ;
        RECT 328.725 36.505 329.245 38.495 ;
        RECT 328.180 34.895 329.790 36.505 ;
        RECT 328.725 32.905 329.245 34.895 ;
        RECT 328.180 31.295 329.790 32.905 ;
        RECT 328.725 29.305 329.245 31.295 ;
        RECT 328.180 27.695 329.790 29.305 ;
        RECT 328.725 25.705 329.245 27.695 ;
        RECT 328.180 24.095 329.790 25.705 ;
        RECT 328.725 22.105 329.245 24.095 ;
        RECT 328.180 20.495 329.790 22.105 ;
        RECT 328.725 18.505 329.245 20.495 ;
        RECT 328.180 16.895 329.790 18.505 ;
        RECT 328.725 14.905 329.245 16.895 ;
        RECT 328.180 13.295 329.790 14.905 ;
        RECT 328.725 11.305 329.245 13.295 ;
        RECT 328.180 9.695 329.790 11.305 ;
        RECT 328.725 7.705 329.245 9.695 ;
        RECT 328.180 6.095 329.790 7.705 ;
        RECT 328.725 4.580 329.245 6.095 ;
        RECT 165.215 4.060 330.185 4.580 ;
        RECT 167.210 4.055 167.740 4.060 ;
        RECT 317.525 3.910 318.045 4.060 ;
        RECT 134.575 -5.170 135.065 -5.165 ;
        RECT 134.575 -5.650 136.440 -5.170 ;
        RECT 134.575 -5.655 135.065 -5.650 ;
  END
END tt_um_tsar_adc
END LIBRARY

