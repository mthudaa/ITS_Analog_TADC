magic
tech sky130A
magscale 1 2
timestamp 1757834164
<< dnwell >>
rect 12318 3709 14718 6109
rect 16941 3702 19353 6114
<< nwell >>
rect 12238 5903 14798 6189
rect 12238 3915 12524 5903
rect 14512 3915 14798 5903
rect 12238 3629 14798 3915
rect 16861 5908 19433 6194
rect 16861 3908 17147 5908
rect 19147 3908 19433 5908
rect 16861 3622 19433 3908
<< nsubdiff >>
rect 12275 6132 14761 6152
rect 12275 6098 12355 6132
rect 14681 6098 14761 6132
rect 12275 6078 14761 6098
rect 12275 6072 12349 6078
rect 12275 3746 12295 6072
rect 12329 3746 12349 6072
rect 12275 3740 12349 3746
rect 14687 6072 14761 6078
rect 14687 3746 14707 6072
rect 14741 3746 14761 6072
rect 14687 3740 14761 3746
rect 12275 3720 14761 3740
rect 12275 3686 12355 3720
rect 14681 3686 14761 3720
rect 12275 3666 14761 3686
rect 16898 6137 19396 6157
rect 16898 6103 16978 6137
rect 19316 6103 19396 6137
rect 16898 6083 19396 6103
rect 16898 6077 16972 6083
rect 16898 3739 16918 6077
rect 16952 3739 16972 6077
rect 16898 3733 16972 3739
rect 19322 6077 19396 6083
rect 19322 3739 19342 6077
rect 19376 3739 19396 6077
rect 19322 3733 19396 3739
rect 16898 3713 19396 3733
rect 16898 3679 16978 3713
rect 19316 3679 19396 3713
rect 16898 3659 19396 3679
<< nsubdiffcont >>
rect 12355 6098 14681 6132
rect 12295 3746 12329 6072
rect 14707 3746 14741 6072
rect 12355 3686 14681 3720
rect 16978 6103 19316 6137
rect 16918 3739 16952 6077
rect 19342 3739 19376 6077
rect 16978 3679 19316 3713
<< locali >>
rect 12295 6098 12355 6132
rect 14681 6098 14741 6132
rect 12295 6072 12329 6098
rect 12295 3720 12329 3746
rect 14707 6072 14741 6098
rect 14707 3720 14741 3746
rect 12295 3686 12355 3720
rect 14681 3686 14741 3720
rect 16918 6103 16978 6137
rect 19316 6103 19376 6137
rect 16918 6077 16952 6103
rect 16918 3713 16952 3739
rect 19342 6077 19376 6103
rect 19342 3713 19376 3739
rect 16918 3679 16978 3713
rect 19316 3679 19376 3713
<< viali >>
rect 8835 -8 8869 26
rect 10702 21 10736 55
rect 20924 2 20958 36
rect 22791 -8 22825 26
<< metal1 >>
rect 11328 6352 20483 6374
rect 11328 6300 15804 6352
rect 15856 6300 20483 6352
rect 11328 6278 20483 6300
rect 11318 338 11434 360
rect 11318 286 11350 338
rect 11402 286 11434 338
rect 11318 264 11434 286
rect 12158 264 14974 520
rect 16686 264 19502 520
rect 20226 338 20342 360
rect 20226 286 20258 338
rect 20310 286 20342 338
rect 20226 264 20342 286
rect 20754 116 20764 168
rect 20816 116 20826 168
rect 10685 55 11048 64
rect 8823 26 8881 32
rect 3079 -8 8835 26
rect 8869 -8 8881 26
rect 10685 21 10702 55
rect 10736 21 11048 55
rect 10685 12 11048 21
rect 11100 12 11110 64
rect 20754 -7 20764 45
rect 20816 36 20975 45
rect 20816 2 20924 36
rect 20958 2 20975 36
rect 20816 -7 20975 2
rect 22779 26 22837 32
rect 8823 -14 8881 -8
rect 22779 -8 22791 26
rect 22825 -8 28581 26
rect 22779 -14 22837 -8
rect 10838 -328 10956 -305
rect 10838 -380 10871 -328
rect 10923 -380 10956 -328
rect 10838 -403 10956 -380
rect 20704 -328 20822 -305
rect 20704 -380 20737 -328
rect 20789 -380 20822 -328
rect 20704 -403 20822 -380
<< via1 >>
rect 15804 6300 15856 6352
rect 11350 286 11402 338
rect 20258 286 20310 338
rect 20764 116 20816 168
rect 11048 12 11100 64
rect 20764 -7 20816 45
rect 10871 -380 10923 -328
rect 20737 -380 20789 -328
<< metal2 >>
rect 15782 6354 15878 6384
rect 15782 6298 15802 6354
rect 15858 6298 15878 6354
rect 15782 6268 15878 6298
rect 11328 340 11424 370
rect 11328 284 11348 340
rect 11404 284 11424 340
rect 11328 254 11424 284
rect 20236 340 20332 370
rect 20236 284 20256 340
rect 20312 284 20332 340
rect 20236 254 20332 284
rect 20764 168 20816 178
rect 20340 116 20764 168
rect 11048 64 11100 74
rect 11100 12 11353 64
rect 20764 45 20816 116
rect 11048 2 11100 12
rect 20764 -17 20816 -7
rect 10848 -326 10946 -295
rect 10848 -382 10869 -326
rect 10925 -382 10946 -326
rect 10848 -413 10946 -382
rect 20714 -326 20812 -295
rect 20714 -382 20735 -326
rect 20791 -382 20812 -326
rect 20714 -413 20812 -382
<< via2 >>
rect 15802 6352 15858 6354
rect 15802 6300 15804 6352
rect 15804 6300 15856 6352
rect 15856 6300 15858 6352
rect 15802 6298 15858 6300
rect 11348 338 11404 340
rect 11348 286 11350 338
rect 11350 286 11402 338
rect 11402 286 11404 338
rect 11348 284 11404 286
rect 20256 338 20312 340
rect 20256 286 20258 338
rect 20258 286 20310 338
rect 20310 286 20312 338
rect 20256 284 20312 286
rect 10869 -328 10925 -326
rect 10869 -380 10871 -328
rect 10871 -380 10923 -328
rect 10923 -380 10925 -328
rect 10869 -382 10925 -380
rect 20735 -328 20791 -326
rect 20735 -380 20737 -328
rect 20737 -380 20789 -328
rect 20789 -380 20791 -328
rect 20735 -382 20791 -380
<< metal3 >>
rect 13172 6114 14984 6380
rect 15772 6354 15888 6379
rect 15772 6298 15802 6354
rect 15858 6298 15888 6354
rect 15772 6273 15888 6298
rect 15782 744 15878 6273
rect 16686 6119 18478 6375
rect 15772 728 15888 744
rect 15772 664 15798 728
rect 15862 664 15888 728
rect 15772 648 15888 664
rect 11318 360 11434 365
rect 20226 360 20342 365
rect 11318 340 20342 360
rect 11318 284 11348 340
rect 11404 284 20256 340
rect 20312 284 20342 340
rect 11318 264 20342 284
rect 11318 259 11434 264
rect 20226 259 20342 264
rect 10838 -305 10956 -300
rect 20704 -305 20822 -300
rect 10838 -323 20822 -305
rect 10838 -326 15798 -323
rect 10838 -382 10869 -326
rect 10925 -382 15798 -326
rect 10838 -387 15798 -382
rect 15862 -326 20822 -323
rect 15862 -382 20735 -326
rect 20791 -382 20822 -326
rect 15862 -387 20822 -382
rect 10838 -403 20822 -387
rect 10838 -408 10956 -403
rect 20704 -408 20822 -403
<< via3 >>
rect 15798 664 15862 728
rect 15798 -387 15862 -323
<< metal4 >>
rect 15781 728 15879 745
rect 15781 664 15798 728
rect 15862 664 15879 728
rect 15781 647 15879 664
rect 15782 -306 15878 647
rect 15781 -323 15879 -306
rect 15781 -387 15798 -323
rect 15862 -387 15879 -323
rect 15781 -404 15879 -387
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_0
timestamp 1750100919
transform -1 0 10848 0 -1 312
box -38 -49 2150 715
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_1
timestamp 1750100919
transform 1 0 20812 0 -1 312
box -38 -49 2150 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1750100919
transform -1 0 8736 0 -1 312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1750100919
transform -1 0 23020 0 -1 312
box -38 -49 134 715
use th_sw  th_sw_0
timestamp 1757834164
transform 1 0 369 0 1 132
box 2710 -132 15509 6253
use th_sw  th_sw_1
timestamp 1757834164
transform -1 0 31291 0 1 132
box 2710 -132 15509 6253
<< labels >>
flabel metal3 s 15706 294 15740 328 0 FreeSans 500 0 0 0 VSS
port 3 nsew
flabel metal1 s 13533 411 13567 445 0 FreeSans 500 0 0 0 VCN
port 4 nsew
flabel metal1 s 18092 413 18126 447 0 FreeSans 500 0 0 0 VCP
port 5 nsew
flabel metal3 s 15782 6278 15878 6374 0 FreeSans 1000 0 0 0 VDD
port 6 nsew
flabel metal3 s 14013 6246 14043 6276 0 FreeSans 1000 0 0 0 VIN
port 7 nsew
flabel metal3 s 17579 6243 17609 6273 0 FreeSans 1000 0 0 0 VIP
port 8 nsew
flabel metal1 28547 -8 28581 26 0 FreeSans 320 0 0 0 CK
port 11 nsew
flabel metal1 3087 -8 3121 26 0 FreeSans 320 0 0 0 CKB
port 13 nsew
<< end >>
