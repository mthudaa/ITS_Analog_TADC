magic
tech sky130A
magscale 1 2
timestamp 1757893939
<< locali >>
rect -351 -3654 -291 -3641
rect -351 -3688 -338 -3654
rect -304 -3688 -291 -3654
rect -351 -3701 -291 -3688
rect -171 -3653 -111 -3640
rect -171 -3687 -158 -3653
rect -124 -3687 -111 -3653
rect -171 -3700 -111 -3687
rect 23 -3670 63 -3667
rect 23 -3704 26 -3670
rect 60 -3704 63 -3670
rect 23 -3707 63 -3704
rect 151 -3707 379 -3667
rect 536 -3717 657 -3677
rect 882 -3681 942 -3668
rect 882 -3715 895 -3681
rect 929 -3715 942 -3681
rect 882 -3728 942 -3715
rect 1009 -3716 1326 -3676
rect 2415 -3677 2475 -3664
rect 1976 -3717 2190 -3677
rect 2415 -3711 2428 -3677
rect 2462 -3711 2475 -3677
rect 2415 -3724 2475 -3711
rect 2824 -3681 2864 -3678
rect 2824 -3715 2827 -3681
rect 2861 -3715 2864 -3681
rect 2824 -3718 2864 -3715
rect -251 -3857 -211 -3854
rect -251 -3891 -248 -3857
rect -214 -3891 -211 -3857
rect -251 -3894 -211 -3891
rect -251 -4229 -211 -4226
rect -251 -4263 -248 -4229
rect -214 -4263 -211 -4229
rect -251 -4266 -211 -4263
rect -631 -4415 -571 -4402
rect -631 -4449 -618 -4415
rect -584 -4449 -571 -4415
rect 13 -4416 73 -4403
rect -631 -4462 -571 -4449
rect -435 -4469 -301 -4429
rect -171 -4431 -111 -4418
rect -171 -4465 -158 -4431
rect -124 -4465 -111 -4431
rect 13 -4450 26 -4416
rect 60 -4450 73 -4416
rect 13 -4463 73 -4450
rect 126 -4453 379 -4413
rect 532 -4443 628 -4403
rect 678 -4406 738 -4393
rect 678 -4440 691 -4406
rect 725 -4440 738 -4406
rect 678 -4453 738 -4440
rect 1009 -4443 1326 -4403
rect 1972 -4443 2190 -4403
rect 2415 -4409 2475 -4396
rect 2415 -4443 2428 -4409
rect 2462 -4443 2475 -4409
rect 2824 -4405 2864 -4402
rect 2824 -4439 2827 -4405
rect 2861 -4439 2864 -4405
rect 2824 -4442 2864 -4439
rect 2415 -4456 2475 -4443
rect -171 -4478 -111 -4465
<< viali >>
rect -338 -3688 -304 -3654
rect -158 -3687 -124 -3653
rect 26 -3704 60 -3670
rect 895 -3715 929 -3681
rect 2428 -3711 2462 -3677
rect 2827 -3715 2861 -3681
rect -248 -3891 -214 -3857
rect -248 -4263 -214 -4229
rect -618 -4449 -584 -4415
rect -158 -4465 -124 -4431
rect 26 -4450 60 -4416
rect 691 -4440 725 -4406
rect 2428 -4443 2462 -4409
rect 2827 -4439 2861 -4405
<< metal1 >>
rect 1060 -3367 1140 -3363
rect 1060 -3419 1074 -3367
rect 1126 -3419 1140 -3367
rect 1060 -3423 1140 -3419
rect -181 -3511 748 -3507
rect -181 -3563 -167 -3511
rect -115 -3563 682 -3511
rect 734 -3563 748 -3511
rect -181 -3567 748 -3563
rect 2578 -3511 2678 -3497
rect 2578 -3563 2602 -3511
rect 2654 -3517 2678 -3511
rect 2654 -3563 2927 -3517
rect 2578 -3577 2927 -3563
rect -363 -3641 -279 -3635
rect -641 -3645 -279 -3641
rect -641 -3697 -627 -3645
rect -575 -3654 -279 -3645
rect -575 -3688 -338 -3654
rect -304 -3688 -279 -3654
rect -575 -3697 -279 -3688
rect -641 -3701 -279 -3697
rect -363 -3707 -279 -3701
rect -183 -3644 -99 -3634
rect -183 -3696 -167 -3644
rect -115 -3696 -99 -3644
rect -183 -3706 -99 -3696
rect 3 -3661 83 -3657
rect 3 -3713 17 -3661
rect 69 -3713 83 -3661
rect 3 -3717 83 -3713
rect 870 -3672 954 -3662
rect 870 -3724 886 -3672
rect 938 -3724 954 -3672
rect 870 -3734 954 -3724
rect 2403 -3668 2487 -3658
rect 2403 -3720 2419 -3668
rect 2471 -3720 2487 -3668
rect 2403 -3730 2487 -3720
rect 2812 -3681 2927 -3668
rect 2812 -3715 2827 -3681
rect 2861 -3715 2927 -3681
rect 2812 -3728 2927 -3715
rect -263 -3848 83 -3844
rect -263 -3857 17 -3848
rect -263 -3891 -248 -3857
rect -214 -3891 17 -3857
rect -263 -3900 17 -3891
rect 69 -3900 83 -3848
rect -263 -3904 83 -3900
rect 2405 -3848 2927 -3844
rect 2405 -3900 2419 -3848
rect 2471 -3900 2927 -3848
rect 2405 -3904 2927 -3900
rect 2791 -4100 2873 -4026
rect -263 -4220 83 -4216
rect -263 -4229 17 -4220
rect -263 -4263 -248 -4229
rect -214 -4263 17 -4229
rect -263 -4272 17 -4263
rect 69 -4272 83 -4220
rect -263 -4276 83 -4272
rect -643 -4406 -559 -4396
rect 666 -4397 750 -4387
rect -643 -4458 -627 -4406
rect -575 -4458 -559 -4406
rect 1 -4407 85 -4397
rect -643 -4468 -559 -4458
rect -183 -4422 -99 -4412
rect -183 -4474 -167 -4422
rect -115 -4474 -99 -4422
rect 1 -4459 17 -4407
rect 69 -4459 85 -4407
rect 666 -4449 682 -4397
rect 734 -4449 750 -4397
rect 666 -4459 750 -4449
rect 2403 -4400 2487 -4390
rect 2403 -4452 2419 -4400
rect 2471 -4452 2487 -4400
rect 2812 -4405 2927 -4392
rect 2812 -4439 2827 -4405
rect 2861 -4439 2927 -4405
rect 2812 -4452 2927 -4439
rect 1 -4469 85 -4459
rect 2403 -4462 2487 -4452
rect -183 -4484 -99 -4474
rect 2405 -4551 2927 -4547
rect 2405 -4603 2419 -4551
rect 2471 -4603 2927 -4551
rect 2405 -4607 2927 -4603
rect 1060 -4700 1140 -4696
rect 1060 -4752 1074 -4700
rect 1126 -4752 1140 -4700
rect 1060 -4756 1140 -4752
rect 2783 -4764 2865 -4690
<< via1 >>
rect 1074 -3419 1126 -3367
rect -167 -3563 -115 -3511
rect 682 -3563 734 -3511
rect 2602 -3563 2654 -3511
rect -627 -3697 -575 -3645
rect -167 -3653 -115 -3644
rect -167 -3687 -158 -3653
rect -158 -3687 -124 -3653
rect -124 -3687 -115 -3653
rect -167 -3696 -115 -3687
rect 17 -3670 69 -3661
rect 17 -3704 26 -3670
rect 26 -3704 60 -3670
rect 60 -3704 69 -3670
rect 17 -3713 69 -3704
rect 886 -3681 938 -3672
rect 886 -3715 895 -3681
rect 895 -3715 929 -3681
rect 929 -3715 938 -3681
rect 886 -3724 938 -3715
rect 2419 -3677 2471 -3668
rect 2419 -3711 2428 -3677
rect 2428 -3711 2462 -3677
rect 2462 -3711 2471 -3677
rect 2419 -3720 2471 -3711
rect 17 -3900 69 -3848
rect 2419 -3900 2471 -3848
rect 17 -4272 69 -4220
rect -627 -4415 -575 -4406
rect -627 -4449 -618 -4415
rect -618 -4449 -584 -4415
rect -584 -4449 -575 -4415
rect -627 -4458 -575 -4449
rect -167 -4431 -115 -4422
rect -167 -4465 -158 -4431
rect -158 -4465 -124 -4431
rect -124 -4465 -115 -4431
rect -167 -4474 -115 -4465
rect 17 -4416 69 -4407
rect 17 -4450 26 -4416
rect 26 -4450 60 -4416
rect 60 -4450 69 -4416
rect 17 -4459 69 -4450
rect 682 -4406 734 -4397
rect 682 -4440 691 -4406
rect 691 -4440 725 -4406
rect 725 -4440 734 -4406
rect 682 -4449 734 -4440
rect 2419 -4409 2471 -4400
rect 2419 -4443 2428 -4409
rect 2428 -4443 2462 -4409
rect 2462 -4443 2471 -4409
rect 2419 -4452 2471 -4443
rect 2419 -4603 2471 -4551
rect 1074 -4752 1126 -4700
<< metal2 >>
rect 1070 -3367 1130 -3353
rect 1070 -3419 1074 -3367
rect 1126 -3419 1130 -3367
rect -631 -3509 -571 -3497
rect -631 -3565 -629 -3509
rect -573 -3565 -571 -3509
rect -631 -3645 -571 -3565
rect -631 -3697 -627 -3645
rect -575 -3697 -571 -3645
rect -631 -4406 -571 -3697
rect -171 -3511 -111 -3497
rect -171 -3563 -167 -3511
rect -115 -3563 -111 -3511
rect -171 -3644 -111 -3563
rect -171 -3696 -167 -3644
rect -115 -3696 -111 -3644
rect 678 -3511 738 -3497
rect 678 -3563 682 -3511
rect 734 -3563 738 -3511
rect -171 -3710 -111 -3696
rect 13 -3661 73 -3647
rect 13 -3713 17 -3661
rect 69 -3713 73 -3661
rect 13 -3848 73 -3713
rect 13 -3900 17 -3848
rect 69 -3900 73 -3848
rect 13 -3914 73 -3900
rect -631 -4458 -627 -4406
rect -575 -4458 -571 -4406
rect 13 -4220 73 -4206
rect 13 -4272 17 -4220
rect 69 -4272 73 -4220
rect 13 -4407 73 -4272
rect -631 -4472 -571 -4458
rect -171 -4422 -111 -4408
rect -171 -4474 -167 -4422
rect -115 -4474 -111 -4422
rect 13 -4459 17 -4407
rect 69 -4459 73 -4407
rect 13 -4473 73 -4459
rect 678 -4397 738 -3563
rect 678 -4449 682 -4397
rect 734 -4449 738 -4397
rect 678 -4463 738 -4449
rect 882 -3672 942 -3658
rect 882 -3724 886 -3672
rect 938 -3724 942 -3672
rect -171 -4551 -111 -4474
rect 882 -4551 942 -3724
rect -171 -4611 942 -4551
rect 1070 -4700 1130 -3419
rect 2588 -3509 2668 -3487
rect 2588 -3565 2600 -3509
rect 2656 -3565 2668 -3509
rect 2588 -3587 2668 -3565
rect 2415 -3668 2475 -3654
rect 2415 -3720 2419 -3668
rect 2471 -3720 2475 -3668
rect 2415 -3848 2475 -3720
rect 2415 -3900 2419 -3848
rect 2471 -3900 2475 -3848
rect 2415 -3914 2475 -3900
rect 2415 -4400 2475 -4386
rect 2415 -4452 2419 -4400
rect 2471 -4452 2475 -4400
rect 2415 -4551 2475 -4452
rect 2415 -4603 2419 -4551
rect 2471 -4603 2475 -4551
rect 2415 -4617 2475 -4603
rect 1070 -4752 1074 -4700
rect 1126 -4752 1130 -4700
rect 1070 -4766 1130 -4752
<< via2 >>
rect -629 -3565 -573 -3509
rect 2600 -3511 2656 -3509
rect 2600 -3563 2602 -3511
rect 2602 -3563 2654 -3511
rect 2654 -3563 2656 -3511
rect 2600 -3565 2656 -3563
<< metal3 >>
rect 2578 -3497 2678 -3492
rect -641 -3509 2678 -3497
rect -641 -3565 -629 -3509
rect -573 -3565 2600 -3509
rect 2656 -3565 2678 -3509
rect -641 -3577 2678 -3565
rect 2578 -3582 2678 -3577
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_0
timestamp 1750100919
transform 1 0 -87 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_1
timestamp 1750100919
transform 1 0 297 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0
timestamp 1750100919
transform 1 0 585 0 -1 -3394
box -38 -49 518 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_0
timestamp 1750100919
transform 1 0 1161 0 -1 -3394
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_1
timestamp 1750100919
transform 1 0 2025 0 -1 -3394
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 -87 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 201 0 1 -4726
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1723858470
transform 1 0 1065 0 1 -4726
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1723858470
transform 1 0 201 0 -1 -3394
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1723858470
transform 1 0 1065 0 -1 -3394
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  x1
timestamp 1723858470
transform 1 0 -375 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x3
timestamp 1750100919
transform 1 0 -663 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x4
timestamp 1750100919
transform 1 0 -87 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x6
timestamp 1750100919
transform 1 0 297 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  x8
timestamp 1750100919
transform 1 0 585 0 1 -4726
box -38 -49 518 715
use sky130_fd_sc_hs__inv_8  x10
timestamp 1750100919
transform 1 0 1161 0 1 -4726
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  x12
timestamp 1750100919
transform 1 0 2025 0 1 -4726
box -38 -49 902 715
<< labels >>
flabel metal1 s 2878 -3567 2918 -3527 0 FreeSans 500 0 0 0 IN
port 1 nsew
flabel metal1 s 2878 -3717 2918 -3677 0 FreeSans 500 0 0 0 CLK0
port 2 nsew
flabel metal1 s 2876 -3894 2916 -3854 0 FreeSans 500 0 0 0 CLKB0
port 3 nsew
flabel metal1 s 2876 -4443 2916 -4403 0 FreeSans 500 0 0 0 CLK1
port 4 nsew
flabel metal1 s 2877 -4597 2917 -4557 0 FreeSans 500 0 0 0 CLKB1
port 5 nsew
flabel metal1 s 2820 -4082 2860 -4042 0 FreeSans 500 0 0 0 VDD
port 6 nsew
flabel metal1 s 2807 -4748 2847 -4708 0 FreeSans 500 0 0 0 VSS
port 7 nsew
<< end >>
