magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -246 -1011 246 1011
<< pmos >>
rect -50 492 50 792
rect -50 64 50 364
rect -50 -364 50 -64
rect -50 -792 50 -492
<< pdiff >>
rect -108 761 -50 792
rect -108 727 -96 761
rect -62 727 -50 761
rect -108 693 -50 727
rect -108 659 -96 693
rect -62 659 -50 693
rect -108 625 -50 659
rect -108 591 -96 625
rect -62 591 -50 625
rect -108 557 -50 591
rect -108 523 -96 557
rect -62 523 -50 557
rect -108 492 -50 523
rect 50 761 108 792
rect 50 727 62 761
rect 96 727 108 761
rect 50 693 108 727
rect 50 659 62 693
rect 96 659 108 693
rect 50 625 108 659
rect 50 591 62 625
rect 96 591 108 625
rect 50 557 108 591
rect 50 523 62 557
rect 96 523 108 557
rect 50 492 108 523
rect -108 333 -50 364
rect -108 299 -96 333
rect -62 299 -50 333
rect -108 265 -50 299
rect -108 231 -96 265
rect -62 231 -50 265
rect -108 197 -50 231
rect -108 163 -96 197
rect -62 163 -50 197
rect -108 129 -50 163
rect -108 95 -96 129
rect -62 95 -50 129
rect -108 64 -50 95
rect 50 333 108 364
rect 50 299 62 333
rect 96 299 108 333
rect 50 265 108 299
rect 50 231 62 265
rect 96 231 108 265
rect 50 197 108 231
rect 50 163 62 197
rect 96 163 108 197
rect 50 129 108 163
rect 50 95 62 129
rect 96 95 108 129
rect 50 64 108 95
rect -108 -95 -50 -64
rect -108 -129 -96 -95
rect -62 -129 -50 -95
rect -108 -163 -50 -129
rect -108 -197 -96 -163
rect -62 -197 -50 -163
rect -108 -231 -50 -197
rect -108 -265 -96 -231
rect -62 -265 -50 -231
rect -108 -299 -50 -265
rect -108 -333 -96 -299
rect -62 -333 -50 -299
rect -108 -364 -50 -333
rect 50 -95 108 -64
rect 50 -129 62 -95
rect 96 -129 108 -95
rect 50 -163 108 -129
rect 50 -197 62 -163
rect 96 -197 108 -163
rect 50 -231 108 -197
rect 50 -265 62 -231
rect 96 -265 108 -231
rect 50 -299 108 -265
rect 50 -333 62 -299
rect 96 -333 108 -299
rect 50 -364 108 -333
rect -108 -523 -50 -492
rect -108 -557 -96 -523
rect -62 -557 -50 -523
rect -108 -591 -50 -557
rect -108 -625 -96 -591
rect -62 -625 -50 -591
rect -108 -659 -50 -625
rect -108 -693 -96 -659
rect -62 -693 -50 -659
rect -108 -727 -50 -693
rect -108 -761 -96 -727
rect -62 -761 -50 -727
rect -108 -792 -50 -761
rect 50 -523 108 -492
rect 50 -557 62 -523
rect 96 -557 108 -523
rect 50 -591 108 -557
rect 50 -625 62 -591
rect 96 -625 108 -591
rect 50 -659 108 -625
rect 50 -693 62 -659
rect 96 -693 108 -659
rect 50 -727 108 -693
rect 50 -761 62 -727
rect 96 -761 108 -727
rect 50 -792 108 -761
<< pdiffc >>
rect -96 727 -62 761
rect -96 659 -62 693
rect -96 591 -62 625
rect -96 523 -62 557
rect 62 727 96 761
rect 62 659 96 693
rect 62 591 96 625
rect 62 523 96 557
rect -96 299 -62 333
rect -96 231 -62 265
rect -96 163 -62 197
rect -96 95 -62 129
rect 62 299 96 333
rect 62 231 96 265
rect 62 163 96 197
rect 62 95 96 129
rect -96 -129 -62 -95
rect -96 -197 -62 -163
rect -96 -265 -62 -231
rect -96 -333 -62 -299
rect 62 -129 96 -95
rect 62 -197 96 -163
rect 62 -265 96 -231
rect 62 -333 96 -299
rect -96 -557 -62 -523
rect -96 -625 -62 -591
rect -96 -693 -62 -659
rect -96 -761 -62 -727
rect 62 -557 96 -523
rect 62 -625 96 -591
rect 62 -693 96 -659
rect 62 -761 96 -727
<< nsubdiff >>
rect -210 941 -85 975
rect -51 941 -17 975
rect 17 941 51 975
rect 85 941 210 975
rect -210 867 -176 941
rect -210 799 -176 833
rect 176 867 210 941
rect 176 799 210 833
rect -210 731 -176 765
rect -210 663 -176 697
rect -210 595 -176 629
rect -210 527 -176 561
rect -210 459 -176 493
rect 176 731 210 765
rect 176 663 210 697
rect 176 595 210 629
rect 176 527 210 561
rect -210 391 -176 425
rect 176 459 210 493
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect -210 -493 -176 -459
rect 176 -425 210 -391
rect -210 -561 -176 -527
rect -210 -629 -176 -595
rect -210 -697 -176 -663
rect -210 -765 -176 -731
rect 176 -493 210 -459
rect 176 -561 210 -527
rect 176 -629 210 -595
rect 176 -697 210 -663
rect 176 -765 210 -731
rect -210 -833 -176 -799
rect -210 -941 -176 -867
rect 176 -833 210 -799
rect 176 -941 210 -867
rect -210 -975 -85 -941
rect -51 -975 -17 -941
rect 17 -975 51 -941
rect 85 -975 210 -941
<< nsubdiffcont >>
rect -85 941 -51 975
rect -17 941 17 975
rect 51 941 85 975
rect -210 833 -176 867
rect -210 765 -176 799
rect 176 833 210 867
rect -210 697 -176 731
rect -210 629 -176 663
rect -210 561 -176 595
rect -210 493 -176 527
rect 176 765 210 799
rect 176 697 210 731
rect 176 629 210 663
rect 176 561 210 595
rect 176 493 210 527
rect -210 425 -176 459
rect -210 357 -176 391
rect 176 425 210 459
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect -210 -459 -176 -425
rect 176 -391 210 -357
rect 176 -459 210 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -210 -663 -176 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect 176 -527 210 -493
rect 176 -595 210 -561
rect 176 -663 210 -629
rect 176 -731 210 -697
rect -210 -867 -176 -833
rect 176 -799 210 -765
rect 176 -867 210 -833
rect -85 -975 -51 -941
rect -17 -975 17 -941
rect 51 -975 85 -941
<< poly >>
rect -50 873 50 889
rect -50 839 -17 873
rect 17 839 50 873
rect -50 792 50 839
rect -50 445 50 492
rect -50 411 -17 445
rect 17 411 50 445
rect -50 364 50 411
rect -50 17 50 64
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -64 50 -17
rect -50 -411 50 -364
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect -50 -492 50 -445
rect -50 -839 50 -792
rect -50 -873 -17 -839
rect 17 -873 50 -839
rect -50 -889 50 -873
<< polycont >>
rect -17 839 17 873
rect -17 411 17 445
rect -17 -17 17 17
rect -17 -445 17 -411
rect -17 -873 17 -839
<< locali >>
rect -210 941 -85 975
rect -51 941 -17 975
rect 17 941 51 975
rect 85 941 210 975
rect -210 867 -176 941
rect -50 839 -17 873
rect 17 839 50 873
rect 176 867 210 941
rect -210 799 -176 833
rect 176 799 210 833
rect -210 731 -176 765
rect -210 663 -176 697
rect -210 595 -176 629
rect -210 527 -176 561
rect -210 459 -176 493
rect -96 767 -62 796
rect -96 695 -62 727
rect -96 625 -62 659
rect -96 557 -62 589
rect -96 488 -62 517
rect 62 767 96 796
rect 62 695 96 727
rect 62 625 96 659
rect 62 557 96 589
rect 62 488 96 517
rect 176 731 210 765
rect 176 663 210 697
rect 176 595 210 629
rect 176 527 210 561
rect 176 459 210 493
rect -210 391 -176 425
rect -50 411 -17 445
rect 17 411 50 445
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -96 339 -62 368
rect -96 267 -62 299
rect -96 197 -62 231
rect -96 129 -62 161
rect -96 60 -62 89
rect 62 339 96 368
rect 62 267 96 299
rect 62 197 96 231
rect 62 129 96 161
rect 62 60 96 89
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect 176 51 210 85
rect -210 -17 -176 17
rect -50 -17 -17 17
rect 17 -17 50 17
rect 176 -17 210 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect -96 -89 -62 -60
rect -96 -161 -62 -129
rect -96 -231 -62 -197
rect -96 -299 -62 -267
rect -96 -368 -62 -339
rect 62 -89 96 -60
rect 62 -161 96 -129
rect 62 -231 96 -197
rect 62 -299 96 -267
rect 62 -368 96 -339
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect 176 -425 210 -391
rect -210 -493 -176 -459
rect -210 -561 -176 -527
rect -210 -629 -176 -595
rect -210 -697 -176 -663
rect -210 -765 -176 -731
rect -96 -517 -62 -488
rect -96 -589 -62 -557
rect -96 -659 -62 -625
rect -96 -727 -62 -695
rect -96 -796 -62 -767
rect 62 -517 96 -488
rect 62 -589 96 -557
rect 62 -659 96 -625
rect 62 -727 96 -695
rect 62 -796 96 -767
rect 176 -493 210 -459
rect 176 -561 210 -527
rect 176 -629 210 -595
rect 176 -697 210 -663
rect 176 -765 210 -731
rect -210 -833 -176 -799
rect 176 -833 210 -799
rect -210 -941 -176 -867
rect -50 -873 -17 -839
rect 17 -873 50 -839
rect 176 -941 210 -867
rect -210 -975 -85 -941
rect -51 -975 -17 -941
rect 17 -975 51 -941
rect 85 -975 210 -941
<< viali >>
rect -17 839 17 873
rect -96 761 -62 767
rect -96 733 -62 761
rect -96 693 -62 695
rect -96 661 -62 693
rect -96 591 -62 623
rect -96 589 -62 591
rect -96 523 -62 551
rect -96 517 -62 523
rect 62 761 96 767
rect 62 733 96 761
rect 62 693 96 695
rect 62 661 96 693
rect 62 591 96 623
rect 62 589 96 591
rect 62 523 96 551
rect 62 517 96 523
rect -17 411 17 445
rect -96 333 -62 339
rect -96 305 -62 333
rect -96 265 -62 267
rect -96 233 -62 265
rect -96 163 -62 195
rect -96 161 -62 163
rect -96 95 -62 123
rect -96 89 -62 95
rect 62 333 96 339
rect 62 305 96 333
rect 62 265 96 267
rect 62 233 96 265
rect 62 163 96 195
rect 62 161 96 163
rect 62 95 96 123
rect 62 89 96 95
rect -17 -17 17 17
rect -96 -95 -62 -89
rect -96 -123 -62 -95
rect -96 -163 -62 -161
rect -96 -195 -62 -163
rect -96 -265 -62 -233
rect -96 -267 -62 -265
rect -96 -333 -62 -305
rect -96 -339 -62 -333
rect 62 -95 96 -89
rect 62 -123 96 -95
rect 62 -163 96 -161
rect 62 -195 96 -163
rect 62 -265 96 -233
rect 62 -267 96 -265
rect 62 -333 96 -305
rect 62 -339 96 -333
rect -17 -445 17 -411
rect -96 -523 -62 -517
rect -96 -551 -62 -523
rect -96 -591 -62 -589
rect -96 -623 -62 -591
rect -96 -693 -62 -661
rect -96 -695 -62 -693
rect -96 -761 -62 -733
rect -96 -767 -62 -761
rect 62 -523 96 -517
rect 62 -551 96 -523
rect 62 -591 96 -589
rect 62 -623 96 -591
rect 62 -693 96 -661
rect 62 -695 96 -693
rect 62 -761 96 -733
rect 62 -767 96 -761
rect -17 -873 17 -839
<< metal1 >>
rect -46 873 46 879
rect -46 839 -17 873
rect 17 839 46 873
rect -46 833 46 839
rect -102 767 -56 792
rect -102 733 -96 767
rect -62 733 -56 767
rect -102 695 -56 733
rect -102 661 -96 695
rect -62 661 -56 695
rect -102 623 -56 661
rect -102 589 -96 623
rect -62 589 -56 623
rect -102 551 -56 589
rect -102 517 -96 551
rect -62 517 -56 551
rect -102 492 -56 517
rect 56 767 102 792
rect 56 733 62 767
rect 96 733 102 767
rect 56 695 102 733
rect 56 661 62 695
rect 96 661 102 695
rect 56 623 102 661
rect 56 589 62 623
rect 96 589 102 623
rect 56 551 102 589
rect 56 517 62 551
rect 96 517 102 551
rect 56 492 102 517
rect -46 445 46 451
rect -46 411 -17 445
rect 17 411 46 445
rect -46 405 46 411
rect -102 339 -56 364
rect -102 305 -96 339
rect -62 305 -56 339
rect -102 267 -56 305
rect -102 233 -96 267
rect -62 233 -56 267
rect -102 195 -56 233
rect -102 161 -96 195
rect -62 161 -56 195
rect -102 123 -56 161
rect -102 89 -96 123
rect -62 89 -56 123
rect -102 64 -56 89
rect 56 339 102 364
rect 56 305 62 339
rect 96 305 102 339
rect 56 267 102 305
rect 56 233 62 267
rect 96 233 102 267
rect 56 195 102 233
rect 56 161 62 195
rect 96 161 102 195
rect 56 123 102 161
rect 56 89 62 123
rect 96 89 102 123
rect 56 64 102 89
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -89 -56 -64
rect -102 -123 -96 -89
rect -62 -123 -56 -89
rect -102 -161 -56 -123
rect -102 -195 -96 -161
rect -62 -195 -56 -161
rect -102 -233 -56 -195
rect -102 -267 -96 -233
rect -62 -267 -56 -233
rect -102 -305 -56 -267
rect -102 -339 -96 -305
rect -62 -339 -56 -305
rect -102 -364 -56 -339
rect 56 -89 102 -64
rect 56 -123 62 -89
rect 96 -123 102 -89
rect 56 -161 102 -123
rect 56 -195 62 -161
rect 96 -195 102 -161
rect 56 -233 102 -195
rect 56 -267 62 -233
rect 96 -267 102 -233
rect 56 -305 102 -267
rect 56 -339 62 -305
rect 96 -339 102 -305
rect 56 -364 102 -339
rect -46 -411 46 -405
rect -46 -445 -17 -411
rect 17 -445 46 -411
rect -46 -451 46 -445
rect -102 -517 -56 -492
rect -102 -551 -96 -517
rect -62 -551 -56 -517
rect -102 -589 -56 -551
rect -102 -623 -96 -589
rect -62 -623 -56 -589
rect -102 -661 -56 -623
rect -102 -695 -96 -661
rect -62 -695 -56 -661
rect -102 -733 -56 -695
rect -102 -767 -96 -733
rect -62 -767 -56 -733
rect -102 -792 -56 -767
rect 56 -517 102 -492
rect 56 -551 62 -517
rect 96 -551 102 -517
rect 56 -589 102 -551
rect 56 -623 62 -589
rect 96 -623 102 -589
rect 56 -661 102 -623
rect 56 -695 62 -661
rect 96 -695 102 -661
rect 56 -733 102 -695
rect 56 -767 62 -733
rect 96 -767 102 -733
rect 56 -792 102 -767
rect -46 -839 46 -833
rect -46 -873 -17 -839
rect 17 -873 46 -839
rect -46 -879 46 -873
<< properties >>
string FIXED_BBOX -193 -958 193 958
<< end >>
