magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< error_p >>
rect -29 791 29 797
rect -29 757 -17 791
rect -29 751 29 757
<< pwell >>
rect -201 -919 201 919
<< nmos >>
rect -15 -781 15 719
<< ndiff >>
rect -73 700 -15 719
rect -73 666 -61 700
rect -27 666 -15 700
rect -73 632 -15 666
rect -73 598 -61 632
rect -27 598 -15 632
rect -73 564 -15 598
rect -73 530 -61 564
rect -27 530 -15 564
rect -73 496 -15 530
rect -73 462 -61 496
rect -27 462 -15 496
rect -73 428 -15 462
rect -73 394 -61 428
rect -27 394 -15 428
rect -73 360 -15 394
rect -73 326 -61 360
rect -27 326 -15 360
rect -73 292 -15 326
rect -73 258 -61 292
rect -27 258 -15 292
rect -73 224 -15 258
rect -73 190 -61 224
rect -27 190 -15 224
rect -73 156 -15 190
rect -73 122 -61 156
rect -27 122 -15 156
rect -73 88 -15 122
rect -73 54 -61 88
rect -27 54 -15 88
rect -73 20 -15 54
rect -73 -14 -61 20
rect -27 -14 -15 20
rect -73 -48 -15 -14
rect -73 -82 -61 -48
rect -27 -82 -15 -48
rect -73 -116 -15 -82
rect -73 -150 -61 -116
rect -27 -150 -15 -116
rect -73 -184 -15 -150
rect -73 -218 -61 -184
rect -27 -218 -15 -184
rect -73 -252 -15 -218
rect -73 -286 -61 -252
rect -27 -286 -15 -252
rect -73 -320 -15 -286
rect -73 -354 -61 -320
rect -27 -354 -15 -320
rect -73 -388 -15 -354
rect -73 -422 -61 -388
rect -27 -422 -15 -388
rect -73 -456 -15 -422
rect -73 -490 -61 -456
rect -27 -490 -15 -456
rect -73 -524 -15 -490
rect -73 -558 -61 -524
rect -27 -558 -15 -524
rect -73 -592 -15 -558
rect -73 -626 -61 -592
rect -27 -626 -15 -592
rect -73 -660 -15 -626
rect -73 -694 -61 -660
rect -27 -694 -15 -660
rect -73 -728 -15 -694
rect -73 -762 -61 -728
rect -27 -762 -15 -728
rect -73 -781 -15 -762
rect 15 700 73 719
rect 15 666 27 700
rect 61 666 73 700
rect 15 632 73 666
rect 15 598 27 632
rect 61 598 73 632
rect 15 564 73 598
rect 15 530 27 564
rect 61 530 73 564
rect 15 496 73 530
rect 15 462 27 496
rect 61 462 73 496
rect 15 428 73 462
rect 15 394 27 428
rect 61 394 73 428
rect 15 360 73 394
rect 15 326 27 360
rect 61 326 73 360
rect 15 292 73 326
rect 15 258 27 292
rect 61 258 73 292
rect 15 224 73 258
rect 15 190 27 224
rect 61 190 73 224
rect 15 156 73 190
rect 15 122 27 156
rect 61 122 73 156
rect 15 88 73 122
rect 15 54 27 88
rect 61 54 73 88
rect 15 20 73 54
rect 15 -14 27 20
rect 61 -14 73 20
rect 15 -48 73 -14
rect 15 -82 27 -48
rect 61 -82 73 -48
rect 15 -116 73 -82
rect 15 -150 27 -116
rect 61 -150 73 -116
rect 15 -184 73 -150
rect 15 -218 27 -184
rect 61 -218 73 -184
rect 15 -252 73 -218
rect 15 -286 27 -252
rect 61 -286 73 -252
rect 15 -320 73 -286
rect 15 -354 27 -320
rect 61 -354 73 -320
rect 15 -388 73 -354
rect 15 -422 27 -388
rect 61 -422 73 -388
rect 15 -456 73 -422
rect 15 -490 27 -456
rect 61 -490 73 -456
rect 15 -524 73 -490
rect 15 -558 27 -524
rect 61 -558 73 -524
rect 15 -592 73 -558
rect 15 -626 27 -592
rect 61 -626 73 -592
rect 15 -660 73 -626
rect 15 -694 27 -660
rect 61 -694 73 -660
rect 15 -728 73 -694
rect 15 -762 27 -728
rect 61 -762 73 -728
rect 15 -781 73 -762
<< ndiffc >>
rect -61 666 -27 700
rect -61 598 -27 632
rect -61 530 -27 564
rect -61 462 -27 496
rect -61 394 -27 428
rect -61 326 -27 360
rect -61 258 -27 292
rect -61 190 -27 224
rect -61 122 -27 156
rect -61 54 -27 88
rect -61 -14 -27 20
rect -61 -82 -27 -48
rect -61 -150 -27 -116
rect -61 -218 -27 -184
rect -61 -286 -27 -252
rect -61 -354 -27 -320
rect -61 -422 -27 -388
rect -61 -490 -27 -456
rect -61 -558 -27 -524
rect -61 -626 -27 -592
rect -61 -694 -27 -660
rect -61 -762 -27 -728
rect 27 666 61 700
rect 27 598 61 632
rect 27 530 61 564
rect 27 462 61 496
rect 27 394 61 428
rect 27 326 61 360
rect 27 258 61 292
rect 27 190 61 224
rect 27 122 61 156
rect 27 54 61 88
rect 27 -14 61 20
rect 27 -82 61 -48
rect 27 -150 61 -116
rect 27 -218 61 -184
rect 27 -286 61 -252
rect 27 -354 61 -320
rect 27 -422 61 -388
rect 27 -490 61 -456
rect 27 -558 61 -524
rect 27 -626 61 -592
rect 27 -694 61 -660
rect 27 -762 61 -728
<< psubdiff >>
rect -175 859 -51 893
rect -17 859 17 893
rect 51 859 175 893
rect -175 765 -141 859
rect 141 765 175 859
rect -175 697 -141 731
rect -175 629 -141 663
rect -175 561 -141 595
rect -175 493 -141 527
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -175 -527 -141 -493
rect -175 -595 -141 -561
rect -175 -663 -141 -629
rect -175 -731 -141 -697
rect -175 -859 -141 -765
rect 141 697 175 731
rect 141 629 175 663
rect 141 561 175 595
rect 141 493 175 527
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 141 -527 175 -493
rect 141 -595 175 -561
rect 141 -663 175 -629
rect 141 -731 175 -697
rect 141 -859 175 -765
rect -175 -893 -51 -859
rect -17 -893 17 -859
rect 51 -893 175 -859
<< psubdiffcont >>
rect -51 859 -17 893
rect 17 859 51 893
rect -175 731 -141 765
rect 141 731 175 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect 141 663 175 697
rect 141 595 175 629
rect 141 527 175 561
rect 141 459 175 493
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect 141 -493 175 -459
rect 141 -561 175 -527
rect 141 -629 175 -595
rect 141 -697 175 -663
rect 141 -765 175 -731
rect -51 -893 -17 -859
rect 17 -893 51 -859
<< poly >>
rect -33 791 33 807
rect -33 757 -17 791
rect 17 757 33 791
rect -33 741 33 757
rect -15 719 15 741
rect -15 -807 15 -781
<< polycont >>
rect -17 757 17 791
<< locali >>
rect -175 859 -51 893
rect -17 859 17 893
rect 51 859 175 893
rect -175 765 -141 859
rect -33 757 -17 791
rect 17 757 33 791
rect 141 765 175 859
rect -175 697 -141 731
rect -175 629 -141 663
rect -175 561 -141 595
rect -175 493 -141 527
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -175 -527 -141 -493
rect -175 -595 -141 -561
rect -175 -663 -141 -629
rect -175 -731 -141 -697
rect -175 -859 -141 -765
rect -61 706 -27 723
rect -61 634 -27 666
rect -61 564 -27 598
rect -61 496 -27 528
rect -61 428 -27 456
rect -61 360 -27 384
rect -61 292 -27 312
rect -61 224 -27 240
rect -61 156 -27 168
rect -61 88 -27 96
rect -61 20 -27 24
rect -61 -86 -27 -82
rect -61 -158 -27 -150
rect -61 -230 -27 -218
rect -61 -302 -27 -286
rect -61 -374 -27 -354
rect -61 -446 -27 -422
rect -61 -518 -27 -490
rect -61 -590 -27 -558
rect -61 -660 -27 -626
rect -61 -728 -27 -696
rect -61 -785 -27 -768
rect 27 706 61 723
rect 27 634 61 666
rect 27 564 61 598
rect 27 496 61 528
rect 27 428 61 456
rect 27 360 61 384
rect 27 292 61 312
rect 27 224 61 240
rect 27 156 61 168
rect 27 88 61 96
rect 27 20 61 24
rect 27 -86 61 -82
rect 27 -158 61 -150
rect 27 -230 61 -218
rect 27 -302 61 -286
rect 27 -374 61 -354
rect 27 -446 61 -422
rect 27 -518 61 -490
rect 27 -590 61 -558
rect 27 -660 61 -626
rect 27 -728 61 -696
rect 27 -785 61 -768
rect 141 697 175 731
rect 141 629 175 663
rect 141 561 175 595
rect 141 493 175 527
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 141 -527 175 -493
rect 141 -595 175 -561
rect 141 -663 175 -629
rect 141 -731 175 -697
rect 141 -859 175 -765
rect -175 -893 -51 -859
rect -17 -893 17 -859
rect 51 -893 175 -859
<< viali >>
rect -17 757 17 791
rect -61 700 -27 706
rect -61 672 -27 700
rect -61 632 -27 634
rect -61 600 -27 632
rect -61 530 -27 562
rect -61 528 -27 530
rect -61 462 -27 490
rect -61 456 -27 462
rect -61 394 -27 418
rect -61 384 -27 394
rect -61 326 -27 346
rect -61 312 -27 326
rect -61 258 -27 274
rect -61 240 -27 258
rect -61 190 -27 202
rect -61 168 -27 190
rect -61 122 -27 130
rect -61 96 -27 122
rect -61 54 -27 58
rect -61 24 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -86
rect -61 -120 -27 -116
rect -61 -184 -27 -158
rect -61 -192 -27 -184
rect -61 -252 -27 -230
rect -61 -264 -27 -252
rect -61 -320 -27 -302
rect -61 -336 -27 -320
rect -61 -388 -27 -374
rect -61 -408 -27 -388
rect -61 -456 -27 -446
rect -61 -480 -27 -456
rect -61 -524 -27 -518
rect -61 -552 -27 -524
rect -61 -592 -27 -590
rect -61 -624 -27 -592
rect -61 -694 -27 -662
rect -61 -696 -27 -694
rect -61 -762 -27 -734
rect -61 -768 -27 -762
rect 27 700 61 706
rect 27 672 61 700
rect 27 632 61 634
rect 27 600 61 632
rect 27 530 61 562
rect 27 528 61 530
rect 27 462 61 490
rect 27 456 61 462
rect 27 394 61 418
rect 27 384 61 394
rect 27 326 61 346
rect 27 312 61 326
rect 27 258 61 274
rect 27 240 61 258
rect 27 190 61 202
rect 27 168 61 190
rect 27 122 61 130
rect 27 96 61 122
rect 27 54 61 58
rect 27 24 61 54
rect 27 -48 61 -14
rect 27 -116 61 -86
rect 27 -120 61 -116
rect 27 -184 61 -158
rect 27 -192 61 -184
rect 27 -252 61 -230
rect 27 -264 61 -252
rect 27 -320 61 -302
rect 27 -336 61 -320
rect 27 -388 61 -374
rect 27 -408 61 -388
rect 27 -456 61 -446
rect 27 -480 61 -456
rect 27 -524 61 -518
rect 27 -552 61 -524
rect 27 -592 61 -590
rect 27 -624 61 -592
rect 27 -694 61 -662
rect 27 -696 61 -694
rect 27 -762 61 -734
rect 27 -768 61 -762
<< metal1 >>
rect -29 791 29 797
rect -29 757 -17 791
rect 17 757 29 791
rect -29 751 29 757
rect -67 706 -21 719
rect -67 672 -61 706
rect -27 672 -21 706
rect -67 634 -21 672
rect -67 600 -61 634
rect -27 600 -21 634
rect -67 562 -21 600
rect -67 528 -61 562
rect -27 528 -21 562
rect -67 490 -21 528
rect -67 456 -61 490
rect -27 456 -21 490
rect -67 418 -21 456
rect -67 384 -61 418
rect -27 384 -21 418
rect -67 346 -21 384
rect -67 312 -61 346
rect -27 312 -21 346
rect -67 274 -21 312
rect -67 240 -61 274
rect -27 240 -21 274
rect -67 202 -21 240
rect -67 168 -61 202
rect -27 168 -21 202
rect -67 130 -21 168
rect -67 96 -61 130
rect -27 96 -21 130
rect -67 58 -21 96
rect -67 24 -61 58
rect -27 24 -21 58
rect -67 -14 -21 24
rect -67 -48 -61 -14
rect -27 -48 -21 -14
rect -67 -86 -21 -48
rect -67 -120 -61 -86
rect -27 -120 -21 -86
rect -67 -158 -21 -120
rect -67 -192 -61 -158
rect -27 -192 -21 -158
rect -67 -230 -21 -192
rect -67 -264 -61 -230
rect -27 -264 -21 -230
rect -67 -302 -21 -264
rect -67 -336 -61 -302
rect -27 -336 -21 -302
rect -67 -374 -21 -336
rect -67 -408 -61 -374
rect -27 -408 -21 -374
rect -67 -446 -21 -408
rect -67 -480 -61 -446
rect -27 -480 -21 -446
rect -67 -518 -21 -480
rect -67 -552 -61 -518
rect -27 -552 -21 -518
rect -67 -590 -21 -552
rect -67 -624 -61 -590
rect -27 -624 -21 -590
rect -67 -662 -21 -624
rect -67 -696 -61 -662
rect -27 -696 -21 -662
rect -67 -734 -21 -696
rect -67 -768 -61 -734
rect -27 -768 -21 -734
rect -67 -781 -21 -768
rect 21 706 67 719
rect 21 672 27 706
rect 61 672 67 706
rect 21 634 67 672
rect 21 600 27 634
rect 61 600 67 634
rect 21 562 67 600
rect 21 528 27 562
rect 61 528 67 562
rect 21 490 67 528
rect 21 456 27 490
rect 61 456 67 490
rect 21 418 67 456
rect 21 384 27 418
rect 61 384 67 418
rect 21 346 67 384
rect 21 312 27 346
rect 61 312 67 346
rect 21 274 67 312
rect 21 240 27 274
rect 61 240 67 274
rect 21 202 67 240
rect 21 168 27 202
rect 61 168 67 202
rect 21 130 67 168
rect 21 96 27 130
rect 61 96 67 130
rect 21 58 67 96
rect 21 24 27 58
rect 61 24 67 58
rect 21 -14 67 24
rect 21 -48 27 -14
rect 61 -48 67 -14
rect 21 -86 67 -48
rect 21 -120 27 -86
rect 61 -120 67 -86
rect 21 -158 67 -120
rect 21 -192 27 -158
rect 61 -192 67 -158
rect 21 -230 67 -192
rect 21 -264 27 -230
rect 61 -264 67 -230
rect 21 -302 67 -264
rect 21 -336 27 -302
rect 61 -336 67 -302
rect 21 -374 67 -336
rect 21 -408 27 -374
rect 61 -408 67 -374
rect 21 -446 67 -408
rect 21 -480 27 -446
rect 61 -480 67 -446
rect 21 -518 67 -480
rect 21 -552 27 -518
rect 61 -552 67 -518
rect 21 -590 67 -552
rect 21 -624 27 -590
rect 61 -624 67 -590
rect 21 -662 67 -624
rect 21 -696 27 -662
rect 61 -696 67 -662
rect 21 -734 67 -696
rect 21 -768 27 -734
rect 61 -768 67 -734
rect 21 -781 67 -768
<< properties >>
string FIXED_BBOX -158 -876 158 876
<< end >>
