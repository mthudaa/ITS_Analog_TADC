magic
tech sky130A
magscale 1 2
timestamp 1757871483
<< metal1 >>
rect -32202 -960 -32192 -864
rect -32096 -960 -31492 -864
rect -31412 -960 -31180 -864
rect -31084 -960 -31074 -864
rect -32202 -3120 -32192 -3024
rect -32096 -3120 -31652 -3024
rect -31572 -3120 -31180 -3024
rect -31084 -3120 -31074 -3024
rect -32202 -3840 -32192 -3744
rect -32096 -3840 -31812 -3744
rect -31732 -3840 -31180 -3744
rect -31084 -3840 -31074 -3744
rect -32834 -4668 -32824 -4572
rect -32744 -4668 -32192 -4572
rect -32096 -4668 -32086 -4572
rect -32514 -5028 -32504 -4932
rect -32424 -5028 -31180 -4932
rect -31084 -5028 -31074 -4932
rect -32674 -5388 -32664 -5292
rect -32584 -5388 -31180 -5292
rect -31084 -5388 -31074 -5292
rect -32514 -5748 -32504 -5652
rect -32424 -5748 -32192 -5652
rect -32096 -5748 -32086 -5652
rect -32202 -6000 -32192 -5904
rect -32096 -6000 -31812 -5904
rect -31732 -6000 -31180 -5904
rect -31084 -6000 -31074 -5904
rect -32202 -7440 -32192 -7344
rect -32096 -7440 -31652 -7344
rect -31572 -7440 -31180 -7344
rect -31084 -7440 -31074 -7344
rect -32202 -9600 -32192 -9504
rect -32096 -9600 -31492 -9504
rect -31412 -9600 -31180 -9504
rect -31084 -9600 -31074 -9504
rect -48044 -11304 -40292 -11200
rect -40188 -11304 -23088 -11200
rect -22984 -11304 -15900 -11200
rect -48044 -11512 -36244 -11408
rect -36140 -11512 -27136 -11408
rect -27032 -11512 -15900 -11408
rect -48044 -11720 -34220 -11616
rect -34116 -11720 -29160 -11616
rect -29056 -11720 -15900 -11616
rect -48044 -11928 -33208 -11824
rect -33104 -11928 -30172 -11824
rect -30068 -11928 -15900 -11824
rect -48044 -12136 -31492 -12032
rect -31412 -12136 -15900 -12032
rect -48044 -12344 -31652 -12240
rect -31572 -12344 -15900 -12240
rect -48044 -12552 -31812 -12448
rect -31732 -12552 -15900 -12448
rect -48044 -12760 -32504 -12656
rect -32424 -12760 -15900 -12656
rect -48044 -12968 -32664 -12864
rect -32584 -12968 -15900 -12864
rect -48044 -13176 -32824 -13072
rect -32744 -13176 -15900 -13072
<< via1 >>
rect -32192 -960 -32096 -864
rect -31492 -960 -31412 -864
rect -31180 -960 -31084 -864
rect -32192 -3120 -32096 -3024
rect -31652 -3120 -31572 -3024
rect -31180 -3120 -31084 -3024
rect -32192 -3840 -32096 -3744
rect -31812 -3840 -31732 -3744
rect -31180 -3840 -31084 -3744
rect -32824 -4668 -32744 -4572
rect -32192 -4668 -32096 -4572
rect -32504 -5028 -32424 -4932
rect -31180 -5028 -31084 -4932
rect -32664 -5388 -32584 -5292
rect -31180 -5388 -31084 -5292
rect -32504 -5748 -32424 -5652
rect -32192 -5748 -32096 -5652
rect -32192 -6000 -32096 -5904
rect -31812 -6000 -31732 -5904
rect -31180 -6000 -31084 -5904
rect -32192 -7440 -32096 -7344
rect -31652 -7440 -31572 -7344
rect -31180 -7440 -31084 -7344
rect -32192 -9600 -32096 -9504
rect -31492 -9600 -31412 -9504
rect -31180 -9600 -31084 -9504
rect -40292 -11304 -40188 -11200
rect -23088 -11304 -22984 -11200
rect -36244 -11512 -36140 -11408
rect -27136 -11512 -27032 -11408
rect -34220 -11720 -34116 -11616
rect -29160 -11720 -29056 -11616
rect -33208 -11928 -33104 -11824
rect -30172 -11928 -30068 -11824
rect -31492 -12136 -31412 -12032
rect -31652 -12344 -31572 -12240
rect -31812 -12552 -31732 -12448
rect -32504 -12760 -32424 -12656
rect -32664 -12968 -32584 -12864
rect -32824 -13176 -32744 -13072
<< metal2 >>
rect -32192 -864 -32096 -854
rect -32192 -970 -32096 -960
rect -31492 -864 -31412 -858
rect -32192 -3024 -32096 -3014
rect -32192 -3130 -32096 -3120
rect -31652 -3024 -31572 -3018
rect -32192 -3744 -32096 -3734
rect -32192 -3850 -32096 -3840
rect -31812 -3744 -31732 -3738
rect -32824 -4572 -32744 -4566
rect -40292 -11200 -40188 -11190
rect -40292 -11314 -40188 -11304
rect -36244 -11408 -36140 -11398
rect -36244 -11522 -36140 -11512
rect -34220 -11616 -34116 -11606
rect -34220 -11730 -34116 -11720
rect -33208 -11824 -33104 -11814
rect -33208 -11938 -33104 -11928
rect -32824 -13072 -32744 -4668
rect -32192 -4572 -32096 -4562
rect -32192 -4678 -32096 -4668
rect -32504 -4932 -32424 -4926
rect -32664 -5292 -32584 -5286
rect -32664 -12864 -32584 -5388
rect -32504 -5652 -32424 -5028
rect -32504 -12656 -32424 -5748
rect -32192 -5652 -32096 -5642
rect -32192 -5758 -32096 -5748
rect -32192 -5904 -32096 -5894
rect -32192 -6010 -32096 -6000
rect -31812 -5904 -31732 -3840
rect -32192 -7344 -32096 -7334
rect -32192 -7450 -32096 -7440
rect -32192 -9504 -32096 -9494
rect -32192 -9610 -32096 -9600
rect -31812 -12448 -31732 -6000
rect -31652 -7344 -31572 -3120
rect -31652 -12240 -31572 -7440
rect -31492 -9504 -31412 -960
rect -31180 -864 -31084 -854
rect -31180 -970 -31084 -960
rect -31180 -3024 -31084 -3014
rect -31180 -3130 -31084 -3120
rect -31180 -3744 -31084 -3734
rect -31180 -3850 -31084 -3840
rect -31180 -4932 -31084 -4922
rect -31180 -5038 -31084 -5028
rect -31180 -5292 -31084 -5282
rect -31180 -5398 -31084 -5388
rect -31180 -5904 -31084 -5894
rect -31180 -6010 -31084 -6000
rect -31180 -7344 -31084 -7334
rect -31180 -7450 -31084 -7440
rect -31492 -12032 -31412 -9600
rect -31180 -9504 -31084 -9494
rect -31180 -9610 -31084 -9600
rect -23088 -11200 -22984 -11190
rect -23088 -11314 -22984 -11304
rect -27136 -11408 -27032 -11398
rect -27136 -11522 -27032 -11512
rect -29160 -11616 -29056 -11606
rect -29160 -11730 -29056 -11720
rect -30172 -11824 -30068 -11814
rect -30172 -11938 -30068 -11928
rect -31492 -12146 -31412 -12136
rect -31652 -12354 -31572 -12344
rect -31812 -12562 -31732 -12552
rect -32504 -12770 -32424 -12760
rect -32664 -12978 -32584 -12968
rect -32824 -13186 -32744 -13176
<< via2 >>
rect -32192 -960 -32096 -864
rect -32192 -3120 -32096 -3024
rect -32192 -3840 -32096 -3744
rect -40292 -11304 -40188 -11200
rect -36244 -11512 -36140 -11408
rect -34220 -11720 -34116 -11616
rect -33208 -11928 -33104 -11824
rect -32192 -4668 -32096 -4572
rect -32192 -5748 -32096 -5652
rect -32192 -6000 -32096 -5904
rect -32192 -7440 -32096 -7344
rect -32192 -9600 -32096 -9504
rect -31180 -960 -31084 -864
rect -31180 -3120 -31084 -3024
rect -31180 -3840 -31084 -3744
rect -31180 -5028 -31084 -4932
rect -31180 -5388 -31084 -5292
rect -31180 -6000 -31084 -5904
rect -31180 -7440 -31084 -7344
rect -31180 -9600 -31084 -9504
rect -23088 -11304 -22984 -11200
rect -27136 -11512 -27032 -11408
rect -29160 -11720 -29056 -11616
rect -30172 -11928 -30068 -11824
<< metal3 >>
rect -32202 -864 -32086 -859
rect -32202 -960 -32192 -864
rect -32096 -960 -32086 -864
rect -32202 -965 -32086 -960
rect -31190 -864 -31074 -859
rect -31190 -960 -31180 -864
rect -31084 -960 -31074 -864
rect -31190 -965 -31074 -960
rect -32202 -3024 -32086 -3019
rect -32202 -3120 -32192 -3024
rect -32096 -3120 -32086 -3024
rect -32202 -3125 -32086 -3120
rect -31190 -3024 -31074 -3019
rect -31190 -3120 -31180 -3024
rect -31084 -3120 -31074 -3024
rect -31190 -3125 -31074 -3120
rect -32202 -3744 -32086 -3739
rect -32202 -3840 -32192 -3744
rect -32096 -3840 -32086 -3744
rect -32202 -3845 -32086 -3840
rect -31190 -3744 -31074 -3739
rect -31190 -3840 -31180 -3744
rect -31084 -3840 -31074 -3744
rect -31190 -3845 -31074 -3840
rect -32202 -4572 -32086 -4567
rect -32202 -4668 -32192 -4572
rect -32096 -4668 -32086 -4572
rect -32202 -4673 -32086 -4668
rect -31190 -4932 -31074 -4927
rect -31190 -5028 -31180 -4932
rect -31084 -5028 -31074 -4932
rect -31190 -5033 -31074 -5028
rect -31190 -5292 -31074 -5287
rect -31190 -5388 -31180 -5292
rect -31084 -5388 -31074 -5292
rect -31190 -5393 -31074 -5388
rect -32202 -5652 -32086 -5647
rect -32202 -5748 -32192 -5652
rect -32096 -5748 -32086 -5652
rect -32202 -5753 -32086 -5748
rect -32202 -5904 -32086 -5899
rect -32202 -6000 -32192 -5904
rect -32096 -6000 -32086 -5904
rect -32202 -6005 -32086 -6000
rect -31190 -5904 -31074 -5899
rect -31190 -6000 -31180 -5904
rect -31084 -6000 -31074 -5904
rect -31190 -6005 -31074 -6000
rect -32202 -7344 -32086 -7339
rect -32202 -7440 -32192 -7344
rect -32096 -7440 -32086 -7344
rect -32202 -7445 -32086 -7440
rect -31190 -7344 -31074 -7339
rect -31190 -7440 -31180 -7344
rect -31084 -7440 -31074 -7344
rect -31190 -7445 -31074 -7440
rect -32202 -9504 -32086 -9499
rect -32202 -9600 -32192 -9504
rect -32096 -9600 -32086 -9504
rect -32202 -9605 -32086 -9600
rect -31190 -9504 -31074 -9499
rect -31190 -9600 -31180 -9504
rect -31084 -9600 -31074 -9504
rect -31190 -9605 -31074 -9600
rect -40302 -11200 -40178 -11195
rect -40302 -11304 -40292 -11200
rect -40188 -11304 -40178 -11200
rect -40302 -11309 -40178 -11304
rect -23098 -11200 -22974 -11195
rect -23098 -11304 -23088 -11200
rect -22984 -11304 -22974 -11200
rect -23098 -11309 -22974 -11304
rect -36254 -11408 -36130 -11403
rect -36254 -11512 -36244 -11408
rect -36140 -11512 -36130 -11408
rect -36254 -11517 -36130 -11512
rect -27146 -11408 -27022 -11403
rect -27146 -11512 -27136 -11408
rect -27032 -11512 -27022 -11408
rect -27146 -11517 -27022 -11512
rect -34230 -11616 -34106 -11611
rect -34230 -11720 -34220 -11616
rect -34116 -11720 -34106 -11616
rect -34230 -11725 -34106 -11720
rect -29170 -11616 -29046 -11611
rect -29170 -11720 -29160 -11616
rect -29056 -11720 -29046 -11616
rect -29170 -11725 -29046 -11720
rect -33218 -11824 -33094 -11819
rect -33218 -11928 -33208 -11824
rect -33104 -11928 -33094 -11824
rect -33218 -11933 -33094 -11928
rect -30182 -11824 -30058 -11819
rect -30182 -11928 -30172 -11824
rect -30068 -11928 -30058 -11824
rect -30182 -11933 -30058 -11928
<< via3 >>
rect -32192 -960 -32096 -864
rect -31180 -960 -31084 -864
rect -32192 -3120 -32096 -3024
rect -31180 -3120 -31084 -3024
rect -32192 -3840 -32096 -3744
rect -31180 -3840 -31084 -3744
rect -32192 -6000 -32096 -5904
rect -31180 -6000 -31084 -5904
rect -32192 -7440 -32096 -7344
rect -31180 -7440 -31084 -7344
rect -32192 -9600 -32096 -9504
rect -31180 -9600 -31084 -9504
rect -40292 -11304 -40188 -11200
rect -23088 -11304 -22984 -11200
rect -36244 -11512 -36140 -11408
rect -27136 -11512 -27032 -11408
rect -34220 -11720 -34116 -11616
rect -29160 -11720 -29056 -11616
rect -33208 -11928 -33104 -11824
rect -30172 -11928 -30068 -11824
<< metal4 >>
rect -48044 704 -15850 808
rect -47856 600 -47752 704
rect -46844 600 -46740 704
rect -45832 600 -45728 704
rect -44820 600 -44716 704
rect -43808 600 -43704 704
rect -42796 600 -42692 704
rect -41784 600 -41680 704
rect -40772 600 -40668 704
rect -39760 600 -39656 704
rect -38748 600 -38644 704
rect -37736 600 -37632 704
rect -36724 600 -36620 704
rect -35712 600 -35608 704
rect -34700 600 -34596 704
rect -33688 600 -33584 704
rect -32676 600 -32572 704
rect -31664 600 -31560 704
rect -30652 455 -30548 704
rect -29640 463 -29536 704
rect -28628 600 -28524 704
rect -27616 600 -27512 704
rect -26604 600 -26500 704
rect -25592 600 -25488 704
rect -24580 600 -24476 704
rect -23568 600 -23464 704
rect -22556 600 -22452 704
rect -21544 600 -21440 704
rect -20532 600 -20428 704
rect -19520 600 -19416 704
rect -18508 600 -18404 704
rect -17496 600 -17392 704
rect -16484 600 -16380 704
rect -32192 -863 -32096 12
rect -31180 -863 -31084 12
rect -32193 -864 -32095 -863
rect -32193 -960 -32192 -864
rect -32096 -960 -32095 -864
rect -32193 -961 -32095 -960
rect -31181 -864 -31083 -863
rect -31181 -960 -31180 -864
rect -31084 -960 -31083 -864
rect -31181 -961 -31083 -960
rect -32192 -1692 -32096 -961
rect -31180 -1692 -31084 -961
rect -32192 -3023 -32096 -2868
rect -31180 -3023 -31084 -2868
rect -32193 -3024 -32095 -3023
rect -32193 -3120 -32192 -3024
rect -32096 -3120 -32095 -3024
rect -32193 -3121 -32095 -3120
rect -31181 -3024 -31083 -3023
rect -31181 -3120 -31180 -3024
rect -31084 -3120 -31083 -3024
rect -31181 -3121 -31083 -3120
rect -32192 -3132 -32096 -3121
rect -31180 -3132 -31084 -3121
rect -32193 -3744 -32095 -3743
rect -32193 -3840 -32192 -3744
rect -32096 -3840 -32095 -3744
rect -32193 -3841 -32095 -3840
rect -31181 -3744 -31083 -3743
rect -31181 -3840 -31180 -3744
rect -31084 -3840 -31083 -3744
rect -31181 -3841 -31083 -3840
rect -32192 -3854 -32096 -3841
rect -31180 -3852 -31084 -3841
rect -32193 -5904 -32095 -5903
rect -32193 -6000 -32192 -5904
rect -32096 -6000 -32095 -5904
rect -32193 -6001 -32095 -6000
rect -31181 -5904 -31083 -5903
rect -31181 -6000 -31180 -5904
rect -31084 -6000 -31083 -5904
rect -31181 -6001 -31083 -6000
rect -32192 -6012 -32096 -6001
rect -31180 -6012 -31084 -6001
rect -32192 -7343 -32096 -7188
rect -31180 -7343 -31084 -7188
rect -32193 -7344 -32095 -7343
rect -32193 -7440 -32192 -7344
rect -32096 -7440 -32095 -7344
rect -32193 -7441 -32095 -7440
rect -31181 -7344 -31083 -7343
rect -31181 -7440 -31180 -7344
rect -31084 -7440 -31083 -7344
rect -31181 -7441 -31083 -7440
rect -32192 -7452 -32096 -7441
rect -31180 -7452 -31084 -7441
rect -32192 -9503 -32096 -8628
rect -31180 -9503 -31084 -8628
rect -32193 -9504 -32095 -9503
rect -32193 -9600 -32192 -9504
rect -32096 -9600 -32095 -9504
rect -32193 -9601 -32095 -9600
rect -31181 -9504 -31083 -9503
rect -31181 -9600 -31180 -9504
rect -31084 -9600 -31083 -9504
rect -31181 -9601 -31083 -9600
rect -32192 -10332 -32096 -9601
rect -31180 -10332 -31084 -9601
rect -47376 -11024 -47272 -10920
rect -46364 -11024 -46260 -10920
rect -45352 -11024 -45248 -10920
rect -44340 -11024 -44236 -10920
rect -43328 -11024 -43224 -10920
rect -42316 -11024 -42212 -10920
rect -41304 -11024 -41200 -10920
rect -40292 -11024 -40188 -10920
rect -47376 -11128 -40188 -11024
rect -39280 -11024 -39176 -10920
rect -38268 -11024 -38164 -10920
rect -37256 -11024 -37152 -10920
rect -36244 -11024 -36140 -10920
rect -39280 -11128 -36140 -11024
rect -35232 -11024 -35128 -10920
rect -34220 -11024 -34116 -10920
rect -35232 -11128 -34116 -11024
rect -40292 -11199 -40188 -11128
rect -40293 -11200 -40187 -11199
rect -40293 -11304 -40292 -11200
rect -40188 -11304 -40187 -11200
rect -40293 -11305 -40187 -11304
rect -36244 -11407 -36140 -11128
rect -36245 -11408 -36139 -11407
rect -36245 -11512 -36244 -11408
rect -36140 -11512 -36139 -11408
rect -36245 -11513 -36139 -11512
rect -34220 -11615 -34116 -11128
rect -34221 -11616 -34115 -11615
rect -34221 -11720 -34220 -11616
rect -34116 -11720 -34115 -11616
rect -34221 -11721 -34115 -11720
rect -33208 -11823 -33104 -10920
rect -30172 -11823 -30068 -10857
rect -29160 -11024 -29056 -10920
rect -28148 -11024 -28044 -10816
rect -29160 -11128 -28044 -11024
rect -27136 -11024 -27032 -10920
rect -26124 -11024 -26020 -10816
rect -25112 -11024 -25008 -10810
rect -24100 -11024 -23996 -10816
rect -27136 -11128 -23996 -11024
rect -23088 -11024 -22984 -10920
rect -22076 -11024 -21972 -10816
rect -21064 -11024 -20960 -10816
rect -20052 -11024 -19948 -10811
rect -19040 -11024 -18936 -10816
rect -18028 -11024 -17924 -10811
rect -17016 -11024 -16912 -10816
rect -16004 -11024 -15900 -10816
rect -23088 -11128 -15900 -11024
rect -29160 -11615 -29056 -11128
rect -27136 -11407 -27032 -11128
rect -23088 -11199 -22984 -11128
rect -23089 -11200 -22983 -11199
rect -23089 -11304 -23088 -11200
rect -22984 -11304 -22983 -11200
rect -23089 -11305 -22983 -11304
rect -27137 -11408 -27031 -11407
rect -27137 -11512 -27136 -11408
rect -27032 -11512 -27031 -11408
rect -27137 -11513 -27031 -11512
rect -29161 -11616 -29055 -11615
rect -29161 -11720 -29160 -11616
rect -29056 -11720 -29055 -11616
rect -29161 -11721 -29055 -11720
rect -33209 -11824 -33103 -11823
rect -33209 -11928 -33208 -11824
rect -33104 -11928 -33103 -11824
rect -33209 -11929 -33103 -11928
rect -30173 -11824 -30067 -11823
rect -30173 -11928 -30172 -11824
rect -30068 -11928 -30067 -11824
rect -30173 -11929 -30067 -11928
use sky130_fd_pr__cap_mim_m3_1_NLQ4WR  sky130_fd_pr__cap_mim_m3_1_NLQ4WR_0
timestamp 1757810374
transform 1 0 -31972 0 1 -5160
box -892 -5760 892 5760
use sky130_fd_pr__cap_mim_m3_1_TE2UD4  sky130_fd_pr__cap_mim_m3_1_TE2UD4_0
timestamp 1757858808
transform 1 0 -40574 0 1 -5160
box -7470 -5760 7470 5760
use sky130_fd_pr__cap_mim_m3_1_TE2UD4  sky130_fd_pr__cap_mim_m3_1_TE2UD4_1
timestamp 1757858808
transform 1 0 -23370 0 1 -5160
box -7470 -5760 7470 5760
<< labels >>
flabel metal1 -16004 -13176 -15900 -13072 0 FreeSans 320 0 0 0 VCM
port 10 nsew
flabel metal1 -16004 -11304 -15900 -11200 0 FreeSans 320 0 0 0 S[0]
port 9 nsew
flabel metal1 -16004 -11512 -15900 -11408 0 FreeSans 320 0 0 0 S[1]
port 8 nsew
flabel metal1 -16004 -11720 -15900 -11616 0 FreeSans 320 0 0 0 S[2]
port 7 nsew
flabel metal1 -16004 -11928 -15900 -11824 0 FreeSans 320 0 0 0 S[3]
port 6 nsew
flabel metal1 -16004 -12136 -15900 -12032 0 FreeSans 320 0 0 0 S[4]
port 5 nsew
flabel metal1 -16004 -12344 -15900 -12240 0 FreeSans 320 0 0 0 S[5]
port 4 nsew
flabel metal1 -16004 -12552 -15900 -12448 0 FreeSans 320 0 0 0 S[6]
port 3 nsew
flabel metal1 -16004 -12760 -15900 -12656 0 FreeSans 320 0 0 0 S[7]
port 2 nsew
flabel metal1 -16004 -12968 -15900 -12864 0 FreeSans 320 0 0 0 S[8]
port 1 nsew
<< end >>
