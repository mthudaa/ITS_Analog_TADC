magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -38 332 2150 704
<< pwell >>
rect 4 49 2111 248
rect 0 0 2112 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 456 368 486 592
rect 546 368 576 592
rect 636 368 666 592
rect 726 368 756 592
rect 816 368 846 592
rect 906 368 936 592
rect 996 368 1026 592
rect 1086 368 1116 592
rect 1176 368 1206 592
rect 1266 368 1296 592
rect 1356 368 1386 592
rect 1446 368 1476 592
rect 1546 368 1576 592
rect 1636 368 1666 592
rect 1726 368 1756 592
rect 1816 368 1846 592
rect 1906 368 1936 592
rect 1996 368 2026 592
<< nmoslvt >>
rect 87 74 117 222
rect 173 74 203 222
rect 259 74 289 222
rect 345 74 375 222
rect 431 74 461 222
rect 517 74 547 222
rect 603 74 633 222
rect 689 74 719 222
rect 775 74 805 222
rect 861 74 891 222
rect 975 74 1005 222
rect 1061 74 1091 222
rect 1175 74 1205 222
rect 1261 74 1291 222
rect 1375 74 1405 222
rect 1461 74 1491 222
rect 1547 74 1577 222
rect 1633 74 1663 222
rect 1719 74 1749 222
rect 1805 74 1835 222
rect 1898 74 1928 222
rect 1998 74 2028 222
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 210 173 222
rect 117 176 128 210
rect 162 176 173 210
rect 117 120 173 176
rect 117 86 128 120
rect 162 86 173 120
rect 117 74 173 86
rect 203 210 259 222
rect 203 176 214 210
rect 248 176 259 210
rect 203 116 259 176
rect 203 82 214 116
rect 248 82 259 116
rect 203 74 259 82
rect 289 210 345 222
rect 289 176 300 210
rect 334 176 345 210
rect 289 120 345 176
rect 289 86 300 120
rect 334 86 345 120
rect 289 74 345 86
rect 375 210 431 222
rect 375 176 386 210
rect 420 176 431 210
rect 375 116 431 176
rect 375 82 386 116
rect 420 82 431 116
rect 375 74 431 82
rect 461 210 517 222
rect 461 176 472 210
rect 506 176 517 210
rect 461 120 517 176
rect 461 86 472 120
rect 506 86 517 120
rect 461 74 517 86
rect 547 187 603 222
rect 547 153 558 187
rect 592 153 603 187
rect 547 116 603 153
rect 547 82 558 116
rect 592 82 603 116
rect 547 74 603 82
rect 633 210 689 222
rect 633 176 644 210
rect 678 176 689 210
rect 633 120 689 176
rect 633 86 644 120
rect 678 86 689 120
rect 633 74 689 86
rect 719 210 775 222
rect 719 176 730 210
rect 764 176 775 210
rect 719 116 775 176
rect 719 82 730 116
rect 764 82 775 116
rect 719 74 775 82
rect 805 210 861 222
rect 805 176 816 210
rect 850 176 861 210
rect 805 120 861 176
rect 805 86 816 120
rect 850 86 861 120
rect 805 74 861 86
rect 891 210 975 222
rect 891 176 916 210
rect 950 176 975 210
rect 891 116 975 176
rect 891 82 916 116
rect 950 82 975 116
rect 891 74 975 82
rect 1005 210 1061 222
rect 1005 176 1016 210
rect 1050 176 1061 210
rect 1005 120 1061 176
rect 1005 86 1016 120
rect 1050 86 1061 120
rect 1005 74 1061 86
rect 1091 191 1175 222
rect 1091 157 1116 191
rect 1150 157 1175 191
rect 1091 116 1175 157
rect 1091 82 1116 116
rect 1150 82 1175 116
rect 1091 74 1175 82
rect 1205 210 1261 222
rect 1205 176 1216 210
rect 1250 176 1261 210
rect 1205 120 1261 176
rect 1205 86 1216 120
rect 1250 86 1261 120
rect 1205 74 1261 86
rect 1291 210 1375 222
rect 1291 176 1316 210
rect 1350 176 1375 210
rect 1291 116 1375 176
rect 1291 82 1316 116
rect 1350 82 1375 116
rect 1291 74 1375 82
rect 1405 210 1461 222
rect 1405 176 1416 210
rect 1450 176 1461 210
rect 1405 120 1461 176
rect 1405 86 1416 120
rect 1450 86 1461 120
rect 1405 74 1461 86
rect 1491 152 1547 222
rect 1491 118 1502 152
rect 1536 118 1547 152
rect 1491 74 1547 118
rect 1577 210 1633 222
rect 1577 176 1588 210
rect 1622 176 1633 210
rect 1577 120 1633 176
rect 1577 86 1588 120
rect 1622 86 1633 120
rect 1577 74 1633 86
rect 1663 152 1719 222
rect 1663 118 1674 152
rect 1708 118 1719 152
rect 1663 74 1719 118
rect 1749 210 1805 222
rect 1749 176 1760 210
rect 1794 176 1805 210
rect 1749 120 1805 176
rect 1749 86 1760 120
rect 1794 86 1805 120
rect 1749 74 1805 86
rect 1835 152 1898 222
rect 1835 118 1846 152
rect 1880 118 1898 152
rect 1835 74 1898 118
rect 1928 210 1998 222
rect 1928 176 1939 210
rect 1973 176 1998 210
rect 1928 120 1998 176
rect 1928 86 1939 120
rect 1973 86 1998 120
rect 1928 74 1998 86
rect 2028 210 2085 222
rect 2028 176 2039 210
rect 2073 176 2085 210
rect 2028 120 2085 176
rect 2028 86 2039 120
rect 2073 86 2085 120
rect 2028 74 2085 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 497 176 546
rect 116 463 129 497
rect 163 463 176 497
rect 116 414 176 463
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 579 266 592
rect 206 545 219 579
rect 253 545 266 579
rect 206 511 266 545
rect 206 477 219 511
rect 253 477 266 511
rect 206 443 266 477
rect 206 409 219 443
rect 253 409 266 443
rect 206 368 266 409
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 497 356 546
rect 296 463 309 497
rect 343 463 356 497
rect 296 414 356 463
rect 296 380 309 414
rect 343 380 356 414
rect 296 368 356 380
rect 386 579 456 592
rect 386 545 409 579
rect 443 545 456 579
rect 386 511 456 545
rect 386 477 409 511
rect 443 477 456 511
rect 386 443 456 477
rect 386 409 409 443
rect 443 409 456 443
rect 386 368 456 409
rect 486 580 546 592
rect 486 546 499 580
rect 533 546 546 580
rect 486 497 546 546
rect 486 463 499 497
rect 533 463 546 497
rect 486 414 546 463
rect 486 380 499 414
rect 533 380 546 414
rect 486 368 546 380
rect 576 580 636 592
rect 576 546 589 580
rect 623 546 636 580
rect 576 512 636 546
rect 576 478 589 512
rect 623 478 636 512
rect 576 443 636 478
rect 576 409 589 443
rect 623 409 636 443
rect 576 368 636 409
rect 666 580 726 592
rect 666 546 679 580
rect 713 546 726 580
rect 666 497 726 546
rect 666 463 679 497
rect 713 463 726 497
rect 666 414 726 463
rect 666 380 679 414
rect 713 380 726 414
rect 666 368 726 380
rect 756 579 816 592
rect 756 545 769 579
rect 803 545 816 579
rect 756 511 816 545
rect 756 477 769 511
rect 803 477 816 511
rect 756 443 816 477
rect 756 409 769 443
rect 803 409 816 443
rect 756 368 816 409
rect 846 580 906 592
rect 846 546 859 580
rect 893 546 906 580
rect 846 497 906 546
rect 846 463 859 497
rect 893 463 906 497
rect 846 414 906 463
rect 846 380 859 414
rect 893 380 906 414
rect 846 368 906 380
rect 936 580 996 592
rect 936 546 949 580
rect 983 546 996 580
rect 936 511 996 546
rect 936 477 949 511
rect 983 477 996 511
rect 936 443 996 477
rect 936 409 949 443
rect 983 409 996 443
rect 936 368 996 409
rect 1026 580 1086 592
rect 1026 546 1039 580
rect 1073 546 1086 580
rect 1026 497 1086 546
rect 1026 463 1039 497
rect 1073 463 1086 497
rect 1026 414 1086 463
rect 1026 380 1039 414
rect 1073 380 1086 414
rect 1026 368 1086 380
rect 1116 579 1176 592
rect 1116 545 1129 579
rect 1163 545 1176 579
rect 1116 511 1176 545
rect 1116 477 1129 511
rect 1163 477 1176 511
rect 1116 443 1176 477
rect 1116 409 1129 443
rect 1163 409 1176 443
rect 1116 368 1176 409
rect 1206 580 1266 592
rect 1206 546 1219 580
rect 1253 546 1266 580
rect 1206 497 1266 546
rect 1206 463 1219 497
rect 1253 463 1266 497
rect 1206 414 1266 463
rect 1206 380 1219 414
rect 1253 380 1266 414
rect 1206 368 1266 380
rect 1296 580 1356 592
rect 1296 546 1309 580
rect 1343 546 1356 580
rect 1296 511 1356 546
rect 1296 477 1309 511
rect 1343 477 1356 511
rect 1296 443 1356 477
rect 1296 409 1309 443
rect 1343 409 1356 443
rect 1296 368 1356 409
rect 1386 580 1446 592
rect 1386 546 1399 580
rect 1433 546 1446 580
rect 1386 497 1446 546
rect 1386 463 1399 497
rect 1433 463 1446 497
rect 1386 414 1446 463
rect 1386 380 1399 414
rect 1433 380 1446 414
rect 1386 368 1446 380
rect 1476 580 1546 592
rect 1476 546 1489 580
rect 1523 546 1546 580
rect 1476 508 1546 546
rect 1476 474 1489 508
rect 1523 474 1546 508
rect 1476 368 1546 474
rect 1576 580 1636 592
rect 1576 546 1589 580
rect 1623 546 1636 580
rect 1576 510 1636 546
rect 1576 476 1589 510
rect 1623 476 1636 510
rect 1576 440 1636 476
rect 1576 406 1589 440
rect 1623 406 1636 440
rect 1576 368 1636 406
rect 1666 580 1726 592
rect 1666 546 1679 580
rect 1713 546 1726 580
rect 1666 508 1726 546
rect 1666 474 1679 508
rect 1713 474 1726 508
rect 1666 368 1726 474
rect 1756 580 1816 592
rect 1756 546 1769 580
rect 1803 546 1816 580
rect 1756 510 1816 546
rect 1756 476 1769 510
rect 1803 476 1816 510
rect 1756 440 1816 476
rect 1756 406 1769 440
rect 1803 406 1816 440
rect 1756 368 1816 406
rect 1846 580 1906 592
rect 1846 546 1859 580
rect 1893 546 1906 580
rect 1846 508 1906 546
rect 1846 474 1859 508
rect 1893 474 1906 508
rect 1846 368 1906 474
rect 1936 580 1996 592
rect 1936 546 1949 580
rect 1983 546 1996 580
rect 1936 510 1996 546
rect 1936 476 1949 510
rect 1983 476 1996 510
rect 1936 440 1996 476
rect 1936 406 1949 440
rect 1983 406 1996 440
rect 1936 368 1996 406
rect 2026 580 2085 592
rect 2026 546 2039 580
rect 2073 546 2085 580
rect 2026 510 2085 546
rect 2026 476 2039 510
rect 2073 476 2085 510
rect 2026 440 2085 476
rect 2026 406 2039 440
rect 2073 406 2085 440
rect 2026 368 2085 406
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 176 162 210
rect 128 86 162 120
rect 214 176 248 210
rect 214 82 248 116
rect 300 176 334 210
rect 300 86 334 120
rect 386 176 420 210
rect 386 82 420 116
rect 472 176 506 210
rect 472 86 506 120
rect 558 153 592 187
rect 558 82 592 116
rect 644 176 678 210
rect 644 86 678 120
rect 730 176 764 210
rect 730 82 764 116
rect 816 176 850 210
rect 816 86 850 120
rect 916 176 950 210
rect 916 82 950 116
rect 1016 176 1050 210
rect 1016 86 1050 120
rect 1116 157 1150 191
rect 1116 82 1150 116
rect 1216 176 1250 210
rect 1216 86 1250 120
rect 1316 176 1350 210
rect 1316 82 1350 116
rect 1416 176 1450 210
rect 1416 86 1450 120
rect 1502 118 1536 152
rect 1588 176 1622 210
rect 1588 86 1622 120
rect 1674 118 1708 152
rect 1760 176 1794 210
rect 1760 86 1794 120
rect 1846 118 1880 152
rect 1939 176 1973 210
rect 1939 86 1973 120
rect 2039 176 2073 210
rect 2039 86 2073 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 545 253 579
rect 219 477 253 511
rect 219 409 253 443
rect 309 546 343 580
rect 309 463 343 497
rect 309 380 343 414
rect 409 545 443 579
rect 409 477 443 511
rect 409 409 443 443
rect 499 546 533 580
rect 499 463 533 497
rect 499 380 533 414
rect 589 546 623 580
rect 589 478 623 512
rect 589 409 623 443
rect 679 546 713 580
rect 679 463 713 497
rect 679 380 713 414
rect 769 545 803 579
rect 769 477 803 511
rect 769 409 803 443
rect 859 546 893 580
rect 859 463 893 497
rect 859 380 893 414
rect 949 546 983 580
rect 949 477 983 511
rect 949 409 983 443
rect 1039 546 1073 580
rect 1039 463 1073 497
rect 1039 380 1073 414
rect 1129 545 1163 579
rect 1129 477 1163 511
rect 1129 409 1163 443
rect 1219 546 1253 580
rect 1219 463 1253 497
rect 1219 380 1253 414
rect 1309 546 1343 580
rect 1309 477 1343 511
rect 1309 409 1343 443
rect 1399 546 1433 580
rect 1399 463 1433 497
rect 1399 380 1433 414
rect 1489 546 1523 580
rect 1489 474 1523 508
rect 1589 546 1623 580
rect 1589 476 1623 510
rect 1589 406 1623 440
rect 1679 546 1713 580
rect 1679 474 1713 508
rect 1769 546 1803 580
rect 1769 476 1803 510
rect 1769 406 1803 440
rect 1859 546 1893 580
rect 1859 474 1893 508
rect 1949 546 1983 580
rect 1949 476 1983 510
rect 1949 406 1983 440
rect 2039 546 2073 580
rect 2039 476 2073 510
rect 2039 406 2073 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 456 592 486 618
rect 546 592 576 618
rect 636 592 666 618
rect 726 592 756 618
rect 816 592 846 618
rect 906 592 936 618
rect 996 592 1026 618
rect 1086 592 1116 618
rect 1176 592 1206 618
rect 1266 592 1296 618
rect 1356 592 1386 618
rect 1446 592 1476 618
rect 1546 592 1576 618
rect 1636 592 1666 618
rect 1726 592 1756 618
rect 1816 592 1846 618
rect 1906 592 1936 618
rect 1996 592 2026 618
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 456 353 486 368
rect 546 353 576 368
rect 636 353 666 368
rect 726 353 756 368
rect 816 353 846 368
rect 906 353 936 368
rect 996 353 1026 368
rect 1086 353 1116 368
rect 1176 353 1206 368
rect 1266 353 1296 368
rect 1356 353 1386 368
rect 1446 353 1476 368
rect 1546 353 1576 368
rect 1636 353 1666 368
rect 1726 353 1756 368
rect 1816 353 1846 368
rect 1906 353 1936 368
rect 1996 353 2026 368
rect 83 326 119 353
rect 173 326 209 353
rect 263 326 299 353
rect 353 326 389 353
rect 453 326 489 353
rect 543 326 579 353
rect 633 326 669 353
rect 723 326 759 353
rect 813 326 849 353
rect 903 326 939 353
rect 993 326 1029 353
rect 1083 326 1119 353
rect 1173 326 1209 353
rect 1263 326 1299 353
rect 1353 326 1389 353
rect 1443 326 1479 353
rect 1543 336 1579 353
rect 1633 336 1669 353
rect 1723 336 1759 353
rect 1813 336 1849 353
rect 1903 336 1939 353
rect 1993 336 2029 353
rect 83 310 1491 326
rect 83 276 213 310
rect 247 276 390 310
rect 424 276 582 310
rect 616 276 755 310
rect 789 276 927 310
rect 961 276 1131 310
rect 1165 276 1316 310
rect 1350 276 1491 310
rect 83 260 1491 276
rect 1543 320 2029 336
rect 1543 286 1571 320
rect 1605 286 1639 320
rect 1673 286 1707 320
rect 1741 286 1775 320
rect 1809 286 1843 320
rect 1877 286 1911 320
rect 1945 286 1979 320
rect 2013 286 2029 320
rect 1543 270 2029 286
rect 87 222 117 260
rect 173 222 203 260
rect 259 222 289 260
rect 345 222 375 260
rect 431 222 461 260
rect 517 222 547 260
rect 603 222 633 260
rect 689 222 719 260
rect 775 222 805 260
rect 861 222 891 260
rect 975 222 1005 260
rect 1061 222 1091 260
rect 1175 222 1205 260
rect 1261 222 1291 260
rect 1375 222 1405 260
rect 1461 222 1491 260
rect 1547 222 1577 270
rect 1633 222 1663 270
rect 1719 222 1749 270
rect 1805 222 1835 270
rect 1898 222 1928 270
rect 1998 222 2028 270
rect 87 48 117 74
rect 173 48 203 74
rect 259 48 289 74
rect 345 48 375 74
rect 431 48 461 74
rect 517 48 547 74
rect 603 48 633 74
rect 689 48 719 74
rect 775 48 805 74
rect 861 48 891 74
rect 975 48 1005 74
rect 1061 48 1091 74
rect 1175 48 1205 74
rect 1261 48 1291 74
rect 1375 48 1405 74
rect 1461 48 1491 74
rect 1547 48 1577 74
rect 1633 48 1663 74
rect 1719 48 1749 74
rect 1805 48 1835 74
rect 1898 48 1928 74
rect 1998 48 2028 74
<< polycont >>
rect 213 276 247 310
rect 390 276 424 310
rect 582 276 616 310
rect 755 276 789 310
rect 927 276 961 310
rect 1131 276 1165 310
rect 1316 276 1350 310
rect 1571 286 1605 320
rect 1639 286 1673 320
rect 1707 286 1741 320
rect 1775 286 1809 320
rect 1843 286 1877 320
rect 1911 286 1945 320
rect 1979 286 2013 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 112 580 163 596
rect 112 546 129 580
rect 112 497 163 546
rect 112 463 129 497
rect 112 424 163 463
rect 112 390 127 424
rect 161 414 163 424
rect 219 579 253 649
rect 219 511 253 545
rect 219 443 253 477
rect 219 393 253 409
rect 293 580 344 596
rect 293 546 309 580
rect 343 546 344 580
rect 293 497 344 546
rect 293 463 309 497
rect 343 463 344 497
rect 293 424 344 463
rect 112 380 129 390
rect 26 210 76 226
rect 26 176 42 210
rect 26 120 76 176
rect 26 86 42 120
rect 26 17 76 86
rect 112 210 163 380
rect 293 390 303 424
rect 337 414 344 424
rect 293 380 309 390
rect 343 380 344 414
rect 393 579 443 649
rect 393 545 409 579
rect 393 511 443 545
rect 393 477 409 511
rect 393 443 443 477
rect 393 409 409 443
rect 393 393 443 409
rect 483 580 535 596
rect 483 546 499 580
rect 533 546 535 580
rect 483 497 535 546
rect 483 463 499 497
rect 533 463 535 497
rect 483 424 535 463
rect 197 350 259 356
rect 197 316 211 350
rect 245 316 259 350
rect 197 310 259 316
rect 197 276 213 310
rect 247 276 259 310
rect 197 260 259 276
rect 112 176 128 210
rect 162 176 163 210
rect 112 120 163 176
rect 112 86 128 120
rect 162 86 163 120
rect 112 70 163 86
rect 198 210 257 226
rect 198 176 214 210
rect 248 176 257 210
rect 198 116 257 176
rect 198 82 214 116
rect 248 82 257 116
rect 198 17 257 82
rect 293 210 344 380
rect 483 390 494 424
rect 528 414 535 424
rect 483 380 499 390
rect 533 380 535 414
rect 589 580 623 649
rect 589 512 623 546
rect 589 443 623 478
rect 589 393 623 409
rect 662 580 713 596
rect 662 546 679 580
rect 662 497 713 546
rect 662 463 679 497
rect 662 424 713 463
rect 378 350 435 356
rect 378 316 390 350
rect 424 316 435 350
rect 378 310 435 316
rect 378 276 390 310
rect 424 276 435 310
rect 378 260 435 276
rect 483 271 535 380
rect 662 390 672 424
rect 706 414 713 424
rect 769 579 803 649
rect 769 511 803 545
rect 769 443 803 477
rect 769 393 803 409
rect 843 580 909 596
rect 843 546 859 580
rect 893 546 909 580
rect 843 497 909 546
rect 843 463 859 497
rect 893 463 909 497
rect 843 424 909 463
rect 843 414 860 424
rect 662 380 679 390
rect 662 364 713 380
rect 843 380 859 414
rect 894 390 909 424
rect 949 580 983 649
rect 949 511 983 546
rect 949 443 983 477
rect 949 393 983 409
rect 1023 580 1082 596
rect 1023 546 1039 580
rect 1073 546 1082 580
rect 1023 497 1082 546
rect 1023 463 1039 497
rect 1073 463 1082 497
rect 1023 424 1082 463
rect 893 380 909 390
rect 1023 380 1039 424
rect 1073 380 1082 424
rect 1129 579 1163 649
rect 1129 511 1163 545
rect 1129 443 1163 477
rect 1129 393 1163 409
rect 1212 580 1266 596
rect 1212 546 1219 580
rect 1253 546 1266 580
rect 1212 497 1266 546
rect 1212 463 1219 497
rect 1253 463 1266 497
rect 1212 424 1266 463
rect 469 237 535 271
rect 569 350 628 356
rect 569 316 582 350
rect 616 316 628 350
rect 569 310 628 316
rect 569 276 582 310
rect 616 276 628 310
rect 569 260 628 276
rect 293 176 300 210
rect 334 176 344 210
rect 293 120 344 176
rect 293 86 300 120
rect 334 86 344 120
rect 293 70 344 86
rect 379 210 420 226
rect 379 176 386 210
rect 379 116 420 176
rect 379 82 386 116
rect 379 17 420 82
rect 469 210 522 237
rect 662 226 696 364
rect 747 350 809 356
rect 747 331 760 350
rect 731 316 760 331
rect 794 316 809 350
rect 731 310 809 316
rect 731 276 755 310
rect 789 276 809 310
rect 731 260 809 276
rect 843 226 877 380
rect 935 350 973 356
rect 935 346 936 350
rect 911 316 936 346
rect 970 316 973 350
rect 911 310 973 316
rect 911 276 927 310
rect 961 276 973 310
rect 911 260 973 276
rect 1023 275 1082 380
rect 1212 380 1219 424
rect 1253 380 1266 424
rect 1309 580 1343 649
rect 1309 511 1343 546
rect 1309 443 1343 477
rect 1309 393 1343 409
rect 1396 580 1449 596
rect 1396 546 1399 580
rect 1433 546 1449 580
rect 1396 497 1449 546
rect 1396 463 1399 497
rect 1433 463 1449 497
rect 1396 424 1449 463
rect 1489 580 1539 649
rect 1523 546 1539 580
rect 1489 508 1539 546
rect 1523 474 1539 508
rect 1489 458 1539 474
rect 1573 580 1639 596
rect 1573 546 1589 580
rect 1623 546 1639 580
rect 1573 510 1639 546
rect 1573 476 1589 510
rect 1623 476 1639 510
rect 1573 440 1639 476
rect 1679 580 1713 649
rect 1679 508 1713 546
rect 1679 458 1713 474
rect 1753 580 1819 596
rect 1753 546 1769 580
rect 1803 546 1819 580
rect 1753 510 1819 546
rect 1753 476 1769 510
rect 1803 476 1819 510
rect 1573 424 1589 440
rect 1396 414 1405 424
rect 1007 241 1082 275
rect 1116 350 1178 356
rect 1116 316 1130 350
rect 1164 316 1178 350
rect 1116 310 1178 316
rect 1116 276 1131 310
rect 1165 276 1178 310
rect 1116 260 1178 276
rect 469 176 472 210
rect 506 176 522 210
rect 644 210 696 226
rect 469 120 522 176
rect 469 86 472 120
rect 506 86 522 120
rect 469 70 522 86
rect 558 187 592 203
rect 558 116 592 153
rect 558 17 592 82
rect 678 176 696 210
rect 644 120 696 176
rect 678 86 696 120
rect 644 70 696 86
rect 730 210 764 226
rect 730 116 764 176
rect 730 17 764 82
rect 800 210 877 226
rect 800 176 816 210
rect 850 176 877 210
rect 800 120 877 176
rect 800 86 816 120
rect 850 86 877 120
rect 800 70 877 86
rect 911 210 966 226
rect 911 176 916 210
rect 950 176 966 210
rect 911 116 966 176
rect 911 82 916 116
rect 950 82 966 116
rect 911 17 966 82
rect 1007 210 1066 241
rect 1212 226 1266 380
rect 1396 380 1399 414
rect 1439 390 1449 424
rect 1433 380 1449 390
rect 1300 350 1362 356
rect 1300 316 1313 350
rect 1347 316 1362 350
rect 1300 310 1362 316
rect 1300 276 1316 310
rect 1350 276 1362 310
rect 1300 260 1362 276
rect 1396 250 1449 380
rect 1484 406 1589 424
rect 1623 424 1639 440
rect 1753 440 1819 476
rect 1859 580 1893 649
rect 1859 508 1893 546
rect 1859 458 1893 474
rect 1933 580 1999 596
rect 1933 546 1949 580
rect 1983 546 1999 580
rect 1933 510 1999 546
rect 1933 476 1949 510
rect 1983 476 1999 510
rect 1753 424 1769 440
rect 1623 406 1769 424
rect 1803 424 1819 440
rect 1933 440 1999 476
rect 1933 424 1949 440
rect 1803 406 1949 424
rect 1983 406 1999 440
rect 1484 390 1999 406
rect 2039 580 2089 649
rect 2073 546 2089 580
rect 2039 510 2089 546
rect 2073 476 2089 510
rect 2039 440 2089 476
rect 2073 406 2089 440
rect 2039 390 2089 406
rect 1484 350 1518 390
rect 1007 176 1016 210
rect 1050 176 1066 210
rect 1200 210 1266 226
rect 1007 120 1066 176
rect 1007 86 1016 120
rect 1050 86 1066 120
rect 1007 70 1066 86
rect 1100 191 1166 207
rect 1100 157 1116 191
rect 1150 157 1166 191
rect 1100 116 1166 157
rect 1100 82 1116 116
rect 1150 82 1166 116
rect 1100 17 1166 82
rect 1200 176 1216 210
rect 1250 176 1266 210
rect 1200 120 1266 176
rect 1200 86 1216 120
rect 1250 86 1266 120
rect 1200 70 1266 86
rect 1300 210 1366 226
rect 1300 176 1316 210
rect 1350 176 1366 210
rect 1300 116 1366 176
rect 1300 82 1316 116
rect 1350 82 1366 116
rect 1300 17 1366 82
rect 1400 210 1450 250
rect 1400 176 1416 210
rect 1484 236 1518 316
rect 1555 320 2087 356
rect 1555 286 1571 320
rect 1605 286 1639 320
rect 1673 286 1707 320
rect 1741 286 1775 320
rect 1809 286 1843 320
rect 1877 286 1911 320
rect 1945 286 1979 320
rect 2013 286 2087 320
rect 1555 270 2087 286
rect 1484 210 1989 236
rect 1484 202 1588 210
rect 1400 120 1450 176
rect 1622 202 1760 210
rect 1400 86 1416 120
rect 1400 70 1450 86
rect 1486 152 1552 168
rect 1486 118 1502 152
rect 1536 118 1552 152
rect 1486 17 1552 118
rect 1588 120 1622 176
rect 1794 202 1939 210
rect 1588 70 1622 86
rect 1658 152 1724 168
rect 1658 118 1674 152
rect 1708 118 1724 152
rect 1658 17 1724 118
rect 1760 120 1794 176
rect 1973 176 1989 210
rect 1760 70 1794 86
rect 1830 152 1896 168
rect 1830 118 1846 152
rect 1880 118 1896 152
rect 1830 17 1896 118
rect 1939 120 1989 176
rect 1973 86 1989 120
rect 1939 70 1989 86
rect 2023 210 2089 226
rect 2023 176 2039 210
rect 2073 176 2089 210
rect 2023 120 2089 176
rect 2023 86 2039 120
rect 2073 86 2089 120
rect 2023 17 2089 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 127 414 161 424
rect 127 390 129 414
rect 129 390 161 414
rect 303 414 337 424
rect 303 390 309 414
rect 309 390 337 414
rect 211 316 245 350
rect 494 414 528 424
rect 494 390 499 414
rect 499 390 528 414
rect 390 316 424 350
rect 672 414 706 424
rect 672 390 679 414
rect 679 390 706 414
rect 860 414 894 424
rect 860 390 893 414
rect 893 390 894 414
rect 1039 414 1073 424
rect 1039 390 1073 414
rect 582 316 616 350
rect 760 316 794 350
rect 936 316 970 350
rect 1219 414 1253 424
rect 1219 390 1253 414
rect 1405 414 1439 424
rect 1130 316 1164 350
rect 1405 390 1433 414
rect 1433 390 1439 414
rect 1313 316 1347 350
rect 1484 316 1518 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 115 424 1451 430
rect 115 390 127 424
rect 161 390 303 424
rect 337 390 494 424
rect 528 390 672 424
rect 706 390 860 424
rect 894 390 1039 424
rect 1073 390 1219 424
rect 1253 390 1405 424
rect 1439 390 1451 424
rect 115 384 1451 390
rect 197 350 1530 356
rect 197 316 211 350
rect 245 316 390 350
rect 424 316 582 350
rect 616 316 760 350
rect 794 316 936 350
rect 970 316 1130 350
rect 1164 316 1313 350
rect 1347 316 1484 350
rect 1518 316 1530 350
rect 197 310 1530 316
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_16
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 1 nsew
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 2 nsew
flabel metal1 s 115 384 1451 430 0 FreeSans 400 0 0 0 X
port 4 nsew
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 3 nsew
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A
port 7 nsew
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A
port 7 nsew
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A
port 7 nsew
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A
port 7 nsew
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2112 666
<< end >>
