* PEX produced on Tue Sep 16 01:29:14 AM CST 2025 using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from tt_um_tsar_adc.ext - technology: sky130A

.subckt tt_um_tsar_adc clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_out[0]
+ uio_out[1] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] VDPWR VGND
X0 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_8403_19478# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_13164_28398# sar9b_0._06_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4 VGND sar9b_0.net5 a_7914_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 VDPWR a_10098_19171# a_9900_19047# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X8 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDPWR a_4749_27652# sar9b_0.net58 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X13 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X14 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X15 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 a_7926_23234# sar9b_0.net62 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X19 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=31.32 ps=341.28 w=0.5 l=0.5
X20 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X22 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X23 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X24 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X26 a_5896_22188# a_4755_22138# a_5739_22488# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X27 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X28 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X30 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X31 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X33 a_40321_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X34 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X35 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X37 VGND a_13011_24802# single_9b_cdac_0.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X38 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B a_16970_11404# VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X39 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X40 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X41 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X43 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X44 a_12047_26517# a_11842_26426# a_11382_26138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X45 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X46 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X48 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X49 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 a_8438_18958# a_8303_18859# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X53 a_3855_25792# a_4125_25958# a_4083_25852# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.05565 ps=0.685 w=0.42 l=0.15
X54 VGND a_12870_22267# a_12828_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X55 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X56 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X57 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X58 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X59 VGND sar9b_0.net52 a_12246_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X60 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VGND sar9b_0.clknet_1_1__leaf_CLK a_2835_24136# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X62 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X63 VGND a_13011_23238# single_9b_cdac_1.CF[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X64 a_5182_22567# sar9b_0.net64 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X65 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X66 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X67 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X68 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X69 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=282.12262 ps=2.58843k w=0.42 l=1
X70 a_12047_22521# a_11658_22138# a_11382_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X71 a_5196_19448# sar9b_0.net16 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X72 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X73 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X75 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X77 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X78 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X80 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X81 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X82 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X83 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X84 sar9b_0.net34 a_10284_25707# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X85 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X86 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X87 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VGND sar9b_0.net47 a_7062_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VGND a_11915_28371# uo_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X92 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X93 a_7890_26108# a_8345_26455# a_8294_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X94 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X96 VDPWR sar9b_0.net59 a_2847_26141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X97 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X98 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X99 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X100 a_12828_22145# a_11658_22138# a_12618_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X101 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X102 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X103 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 a_2918_20140# a_2739_20140# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X105 a_7343_27849# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X106 VDPWR a_11178_24802# a_11430_24931# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X107 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X108 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X109 VDPWR a_4771_18260# sar9b_0.net56 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X110 a_6634_18206# sar9b_0.net73 a_7155_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X111 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X112 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X113 a_10895_22855# a_10690_22806# a_10230_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X114 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X115 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10254_2858# dw_12589_1395# dw_12589_1395# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X116 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X117 a_26951_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X118 VGND a_6880_26815# sar9b_0.net21 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X119 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X120 single_9b_cdac_0.SW[7] a_10859_26330# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X121 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X122 a_2706_26108# a_3161_26455# a_3110_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X124 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X125 a_6534_27123# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X126 a_7978_22202# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X127 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X130 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 a_11842_19766# a_11658_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X132 VDPWR sar9b_0.net17 a_2931_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X133 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X135 a_11436_17742# sar9b_0.net2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X136 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X137 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 a_7155_18146# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X140 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X141 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X142 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 uo_out[0] a_11915_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X145 VGND a_4044_24776# sar9b_0.net72 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X146 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X147 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X148 sar9b_0.net40 a_6444_19448# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X149 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X153 VDPWR a_13216_23805# sar9b_0.net32 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X154 single_9b_cdac_1.SW[6] a_13011_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X155 VGND a_9588_27045# a_9593_26914# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X156 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X159 VGND sar9b_0.net52 a_10710_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X161 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X162 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=486.22675 ps=3.99183k w=1 l=1
X165 sar9b_0.net1 a_6867_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X166 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X167 a_5962_24151# a_5753_24250# a_5298_24499# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X168 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X169 VDPWR a_6834_20780# a_6636_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X170 a_10098_19171# a_10548_19053# a_10500_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X171 a_3561_22527# a_3027_22138# a_3454_22567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X172 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X176 a_12618_18142# a_11842_18434# a_12182_18427# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X177 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X178 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X179 a_8006_17229# a_7743_16817# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X180 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[1] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X182 a_9414_23127# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X183 a_6444_21738# sar9b_0._02_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X187 a_7404_17715# sar9b_0.net1 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24915 pd=2.37 as=0.15198 ps=1.17 w=0.55 l=0.15
X188 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VDPWR sar9b_0.net58 a_5046_27230# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X190 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X191 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X192 a_11568_24809# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X193 a_7831_22521# a_7402_22441# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X194 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X196 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X197 a_4072_19474# sar9b_0.net46 a_3994_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.20165 pd=1.285 as=0.0888 ps=0.98 w=0.74 l=0.15
X198 VGND a_8166_27595# a_8124_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X199 a_8842_16874# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X200 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X201 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 single_9b_cdac_0.SW[3] a_12491_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X204 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X205 sar9b_0.net18 a_2508_27440# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X206 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X207 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=93.96 ps=773.28003 w=1.5 l=0.5
X208 VDPWR sar9b_0._10_ a_4496_20468# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 th_dif_sw_0.CK a_10227_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X212 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X214 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X215 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X216 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X219 a_5459_22165# a_4934_22432# a_5289_22527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X220 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X222 VDPWR a_10932_25713# a_10937_25582# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X224 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X225 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X226 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X227 a_5506_17478# a_5322_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X228 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 a_8124_27473# a_6954_27466# a_7914_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X231 VDPWR a_7590_24931# a_7540_25221# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X232 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X233 a_10830_19068# a_10548_19053# a_11191_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X234 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDPWR a_5235_27466# uo_out[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X236 VGND a_4210_22378# a_4168_22188# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X237 a_6038_20140# a_5126_20140# a_5931_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X238 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X239 VDPWR sar9b_0.net22 a_8691_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X240 a_4011_22488# a_3206_22432# a_3713_22522# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X241 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X242 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X243 VDPWR sar9b_0.net35 a_3946_26198# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X244 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VDPWR sar9b_0.net54 a_7926_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X246 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X251 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X252 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X255 a_10926_17021# a_10649_17131# a_11256_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X256 a_11915_27039# sar9b_0.net30 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X257 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X258 sar9b_0.net36 a_9996_16784# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X259 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X260 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X261 a_2508_20780# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X262 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X266 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X267 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X268 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X270 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X271 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X272 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X273 a_5481_20185# a_5126_20140# a_5374_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X274 a_11382_18146# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X275 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X276 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X277 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X278 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X280 a_13216_19809# a_12618_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X281 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X282 a_7542_27530# a_7478_27751# a_7464_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X283 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VGND sar9b_0.net45 a_12647_27128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X285 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X286 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X287 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X288 VDPWR a_11030_22954# a_10985_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X289 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X290 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X291 a_11256_16874# a_10858_17113# a_11178_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X292 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X294 VGND sar9b_0.net68 a_3073_24815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X295 a_5289_22527# a_4934_22432# a_5182_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X296 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X297 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X298 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X299 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X301 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X302 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X303 VGND a_13011_24570# single_9b_cdac_1.CF[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X304 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 a_8303_23853# a_8098_23762# a_7638_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X306 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X307 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X308 a_12618_26134# a_11658_26134# a_12182_26419# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X309 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X310 VDPWR a_6579_18832# sar9b_0.net46 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X311 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X312 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A a_50962_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X313 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X316 a_11842_23762# a_11658_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X317 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 a_7464_27530# a_7138_27758# a_7343_27849# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X319 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X320 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X321 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X322 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X323 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X324 VGND sar9b_0.clknet_1_0__leaf_CLK a_4947_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X325 a_12870_19603# a_12618_19474# a_13008_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X326 VDPWR sar9b_0.net59 a_9279_27227# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 single_9b_cdac_0.SW[2] a_13067_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X329 VGND sar9b_0.net63 a_4811_23656# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2695 pd=2.08 as=0.13062 ps=1.025 w=0.55 l=0.15
X330 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X331 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A a_59529_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X332 a_11178_16874# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X333 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X334 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X335 a_3073_24815# sar9b_0._14_ sar9b_0._16_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X336 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X337 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X338 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X339 VGND a_7890_26108# a_7692_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X340 a_9935_24187# a_9730_24138# a_9270_24566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X341 VDPWR a_8595_17910# single_9b_cdac_1.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X342 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X343 VGND a_11776_27801# sar9b_0.net25 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X344 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X345 VDPWR a_10506_24506# a_10758_24459# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X346 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X347 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X348 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X349 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X351 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X352 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X353 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X354 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X355 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X356 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 a_21368_4076# th_dif_sw_0.th_sw_1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X358 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X359 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X360 a_9974_17626# a_9839_17527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X361 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X362 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X363 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X364 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X365 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X366 a_5151_28559# a_5010_28495# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X367 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X368 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X369 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X370 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X371 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X374 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X375 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X376 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDPWR tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X378 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 single_9b_cdac_1.SW[5] a_13011_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X380 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VGND a_7590_24931# a_7548_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X383 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X384 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X385 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X386 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X387 a_9634_17478# a_9450_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X388 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X391 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X392 VGND a_4811_23656# sar9b_0._13_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X393 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X394 a_12870_18271# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X396 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X397 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 a_9174_17906# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X400 VGND a_7347_24160# sar9b_0.net54 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X401 VDPWR a_12588_16784# sar9b_0.net2 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X402 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X403 a_16185_12837# tdc_0.phase_detector_0.pd_out_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X404 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X405 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X406 sar9b_0.net39 a_6540_22112# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X407 VGND a_12870_19603# a_12828_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X408 a_3454_22567# sar9b_0.net67 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X409 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X410 a_5832_27170# a_5506_26802# a_5711_26851# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X411 a_11466_23174# a_10690_22806# a_11030_22954# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X412 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X413 VGND a_8691_28566# uo_out[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X414 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X415 sar9b_0.clk_div_0.COUNT\[0\] a_5938_22378# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X416 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X419 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X420 VDPWR sar9b_0.net7 a_11658_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X421 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X424 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X425 a_11214_25728# a_10937_25582# a_11544_25838# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X426 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X429 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X430 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X433 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X434 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X435 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X436 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X437 a_9942_27470# sar9b_0.net43 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X438 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X440 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X441 a_11146_25483# a_10932_25713# a_10482_25831# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X442 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X445 a_12828_19481# a_11658_19474# a_12618_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X446 a_10926_17021# a_10644_16791# a_11287_17193# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X447 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X448 VGND sar9b_0.net59 a_8118_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X449 VDPWR a_10035_19474# sar9b_0.net48 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X451 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 a_10932_25713# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X453 a_6922_23534# sar9b_0.net10 a_7443_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X454 VGND sar9b_0.net43 a_11859_20574# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X455 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X456 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X457 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[2] a_55773_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X458 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X459 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X460 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VDPWR single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X462 a_11008_17491# a_10410_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X463 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X464 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X465 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X466 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X467 VGND a_5633_20244# a_5651_20547# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X468 a_64331_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X469 a_4330_27170# a_3545_26914# a_3822_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X470 VDPWR a_6880_26815# sar9b_0.net21 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X471 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X472 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X474 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X475 a_10690_22806# a_10506_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X476 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 sar9b_0.net44 a_6307_27584# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X478 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X479 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X480 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X481 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X482 VDPWR a_9974_17626# a_9929_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X483 VDPWR a_10742_27751# a_10697_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X484 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X485 VDPWR a_7890_26108# a_7692_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X486 VDPWR sar9b_0._07_ a_5628_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X487 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDPWR clk a_4332_23043# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X489 a_11382_22142# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X490 a_10607_21189# a_10402_21098# a_9942_20810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X491 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X492 a_13216_23805# a_12618_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X493 a_11287_17193# a_10858_17113# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X494 VDPWR sar9b_0.net44 a_6954_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X495 VDPWR a_5633_20244# a_5588_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X496 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 a_10098_19171# a_10553_18922# a_10502_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X498 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X499 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X500 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X502 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X503 VGND a_8595_17910# single_9b_cdac_1.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X504 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X505 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X507 a_4293_25852# a_4136_25584# a_3855_25792# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1181 ps=1.035 w=0.55 l=0.15
X508 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X509 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X510 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 a_9929_17527# a_9450_17846# a_9839_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X512 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] a_46159_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X515 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X516 VGND sar9b_0.net46 a_7830_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X517 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VDPWR sar9b_0.cyclic_flag_0.FINAL a_8883_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X519 a_10697_27849# a_10218_27466# a_10607_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X520 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X521 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X522 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X523 single_9b_cdac_1.SW[3] a_10803_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X524 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X525 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X526 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X527 a_7978_22202# a_7193_22459# a_7470_22349# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X528 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X531 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 a_9802_26815# a_9593_26914# a_9138_27163# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X533 a_7638_23474# sar9b_0.net11 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X534 a_9472_23805# a_8874_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X535 a_5588_20145# a_4947_20140# a_5481_20185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X536 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X537 a_11380_27885# a_10402_27758# a_11178_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X538 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X539 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X540 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X541 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X542 a_8842_16874# a_8057_17131# a_8334_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X543 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X544 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VGND sar9b_0.net21 a_7539_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X548 VGND a_10528_20155# sar9b_0.net38 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X549 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X550 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X551 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X552 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X553 single_9b_cdac_1.CF[7] a_12435_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X554 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X555 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X557 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X558 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X559 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 a_2940_25096# a_2893_24992# sar9b_0._16_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X561 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X562 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X563 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X564 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X565 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X567 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X568 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X571 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X573 VDPWR single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X574 VDPWR a_4811_23656# sar9b_0._13_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.3346 pd=1.76 as=0.3304 ps=2.83 w=1.12 l=0.15
X575 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X576 VGND a_5196_24776# sar9b_0.net68 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X577 VDPWR a_13011_16810# single_9b_cdac_1.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X578 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X579 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 single_9b_cdac_0.SW[8] a_9323_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X581 sar9b_0.net39 a_6540_22112# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X582 VDPWR sar9b_0.net47 a_6879_22145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X583 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X584 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X586 VDPWR a_10859_26330# single_9b_cdac_0.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X587 a_3180_19448# sar9b_0._09_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X588 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X589 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X590 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X591 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X592 a_8874_23470# a_7914_23470# a_8438_23755# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X593 a_3725_23194# a_3695_23038# a_3647_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X594 a_3273_20185# a_2739_20140# a_3166_20145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X595 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X598 VDPWR a_6534_27123# a_6484_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X599 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X600 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X601 VDPWR a_10182_20463# a_10132_20155# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X602 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X603 VGND a_3819_24136# a_4018_24235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X604 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X606 VDPWR a_8691_28566# uo_out[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X607 a_6738_22112# a_7193_22459# a_7142_22557# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X608 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X609 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A a_45123_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X610 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X611 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X612 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X614 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X615 VGND a_13011_24570# single_9b_cdac_1.CF[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X616 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X618 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X619 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 a_4236_21738# sar9b_0._05_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X621 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X622 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X623 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X624 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X626 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X627 a_11160_19178# a_10762_18823# a_11082_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X628 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X630 a_3539_24543# a_3014_24136# a_3369_24181# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X631 VDPWR sar9b_0.net10 a_11658_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X632 a_10218_21842# a_9258_21842# a_9782_21622# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X633 single_9b_cdac_1.CF[3] a_13011_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X634 a_8303_18859# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X635 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X637 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VDPWR a_12618_18142# a_12870_18271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X639 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X640 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X641 VDPWR a_12435_20806# single_9b_cdac_1.CF[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X642 VDPWR a_9126_23599# a_9076_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X643 single_9b_cdac_0.SW[1] a_13011_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X644 single_9b_cdac_1.SW[7] a_13011_19242# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X645 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X646 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X647 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X649 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X650 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 sar9b_0.net11 a_5484_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X652 sar9b_0._08_ a_4072_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.20905 ps=1.305 w=0.74 l=0.15
X653 a_6484_17491# a_5506_17478# a_6282_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X654 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X655 VGND a_13011_21906# single_9b_cdac_1.CF[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X656 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X657 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X658 a_11776_25137# a_11178_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X659 VDPWR a_9414_23127# a_9364_22819# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X660 sar9b_0.net35 a_7404_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X661 a_8013_23234# sar9b_0.net62 a_7926_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X662 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X663 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X664 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 a_11082_19178# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X666 a_10662_17799# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X667 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X668 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 a_9366_27227# a_9138_27163# a_9279_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X670 a_7284_20787# sar9b_0.net56 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X671 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X673 a_11842_22430# a_11658_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 VDPWR sar9b_0._07_ a_3795_19512# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2478 ps=2.27 w=0.84 l=0.15
X676 a_10194_16784# a_10649_17131# a_10598_17229# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X677 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X678 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X680 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X681 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X682 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X684 VDPWR a_3822_27060# a_3754_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X685 a_11722_25838# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X686 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X687 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X688 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X689 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X690 VGND sar9b_0.net20 a_8115_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X691 a_13008_23477# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X692 VGND a_10470_21795# a_10428_21899# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X693 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 uo_out[6] a_8115_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X695 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X696 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X697 single_9b_cdac_0.SW[0] a_13011_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X698 uo_out[7] a_5235_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X699 a_9138_27163# a_9588_27045# a_9540_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X700 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X701 VGND sar9b_0.clk_div_0.COUNT\[1\] a_3219_22860# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11312 pd=1.065 as=0.15675 ps=1.67 w=0.55 l=0.15
X702 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X703 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X704 VGND sar9b_0.net51 a_9363_20826# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X705 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X708 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X709 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X711 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X712 VGND sar9b_0.net66 sar9b_0._05_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X713 VDPWR sar9b_0.net8 a_8970_20510# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X714 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X716 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X717 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X718 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X719 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X721 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A a_41357_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X722 uio_out[1] a_2931_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X723 a_6744_23238# a_6484_22845# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X724 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X726 VDPWR single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X727 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X728 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VDPWR single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X730 a_10428_21899# a_9258_21842# a_10218_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X731 a_9323_27662# sar9b_0.net34 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X732 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X733 a_8512_27801# a_7914_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X734 VDPWR sar9b_0.net45 a_10218_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X735 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X736 VDPWR sar9b_0.net47 a_7374_19685# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X737 a_8006_18561# a_7743_18149# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X738 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X739 a_10070_24286# a_9935_24187# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X740 a_2892_23070# sar9b_0._18_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X741 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X743 a_5289_22527# a_4755_22138# a_5182_22567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X744 a_4496_20468# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X745 VDPWR a_3156_27447# a_3161_27787# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X746 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X747 a_2892_23070# sar9b_0._18_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X748 VGND a_5394_18116# a_5196_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X749 VDPWR sar9b_0.net49 a_10227_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X750 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X751 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X752 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X753 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X754 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X755 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X756 a_6538_24506# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X757 a_9494_20290# a_9359_20191# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X758 VGND sar9b_0.net48 a_8502_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X759 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X760 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 a_12243_25898# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X763 VDPWR a_3438_27677# a_3370_27769# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X764 sar9b_0.net45 a_8883_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X765 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X767 a_5046_17906# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X768 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X769 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 a_5506_26802# a_5322_27170# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X771 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X773 a_12182_18427# a_12047_18525# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X774 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X777 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X780 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X783 VGND sar9b_0.net37 a_8019_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X784 single_9b_cdac_1.SW[0] a_8595_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X785 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X786 VDPWR sar9b_0.net60 a_6678_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X787 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X788 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X789 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 VDPWR a_13011_20806# single_9b_cdac_1.CF[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X791 single_9b_cdac_1.SW[8] a_11859_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X792 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X793 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X794 a_15265_9613# th_dif_sw_0.VCP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X795 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X797 VDPWR a_12870_26263# a_12820_26553# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X798 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X799 a_8502_19178# a_8438_18958# a_8424_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X800 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X801 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X802 tdc_0.phase_detector_0.INN a_16527_10454# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X803 VDPWR sar9b_0.net58 a_3438_27677# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X804 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X805 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X806 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X807 a_5414_28147# a_5151_28559# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X808 a_10816_21487# a_10218_21842# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X809 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X810 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X811 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X814 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X816 VDPWR a_3372_25734# sar9b_0.net69 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X817 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X819 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X820 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X822 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X823 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X824 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X826 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X827 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X828 a_7138_27758# a_6954_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X829 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X830 single_9b_cdac_0.SW[7] a_10859_26330# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X831 single_9b_cdac_0.SW[6] a_9323_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X832 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X833 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X834 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X835 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X836 a_8386_22806# a_8202_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X837 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X838 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X839 a_8424_19178# a_8098_18810# a_8303_18859# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X841 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X842 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X843 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X844 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X845 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X846 VGND a_11859_20574# single_9b_cdac_1.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X847 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X849 VDPWR tdc_0.OUTP tdc_0.OUTN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X850 uo_out[4] a_8691_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X851 VDPWR a_13011_24570# single_9b_cdac_1.CF[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X852 VDPWR sar9b_0.net47 a_6783_19481# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X853 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X854 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X855 sar9b_0._07_ a_3371_23106# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.4816 pd=3.1 as=0.203 ps=1.505 w=1.12 l=0.15
X856 single_9b_cdac_1.CF[5] a_13011_23238# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X857 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X858 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X859 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X860 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X861 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 a_5846_22572# a_4934_22432# a_5739_22488# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X863 a_12047_18525# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X864 tdc_0.OUTN tdc_0.phase_detector_0.pd_out_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X865 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X867 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X868 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X869 a_6052_19792# sar9b_0._07_ a_5581_19664# VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X870 a_21368_4076# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_18214_3039# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X871 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X872 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X874 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X875 a_8842_18206# sar9b_0.net5 a_9363_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X876 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X877 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X878 a_6642_19448# a_7097_19795# a_7046_19893# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X879 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X880 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X881 a_4330_27170# a_3540_27045# a_3822_27060# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X882 a_5002_23764# sar9b_0.net72 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.3346 ps=1.76 w=0.84 l=0.15
X883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X884 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X885 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X886 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 a_7343_27849# a_6954_27466# a_6678_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X888 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X889 a_5801_17527# a_5322_17846# a_5711_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X890 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X891 sar9b_0.net48 a_10035_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X892 VDPWR sar9b_0.net48 a_6126_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X893 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X896 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X897 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X898 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X899 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X900 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X901 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X902 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X903 VDPWR a_5394_18116# a_5196_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X904 a_21368_4076# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X905 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X906 VDPWR a_5580_24776# sar9b_0._03_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X907 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X908 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X909 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X910 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X912 a_5812_21028# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3685 pd=2.44 as=0.17462 ps=1.185 w=0.55 l=0.15
X913 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X914 a_3994_19474# sar9b_0._07_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.14457 ps=1.15 w=0.74 l=0.15
X915 a_11214_25728# a_10932_25713# a_11575_25519# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X916 a_9363_18146# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X918 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X919 uo_out[7] a_5235_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X920 VGND sar9b_0.net59 a_9366_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X921 a_9782_21622# a_9647_21523# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X922 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X924 sar9b_0._06_ a_12560_27128# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X925 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X926 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X927 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X928 VDPWR a_2603_17006# th_dif_sw_0.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X929 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X930 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X931 VGND sar9b_0.net52 a_8502_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X932 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X933 sar9b_0._15_ a_4467_24162# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X934 sar9b_0.net44 a_6307_27584# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X935 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X936 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X937 VDPWR tdc_0.phase_detector_0.pd_out_0.A a_16185_13034# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X938 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X939 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X940 VGND a_12491_27662# single_9b_cdac_0.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X941 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X942 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X943 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X944 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X945 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X946 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X947 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X948 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X949 a_11575_25519# a_11146_25483# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X950 a_12137_26517# a_11658_26134# a_12047_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X951 a_2508_23444# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X952 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X953 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 a_8502_23534# a_8438_23755# a_8424_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X955 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X956 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X957 a_9076_23889# a_8098_23762# a_8874_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X958 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X959 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X960 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X961 dw_17224_1400# a_18214_3039# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X962 VGND a_13011_21906# single_9b_cdac_1.CF[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X965 a_5711_26851# a_5322_27170# a_5046_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X966 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X967 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X968 a_12182_22423# a_12047_22521# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X969 a_6252_20780# sar9b_0._11_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X970 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X971 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 VGND sar9b_0.net12 a_12435_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X973 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X974 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X975 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X976 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X977 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X979 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X980 a_7590_24931# a_7338_24802# a_7728_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X981 a_6252_20780# sar9b_0._11_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X983 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X984 a_10598_17229# a_10335_16817# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X985 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X986 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X987 a_44418_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X988 a_8424_23534# a_8098_23762# a_8303_23853# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X989 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X990 a_10623_25895# a_10482_25831# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 a_9552_23231# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X993 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X994 a_10985_22855# a_10506_23174# a_10895_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X995 a_6250_28502# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X996 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X997 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X999 VGND sar9b_0.net9 a_10506_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1000 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1001 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1002 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1003 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1004 VDPWR a_9930_20510# a_10182_20463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1005 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1006 VDPWR a_6282_27170# a_6534_27123# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1007 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1008 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1009 VDPWR sar9b_0.net61 a_7978_22202# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1010 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1011 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1012 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1013 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1014 a_5628_19768# a_5581_19664# sar9b_0._10_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X1015 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1016 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1017 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1018 sar9b_0._18_ sar9b_0._17_ a_5183_20819# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1019 a_9138_27163# a_9593_26914# a_9542_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X1020 VGND a_8622_26345# a_8554_26437# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1021 single_9b_cdac_1.SW[4] a_11859_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1022 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1023 a_9935_24187# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1024 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1025 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1026 a_11842_19766# a_11658_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1027 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1028 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1029 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1030 a_12047_22521# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1031 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1033 sar9b_0.net49 a_9363_20826# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X1034 sar9b_0.net6 a_7404_18116# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1035 th_dif_sw_0.VCN ua[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1036 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1037 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1039 a_11030_22954# a_10895_22855# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1040 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1041 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1043 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1044 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1045 a_7540_25221# a_6562_25094# a_7338_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1046 a_5183_20819# sar9b_0.net65 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X1047 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1048 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 a_10742_27751# a_10607_27849# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1050 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1051 a_5581_20992# a_5812_21028# a_5761_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1052 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1055 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1056 VDPWR a_12064_22819# sar9b_0.net30 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1057 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1058 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1060 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1061 a_7402_22441# a_7188_22119# a_6738_22112# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1062 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1063 VGND a_11915_27039# single_9b_cdac_0.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X1064 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1065 VDPWR a_9162_23174# a_9414_23127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1066 sar9b_0._12_ a_5523_21528# a_5765_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3182 pd=2.34 as=0.0888 ps=0.98 w=0.74 l=0.15
X1067 VGND a_12588_16784# sar9b_0.net2 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X1068 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1069 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1070 sar9b_0.net48 a_10035_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1071 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1072 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1074 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1075 a_6771_28562# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1076 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15182 ps=1.125 w=0.55 l=0.15
X1077 VDPWR sar9b_0.net12 a_12435_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1078 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1079 VDPWR sar9b_0.net61 a_8842_16874# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1080 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1081 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1082 VDPWR a_12491_27662# single_9b_cdac_0.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1083 a_3819_24136# a_3014_24136# a_3521_24240# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X1084 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1085 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1086 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1087 VGND a_9323_27662# single_9b_cdac_0.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X1088 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1089 VDPWR sar9b_0.clk_div_0.COUNT\[1\] sar9b_0._17_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3304 ps=2.83 w=1.12 l=0.15
X1090 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1091 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 VDPWR a_10227_18142# th_dif_sw_0.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1093 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1094 a_8622_26345# a_8340_26115# a_8983_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X1095 VDPWR a_4365_25770# a_4293_25852# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.2331 ps=1.395 w=0.84 l=0.15
X1096 VGND sar9b_0.net26 a_13011_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1097 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1098 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1099 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1100 a_3262_24141# sar9b_0.net70 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X1101 a_5765_21842# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.22412 ps=1.365 w=0.74 l=0.15
X1102 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1103 a_7566_21017# a_7284_20787# a_7927_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X1104 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1105 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1106 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1108 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1109 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1110 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1111 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1112 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1113 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1114 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1115 a_6102_24806# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1116 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1117 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1118 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1119 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1120 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1121 VGND sar9b_0.net10 a_13011_23238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1122 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1123 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1124 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1125 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1126 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1127 a_11338_19178# a_10553_18922# a_10830_19068# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1128 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1129 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1130 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1131 VDPWR a_10528_20155# sar9b_0.net38 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1132 a_5443_19074# sar9b_0.net4 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1133 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1134 uo_out[7] a_5235_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1135 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1136 VDPWR a_2706_27440# a_2508_27440# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1137 VGND a_11339_27039# single_9b_cdac_0.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1138 VDPWR a_10662_17799# a_10612_17491# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1139 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1140 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1141 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1142 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1143 a_8781_20570# sar9b_0.net61 a_8694_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1144 a_8266_17113# a_8052_16791# a_7602_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1145 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1146 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1147 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1148 VDPWR a_13216_18477# sar9b_0.net28 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1149 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1150 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1151 a_9846_21842# a_9782_21622# a_9768_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1152 a_7927_21189# a_7498_21109# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X1153 VDPWR a_11430_20935# a_11380_21225# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1154 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1155 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1156 VGND single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1157 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1158 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A a_65367_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1159 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1160 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1161 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1162 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1163 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1164 VDPWR single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1165 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1166 VDPWR sar9b_0.clknet_0_CLK a_2508_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1167 a_4934_22432# a_4755_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X1168 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1169 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1170 a_10859_26330# sar9b_0.net33 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X1171 VDPWR a_8438_23755# a_8393_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1172 a_4583_20468# sar9b_0.net60 a_4496_20468# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X1173 a_7046_19893# a_6783_19481# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1175 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1176 a_11008_17491# a_10410_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1177 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1178 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1179 VGND single_9b_cdac_0.SW[7] a_30012_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1180 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1181 a_5962_24151# a_5748_24381# a_5298_24499# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1182 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1183 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1184 VDPWR sar9b_0.net50 a_11382_18146# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1185 a_9768_21842# a_9442_21474# a_9647_21523# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1186 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1187 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1188 a_5581_20992# sar9b_0._08_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.19322 ps=1.32 w=0.55 l=0.15
X1189 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1190 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1191 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1192 VGND sar9b_0.net54 a_6966_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1194 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1195 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1196 VGND sar9b_0.net10 a_11658_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1197 single_9b_cdac_1.CF[0] a_13011_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1198 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1199 a_3946_26198# sar9b_0.net35 a_4467_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1200 a_8393_23853# a_7914_23470# a_8303_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1201 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1202 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1203 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1204 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1205 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1206 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 VGND sar9b_0.net68 a_2893_24992# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X1208 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1209 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1210 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1211 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1212 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1213 single_9b_cdac_1.CF[2] a_11859_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1214 VGND sar9b_0.net50 a_11469_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1215 a_10378_27170# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X1216 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1217 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1218 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1219 VDPWR sar9b_0.net26 a_13011_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1220 a_11842_23762# a_11658_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1221 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1222 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1223 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1224 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1225 VDPWR a_13067_27662# single_9b_cdac_0.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1226 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1227 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y a_54737_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1228 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1229 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1230 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1231 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1232 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1234 a_4293_25852# a_4125_25958# a_3855_25792# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.1428 ps=1.225 w=0.84 l=0.15
X1235 single_9b_cdac_1.SW[0] a_8595_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1236 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1237 a_4467_26138# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1238 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1239 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1240 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1241 a_9540_27227# a_9279_27227# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1242 a_12182_22423# a_12047_22521# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1243 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1244 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1245 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1246 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1247 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1248 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1249 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1250 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1251 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1252 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1253 VDPWR a_7566_21017# a_7498_21109# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1254 a_11469_19478# sar9b_0.net73 a_11382_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1255 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1256 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1257 VDPWR a_10926_17021# a_10858_17113# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1258 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1259 VGND a_3603_28156# sar9b_0.net59 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1260 VDPWR a_9323_27662# single_9b_cdac_0.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1261 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1262 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1263 VDPWR sar9b_0.net58 a_5151_28559# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1264 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1266 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1267 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1268 a_10470_21795# a_10218_21842# a_10608_21899# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1269 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1270 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1271 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1272 VGND a_11915_27039# single_9b_cdac_0.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1273 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1274 a_3166_20145# sar9b_0._00_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X1275 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1276 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1277 a_9647_21523# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1278 VGND a_7374_19685# a_7306_19777# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1280 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1281 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1282 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1283 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1284 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1285 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1286 a_5046_27230# sar9b_0.net39 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1287 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1288 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1289 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1290 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[1] a_60565_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1291 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1292 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1293 a_10528_20155# a_9930_20510# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1294 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1295 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1296 single_9b_cdac_1.SW[1] a_10803_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1297 VDPWR sar9b_0.net48 a_9174_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1298 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1299 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1300 VGND a_10098_19171# a_9900_19047# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1301 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1302 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1303 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1304 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1305 a_5238_28559# a_5010_28495# a_5151_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1306 VGND a_9323_27662# single_9b_cdac_0.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1307 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1308 a_9942_20810# sar9b_0.net7 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1309 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1310 a_50962_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1311 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1312 VGND a_13011_19242# single_9b_cdac_1.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1313 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1314 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1315 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1316 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1317 sar9b_0.net47 a_7443_21496# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X1318 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A a_36555_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1319 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1320 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1321 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1322 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1323 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1324 VDPWR single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1325 a_35519_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1326 a_11842_18434# a_11658_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1328 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1329 VDPWR single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1330 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1331 VDPWR a_5196_24776# sar9b_0.net68 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1332 VGND sar9b_0.clknet_0_CLK a_2508_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X1333 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1334 VDPWR a_6642_19448# a_6444_19448# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1335 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1336 a_7092_19455# sar9b_0.net10 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1337 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1338 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1339 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1340 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1341 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1342 VGND a_3438_27677# a_3370_27769# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1343 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1344 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1345 single_9b_cdac_0.SW[4] a_11915_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X1346 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1347 VDPWR sar9b_0.net72 sar9b_0._14_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1348 a_6534_17799# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1349 a_8074_20870# a_7289_21127# a_7566_21017# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1350 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VDPWR a_10482_3438# VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X1351 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1352 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1353 VDPWR a_13216_22473# sar9b_0.net31 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1354 VDPWR a_10742_21091# a_10697_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1355 a_11434_16874# a_10649_17131# a_10926_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1356 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1357 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1358 VGND sar9b_0.net44 a_6954_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1359 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1360 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1361 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1362 a_5481_20185# a_4947_20140# a_5374_20145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X1363 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1364 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1365 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1366 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1367 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1368 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1369 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1370 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1371 uio_out[0] a_4083_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1372 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1373 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1374 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1375 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1376 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1377 VDPWR a_11776_25137# sar9b_0.net13 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1378 a_8303_18859# a_7914_19178# a_7638_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1379 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1380 VGND sar9b_0._04_ a_3027_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1381 a_4811_23656# sar9b_0.net63 a_5002_23764# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1134 ps=1.11 w=0.84 l=0.15
X1382 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1383 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1384 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1385 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1387 a_3425_20244# a_3273_20185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X1388 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1389 VDPWR a_6307_27584# sar9b_0.net44 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1390 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1391 a_12820_23889# a_11842_23762# a_12618_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1392 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1393 a_6444_21738# sar9b_0._02_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1394 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1396 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1397 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1398 a_16555_12124# tdc_0.OUTN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1399 VGND sar9b_0.net17 a_2931_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1400 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1401 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1402 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1403 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1404 a_3156_27447# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1405 a_4332_23043# clk VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1406 VDPWR sar9b_0.net53 a_11382_22142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1407 a_10697_21189# a_10218_20806# a_10607_21189# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1408 VGND a_10803_19474# single_9b_cdac_1.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1409 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1410 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1411 uio_out[1] a_2931_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1412 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1413 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1414 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1415 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1416 a_7138_27758# a_6954_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1418 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1419 sar9b_0.net56 a_4771_18260# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X1420 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1421 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1422 sar9b_0.net17 a_2508_26108# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1423 a_3822_27060# a_3545_26914# a_4152_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X1424 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1425 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1426 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1427 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1428 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1429 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1430 VDPWR th_dif_sw_0.th_sw_1.CKB a_18214_3039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X1431 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1432 a_9760_22819# a_9162_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1433 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1434 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1435 sar9b_0.net51 a_5811_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2051 ps=1.52 w=1.12 l=0.15
X1436 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1437 VGND sar9b_0.net46 a_7830_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1438 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1439 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1440 VGND single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1441 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1442 VGND sar9b_0.net53 a_11469_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1443 a_10132_20155# a_9154_20142# a_9930_20510# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1444 VGND a_6126_18353# a_6058_18445# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1445 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1446 VGND a_4011_22488# a_4210_22378# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X1447 a_4812_21738# sar9b_0.clk_div_0.COUNT\[3\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1448 th_dif_sw_0.VCN th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCN VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X1449 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1450 VDPWR sar9b_0.net52 a_7638_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1451 sar9b_0._05_ sar9b_0.net66 a_2828_22432# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X1452 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1453 VGND sar9b_0.net58 a_2934_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1454 VGND single_9b_cdac_0.SW[4] a_44418_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1455 a_7142_22557# a_6879_22145# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1456 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1457 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1458 a_9279_27227# a_9138_27163# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X1459 a_4152_27170# a_3754_26815# a_4074_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1460 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1461 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1462 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1463 a_3747_25724# a_3855_25792# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1229 ps=1.085 w=0.64 l=0.15
X1464 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 a_21368_4076# th_dif_sw_0.th_sw_1.CKB a_18214_3039# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X1466 VDPWR a_12435_24802# single_9b_cdac_1.CF[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1467 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1468 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1469 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] a_31753_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1470 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1471 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1472 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1474 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1475 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1476 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1477 single_9b_cdac_1.SW[6] a_13011_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1478 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1479 a_11469_23474# sar9b_0.net74 a_11382_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1480 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1481 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1483 VDPWR a_5010_28495# a_4812_28371# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1484 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1485 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1486 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11655 ps=1.055 w=0.74 l=0.15
X1487 a_5526_24563# a_5298_24499# a_5439_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1488 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1489 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1490 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1491 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1492 VDPWR a_9323_27662# single_9b_cdac_0.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1493 a_3443_20547# a_2918_20140# a_3273_20185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X1494 VDPWR a_8595_17910# single_9b_cdac_1.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1495 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1496 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1497 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1498 a_8074_20870# a_7284_20787# a_7566_21017# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1499 a_4074_27170# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X1500 a_10134_24506# a_10070_24286# a_10056_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1501 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1502 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1503 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1504 a_13216_18477# a_12618_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1505 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1506 sar9b_0._14_ sar9b_0.net72 a_2637_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1507 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1508 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1509 a_7478_27751# a_7343_27849# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1510 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1511 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1512 VDPWR a_5844_18123# a_5849_18463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1513 VGND sar9b_0.net22 a_8691_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1514 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1515 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1516 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1517 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1518 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1519 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1520 VDPWR a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
X1521 a_55773_15501# single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1522 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y a_49926_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1523 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1524 VDPWR clk a_15151_10456# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X1525 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1526 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1528 VGND a_9126_19131# a_9084_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1529 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1530 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1531 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1532 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1533 a_10056_24506# a_9730_24138# a_9935_24187# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1534 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1535 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1536 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1537 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1538 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1539 a_8303_23853# a_7914_23470# a_7638_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1540 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1541 a_11842_22430# a_11658_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1542 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1543 uo_out[5] a_7539_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1544 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1545 a_11338_19178# a_10548_19053# a_10830_19068# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1546 a_5506_17478# a_5322_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1547 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1549 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1550 VDPWR a_10803_19474# single_9b_cdac_1.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1551 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1552 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1553 VDPWR a_13011_19242# single_9b_cdac_1.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1554 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1555 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1556 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1557 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1558 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1559 single_9b_cdac_1.CF[8] a_13011_25902# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1560 VGND a_6744_23238# a_6861_22828# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11485 pd=1.085 as=0.2436 ps=2 w=0.42 l=0.18
X1561 VDPWR a_9472_18823# sar9b_0.net26 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1562 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1563 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1564 a_6346_23773# a_6132_23451# a_5682_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X1565 VGND a_7470_22349# a_7402_22441# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1566 VDPWR a_11436_17742# sar9b_0.net61 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1567 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1568 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1570 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1571 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1572 a_3976_24520# a_2835_24136# a_3819_24136# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X1573 a_9084_19235# a_7914_19178# a_8874_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1574 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1575 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1576 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1577 a_5394_18116# a_5844_18123# a_5796_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X1578 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1579 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1580 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1581 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1582 VDPWR a_10410_17846# a_10662_17799# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1583 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1584 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1585 a_6250_28502# a_5460_28377# a_5742_28392# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1586 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1587 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1588 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1589 a_12618_26134# a_11842_26426# a_12182_26419# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1590 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1591 a_46159_15501# single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1592 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1593 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1594 a_9935_24187# a_9546_24506# a_9270_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1595 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1596 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1597 a_6767_25185# a_6562_25094# a_6102_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1598 VGND sar9b_0.net8 a_11658_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1599 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1600 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1601 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1602 uo_out[1] a_12531_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1603 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1604 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1605 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1606 a_13216_19809# a_12618_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1607 VGND sar9b_0.net35 a_8595_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1608 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1609 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1611 a_39616_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1612 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1613 a_10420_21487# a_9442_21474# a_10218_21842# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1614 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1615 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1616 a_4211_19474# sar9b_0.net71 a_4072_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=1.55 as=0.20165 ps=1.285 w=0.74 l=0.15
X1617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1618 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1619 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1620 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1621 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1622 VDPWR a_8115_28566# uo_out[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1623 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1624 VDPWR a_13011_24802# single_9b_cdac_0.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1625 a_7188_22119# sar9b_0.net9 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1626 a_5796_18149# a_5535_18149# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1627 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1628 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1629 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.B a_16185_12837# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1630 a_6880_26815# a_6282_27170# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1631 VDPWR sar9b_0.net56 a_10218_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1632 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1633 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1634 a_11776_27801# a_11178_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1635 a_7882_19538# a_7092_19455# a_7374_19685# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1636 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1637 a_9154_20142# a_8970_20510# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1638 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1639 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1640 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1641 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1642 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1643 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1644 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1645 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1646 VGND a_8340_26115# a_8345_26455# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1647 sar9b_0.net57 a_5443_19074# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1648 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1649 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1650 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1651 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1652 a_12182_19759# a_12047_19857# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1653 VGND a_13011_19242# single_9b_cdac_1.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X1654 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1655 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1656 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1657 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1658 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1659 VDPWR clk a_4332_23043# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1660 VDPWR a_10830_19068# a_10762_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1661 VDPWR a_2931_28566# uio_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1662 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1663 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1664 a_4531_25875# a_4293_25852# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1648 ps=1.245 w=0.42 l=0.15
X1665 a_9839_17527# a_9634_17478# a_9174_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1666 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1667 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1668 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1669 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1670 VDPWR a_3540_27045# a_3545_26914# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1671 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1672 a_11178_24802# a_10218_24802# a_10742_25087# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1673 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1675 a_10402_27758# a_10218_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1676 a_11178_20806# a_10402_21098# a_10742_21091# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1677 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1678 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1679 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1680 a_10895_22855# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1681 VDPWR sar9b_0.net46 a_8334_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X1682 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1683 a_3156_27447# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1684 VDPWR a_7602_18116# a_7404_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1685 a_9126_23599# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1686 tdc_0.phase_detector_0.INP a_15151_10456# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X1687 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1688 VDPWR sar9b_0.net62 a_6538_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1689 a_7602_18116# a_8052_18123# a_8004_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X1690 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1691 a_3521_24240# a_3369_24181# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X1692 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1693 VDPWR a_8883_27466# sar9b_0.net45 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1694 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1695 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1696 single_9b_cdac_1.CF[4] a_13011_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1697 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1698 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1699 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1700 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1701 a_8554_26437# a_8345_26455# a_7890_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X1702 a_5580_24776# sar9b_0._15_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1703 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1704 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1705 VGND a_9939_28566# uo_out[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1706 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1707 VGND sar9b_0.clknet_0_CLK a_2508_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X1708 a_11434_16874# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X1709 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1710 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1711 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1712 a_5126_20140# a_4947_20140# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X1713 VGND a_5443_19074# sar9b_0.net57 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1714 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X1715 uo_out[6] a_8115_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1716 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1717 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1718 VDPWR a_3713_22522# a_3668_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X1719 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1720 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1721 a_11382_26138# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1722 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1723 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1724 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1725 a_6879_22145# a_6738_22112# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X1726 ua[3] th_dif_sw_0.th_sw_1.CK ua[3] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X1727 a_13008_18149# sar9b_0.net50 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1728 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1729 a_10402_21098# a_10218_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1730 VGND a_10803_19474# single_9b_cdac_1.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X1731 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1732 VGND sar9b_0.net11 a_13011_24570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X1733 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1734 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1735 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1736 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1737 a_9634_17478# a_9450_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1738 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1739 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1740 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1741 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1742 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1743 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1744 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1745 a_8118_26141# a_7890_26108# a_8031_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1746 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1747 a_41357_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1748 VGND sar9b_0.net54 a_5526_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1749 VDPWR a_11430_27595# a_11380_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1750 VGND a_9472_23805# sar9b_0.net12 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1751 VDPWR a_10859_26330# single_9b_cdac_0.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1752 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1753 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1754 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1755 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1756 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1757 a_3668_22567# a_3027_22138# a_3561_22527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X1758 sar9b_0._04_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1759 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1760 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1761 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1762 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1763 VDPWR a_11859_17910# single_9b_cdac_1.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1764 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1765 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1766 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1767 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1768 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1769 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1770 a_9647_21523# a_9258_21842# a_8982_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1771 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1772 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1773 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1774 a_3713_22522# a_3561_22527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X1775 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1776 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1777 VDPWR a_8691_28566# uo_out[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1778 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1779 VDPWR sar9b_0.net47 a_6975_20813# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1780 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1781 uo_out[5] a_7539_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1782 VDPWR single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1783 VDPWR a_13011_23238# single_9b_cdac_1.CF[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1784 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1785 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1786 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1787 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1788 a_6252_19074# sar9b_0.net15 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1789 a_2828_22432# sar9b_0._12_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X1790 a_6634_18206# a_5844_18123# a_6126_18353# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1792 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1793 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1794 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1795 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1796 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1797 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1798 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1799 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1800 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1801 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1802 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1803 VDPWR a_13164_28398# sar9b_0.net14 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1804 single_9b_cdac_1.SW[2] a_8019_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1805 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1806 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1807 VGND sar9b_0.net53 a_11094_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1808 a_8842_16874# sar9b_0.net61 a_9363_16814# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1809 VDPWR single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1810 a_59529_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1812 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1813 VGND a_3372_25734# sar9b_0.net69 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X1814 VGND sar9b_0.net11 a_11658_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1815 VGND a_4083_28566# uio_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1816 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1817 VDPWR sar9b_0.clknet_1_1__leaf_CLK a_4755_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1819 a_3946_27530# sar9b_0.net36 a_4467_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1820 a_9323_27662# sar9b_0.net34 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X1821 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1822 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1823 VGND single_9b_cdac_0.SW[8] a_25210_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1824 a_13216_23805# a_12618_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1825 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1826 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1827 single_9b_cdac_0.SW[0] a_13011_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1828 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1829 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1830 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1831 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1832 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1833 a_13164_28398# sar9b_0._06_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1834 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1835 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1836 a_7936_25137# a_7338_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1837 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1838 a_12870_26263# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1839 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1840 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1841 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1842 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1843 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1844 a_11722_25838# a_10937_25582# a_11214_25728# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1845 a_11094_23174# a_11030_22954# a_11016_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1846 single_9b_cdac_1.CF[5] a_13011_23238# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X1847 a_9363_16814# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1848 th_dif_sw_0.CKB a_2603_17006# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1849 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1850 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1851 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1852 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1853 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1854 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1856 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1857 a_4467_27470# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1858 a_8983_26517# a_8554_26437# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X1859 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1860 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1861 a_12182_23755# a_12047_23853# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1862 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1863 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1864 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1865 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1867 VDPWR sar9b_0.net12 a_11658_26134# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1868 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1869 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1870 a_10607_27849# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1871 VDPWR a_6534_17799# a_6484_17491# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1872 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1874 VDPWR a_5682_23444# a_5484_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1875 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1876 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1877 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1878 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1879 VDPWR sar9b_0.net59 a_9942_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1880 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1881 VDPWR a_3723_20140# a_3922_20239# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X1882 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1883 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1884 sar9b_0.net63 a_6861_22828# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.11485 ps=1.085 w=0.74 l=0.15
X1885 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1886 VDPWR sar9b_0.net36 a_10803_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1887 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1888 a_11030_22954# a_10895_22855# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1889 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1890 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1891 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1892 VGND sar9b_0.net58 a_3318_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X1893 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1894 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1895 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1896 a_12064_22819# a_11466_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1897 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1898 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1899 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1900 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1901 a_9542_26815# a_9279_27227# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1902 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1903 a_5812_21028# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2898 ps=2.37 w=0.84 l=0.15
X1904 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1905 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1906 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1907 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[2] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1908 sar9b_0._11_ a_4496_20468# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X1909 VGND a_7092_19455# a_7097_19795# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1910 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1911 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1912 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1913 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1914 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1915 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1916 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1917 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1918 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1919 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1920 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1921 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1922 VGND a_11104_24151# sar9b_0.net42 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1923 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1924 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1925 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1926 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1927 sar9b_0.net34 a_10284_25707# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X1928 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1929 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1930 a_5910_23477# a_5682_23444# a_5823_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1931 a_13008_22145# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1932 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1933 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1935 VDPWR sar9b_0.net52 a_10623_25895# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1936 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1937 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1938 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1939 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1940 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1941 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1942 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1943 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1944 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1945 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1946 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1947 VDPWR sar9b_0.net18 a_4083_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1948 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1949 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1950 VDPWR sar9b_0.net61 a_11434_16874# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1952 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1953 VDPWR sar9b_0.net38 a_6250_28502# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1954 a_6966_24866# a_6902_25087# a_6888_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1955 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1956 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1957 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1958 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1959 VDPWR a_8340_26115# a_8345_26455# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1960 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1961 a_7236_20813# a_6975_20813# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1962 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1964 sar9b_0.net58 a_4749_27652# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1965 VDPWR a_11859_21906# single_9b_cdac_1.CF[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1966 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1967 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1968 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1969 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1970 VGND a_3156_27447# a_3161_27787# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1971 VGND tdc_0.RDY a_5331_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1972 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1973 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1974 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1975 VDPWR a_8622_26345# a_8554_26437# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1976 a_5711_26851# a_5506_26802# a_5046_27230# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1977 VDPWR a_11859_17910# single_9b_cdac_1.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1978 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1979 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1980 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X1981 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1982 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1983 a_5133_27230# sar9b_0.net39 a_5046_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1984 a_10742_21091# a_10607_21189# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1985 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1986 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1987 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1988 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1989 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1990 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1991 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1992 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1993 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1994 VDPWR a_3156_26115# a_3161_26455# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1995 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1996 a_3723_20140# a_2918_20140# a_3425_20244# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X1997 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1998 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1999 a_6888_24866# a_6562_25094# a_6767_25185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2000 VDPWR a_9363_20826# sar9b_0.net49 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X2001 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2002 a_10482_25831# a_10932_25713# a_10884_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2003 single_9b_cdac_1.CF[7] a_12435_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2004 VGND sar9b_0.net50 a_12246_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2005 sar9b_0.net35 a_7404_16784# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2006 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2007 VDPWR a_3438_26345# a_3370_26437# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2008 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2009 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2010 VDPWR sar9b_0.net59 a_8622_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2011 a_4467_24162# sar9b_0._13_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X2012 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2013 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2014 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2015 a_5010_28495# a_5465_28246# a_5414_28147# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2016 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2017 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2018 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2019 a_54032_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2020 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2021 sar9b_0.net53 a_10227_23490# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2022 a_3370_27769# a_3161_27787# a_2706_27440# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2023 VGND sar9b_0.net59 a_10806_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2024 a_5742_28392# a_5460_28377# a_6103_28183# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2025 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2026 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2027 a_9782_21622# a_9647_21523# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X2028 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2030 VGND a_12531_28566# uo_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2031 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2032 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2033 VDPWR sar9b_0.net59 a_3438_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2034 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2035 a_8591_22855# a_8386_22806# a_7926_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2036 single_9b_cdac_0.SW[3] a_12491_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2037 a_10884_25895# a_10623_25895# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2038 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2039 single_9b_cdac_0.SW[1] a_13011_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2040 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2041 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2042 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2043 VDPWR a_2706_26108# a_2508_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2044 a_5931_20140# a_4947_20140# a_5633_20244# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X2045 VDPWR sar9b_0.net41 a_13011_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2046 a_10422_16817# a_10194_16784# a_10335_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2047 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2048 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2049 VGND a_5739_22488# a_5938_22378# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X2050 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2051 a_9130_26198# a_8345_26455# a_8622_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X2052 VGND a_11859_21906# single_9b_cdac_1.CF[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2053 th_dif_sw_0.CK a_10227_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2055 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2056 th_dif_sw_0.CKB a_2603_17006# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2057 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2058 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2059 a_6103_28183# a_5674_28147# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2060 a_10806_27530# a_10742_27751# a_10728_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2061 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2062 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2063 VDPWR sar9b_0.net54 a_6102_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2064 VDPWR sar9b_0.net65 a_5083_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X2065 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2066 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2067 VDPWR sar9b_0.net47 a_6052_19792# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X2068 VDPWR a_12618_26134# a_12870_26263# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2069 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A a_54737_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2070 a_8304_27473# sar9b_0.net60 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2071 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2072 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2074 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2075 a_45123_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2076 VGND single_9b_cdac_0.SW[5] a_39616_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2077 VGND sar9b_0.net9 a_13011_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X2078 a_3180_19448# sar9b_0._09_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2079 VDPWR a_5196_19448# sar9b_0.net71 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2080 VGND a_10830_19068# a_10762_18823# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2081 VDPWR a_5235_27466# uo_out[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2082 a_7374_19685# a_7092_19455# a_7735_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2083 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2084 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2086 VGND a_10816_21487# sar9b_0.net9 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2087 a_9930_20510# a_9154_20142# a_9494_20290# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2088 a_5910_17846# a_5846_17626# a_5832_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2089 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2090 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2091 a_5374_20145# sar9b_0._01_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X2092 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2093 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2094 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2095 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2096 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2097 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2098 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2099 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[8] a_26951_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2100 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2101 a_10728_27530# a_10402_27758# a_10607_27849# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2102 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2103 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2104 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2105 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2106 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2107 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2108 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2109 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2110 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2111 a_7478_27751# a_7343_27849# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2112 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2113 a_5700_24563# a_5439_24563# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2114 a_6058_18445# a_5849_18463# a_5394_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2115 VGND th_dif_sw_0.th_sw_1.CK a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X2116 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2117 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2118 a_10830_19068# a_10553_18922# a_11160_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2119 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2120 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2121 a_2508_23444# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2122 VGND sar9b_0.net56 a_5322_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2123 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2124 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2125 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2126 a_10548_19053# sar9b_0.net7 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2127 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2128 a_15400_11316# tdc_0.phase_detector_0.INP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X2129 VGND a_4083_28566# uio_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2130 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2131 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2132 a_10816_21487# a_10218_21842# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2133 VGND clk a_4332_23043# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X2134 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2135 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2136 a_3438_27677# a_3156_27447# a_3799_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2137 VGND a_8883_27466# sar9b_0.net45 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2138 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2139 a_12246_26198# a_12182_26419# a_12168_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2140 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2141 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2142 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2143 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2144 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2145 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2146 a_5742_28392# a_5465_28246# a_6072_28502# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2147 a_9130_26198# a_8340_26115# a_8622_26345# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2148 a_6922_23534# a_6132_23451# a_6414_23681# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2149 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2150 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2151 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2152 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2153 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2154 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2155 a_35519_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2156 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2157 VDPWR sar9b_0.net25 a_12531_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2158 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2159 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2160 a_5846_17626# a_5711_17527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2161 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2162 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2163 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2164 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2165 VDPWR a_6744_23238# a_6861_22828# VDPWR sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.475 as=0.51 ps=3.02 w=1 l=0.25
X2166 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2167 VGND sar9b_0.net54 a_5910_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2168 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2169 a_10182_20463# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2170 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2171 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2172 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2173 a_10620_17903# a_9450_17846# a_10410_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2175 a_3799_27849# a_3370_27769# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2176 a_11339_27039# sar9b_0.net31 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X2177 VDPWR sar9b_0.net42 a_10378_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X2178 VDPWR a_11859_21906# single_9b_cdac_1.CF[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2180 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2182 a_2940_25096# sar9b_0.net68 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X2183 VGND a_7188_22119# a_7193_22459# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2185 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2186 a_12168_26198# a_11842_26426# a_12047_26517# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2187 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2188 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2189 a_6072_28502# a_5674_28147# a_5994_28502# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2190 single_9b_cdac_0.SW[2] a_13067_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2191 VDPWR a_7338_24802# a_7590_24931# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2192 a_5633_20244# a_5481_20185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X2193 a_5844_18123# sar9b_0.net6 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2194 VGND sar9b_0.net48 a_10038_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2195 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2196 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2197 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2198 a_7374_19685# a_7097_19795# a_7704_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2199 th_dif_sw_0.CKB a_2603_17006# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X2200 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2201 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2202 a_65367_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2203 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2204 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2205 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2206 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2207 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2208 sar9b_0.net43 a_5100_24375# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2210 VDPWR a_9870_27060# a_9802_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2211 a_12182_26419# a_12047_26517# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X2212 VGND sar9b_0.net53 a_12246_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2213 VDPWR a_4011_22488# a_4210_22378# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2214 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2215 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2216 VGND single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2217 VDPWR a_9939_28566# uo_out[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2218 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2219 single_9b_cdac_1.CF[7] a_12435_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2220 a_11430_20935# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2221 sar9b_0.net16 a_3922_20239# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X2222 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2223 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2224 VDPWR th_dif_sw_0.CKB a_21177_7457# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2225 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2226 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2227 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2228 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2229 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2230 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2231 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2232 a_2603_17006# sar9b_0.net16 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2235 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2236 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2237 uo_out[4] a_8691_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2238 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2239 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2240 a_5711_17527# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2241 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2242 VDPWR a_7092_19455# a_7097_19795# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2243 a_6126_18353# a_5844_18123# a_6487_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2244 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2245 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2246 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2247 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2248 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2249 a_7704_19538# a_7306_19777# a_7626_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2250 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2251 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2252 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2253 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2254 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2255 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2256 VDPWR a_7374_19685# a_7306_19777# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2257 VGND a_8334_18353# a_8266_18445# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2258 single_9b_cdac_1.SW[5] a_13011_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2259 VGND single_9b_cdac_0.SW[2] a_54032_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2260 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2261 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2262 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2263 VGND clk a_15197_10290# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X2264 VGND a_12064_22819# sar9b_0.net30 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2266 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2267 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2268 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2269 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2270 VDPWR sar9b_0.net9 a_13011_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2271 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2272 VGND a_2603_17006# th_dif_sw_0.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2273 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2274 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2275 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2276 sar9b_0.net23 a_7692_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X2277 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2278 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2279 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2280 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2281 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2282 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2283 a_6487_18525# a_6058_18445# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2284 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2286 VGND a_13011_17910# single_9b_cdac_1.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2287 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2288 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2289 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2290 VDPWR a_7443_21496# sar9b_0.net47 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X2291 a_7626_19538# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2292 VDPWR a_12182_19759# a_12137_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2293 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2294 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2295 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2296 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2297 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2298 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2299 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2300 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2301 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2302 a_7728_24809# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2303 a_2508_23444# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X2304 a_7483_23174# sar9b_0.clk_div_0.COUNT\[1\] sar9b_0._17_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X2305 VGND sar9b_0.net56 a_10218_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2306 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2307 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2308 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2309 a_10506_24506# a_9546_24506# a_10070_24286# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2310 a_8052_18123# sar9b_0.net56 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2311 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2312 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2313 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2314 a_11842_18434# a_11658_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2315 VDPWR sar9b_0.net39 a_11859_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2316 VGND sar9b_0.net48 a_10422_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2317 VGND single_9b_cdac_1.SW[7] a_30012_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2318 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2319 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2320 VGND sar9b_0.net56 a_9450_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2321 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2322 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2323 a_12047_26517# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2324 a_5651_20547# a_5126_20140# a_5481_20185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X2325 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2326 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y a_30717_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2327 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2328 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2329 a_6282_27170# a_5506_26802# a_5846_26950# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2330 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2331 VDPWR sar9b_0.clk_div_0.COUNT\[1\] a_3219_22860# VDPWR sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X2332 VDPWR a_6282_17846# a_6534_17799# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2333 a_9960_17846# a_9634_17478# a_9839_17527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2334 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2335 a_15197_10290# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_15151_10456# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X2336 a_13008_19481# sar9b_0.net50 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2337 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2338 a_7890_26108# a_8340_26115# a_8292_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2339 VDPWR a_5441_22522# a_5396_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X2340 VDPWR sar9b_0.net51 a_6579_18832# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X2341 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2342 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2344 VDPWR a_4083_28566# uio_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2345 a_7404_17715# sar9b_0.net1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2051 ps=1.52 w=0.84 l=0.15
X2346 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2347 a_8166_27595# a_7914_27466# a_8304_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X2348 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2349 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2350 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2352 a_6538_24506# sar9b_0.net62 a_7059_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2353 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2354 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2355 single_9b_cdac_1.CF[2] a_11859_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2356 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2357 a_6307_27584# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X2358 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2359 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2360 dw_12589_1395# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VDPWR dw_12589_1395# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X2361 a_6126_18353# a_5849_18463# a_6456_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2362 a_8694_20570# sar9b_0.net61 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2363 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2364 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2365 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2366 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2367 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2368 a_8292_26141# a_8031_26141# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2369 VGND a_10758_24459# a_10716_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2370 a_7830_18149# a_7602_18116# a_7743_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2371 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2373 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2374 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2375 VGND a_12531_28566# uo_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2376 a_5396_22567# a_4755_22138# a_5289_22527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X2377 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A a_49926_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2378 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2380 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2381 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2382 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2383 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2384 VGND th_dif_sw_0.th_sw_1.CK a_10482_3438# VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X2385 a_36555_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2387 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2388 VGND a_3713_22522# a_3731_22165# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X2389 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2390 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2391 a_9162_23174# a_8386_22806# a_8726_22954# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2392 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2393 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2394 a_7059_24566# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2395 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2396 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2397 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2398 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2399 a_3713_22522# a_3561_22527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2400 sar9b_0.net46 a_6579_18832# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2401 sar9b_0.net4 a_5331_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2402 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2403 a_6456_18206# a_6058_18445# a_6378_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2404 VDPWR a_5846_17626# a_5801_17527# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2405 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2406 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2407 VDPWR a_6126_18353# a_6058_18445# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2408 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2410 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2411 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2412 a_10716_24563# a_9546_24506# a_10506_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2413 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2414 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2415 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2416 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2417 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2418 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2419 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2420 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2421 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2423 a_60565_15501# single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2424 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2425 single_9b_cdac_1.CF[7] a_12435_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2426 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2427 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2428 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2429 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2430 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2431 a_12491_27662# sar9b_0.net29 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2432 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2433 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2434 a_8004_18149# a_7743_18149# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2435 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2436 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2437 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2438 a_6378_18206# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2439 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2440 VDPWR a_13011_17910# single_9b_cdac_1.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2441 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2442 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2443 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2444 single_9b_cdac_1.CF[6] a_13011_24570# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2445 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2446 VDPWR a_2547_28132# sar9b_0.net60 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2447 a_7638_19238# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2448 VGND a_16159_13315# tdc_0.RDY VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X2449 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2450 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X2451 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2454 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2455 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2456 single_9b_cdac_0.SW[8] a_9323_27662# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2457 a_6282_27170# a_5322_27170# a_5846_26950# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2458 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2459 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2460 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2461 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2462 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2463 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2464 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2465 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2467 a_4365_25770# a_4125_25958# a_4588_25473# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.0504 ps=0.66 w=0.42 l=0.15
X2468 VDPWR sar9b_0.net59 a_9870_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2469 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2470 VDPWR sar9b_0.net51 a_7443_21496# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X2471 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2472 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2473 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2474 VGND a_13216_22473# sar9b_0.net31 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2475 a_5844_18123# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2476 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2477 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2478 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2479 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2480 a_4771_18260# sar9b_0.net57 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2481 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2483 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2484 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2485 VGND sar9b_0.net1 a_10707_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2486 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2487 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2488 a_3880_20524# a_2739_20140# a_3723_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X2489 a_24332_16877# single_9b_cdac_1.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2490 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2491 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2492 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2493 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2494 sar9b_0.net20 a_4812_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2495 a_3369_24181# a_2835_24136# a_3262_24141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X2496 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2497 sar9b_0._10_ a_5581_19664# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X2498 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2499 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2500 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2501 a_4588_25473# a_4293_25852# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.18985 ps=1.545 w=0.42 l=0.15
X2502 VDPWR a_12182_23755# a_12137_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2503 single_9b_cdac_1.SW[8] a_11859_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2504 VGND sar9b_0.net50 a_11469_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2505 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2506 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2507 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2508 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2509 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2510 a_6391_24187# a_5962_24151# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2511 VDPWR a_6902_25087# a_6857_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2512 a_6834_20780# a_7289_21127# a_7238_21225# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2513 VGND a_7404_17715# sar9b_0.net73 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X2514 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2515 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2516 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2517 a_7548_24809# a_6378_24802# a_7338_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2518 VGND a_8940_24402# sar9b_0.net62 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2519 VDPWR sar9b_0.net7 a_11859_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2520 single_9b_cdac_1.SW[1] a_10803_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2521 VGND tdc_0.OUTN a_6867_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2522 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2523 a_9162_23174# a_8202_23174# a_8726_22954# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2524 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2525 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2526 a_6307_27584# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2527 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2528 VGND a_10227_18142# th_dif_sw_0.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2529 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2530 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2531 sar9b_0._14_ sar9b_0.net63 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2532 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2533 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2534 sar9b_0.net52 a_9165_24988# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2535 VGND a_11776_25137# sar9b_0.net13 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2536 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2537 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2538 a_15052_11404# tdc_0.phase_detector_0.INN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X2539 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2540 VGND single_9b_cdac_0.SW[3] a_49221_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2541 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2542 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2543 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2544 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2545 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2546 sar9b_0.net16 a_3922_20239# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X2547 a_11469_18146# sar9b_0.net73 a_11382_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2550 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2551 VDPWR sar9b_0.net9 a_10506_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2552 a_11776_21141# a_11178_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2553 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2554 a_6857_25185# a_6378_24802# a_6767_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2555 VDPWR a_11104_24151# sar9b_0.net42 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2556 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2557 VDPWR a_12531_28566# uo_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2558 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2559 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2560 a_11544_25838# a_11146_25483# a_11466_25838# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2561 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2562 VDPWR clk a_16527_10454# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X2563 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2564 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2565 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2566 a_11178_27466# a_10402_27758# a_10742_27751# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2567 a_6767_25185# a_6378_24802# a_6102_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2568 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2569 VGND single_9b_cdac_1.SW[4] a_44418_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2570 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2571 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2572 VGND a_6252_19074# sar9b_0.net55 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2573 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2574 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2575 VGND tdc_0.phase_detector_0.pd_out_0.B a_16159_13315# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X2576 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2577 single_9b_cdac_0.SW[0] a_13011_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2578 sar9b_0.net47 a_7443_21496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2579 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2580 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2581 VGND sar9b_0.net47 a_5581_19664# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X2582 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2583 a_13067_27662# sar9b_0.net28 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2584 a_10402_21098# a_10218_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2585 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2586 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2587 a_9942_24806# sar9b_0.net12 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2588 a_7443_23474# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2589 sar9b_0.net74 a_10707_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2590 VGND sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X2591 single_9b_cdac_1.SW[3] a_10803_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2592 a_31753_15501# single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2593 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2594 a_3425_20244# a_3273_20185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2595 a_8842_18206# a_8052_18123# a_8334_18353# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X2596 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2597 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2598 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2599 a_11016_23174# a_10690_22806# a_10895_22855# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2600 VDPWR a_5443_19074# sar9b_0.net57 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2601 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2602 a_6642_19448# a_7092_19455# a_7044_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2603 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2604 a_3747_25724# a_3855_25792# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1862 ps=1.475 w=0.84 l=0.15
X2605 VGND a_9165_24988# sar9b_0.net52 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X2606 a_8303_23853# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2607 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2608 a_11466_25838# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2609 a_3754_26815# a_3540_27045# a_3090_27163# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2610 VGND a_13011_17910# single_9b_cdac_1.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2611 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2612 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2613 a_16222_11316# tdc_0.phase_detector_0.INN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X2614 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2615 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2616 a_6250_28502# sar9b_0.net38 a_6771_28562# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2617 a_3540_27045# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2618 VDPWR single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2619 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2620 a_10608_21899# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2621 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2622 a_6880_17491# a_6282_17846# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2623 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2624 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2625 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2626 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2627 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2628 VDPWR sar9b_0.net27 a_13011_27234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2629 a_3819_24136# a_2835_24136# a_3521_24240# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X2630 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2631 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2632 VDPWR a_9138_27163# a_8940_27039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2633 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2634 a_10402_27758# a_10218_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2635 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2636 VGND a_3438_26345# a_3370_26437# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2637 VDPWR a_13216_26469# sar9b_0.net33 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2638 sar9b_0.net51 a_5811_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15198 ps=1.17 w=0.74 l=0.15
X2639 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2640 a_5439_24563# a_5298_24499# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2641 VDPWR a_8874_23470# a_9126_23599# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X2642 VGND a_12435_20806# single_9b_cdac_1.CF[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2643 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2644 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2645 a_6360_24506# a_5962_24151# a_6282_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2646 VGND sar9b_0.net49 a_10806_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2647 a_3690_27530# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2648 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2649 VDPWR a_12870_23599# a_12820_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2650 a_59529_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2651 VGND a_13067_27662# single_9b_cdac_0.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2652 a_7602_16784# a_8052_16791# a_8004_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2653 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2654 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2655 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2656 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2657 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2658 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2659 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2660 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2661 VDPWR a_13011_21906# single_9b_cdac_1.CF[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2662 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2663 a_2706_27440# a_3156_27447# a_3108_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2664 a_2508_20780# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X2665 VDPWR a_10548_19053# a_10553_18922# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2666 single_9b_cdac_1.SW[0] a_8595_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2667 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2668 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2670 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2671 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2672 VDPWR sar9b_0.net54 a_6030_24396# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2673 a_11434_16874# sar9b_0.net61 a_11955_16814# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2674 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2675 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2676 VDPWR sar9b_0.net3 a_2547_28132# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X2677 a_12820_22557# a_11842_22430# a_12618_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X2678 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2679 VDPWR sar9b_0.net52 a_11382_26138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2680 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2681 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2682 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2683 a_10482_25831# a_10937_25582# a_10886_25483# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2684 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2685 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2686 a_3156_26115# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2687 a_6282_24506# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2688 VGND a_10803_18142# single_9b_cdac_1.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2689 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2690 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2691 th_dif_sw_0.VCN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X2692 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2693 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2694 a_10806_20870# a_10742_21091# a_10728_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2695 a_7882_19538# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X2696 a_10607_27849# a_10218_27466# a_9942_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2697 VGND sar9b_0.net49 a_8781_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2698 VDPWR a_5931_20140# a_6130_20239# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2699 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2700 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2701 VDPWR a_4236_21738# sar9b_0.net67 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2702 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2703 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2704 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2705 a_12588_16784# tdc_0.OUTP VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2707 a_3108_27473# a_2847_27473# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2708 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2709 sar9b_0.net27 a_5196_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X2710 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2711 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2712 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2713 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2714 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2715 VGND a_6642_19448# a_6444_19448# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2716 a_9472_18823# a_8874_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2717 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2718 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2719 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X2720 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2721 VGND a_10548_19053# a_10553_18922# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2722 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2723 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2724 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2725 a_7498_21109# a_7284_20787# a_6834_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2726 VGND sar9b_0.net53 a_11469_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2727 a_10728_20870# a_10402_21098# a_10607_21189# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2728 a_10858_17113# a_10644_16791# a_10194_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2729 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2730 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2731 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2732 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2733 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2734 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2735 a_3371_23106# sar9b_0.clk_div_0.COUNT\[2\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X2736 VDPWR a_10816_21487# sar9b_0.net9 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2737 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2738 VGND sar9b_0.net59 a_2934_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2739 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2741 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2742 a_8622_26345# a_8345_26455# a_8952_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2743 a_3647_23194# a_3219_22860# a_3371_23106# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X2744 a_6414_23681# a_6137_23791# a_6744_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2746 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2747 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2748 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2749 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2750 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2751 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2752 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2753 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2754 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2755 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2756 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2757 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2758 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2759 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# a_16357_9613# VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X2760 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2761 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2762 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2763 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2764 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2765 sar9b_0.clk_div_0.COUNT\[3\] a_4210_22378# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X2766 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2767 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2768 a_11469_22142# sar9b_0.net73 a_11382_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2769 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2770 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2771 VGND a_2706_27440# a_2508_27440# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2772 VDPWR a_7478_27751# a_7433_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2773 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2774 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2775 VGND sar9b_0.net49 a_9069_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2776 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCP VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X2777 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2778 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2779 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2780 a_12047_26517# a_11658_26134# a_11382_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2781 a_4934_22432# a_4755_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2782 VGND a_5844_18123# a_5849_18463# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2783 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2784 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2785 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2786 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2787 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2788 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2789 VDPWR sar9b_0.net4 a_6378_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2790 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X2791 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2792 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2793 a_7566_21017# a_7289_21127# a_7896_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2794 a_10607_21189# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2795 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2796 VGND a_13011_20806# single_9b_cdac_1.CF[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2797 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2798 VGND sar9b_0.net42 a_13011_19242# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X2799 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2800 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2801 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2802 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2803 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2804 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2805 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2806 a_2893_24992# sar9b_0._14_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X2807 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2808 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2809 a_7936_25137# a_7338_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2810 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2812 VDPWR sar9b_0.net49 a_9942_20810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2814 VGND a_13011_27234# single_9b_cdac_0.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2815 VDPWR a_2603_17006# th_dif_sw_0.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2816 a_9069_21902# sar9b_0.net8 a_8982_21902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2817 single_9b_cdac_1.CF[4] a_13011_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X2818 a_5931_20140# a_5126_20140# a_5633_20244# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X2819 VDPWR sar9b_0.net12 a_9546_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2820 a_2918_20140# a_2739_20140# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2821 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2822 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2823 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2824 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2825 a_11430_27595# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2826 a_7338_24802# a_6562_25094# a_6902_25087# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2827 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2828 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2829 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2830 a_11842_26426# a_11658_26134# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2831 VGND a_12491_27662# single_9b_cdac_0.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X2832 a_7896_20870# a_7498_21109# a_7818_20870# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2833 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2834 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2835 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2836 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2837 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2838 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2839 a_3014_24136# a_2835_24136# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X2840 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2841 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2842 VDPWR a_5739_22488# a_5938_22378# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X2843 VDPWR a_3795_19512# a_4292_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2557 pd=1.59 as=0.21 ps=1.42 w=1 l=0.15
X2844 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2845 VDPWR a_10803_18142# single_9b_cdac_1.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2846 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2847 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2848 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2849 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2850 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2851 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2852 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2853 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X2854 VGND a_10227_18142# th_dif_sw_0.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2856 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2857 VGND single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2858 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2859 VGND a_13216_19809# sar9b_0.net29 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2860 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2861 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2862 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2863 VDPWR a_10470_21795# a_10420_21487# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2864 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2865 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2866 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2867 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2868 a_7818_20870# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2869 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2870 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2871 VGND a_6534_17799# a_6492_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2872 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2873 VGND a_8052_18123# a_8057_18463# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2874 VGND sar9b_0.net7 a_11658_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2875 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2876 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2877 a_6562_25094# a_6378_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2878 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2879 sar9b_0.net54 a_7347_24160# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X2880 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2882 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2883 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2884 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2885 a_9839_17527# a_9450_17846# a_9174_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2886 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2887 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2888 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2889 VDPWR single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2890 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2891 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2892 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2893 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2895 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2896 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2897 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2898 sar9b_0.net53 a_10227_23490# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X2899 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2900 a_8940_24402# sar9b_0.net2 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2901 VDPWR sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# VDPWR sky130_fd_pr__pfet_01v8 ad=0.27625 pd=1.625 as=0.1176 ps=1.4 w=0.42 l=0.15
X2902 VDPWR tdc_0.OUTN a_6867_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2903 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2904 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2905 a_5126_20140# a_4947_20140# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2906 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2907 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2908 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2909 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2910 a_6492_17903# a_5322_17846# a_6282_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2911 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2912 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2913 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2914 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2915 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2916 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2918 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2919 a_12182_18427# a_12047_18525# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2920 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2921 a_45123_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2922 a_8266_18445# a_8057_18463# a_7602_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2923 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2924 a_5801_26851# a_5322_27170# a_5711_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2925 a_9839_17527# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2926 single_9b_cdac_1.SW[4] a_11859_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2927 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2928 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2929 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2930 VGND single_9b_cdac_1.SW[8] a_25210_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2931 VDPWR sar9b_0.net58 a_5742_28392# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2932 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y a_25915_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2933 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2934 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2935 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2936 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2937 VGND sar9b_0.net63 sar9b_0._02_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2938 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2939 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2940 a_3156_26115# sar9b_0.net44 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2941 a_6975_20813# a_6834_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2942 VDPWR a_7602_16784# a_7404_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2943 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2944 a_5994_28502# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2945 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2946 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2947 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2948 VGND a_12435_20806# single_9b_cdac_1.CF[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2949 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2950 single_9b_cdac_0.SW[8] a_9323_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X2951 VGND a_9126_23599# a_9084_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2952 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2953 VGND a_3822_27060# a_3754_26815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2954 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2955 single_9b_cdac_1.CF[8] a_13011_25902# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2956 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2957 VDPWR sar9b_0._14_ a_4467_24162# VDPWR sky130_fd_pr__pfet_01v8 ad=0.36323 pd=1.84 as=0.126 ps=1.14 w=0.84 l=0.15
X2958 single_9b_cdac_1.CF[0] a_13011_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2959 VGND single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2960 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2961 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2962 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2963 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2964 VDPWR sar9b_0.net57 a_9258_21842# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2965 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2966 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X2967 a_6250_28502# a_5465_28246# a_5742_28392# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X2968 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X2969 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2970 a_13216_26469# a_12618_26134# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2971 VDPWR a_5523_21528# sar9b_0._12_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.196 ps=1.47 w=1.12 l=0.15
X2972 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2973 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2974 a_8681_22855# a_8202_23174# a_8591_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2975 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2976 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2977 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2978 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2979 VGND a_10803_18142# single_9b_cdac_1.SW[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2980 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2981 VDPWR a_12491_27662# single_9b_cdac_0.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2982 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2983 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2984 a_10886_25483# a_10623_25895# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X2985 a_9084_23477# a_7914_23470# a_8874_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2986 a_5441_22522# a_5289_22527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2987 sar9b_0.net70 a_3027_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2988 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2989 VDPWR a_13011_27234# single_9b_cdac_0.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2990 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2992 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2993 a_3540_27045# sar9b_0.net44 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2994 a_25210_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2995 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2996 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2997 VDPWR a_10227_18142# th_dif_sw_0.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2999 a_9154_20142# a_8970_20510# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3000 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3001 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3002 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3003 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3004 a_4811_23656# sar9b_0.net72 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.13062 pd=1.025 as=0.15198 ps=1.17 w=0.55 l=0.15
X3005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3006 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3007 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3008 a_12870_26263# a_12618_26134# a_13008_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3009 ua[4] th_dif_sw_0.th_sw_1.CK ua[4] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X3010 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3011 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3012 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3013 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3014 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3015 a_11380_25221# a_10402_25094# a_11178_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3016 a_7882_19538# a_7097_19795# a_7374_19685# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3017 a_8334_18353# a_8052_18123# a_8695_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3018 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3019 a_10742_21091# a_10607_21189# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3020 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3021 VGND a_11339_27039# single_9b_cdac_0.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X3022 a_12820_19893# a_11842_19766# a_12618_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3023 VGND a_4771_18260# sar9b_0.net56 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3024 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3025 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3026 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y a_40321_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3027 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3028 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3030 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3031 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3032 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3033 a_4698_25851# a_4136_25584# a_4365_25770# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X3034 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3035 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3036 VGND a_13216_23805# sar9b_0.net32 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3037 VDPWR a_6252_20780# sar9b_0._01_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3039 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3040 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3041 a_5702_24151# a_5439_24563# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3042 VGND a_5938_22378# a_5896_22188# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X3043 VGND sar9b_0.net54 a_6189_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3044 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3045 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3046 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3047 VDPWR sar9b_0.clknet_0_CLK a_2508_23444# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3048 a_5739_22488# a_4934_22432# a_5441_22522# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X3049 VGND sar9b_0.net48 a_7725_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3050 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3051 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3052 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3054 a_8695_18525# a_8266_18445# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X3055 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3056 VGND a_6307_27584# sar9b_0.net44 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3057 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3058 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3059 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3060 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3061 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3062 a_4332_23043# clk VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X3063 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3064 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3065 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3066 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3067 a_3946_27530# a_3161_27787# a_3438_27677# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3068 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3069 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3070 VGND a_13011_20806# single_9b_cdac_1.CF[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3071 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3072 a_5182_22567# sar9b_0.net64 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X3073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3074 VGND a_5196_19448# sar9b_0.net71 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3075 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3076 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3077 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3078 VGND a_12870_26263# a_12828_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3079 a_6189_24806# sar9b_0.net13 a_6102_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3080 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3081 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3082 VGND a_13011_27234# single_9b_cdac_0.SW[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3083 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3084 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 a_48343_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3086 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3087 a_7725_19238# sar9b_0.net73 a_7638_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3088 th_dif_sw_0.CK a_10227_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3089 a_11104_24151# a_10506_24506# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3090 VDPWR clk a_14871_9671# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X3091 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3092 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3093 a_6902_25087# a_6767_25185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3094 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3095 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3096 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3097 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3098 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3099 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3100 a_4083_25852# a_3747_25724# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1197 ps=1.41 w=0.42 l=0.15
X3101 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3102 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3103 single_9b_cdac_1.CF[2] a_11859_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3104 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A a_30717_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3105 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3106 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3108 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3109 single_9b_cdac_0.SW[6] a_9323_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3110 VDPWR a_13067_27662# single_9b_cdac_0.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3111 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3112 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3113 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3114 a_8334_18353# a_8057_18463# a_8664_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X3115 VDPWR sar9b_0.net38 a_10803_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3116 a_10378_27170# sar9b_0.net42 a_10899_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3117 a_12828_26141# a_11658_26134# a_12618_26134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3118 a_10895_22855# a_10506_23174# a_10230_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3119 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3120 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3121 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3122 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3123 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3124 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3125 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3126 uo_out[3] a_9939_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3127 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3128 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3129 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3130 VDPWR a_11178_20806# a_11430_20935# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3131 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3132 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3133 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3134 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3135 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3136 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3137 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3138 single_9b_cdac_1.SW[2] a_8019_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3139 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3140 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3141 uo_out[2] a_10995_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3142 VDPWR sar9b_0._07_ a_5523_21528# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2786 pd=1.64 as=0.2478 ps=2.27 w=0.84 l=0.15
X3143 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3144 VGND a_11430_20935# a_11388_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3145 a_7092_19455# sar9b_0.net10 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3146 a_6634_18206# a_5849_18463# a_6126_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3147 VDPWR a_8052_18123# a_8057_18463# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3148 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3149 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3150 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3151 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3152 VGND sar9b_0.net45 a_10218_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3153 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3154 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3155 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3156 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3157 a_8664_18206# a_8266_18445# a_8586_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3158 VGND single_9b_cdac_1.SW[5] a_39616_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3159 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3160 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3161 a_10899_27230# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3162 sar9b_0.net54 a_7347_24160# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X3163 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3164 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3165 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3166 VDPWR a_8334_18353# a_8266_18445# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3167 VDPWR a_5742_28392# a_5674_28147# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3168 VGND a_8334_17021# a_8266_17113# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3169 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3170 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3171 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3172 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3173 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3174 VGND a_10482_25831# a_10284_25707# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3175 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3176 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3177 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3178 a_26951_15501# single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3180 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3181 a_6767_25185# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3182 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3183 a_3318_27227# a_3090_27163# a_3231_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3184 VDPWR a_11214_25728# a_11146_25483# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3185 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3186 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3187 a_10254_2858# th_dif_sw_0.th_sw_1.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X3188 VGND a_5682_23444# a_5484_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3189 a_11388_20813# a_10218_20806# a_11178_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3190 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3191 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3192 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3193 VDPWR a_9494_20290# a_9449_20191# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3194 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3195 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3196 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3197 VDPWR a_11859_20574# single_9b_cdac_1.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3198 a_8586_18206# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3199 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3200 single_9b_cdac_0.SW[5] a_11339_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3201 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3202 VGND a_3156_26115# a_3161_26455# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3203 single_9b_cdac_0.SW[6] a_9323_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3204 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3205 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3206 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3207 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3208 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3209 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3210 a_8052_16791# sar9b_0.net5 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3211 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3212 VDPWR sar9b_0._03_ a_4698_25851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2972 pd=2.41 as=0.09835 ps=1.005 w=0.42 l=0.15
X3213 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3214 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3215 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3216 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3217 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3218 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3219 a_10254_2858# th_dif_sw_0.th_sw_1.CKB a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X3220 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3221 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3222 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3223 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3224 a_6870_19481# a_6642_19448# a_6783_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3225 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3226 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3227 VGND sar9b_0.net18 a_4083_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3228 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3229 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3230 VGND sar9b_0.net50 a_12246_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3231 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3232 uio_out[0] a_4083_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3233 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3235 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3236 VGND sar9b_0._14_ a_4673_24464# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.111 ps=1.045 w=0.64 l=0.15
X3237 a_10607_21189# a_10218_20806# a_9942_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3238 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3239 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3240 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3241 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3242 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3243 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3244 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3245 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3246 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3247 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3249 a_3370_26437# a_3161_26455# a_2706_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3250 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3251 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3252 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3253 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3254 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3255 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3256 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3257 VDPWR sar9b_0.net49 a_8694_20570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3258 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3259 uio_out[1] a_2931_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3260 sar9b_0.net24 a_8940_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3261 VGND a_9472_18823# sar9b_0.net26 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3262 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3263 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3264 a_9323_28371# sar9b_0.net32 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X3265 VGND a_11718_23127# a_11676_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3266 a_10029_20810# sar9b_0.net7 a_9942_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3267 a_7830_16817# a_7602_16784# a_7743_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3268 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3269 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3270 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3271 VGND a_8512_27801# sar9b_0.net22 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3272 single_9b_cdac_0.SW[5] a_11339_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X3273 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X3274 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3275 VDPWR a_11718_23127# a_11668_22819# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3276 a_2934_27473# a_2706_27440# a_2847_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X3277 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3278 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3279 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3280 VGND a_3723_20140# a_3922_20239# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X3281 VDPWR sar9b_0.net63 a_6286_22804# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X3282 tdc_0.phase_detector_0.INP a_15151_10456# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3283 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3284 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3285 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3286 VGND a_11214_25728# a_11146_25483# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3287 VGND a_10194_16784# a_9996_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3288 a_9132_7271# th_dif_sw_0.CK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3289 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3290 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3291 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3292 sar9b_0.net15 a_6130_20239# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X3293 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3294 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3295 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3296 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3297 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3298 sar9b_0.net70 a_3027_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3299 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3300 a_8098_23762# a_7914_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3301 a_11676_23231# a_10506_23174# a_11466_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3302 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3303 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3304 VDPWR sar9b_0.net54 a_6414_23681# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X3305 sar9b_0.clk_div_0.COUNT\[0\] a_5938_22378# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X3306 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3307 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3308 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3309 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3310 VGND single_9b_cdac_1.SW[2] a_54032_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3312 a_7590_24931# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3313 a_21684_3438# VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X3314 VDPWR a_12435_24802# single_9b_cdac_1.CF[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3315 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3316 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3317 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[3] a_50962_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3318 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3319 a_5682_23444# a_6132_23451# a_6084_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3320 VGND a_6534_27123# a_6492_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3321 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3322 VGND th_dif_sw_0.VCN a_14897_9355# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3323 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3324 a_11718_23127# a_11466_23174# a_11856_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3325 VGND sar9b_0.net69 sar9b_0._04_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3326 VGND sar9b_0.net51 a_7443_21496# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X3327 a_8004_16817# a_7743_16817# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3328 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3329 uo_out[3] a_9939_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3330 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3331 VGND a_5812_21028# a_5581_20992# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17462 pd=1.185 as=0.077 ps=0.83 w=0.55 l=0.15
X3332 single_9b_cdac_1.SW[6] a_13011_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3333 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3334 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3335 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3336 a_10932_25713# sar9b_0.net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3337 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3338 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3339 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3340 VDPWR sar9b_0.net48 a_7638_19238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3341 VGND a_13011_20574# single_9b_cdac_1.CF[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3342 sar9b_0.net24 a_8940_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X3343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3344 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3345 a_11955_16814# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3346 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3347 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3348 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3349 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3350 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3352 VGND a_3521_24240# a_3539_24543# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X3353 VDPWR a_9126_19131# a_9076_18823# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3354 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3355 a_3438_26345# a_3156_26115# a_3799_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3356 VGND a_6030_24396# a_5962_24151# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3357 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3358 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3359 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3360 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3361 a_6084_23477# a_5823_23477# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3362 sar9b_0.net1 a_6867_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X3363 a_6492_27227# a_5322_27170# a_6282_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3364 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3365 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3366 uo_out[4] a_8691_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3367 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3368 VGND single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3369 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3370 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3371 a_6744_23238# a_6484_22845# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.27625 ps=1.625 w=1 l=0.25
X3372 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3373 VGND sar9b_0.net4 a_6378_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3374 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3375 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3376 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3377 VDPWR a_3521_24240# a_3476_24141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X3378 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3379 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3381 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3382 tdc_0.OUTN tdc_0.OUTP a_16555_12412# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3383 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3384 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3385 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3386 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3387 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3388 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3389 a_3799_26517# a_3370_26437# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X3390 VDPWR a_11859_20574# single_9b_cdac_1.SW[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3391 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3392 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3393 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3394 VDPWR a_10803_19474# single_9b_cdac_1.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3395 a_15151_10456# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X3396 a_2508_20780# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X3397 a_12684_20379# sar9b_0.net51 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24915 pd=2.37 as=0.15198 ps=1.17 w=0.55 l=0.15
X3398 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3399 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3400 a_8952_26198# a_8554_26437# a_8874_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3401 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3402 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3403 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3404 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3405 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3406 a_3476_24141# a_2835_24136# a_3369_24181# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X3407 VGND sar9b_0.net53 a_12246_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3408 a_9264_19235# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3409 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3410 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3411 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3412 a_6902_25087# a_6767_25185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3413 VDPWR a_6444_21738# sar9b_0.net64 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3414 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3415 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3416 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3417 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3418 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3419 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3420 a_12047_19857# a_11842_19766# a_11382_19478# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3421 single_9b_cdac_1.SW[7] a_13011_19242# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3422 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3423 VGND sar9b_0.net25 a_12531_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3424 a_10690_22806# a_10506_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3425 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3426 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3427 uo_out[1] a_12531_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3428 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3429 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3430 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3431 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3432 a_10230_23234# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3433 a_8874_26198# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3434 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3435 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3436 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3437 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3438 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3439 VGND sar9b_0.net47 a_6870_19481# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X3440 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3441 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3442 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3443 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3444 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y a_64331_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3445 VDPWR a_2892_23070# sar9b_0.net66 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3446 VDPWR a_13011_24802# single_9b_cdac_0.SW[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3447 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3448 VDPWR sar9b_0.net13 a_13011_25902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3449 a_12491_27662# sar9b_0.net29 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X3450 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3453 VDPWR sar9b_0.net5 a_13011_20574# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3454 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3455 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3456 VDPWR a_7936_25137# sar9b_0.cyclic_flag_0.FINAL VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3457 VDPWR a_4812_21738# sar9b_0.net65 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3458 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3459 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3460 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3461 a_5443_19074# sar9b_0.net4 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X3462 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3463 a_3690_26198# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3464 a_12684_20379# sar9b_0.net51 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2051 ps=1.52 w=0.84 l=0.15
X3465 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X3467 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3468 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3469 a_3946_27530# a_3156_27447# a_3438_27677# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X3470 sar9b_0.net3 a_2451_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3471 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3472 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3473 sar9b_0._12_ sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2786 ps=1.64 w=1.12 l=0.15
X3474 VDPWR a_12182_18427# a_12137_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3475 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3476 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3477 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3478 sar9b_0.net10 a_6636_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3479 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3480 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3481 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3482 a_8074_20870# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3483 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3484 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3485 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3486 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3487 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3488 VGND sar9b_0.net60 a_6765_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3489 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3490 VGND sar9b_0.net36 a_10803_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3491 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3492 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3493 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3494 VGND a_3540_27045# a_3545_26914# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3495 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3496 a_9974_17626# a_9839_17527# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3497 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3498 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3499 a_10607_25185# a_10402_25094# a_9942_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3500 VDPWR sar9b_0.net54 a_5439_24563# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X3501 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3502 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3503 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A a_55773_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3504 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3505 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3506 a_3166_20145# sar9b_0._00_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X3507 VGND sar9b_0.net8 a_8970_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3508 sar9b_0.net4 a_5331_16810# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X3509 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3510 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3511 a_54737_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3512 a_6538_24506# a_5748_24381# a_6030_24396# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X3513 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3514 VGND th_dif_sw_0.VCP a_17125_9355# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3515 VGND a_9939_28566# uo_out[3] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3516 a_9480_20510# a_9154_20142# a_9359_20191# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3517 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3518 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3519 single_9b_cdac_1.CF[4] a_13011_21906# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3520 a_10762_18823# a_10548_19053# a_10098_19171# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X3521 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[8] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3522 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3523 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3524 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3525 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3526 a_10548_19053# sar9b_0.net7 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3527 a_16357_9613# th_dif_sw_0.VCN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3528 a_7978_22202# sar9b_0.net61 a_8499_22142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3529 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3530 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3531 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3532 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3533 sar9b_0.net60 a_2547_28132# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3534 a_6765_27470# sar9b_0.net40 a_6678_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3535 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3536 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3537 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3538 VGND a_10995_28566# uo_out[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3539 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3540 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3541 VDPWR sar9b_0.net45 a_12560_27128# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X3542 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3543 VDPWR sar9b_0.net62 a_7882_19538# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X3544 VGND sar9b_0.net46 a_5910_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3545 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3546 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3547 VGND a_3180_19448# sar9b_0._00_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3548 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3550 a_3754_26815# a_3545_26914# a_3090_27163# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3551 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3552 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3553 tdc_0.RDY a_16159_13315# a_16185_13034# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X3554 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3555 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3556 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3557 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3558 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3559 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3560 VGND single_9b_cdac_1.SW[3] a_49221_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3561 single_9b_cdac_0.SW[5] a_11339_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3562 a_5298_24499# a_5748_24381# a_5700_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3563 a_8499_22142# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3564 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3565 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A a_46159_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3566 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3567 VGND sar9b_0._03_ a_4698_25851# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.23015 pd=2.1 as=0.15563 ps=1.215 w=0.42 l=0.15
X3568 a_4118_22572# a_3206_22432# a_4011_22488# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X3569 VGND a_7602_18116# a_7404_18116# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3570 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3571 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3572 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3573 a_11668_22819# a_10690_22806# a_11466_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3574 VDPWR single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3575 VGND a_10227_23490# sar9b_0.net53 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3576 VDPWR single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3577 a_6286_22804# sar9b_0._12_ sar9b_0._02_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X3578 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3579 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3580 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3581 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3582 VDPWR sar9b_0.net65 a_3371_23106# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.26 as=0.126 ps=1.14 w=0.84 l=0.15
X3583 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3584 th_dif_sw_0.VCP ua[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3585 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3586 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3587 a_3370_27769# a_3156_27447# a_2706_27440# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X3588 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3589 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3590 a_2637_24802# sar9b_0.net63 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3591 sar9b_0._11_ a_4496_20468# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3592 a_13067_27662# sar9b_0.net28 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X3593 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3594 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3595 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3596 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3597 VGND a_5742_28392# a_5674_28147# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3598 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3599 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3600 VDPWR th_dif_sw_0.CK a_9132_7271# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3601 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3602 a_12870_23599# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3603 VGND sar9b_0.net46 a_5133_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3604 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3606 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3607 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3608 a_12047_23853# a_11842_23762# a_11382_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3609 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3610 sar9b_0.net49 a_9363_20826# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X3611 VGND a_10662_17799# a_10620_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X3612 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3613 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3614 VDPWR a_10482_25831# a_10284_25707# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3615 VDPWR sar9b_0.clknet_0_CLK a_2508_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3616 VGND a_11859_17910# single_9b_cdac_1.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3617 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3618 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3619 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3620 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3621 VGND a_13011_20574# single_9b_cdac_1.CF[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3622 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3623 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3624 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3625 single_9b_cdac_0.SW[0] a_13011_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3626 VDPWR sar9b_0.net57 a_7914_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3627 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3628 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X3629 VGND a_12684_20379# sar9b_0.net50 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X3630 a_11382_19478# sar9b_0.net73 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3631 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3632 a_6562_25094# a_6378_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3633 a_9126_19131# a_8874_19178# a_9264_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3634 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3635 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3636 VDPWR single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3637 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3638 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3639 a_5460_28377# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3640 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3641 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3642 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3643 VGND a_7539_28566# uo_out[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3644 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3645 VGND sar9b_0.net41 a_13011_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3646 a_9076_18823# a_8098_18810# a_8874_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3647 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3648 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3649 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3650 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3651 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3652 single_9b_cdac_1.CF[5] a_13011_23238# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3653 VDPWR a_4210_22378# a_4118_22572# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X3654 a_6282_17846# a_5322_17846# a_5846_17626# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3655 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3656 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3657 VDPWR sar9b_0.net24 a_10995_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3658 VGND a_13011_25902# single_9b_cdac_1.CF[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3659 VDPWR sar9b_0.net37 a_8019_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3660 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3661 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3662 a_9730_24138# a_9546_24506# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3663 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3664 VDPWR a_11178_27466# a_11430_27595# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3665 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3666 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3667 a_11776_21141# a_11178_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3668 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3670 VDPWR a_12182_22423# a_12137_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3671 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3672 a_9270_24566# sar9b_0.net62 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3673 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A a_25915_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3675 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3676 a_11842_26426# a_11658_26134# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3677 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3678 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X3679 VDPWR sar9b_0.clknet_1_1__leaf_CLK a_2835_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3680 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3681 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3682 VDPWR sar9b_0.net51 a_9363_20826# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X3683 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3684 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3685 VDPWR sar9b_0.net43 a_11859_20574# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3686 single_9b_cdac_1.SW[3] a_10803_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3687 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3688 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3689 uo_out[0] a_11915_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3690 VDPWR a_5298_24499# a_5100_24375# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3691 a_12618_19474# a_11658_19474# a_12182_19759# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3692 VDPWR a_8512_27801# sar9b_0.net22 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3693 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3694 VGND sar9b_0.net49 a_10029_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3695 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3696 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] a_41357_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3697 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3698 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3699 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3700 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3701 a_3090_27163# a_3540_27045# a_3492_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3702 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3703 VDPWR a_10194_16784# a_9996_16784# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3704 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3705 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3706 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3707 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3708 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3709 a_3110_27885# a_2847_27473# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3710 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3711 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3712 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3713 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3714 VGND a_10859_26330# single_9b_cdac_0.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3715 a_5739_22488# a_4755_22138# a_5441_22522# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X3716 a_11430_20935# a_11178_20806# a_11568_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3717 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3718 a_11776_25137# a_11178_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3719 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3720 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3721 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3722 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3723 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3724 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3725 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3726 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3727 a_7402_22441# a_7193_22459# a_6738_22112# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3728 sar9b_0.net48 a_10035_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3729 VGND a_8052_16791# a_8057_17131# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3730 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3731 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3732 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3733 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3734 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3735 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3736 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3737 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3738 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3739 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3741 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3742 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3743 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3744 a_9870_27060# a_9588_27045# a_10231_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3745 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3746 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3747 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3748 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3749 a_3492_27227# a_3231_27227# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3750 a_4922_20857# sar9b_0._17_ a_4886_21124# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3751 a_11338_19178# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3752 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3753 VDPWR a_10227_23490# sar9b_0.net53 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X3754 sar9b_0.net63 a_6861_22828# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.194 ps=1.475 w=1.12 l=0.15
X3755 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3756 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3757 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3758 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3759 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3760 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3761 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3762 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3763 a_5761_19487# sar9b_0._07_ sar9b_0._10_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X3764 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3765 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3766 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3767 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3768 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X3769 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3770 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3771 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3772 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3773 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3774 a_49926_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3775 VDPWR a_6252_19074# sar9b_0.net55 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3776 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3777 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3778 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3779 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3780 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3781 a_8266_17113# a_8057_17131# a_7602_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3783 VDPWR a_9323_28371# single_9b_cdac_0.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3784 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3785 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3787 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3788 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A a_40321_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3789 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3790 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3791 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3792 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3793 VGND sar9b_0.net52 a_10806_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3794 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3795 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3796 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3797 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3798 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3799 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3800 a_9130_26198# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3801 VDPWR a_12870_22267# a_12820_22557# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3802 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3803 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3804 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3805 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3806 VGND sar9b_0.net7 a_11859_21906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3807 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3808 VDPWR a_13011_25902# single_9b_cdac_1.CF[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3809 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3811 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3812 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3813 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3814 VDPWR a_13011_20574# single_9b_cdac_1.CF[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3815 a_9261_17906# sar9b_0.net6 a_9174_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3816 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3817 a_10470_21795# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3818 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3819 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3820 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3821 a_2706_26108# a_3156_26115# a_3108_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X3822 a_9442_21474# a_9258_21842# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3823 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3824 VGND a_6880_17491# sar9b_0.net5 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3826 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3827 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3828 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3829 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3830 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3831 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3832 th_dif_sw_0.th_sw_1.CKB a_21177_7457# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3833 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3834 a_10806_24866# a_10742_25087# a_10728_24866# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3835 a_8982_21902# sar9b_0.net8 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3836 a_5628_19768# sar9b_0.net47 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X3837 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3838 VDPWR single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3839 VGND a_10995_28566# uo_out[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3840 a_5506_26802# a_5322_27170# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3841 a_11382_23474# sar9b_0.net74 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3842 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3843 a_8512_27801# a_7914_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3844 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3845 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3846 a_10742_27751# a_10607_27849# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3847 VGND a_6414_23681# a_6346_23773# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3848 VDPWR a_12618_23470# a_12870_23599# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3849 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3850 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3851 single_9b_cdac_0.SW[1] a_13011_27234# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3852 a_5441_22522# a_5289_22527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X3853 single_9b_cdac_1.SW[5] a_13011_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3854 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3856 sar9b_0.net23 a_7692_26108# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3857 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3858 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3859 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3860 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3861 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3862 VDPWR sar9b_0.net23 a_9939_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3863 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3864 VGND a_4922_20857# sar9b_0._18_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X3865 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3866 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3867 a_3108_26141# a_2847_26141# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3868 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3869 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3870 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3871 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3872 VGND a_4236_21738# sar9b_0.net67 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3873 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3874 a_7343_27849# a_7138_27758# a_6678_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3875 a_8098_23762# a_7914_23470# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3876 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3877 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3878 VGND sar9b_0.net52 a_11469_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3879 a_10728_24866# a_10402_25094# a_10607_25185# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3880 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3881 VGND a_8019_17910# single_9b_cdac_1.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X3882 VGND sar9b_0.net49 a_10227_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X3883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3884 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3885 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3886 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3887 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.th_sw_main_0.VGS ua[4] VGND sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X3888 uio_out[0] a_4083_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3889 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3890 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3891 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3892 a_3855_25792# a_4136_25584# a_4091_25468# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.09975 ps=0.895 w=0.42 l=0.15
X3893 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3894 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3895 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3896 a_9165_24988# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.2102 ps=1.505 w=1 l=0.15
X3897 VGND a_4018_24235# a_3976_24520# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X3898 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3899 a_6132_23451# sar9b_0.net57 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3900 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3901 a_8842_18206# a_8057_18463# a_8334_18353# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3902 single_9b_cdac_1.SW[4] a_11859_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X3903 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3904 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3905 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3906 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3907 VGND a_9138_27163# a_8940_27039# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3908 a_12618_23470# a_11658_23470# a_12182_23755# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3909 VGND a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.2109 ps=2.05 w=0.74 l=0.15
X3910 a_8874_23470# a_8098_23762# a_8438_23755# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3911 a_8386_22806# a_8202_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3912 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3913 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3914 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3915 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3916 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3917 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3918 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3919 single_9b_cdac_1.CF[1] a_12435_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3920 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3921 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3922 VGND sar9b_0._07_ a_5523_21528# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.22412 pd=1.365 as=0.15675 ps=1.67 w=0.55 l=0.15
X3923 VDPWR a_9782_21622# a_9737_21523# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3924 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3925 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3926 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3928 a_11469_26138# sar9b_0.net74 a_11382_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3929 a_11146_25483# a_10937_25582# a_10482_25831# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3930 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3931 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3932 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3933 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3935 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3936 VGND a_2706_26108# a_2508_26108# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3937 VGND a_6252_20780# sar9b_0._01_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3938 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3939 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3940 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3941 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3942 a_6030_24396# a_5748_24381# a_6391_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3943 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3944 a_3231_27227# a_3090_27163# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X3945 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3946 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3947 sar9b_0._17_ sar9b_0.net63 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2352 ps=1.54 w=1.12 l=0.15
X3948 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3949 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3950 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3952 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3953 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3954 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3955 a_9930_20510# a_8970_20510# a_9494_20290# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3956 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3957 tdc_0.RDY tdc_0.phase_detector_0.pd_out_0.B a_16542_13134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X3958 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3959 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3960 VDPWR sar9b_0.net54 a_10227_23490# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X3961 sar9b_0.net10 a_6636_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X3962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3963 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3964 VDPWR a_8166_27595# a_8116_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3965 VDPWR sar9b_0.net52 a_9942_24806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3966 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3967 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3968 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3969 VGND a_10926_17021# a_10858_17113# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X3970 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3971 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3972 a_2847_27473# a_2706_27440# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X3973 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3974 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3975 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3976 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3977 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3978 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_4947_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3979 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3980 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X3981 VGND a_13011_25902# single_9b_cdac_1.CF[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3983 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3984 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3985 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3986 VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# dw_17224_1400# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X3987 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3988 a_8438_23755# a_8303_23853# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3989 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3990 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3991 VDPWR a_5581_20992# sar9b_0._09_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.3304 ps=2.83 w=1.12 l=0.15
X3992 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3993 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3994 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3995 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3996 a_10800_17903# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3997 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3999 VGND a_11430_27595# a_11388_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4000 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4001 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4002 VGND sar9b_0.net6 a_12435_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4003 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4004 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4005 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4006 VGND sar9b_0.net53 a_9357_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4007 sar9b_0.net74 a_10707_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4008 a_7306_19777# a_7097_19795# a_6642_19448# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4009 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4010 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4011 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4012 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4013 VDPWR a_9323_28371# single_9b_cdac_0.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4014 VDPWR sar9b_0.net58 a_4467_24162# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X4015 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4016 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4017 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4018 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4019 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4020 sar9b_0.net59 a_3603_28156# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X4021 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4022 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4023 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4024 VDPWR a_9939_28566# uo_out[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4025 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4026 VGND a_13216_18477# sar9b_0.net28 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4027 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4028 sar9b_0.net43 a_5100_24375# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4029 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4030 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4031 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4032 a_3438_27677# a_3161_27787# a_3768_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4033 sar9b_0._07_ a_3371_23106# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.11312 ps=1.065 w=0.74 l=0.15
X4034 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4035 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4036 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4037 a_11388_27473# a_10218_27466# a_11178_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4038 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4039 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4040 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4041 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INN a_15400_11316# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4042 VGND sar9b_0.net58 a_5238_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4043 VDPWR a_10995_28566# uo_out[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4044 a_9357_24566# sar9b_0.net62 a_9270_24566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4045 VDPWR a_8019_17910# single_9b_cdac_1.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4046 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4047 a_8052_18123# sar9b_0.net56 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4048 a_10859_26330# sar9b_0.net33 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X4049 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4050 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4051 VDPWR a_7347_24160# sar9b_0.net54 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X4052 VGND sar9b_0.net53 a_10317_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4053 a_6088_20524# a_4947_20140# a_5931_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X4054 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4055 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4056 VDPWR sar9b_0.net10 a_6922_23534# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4057 sar9b_0._04_ sar9b_0.net69 a_2540_22432# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X4058 a_5535_18149# a_5394_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4059 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4060 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4061 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4062 a_9802_26815# a_9588_27045# a_9138_27163# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4063 a_6030_24396# a_5753_24250# a_6360_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4064 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4065 single_9b_cdac_1.CF[3] a_13011_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4066 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4067 a_3768_27530# a_3370_27769# a_3690_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4068 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4069 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4070 a_9359_20191# a_8970_20510# a_8694_20570# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4071 a_12246_19538# a_12182_19759# a_12168_19538# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4072 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4073 a_11915_28371# sar9b_0.net14 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X4074 a_5748_24381# sar9b_0.net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4075 VGND a_2603_17006# th_dif_sw_0.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4076 a_4886_21124# sar9b_0.net65 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4077 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4078 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4079 a_3991_19768# sar9b_0._07_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.4075 pd=1.815 as=0.1853 ps=1.385 w=1 l=0.15
X4080 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4081 VDPWR a_3180_19448# sar9b_0._00_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4082 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4083 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4084 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4086 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4087 a_10506_24506# a_9730_24138# a_10070_24286# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4088 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4089 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4090 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4091 VDPWR a_11339_27039# single_9b_cdac_0.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4092 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4093 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4094 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4095 a_12560_27128# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X4096 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X4097 a_10317_23234# sar9b_0.net74 a_10230_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4098 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4099 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4100 VDPWR single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4101 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4102 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4103 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4104 a_10194_16784# a_10644_16791# a_10596_16817# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X4105 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4106 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4107 VDPWR a_5460_28377# a_5465_28246# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4108 a_12168_19538# a_11842_19766# a_12047_19857# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4109 VGND sar9b_0.net23 a_9939_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4110 uo_out[1] a_12531_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4111 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4112 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4113 a_10029_27470# sar9b_0.net43 a_9942_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4114 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4115 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4116 a_10326_19235# a_10098_19171# a_10239_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X4117 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4118 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4119 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4120 uo_out[2] a_10995_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4121 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4122 single_9b_cdac_1.CF[6] a_13011_24570# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4123 a_16970_11404# tdc_0.phase_detector_0.INP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X4124 VDPWR a_4083_28566# uio_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4125 VDPWR sar9b_0.net55 a_5811_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X4126 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4127 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4128 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4129 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4130 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4131 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4132 VGND sar9b_0.net8 a_13011_20806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4133 a_10596_16817# a_10335_16817# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4134 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4135 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4136 a_3731_22165# a_3206_22432# a_3561_22527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X4137 single_9b_cdac_1.CF[2] a_11859_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4138 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4139 a_10200_27170# a_9802_26815# a_10122_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4140 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4141 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4142 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4143 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4144 a_7735_19857# a_7306_19777# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4145 VDPWR a_7539_28566# uo_out[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4146 a_8438_18958# a_8303_18859# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4147 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4148 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4149 VGND sar9b_0.net27 a_13011_27234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4150 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4151 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4152 a_5832_17846# a_5506_17478# a_5711_17527# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4153 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4154 a_7914_27466# a_6954_27466# a_7478_27751# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4155 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] a_65367_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4156 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4157 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4158 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4159 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4160 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4161 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4162 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4163 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4164 VGND sar9b_0.net52 a_7725_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4165 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4166 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4167 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4168 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4169 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4170 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4171 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4172 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4173 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4174 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4175 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4176 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4177 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4178 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4179 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4180 VDPWR a_11430_24931# a_11380_25221# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4181 single_9b_cdac_1.SW[1] a_10803_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4182 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4183 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4184 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4185 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4186 VDPWR a_12870_19603# a_12820_19893# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4187 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4188 a_10122_27170# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4189 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4190 VGND sar9b_0._10_ a_4583_20468# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X4191 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4192 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4193 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4194 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4195 a_5711_26851# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4196 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4197 VGND a_5460_28377# a_5465_28246# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4198 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4199 a_10896_24563# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4200 a_7725_23474# sar9b_0.net11 a_7638_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4201 VGND a_11859_21906# single_9b_cdac_1.CF[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4202 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4203 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4204 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4205 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4206 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4207 a_5298_24499# a_5753_24250# a_5702_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X4208 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4209 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4210 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4211 a_12820_18561# a_11842_18434# a_12618_18142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4212 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4213 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4214 VDPWR a_3922_20239# a_3830_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4215 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4216 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4217 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4218 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4219 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4220 a_6634_18206# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4221 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4222 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4223 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4224 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4225 VGND sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X4226 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4227 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4228 a_10762_18823# a_10553_18922# a_10098_19171# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4229 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4230 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4231 a_3561_22527# a_3206_22432# a_3454_22567# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X4232 a_10662_17799# a_10410_17846# a_10800_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4233 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4234 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4235 a_4749_27652# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.2102 ps=1.505 w=1 l=0.15
X4236 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4237 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4238 a_9494_20290# a_9359_20191# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4239 VDPWR a_13011_17910# single_9b_cdac_1.SW[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4240 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4241 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4242 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4243 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4244 VGND sar9b_0.net60 a_7542_27530# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4245 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4246 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4247 VGND sar9b_0.net12 a_11658_26134# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4248 single_9b_cdac_1.CF[6] a_13011_24570# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4249 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4250 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4251 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4252 sar9b_0.net60 a_2547_28132# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4253 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4254 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4255 a_10218_21842# a_9442_21474# a_9782_21622# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4256 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4257 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4258 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A a_64331_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4259 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4260 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4261 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4262 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4263 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4264 a_10038_17846# a_9974_17626# a_9960_17846# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4266 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4267 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4268 a_5674_28147# a_5465_28246# a_5010_28495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4269 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4270 a_7743_16817# a_7602_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4271 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4272 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4273 a_3946_26198# a_3161_26455# a_3438_26345# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4274 a_8591_22855# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4275 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4276 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4277 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4278 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4279 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4280 VGND th_dif_sw_0.CK a_9132_7271# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1295 ps=1.09 w=0.74 l=0.15
X4281 a_16881_10256# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16527_10454# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4282 a_12246_23534# a_12182_23755# a_12168_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4283 sar9b_0.net27 a_5196_18116# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4284 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4285 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4286 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4287 VDPWR a_7188_22119# a_7193_22459# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4288 a_13216_18477# a_12618_18142# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4290 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4291 a_21684_3438# th_dif_sw_0.th_sw_1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X4292 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4293 a_3380_20145# a_2739_20140# a_3273_20185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X4294 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4295 a_8116_27885# a_7138_27758# a_7914_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4296 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4297 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4298 a_7800_22202# a_7402_22441# a_7722_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4299 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4300 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4301 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4302 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4303 a_12182_26419# a_12047_26517# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4304 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4305 a_11718_23127# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4306 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4307 VGND clk a_16881_10256# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X4308 VDPWR a_7470_22349# a_7402_22441# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4309 a_5374_20145# sar9b_0._01_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X4310 VDPWR sar9b_0.net49 a_10035_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4312 sar9b_0.net20 a_4812_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4313 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4314 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4315 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4316 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4317 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4318 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4319 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4320 single_9b_cdac_1.SW[8] a_11859_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4321 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4322 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4323 VGND a_2547_28132# sar9b_0.net60 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4324 VDPWR a_6130_20239# a_6038_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4325 a_12168_23534# a_11842_23762# a_12047_23853# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4326 VDPWR a_7404_17715# sar9b_0.net73 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4327 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4328 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4329 sar9b_0.net17 a_2508_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4330 a_54737_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4331 VGND a_5235_27466# uo_out[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4332 a_10231_26851# a_9802_26815# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4333 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] a_36555_29911# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4334 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4335 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4336 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4337 VDPWR sar9b_0.net47 a_7470_22349# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4338 a_7722_22202# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4339 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4340 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4341 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4342 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4343 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4344 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4345 VGND a_21177_7457# th_dif_sw_0.th_sw_1.CKB VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4346 VGND a_13011_16810# single_9b_cdac_1.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4347 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4348 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4349 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4350 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4351 a_6738_22112# a_7188_22119# a_7140_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X4352 sar9b_0._18_ a_4922_20857# a_5083_21100# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X4353 a_9359_20191# a_9154_20142# a_8694_20570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4354 VDPWR sar9b_0.net46 a_8334_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4355 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4356 VDPWR a_9588_27045# a_9593_26914# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4357 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4358 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4359 a_4091_25468# a_3747_25724# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1239 ps=1.43 w=0.42 l=0.15
X4360 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4361 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4362 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4363 a_12137_19857# a_11658_19474# a_12047_19857# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4364 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4365 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4366 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4367 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4368 VGND a_11430_24931# a_11388_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4369 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4370 VDPWR a_10644_16791# a_10649_17131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4371 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4372 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4373 single_9b_cdac_1.SW[6] a_13011_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4374 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4375 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4376 VDPWR a_12531_28566# uo_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4377 VDPWR a_5846_26950# a_5801_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4378 VDPWR a_8052_16791# a_8057_17131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4379 a_3946_26198# a_3156_26115# a_3438_26345# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4381 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4382 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4383 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4384 VDPWR sar9b_0.net53 a_10230_23234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4385 VGND sar9b_0.net48 a_10326_19235# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4386 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4387 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4388 sar9b_0.clk_div_0.COUNT\[2\] a_4018_24235# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X4389 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4390 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4391 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4392 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A a_60565_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4393 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4394 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4395 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4396 a_5910_27170# a_5846_26950# a_5832_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4397 VGND sar9b_0.clknet_0_CLK a_2508_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4398 a_9126_19131# sar9b_0.net48 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4399 VDPWR tdc_0.RDY a_5331_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4400 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4401 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4402 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4403 a_50962_15501# single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4404 a_3494_26815# a_3231_27227# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4405 VDPWR a_9472_23805# sar9b_0.net12 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4406 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4407 VDPWR a_10742_25087# a_10697_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4408 a_11388_24809# a_10218_24802# a_11178_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4409 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4410 a_16527_10454# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X4411 VDPWR a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4412 a_4072_19474# sar9b_0.net71 a_3991_19768# VDPWR sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.4075 ps=1.815 w=1 l=0.15
X4413 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4414 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4415 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4416 VGND a_2892_23070# sar9b_0.net66 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4417 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4418 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4419 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4420 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4421 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4422 VGND sar9b_0.net44 a_5322_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4423 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4424 a_4330_27170# sar9b_0.net37 a_4851_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4425 VGND a_3795_19512# a_4211_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.20905 pd=1.305 as=0.2997 ps=1.55 w=0.74 l=0.15
X4426 VGND a_9870_27060# a_9802_26815# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X4427 VDPWR sar9b_0.net9 a_8074_20870# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4428 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4429 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4430 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4431 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4432 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4433 VDPWR sar9b_0.net40 a_13011_16810# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4434 th_dif_sw_0.th_sw_1.CK a_9132_7271# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4435 VDPWR a_8726_22954# a_8681_22855# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4436 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4437 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4438 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4439 a_10697_25185# a_10218_24802# a_10607_25185# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4440 a_8303_18859# a_8098_18810# a_7638_19238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4441 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 a_24332_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4442 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4443 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A a_15052_11404# VGND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X4444 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4445 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4446 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4447 a_12588_16784# tdc_0.OUTP VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4448 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4449 a_6880_26815# a_6282_27170# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4450 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4451 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4452 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4454 VGND a_13067_27662# single_9b_cdac_0.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4455 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4456 a_8790_23174# a_8726_22954# a_8712_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4457 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4458 a_10607_25185# a_10218_24802# a_9942_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4459 VDPWR a_10758_24459# a_10708_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4460 VGND a_6738_22112# a_6540_22112# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4461 VDPWR a_13011_21906# single_9b_cdac_1.CF[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4462 VDPWR tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4463 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4464 a_5846_26950# a_5711_26851# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4465 a_3364_25120# sar9b_0._14_ a_2893_24992# VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4466 a_10758_24459# a_10506_24506# a_10896_24563# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4467 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4468 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4469 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4470 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4471 tdc_0.OUTP tdc_0.OUTN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4472 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4473 VGND a_6132_23451# a_6137_23791# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4474 VGND clk a_4332_23043# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4475 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4476 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4477 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4478 VGND sar9b_0.net11 a_8202_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4479 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4480 a_10029_24806# sar9b_0.net12 a_9942_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4481 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4482 VGND a_13164_28398# sar9b_0.net14 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4483 a_8712_23174# a_8386_22806# a_8591_22855# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4484 VDPWR sar9b_0.net6 a_12435_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4485 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4486 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4487 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4488 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4489 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4490 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4491 a_13216_22473# a_12618_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4492 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4493 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4494 sar9b_0.net15 a_6130_20239# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X4495 a_3946_27530# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4496 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4497 a_2934_26141# a_2706_26108# a_2847_26141# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X4498 a_8031_26141# a_7890_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4499 VDPWR a_9165_24988# sar9b_0.net52 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X4500 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4501 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4502 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4503 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4504 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4505 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4506 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP a_16222_11316# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4507 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4508 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4509 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4510 a_9760_22819# a_9162_23174# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4511 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4512 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4513 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4514 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4515 VGND a_7602_16784# a_7404_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4516 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4517 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4518 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4519 VGND a_10035_19474# sar9b_0.net48 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4520 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4521 a_6346_23773# a_6137_23791# a_5682_23444# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4522 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4523 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4524 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4525 a_55773_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4526 VDPWR sar9b_0.net55 a_7347_24160# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X4527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4528 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4529 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4530 VGND sar9b_0.net57 a_7914_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4531 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4532 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4533 VDPWR sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4534 VGND a_10182_20463# a_10140_20567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4535 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A a_31753_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4536 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4537 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4538 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4539 VDPWR a_5748_24381# a_5753_24250# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4540 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4541 a_30717_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4542 a_4332_23043# clk VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4543 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4544 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4545 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4546 sar9b_0.net45 a_8883_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4547 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4548 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4549 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4550 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4551 a_12137_23853# a_11658_23470# a_12047_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4552 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4553 VGND sar9b_0.net47 a_6966_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X4554 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4555 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4556 a_11776_27801# a_11178_27466# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4557 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4558 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4559 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4560 VGND a_10932_25713# a_10937_25582# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4561 a_2508_20780# sar9b_0.clknet_0_CLK VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4562 sar9b_0.net40 a_6444_19448# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4563 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4564 single_9b_cdac_0.SW[3] a_12491_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X4565 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4567 VDPWR sar9b_0.net1 a_10707_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4568 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4569 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4570 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4571 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4572 a_8438_23755# a_8303_23853# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4573 VDPWR sar9b_0.net50 a_11382_19478# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4574 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4575 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4576 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4577 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4578 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4579 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4580 VGND single_9b_cdac_0.SW[6] a_34814_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4581 VGND sar9b_0.net59 a_10029_27470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4582 a_46159_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4583 VGND a_7936_25137# sar9b_0.cyclic_flag_0.FINAL VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4584 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4585 a_21177_7457# th_dif_sw_0.CKB VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4586 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4587 VGND sar9b_0.net54 a_10227_23490# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X4588 a_49926_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4589 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4590 single_9b_cdac_1.CF[4] a_13011_21906# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4591 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4592 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4593 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4594 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4595 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4596 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4597 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4598 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4599 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4600 a_11430_27595# a_11178_27466# a_11568_27473# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4601 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4602 uo_out[0] a_11915_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4603 a_4330_27170# sar9b_0.net58 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4604 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4605 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4606 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4607 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4609 VDPWR sar9b_0.net53 a_9270_24566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4610 a_5196_19448# sar9b_0.net16 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4611 VGND a_11436_17742# sar9b_0.net61 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4612 a_12618_22138# a_11842_22430# a_12182_22423# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4613 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4614 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4615 a_3014_24136# a_2835_24136# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4616 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4617 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4618 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4619 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4620 VDPWR sar9b_0.net8 a_13011_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4621 VDPWR a_10803_18142# single_9b_cdac_1.SW[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4622 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4623 a_6414_23681# a_6132_23451# a_6775_23853# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X4624 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4625 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4626 VDPWR a_11915_28371# uo_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4627 VGND a_5748_24381# a_5753_24250# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X4628 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4629 single_9b_cdac_0.SW[4] a_11915_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4630 VGND a_5235_27466# uo_out[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4631 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4632 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4633 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4634 a_63626_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4635 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4636 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4637 a_9165_24988# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X4638 VDPWR sar9b_0.net57 a_10218_24802# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4639 a_7044_19481# a_6783_19481# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4640 VGND a_13011_16810# single_9b_cdac_1.SW[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4641 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4642 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4643 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4644 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4645 VGND a_7443_21496# sar9b_0.net47 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4646 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4647 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4648 VGND a_7566_21017# a_7498_21109# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X4649 VGND sar9b_0.net51 a_6579_18832# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X4650 a_12047_18525# a_11842_18434# a_11382_18146# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4651 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4652 VGND a_5580_24776# sar9b_0._03_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4653 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4654 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4655 VGND a_6444_21738# sar9b_0.net64 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4656 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4657 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4658 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4659 a_3830_20140# a_2918_20140# a_3723_20140# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X4660 VDPWR a_10035_19474# sar9b_0.net48 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4661 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4662 a_12047_19857# a_11658_19474# a_11382_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4663 VGND a_11008_17491# sar9b_0.net7 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4664 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4665 a_6775_23853# a_6346_23773# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4666 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4667 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4668 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4670 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4671 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4672 a_10378_27170# a_9593_26914# a_9870_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4673 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4676 a_11178_24802# a_10402_25094# a_10742_25087# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4677 a_3369_24181# a_3014_24136# a_3262_24141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X4678 a_5823_23477# a_5682_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4679 sar9b_0._08_ a_4072_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2557 ps=1.59 w=1.12 l=0.15
X4680 VDPWR sar9b_0.net11 a_13011_24570# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X4681 a_11178_20806# a_10218_20806# a_10742_21091# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4682 VDPWR sar9b_0.net61 a_11338_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4683 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4684 VDPWR a_6030_24396# a_5962_24151# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4685 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4686 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4687 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4688 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4689 uo_out[0] a_11915_28371# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X4690 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4691 a_6672_17903# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4692 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4693 VDPWR a_3695_23038# a_3371_23106# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.147 ps=1.19 w=0.84 l=0.15
X4694 a_7284_20787# sar9b_0.net56 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4695 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4696 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4697 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4698 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4699 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4700 a_10644_16791# sar9b_0.net6 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4701 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4702 single_9b_cdac_0.SW[2] a_13067_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X4703 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4704 VGND a_4812_21738# sar9b_0.net65 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4705 a_5711_17527# a_5322_17846# a_5046_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4706 a_11722_25838# sar9b_0.net74 a_12243_25898# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4707 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4708 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4709 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4710 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4711 VGND a_11859_20574# single_9b_cdac_1.SW[8] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4712 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4713 a_4561_24464# sar9b_0.net58 a_4467_24162# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1312 pd=1.05 as=0.1824 ps=1.85 w=0.64 l=0.15
X4714 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4715 VGND sar9b_0.clknet_0_CLK a_2508_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4716 a_10500_19235# a_10239_19235# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4717 VGND sar9b_0.net38 a_10803_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4718 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4719 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4720 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4721 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4722 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4723 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4724 a_5581_19664# sar9b_0._07_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X4725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4726 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X4727 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4728 a_10402_25094# a_10218_24802# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4729 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4730 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4731 tdc_0.phase_detector_0.INN a_16527_10454# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X4732 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4733 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4734 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4735 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4736 VDPWR sar9b_0.net41 a_9130_26198# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4737 VGND a_5298_24499# a_5100_24375# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4738 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4739 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4740 single_9b_cdac_1.CF[8] a_13011_25902# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4741 VGND sar9b_0.net5 a_13011_20574# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4742 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4743 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4744 single_9b_cdac_1.CF[0] a_13011_20574# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4746 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4747 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4748 VDPWR a_10218_21842# a_10470_21795# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X4749 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4750 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4751 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4752 VDPWR a_9132_7271# th_dif_sw_0.th_sw_1.CK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4753 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4754 VDPWR a_11776_21141# sar9b_0.net8 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4755 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4756 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4757 a_10708_24151# a_9730_24138# a_10506_24506# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4758 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4759 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4760 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4761 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4762 VDPWR a_6132_23451# a_6137_23791# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4763 a_2603_17006# sar9b_0.net16 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X4764 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4765 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4766 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4767 a_3521_24240# a_3369_24181# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X4768 a_16542_13134# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X4769 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4770 VDPWR sar9b_0.net53 a_11382_23474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4771 VDPWR sar9b_0.net49 a_8982_21902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4772 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4773 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4774 a_6744_23534# a_6346_23773# a_6666_23534# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4775 a_12870_23599# a_12618_23470# a_13008_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4776 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4777 VDPWR a_6414_23681# a_6346_23773# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4778 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4779 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4780 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4781 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4782 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4783 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4784 VDPWR a_13011_27234# single_9b_cdac_0.SW[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4785 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4786 a_9264_23477# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4787 a_4168_22188# a_3027_22138# a_4011_22488# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X4788 VDPWR a_13011_16810# single_9b_cdac_1.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4789 a_43540_16877# single_9b_cdac_1.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4790 a_41357_15501# single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4792 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4793 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4794 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4795 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4796 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4797 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4798 a_11191_18859# a_10762_18823# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4799 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4800 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4801 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4802 a_8554_26437# a_8340_26115# a_7890_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4803 VDPWR sar9b_0.net5 a_7914_19178# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4804 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4805 VGND sar9b_0.net3 a_2547_28132# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4806 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4807 a_7433_27849# a_6954_27466# a_7343_27849# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4808 a_34814_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4809 a_8098_18810# a_7914_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4810 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4812 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4813 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4814 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4815 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4816 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4817 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4818 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4819 a_6666_23534# sar9b_0.net54 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X4820 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4821 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4822 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4823 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4824 a_62748_26999# single_9b_cdac_0.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4825 VGND a_10035_19474# sar9b_0.net48 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X4826 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4827 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4828 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4829 a_3370_26437# a_3156_26115# a_2706_26108# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4830 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4831 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4832 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4833 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4834 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4835 VGND a_4365_25770# a_4293_25852# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.10905 ps=1.025 w=0.55 l=0.15
X4836 a_3372_25734# sar9b_0._16_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4837 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4838 single_9b_cdac_1.CF[3] a_13011_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4839 VDPWR a_11915_28371# uo_out[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4840 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4841 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4842 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4843 VGND a_9760_22819# sar9b_0.net41 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4844 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4845 a_7238_21225# a_6975_20813# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4846 a_5633_20244# a_5481_20185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X4847 a_7743_18149# a_7602_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4848 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4849 a_12647_27128# sar9b_0.net52 a_12560_27128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4850 VDPWR a_12435_20806# single_9b_cdac_1.CF[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4851 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4852 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4853 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4854 a_12870_22267# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4855 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4856 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4857 single_9b_cdac_0.SW[1] a_13011_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X4858 single_9b_cdac_1.SW[7] a_13011_19242# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4859 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4860 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4861 VGND a_5010_28495# a_4812_28371# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4862 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4863 a_12047_22521# a_11842_22430# a_11382_22142# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4864 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4865 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4867 VGND a_12870_23599# a_12828_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4868 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4869 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4870 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4871 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4872 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4874 a_6538_24506# a_5753_24250# a_6030_24396# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4875 a_12047_23853# a_11658_23470# a_11382_23474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4876 VDPWR a_6738_22112# a_6540_22112# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X4877 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4878 single_9b_cdac_0.SW[3] a_12491_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X4879 VDPWR sar9b_0.net58 a_3231_27227# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4880 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4881 a_8940_24402# sar9b_0.net2 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4882 a_12064_22819# a_11466_23174# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4884 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4885 a_3372_25734# sar9b_0._16_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4886 VDPWR sar9b_0.clk_div_0.COUNT\[2\] sar9b_0._17_ VDPWR sky130_fd_pr__pfet_01v8 ad=0.42 pd=2.99 as=0.168 ps=1.42 w=1.12 l=0.15
X4887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4888 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4889 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4890 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4891 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4892 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4893 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4894 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4895 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4896 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X4897 VGND a_10859_26330# single_9b_cdac_0.SW[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X4898 VGND a_3090_27163# a_2892_27039# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4899 a_10320_20567# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4900 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4901 a_5083_21100# sar9b_0._17_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X4902 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4903 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4904 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4905 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4906 sar9b_0.net18 a_2508_27440# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4907 VDPWR sar9b_0.net58 a_2847_27473# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4908 sar9b_0.net3 a_2451_27234# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4909 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4910 VDPWR a_4044_24776# sar9b_0.net72 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4911 a_12828_23477# a_11658_23470# a_12618_23470# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4912 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4913 th_dif_sw_0.CK a_10227_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4914 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4915 uo_out[6] a_8115_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4916 a_29134_26999# single_9b_cdac_0.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4917 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4918 VDPWR a_12182_26419# a_12137_26517# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4919 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4920 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4921 a_3438_26345# a_3161_26455# a_3768_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4922 a_2540_22432# sar9b_0._12_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X4923 a_7140_22145# a_6879_22145# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X4924 a_10239_19235# a_10098_19171# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4925 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4926 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4927 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4928 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4929 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4930 a_8294_26553# a_8031_26141# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4931 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4932 a_2706_27440# a_3161_27787# a_3110_27885# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X4933 a_5580_24776# sar9b_0._15_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4934 a_8842_16874# a_8052_16791# a_8334_17021# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4935 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4936 single_9b_cdac_0.SW[6] a_9323_28371# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4937 VGND sar9b_0.net52 a_10029_24806# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4938 a_12618_18142# a_11658_18142# a_12182_18427# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4939 a_6534_17799# a_6282_17846# a_6672_17903# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4940 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4941 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4942 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4943 uio_out[1] a_2931_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4944 a_4749_27652# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X4945 a_13008_26141# sar9b_0.net52 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4946 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4947 VDPWR a_3603_28156# sar9b_0.net59 VDPWR sky130_fd_pr__pfet_01v8 ad=0.756 pd=3.59 as=0.168 ps=1.42 w=1.12 l=0.15
X4948 VDPWR a_5938_22378# a_5846_22572# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4949 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4950 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4951 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4952 VDPWR sar9b_0.net48 a_10830_19068# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X4953 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4954 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4955 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4956 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4957 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4958 a_11430_24931# a_11178_24802# a_11568_24809# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4959 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4960 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4961 a_3110_26553# a_2847_26141# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X4962 a_3768_26198# a_3370_26437# a_3690_26198# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4963 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4964 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4965 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4966 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4967 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4968 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4969 VGND sar9b_0.net24 a_10995_28566# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4970 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4971 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4972 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4973 a_3262_24141# sar9b_0.net70 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X4974 VGND sar9b_0.net49 a_9558_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4975 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4976 uo_out[2] a_10995_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4977 single_9b_cdac_1.SW[2] a_8019_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4978 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4979 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4980 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4981 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4982 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4983 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4984 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4985 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4986 a_4851_27230# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4987 a_33936_26999# single_9b_cdac_0.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4988 VGND a_5441_22522# a_5459_22165# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X4989 sar9b_0.net36 a_9996_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4990 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4991 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4992 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4993 VDPWR sar9b_0.net48 a_5535_18149# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4994 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4995 a_10742_25087# a_10607_25185# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4996 a_12618_19474# a_11842_19766# a_12182_19759# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4997 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4998 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4999 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 a_62748_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5000 single_9b_cdac_1.SW[8] a_11859_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5001 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5002 VDPWR a_13011_20806# single_9b_cdac_1.CF[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5003 a_8166_27595# sar9b_0.net60 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5004 a_6966_22145# a_6738_22112# a_6879_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5005 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5006 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5007 a_11915_27039# sar9b_0.net30 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X5008 a_9558_20510# a_9494_20290# a_9480_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5009 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5010 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5011 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5012 a_4771_18260# sar9b_0.net57 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X5013 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5014 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5015 a_11568_20813# sar9b_0.net49 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5016 a_8842_18206# sar9b_0.net46 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5017 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5018 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5019 a_9730_24138# a_9546_24506# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5020 single_9b_cdac_1.CF[1] a_12435_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5021 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5022 a_21177_7457# th_dif_sw_0.CKB VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.11655 ps=1.055 w=0.74 l=0.15
X5023 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5024 single_9b_cdac_0.SW[2] a_13067_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5025 single_9b_cdac_0.SW[5] a_11339_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5026 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5027 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5028 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5029 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5030 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5031 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5032 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5033 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5034 a_10410_17846# a_9450_17846# a_9974_17626# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5035 a_9126_23599# a_8874_23470# a_9264_23477# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5036 a_8591_22855# a_8202_23174# a_7926_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5037 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5038 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5039 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5040 a_5674_28147# a_5460_28377# a_5010_28495# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5041 VGND single_9b_cdac_0.SW[1] a_58824_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5042 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5043 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5044 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5045 a_5460_28377# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5046 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5047 a_8098_18810# a_7914_19178# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5048 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5049 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5050 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5051 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5052 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5053 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5054 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5055 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5056 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5057 VGND single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5058 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5059 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5060 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5061 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5062 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5063 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5064 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5065 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5066 VDPWR a_13011_24570# single_9b_cdac_1.CF[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5067 single_9b_cdac_1.CF[5] a_13011_23238# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5068 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5069 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5070 a_5846_17626# a_5711_17527# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5071 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5072 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5073 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5074 VGND sar9b_0.clk_div_0.COUNT\[2\] a_7597_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5075 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5076 a_7306_19777# a_7092_19455# a_6642_19448# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5077 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5078 sar9b_0.net11 a_5484_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5079 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5080 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5081 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5082 a_9359_20191# sar9b_0.net49 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5083 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5084 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5085 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5086 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5087 VDPWR a_3090_27163# a_2892_27039# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X5088 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5089 VGND a_9323_28371# single_9b_cdac_0.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X5090 a_11915_28371# sar9b_0.net14 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X5091 uo_out[5] a_7539_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5092 a_10378_27170# a_9588_27045# a_9870_27060# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5093 a_11466_23174# a_10506_23174# a_11030_22954# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5094 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5095 VGND a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5096 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5097 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5098 VGND sar9b_0.net13 a_13011_25902# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5099 VDPWR a_12618_22138# a_12870_22267# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5100 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5101 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5102 a_8074_20870# sar9b_0.net9 a_8595_20810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5103 a_10335_16817# a_10194_16784# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5104 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5105 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5106 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5107 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5108 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5109 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5110 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5111 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5112 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5113 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5114 VGND single_9b_cdac_0.SW[0] a_63626_26990# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5115 a_7597_23174# sar9b_0.net63 a_7483_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X5116 a_9647_21523# a_9442_21474# a_8982_21902# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5117 a_10140_20567# a_8970_20510# a_9930_20510# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5118 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5119 a_10070_24286# a_9935_24187# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5120 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5121 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5122 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5123 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5124 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5125 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5126 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5127 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5128 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5129 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5130 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5131 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5132 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5133 VDPWR sar9b_0.net60 a_3603_28156# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.32 ps=2.64 w=1 l=0.15
X5134 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5135 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5136 VGND sar9b_0.net55 a_7347_24160# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X5137 VGND sar9b_0.net49 a_9846_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5138 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5139 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5140 sar9b_0.net58 a_4749_27652# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.756 ps=3.59 w=1.12 l=0.15
X5141 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5142 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y a_35519_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5143 a_4673_24464# sar9b_0._13_ a_4561_24464# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.045 as=0.1312 ps=1.05 w=0.64 l=0.15
X5144 a_11856_23231# sar9b_0.net53 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5145 a_10182_20463# a_9930_20510# a_10320_20567# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5146 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5147 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5148 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5149 VDPWR a_21177_7457# th_dif_sw_0.th_sw_1.CKB VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5150 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5151 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5152 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5153 a_8595_20810# sar9b_0.net47 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5154 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5155 a_12618_22138# a_11658_22138# a_12182_22423# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5156 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A a_26951_15501# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5157 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5158 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5159 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5160 VDPWR sar9b_0.net73 a_6634_18206# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5161 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5162 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5163 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5164 a_25915_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5165 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 a_33936_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5166 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X5167 single_9b_cdac_0.SW[7] a_10859_26330# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X5168 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5169 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5170 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5171 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5172 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5173 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5174 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5175 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5176 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5177 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5178 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5179 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5180 a_53154_26999# single_9b_cdac_0.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5181 VDPWR sar9b_0.net48 a_10926_17021# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5182 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5183 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5184 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5185 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5186 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5187 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5188 a_9442_21474# a_9258_21842# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5189 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5190 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5191 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5192 VGND a_9414_23127# a_9372_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5193 sar9b_0._05_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5194 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5195 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5196 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5197 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5198 VDPWR sar9b_0.net46 a_7743_16817# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5199 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5200 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5201 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B a_16555_12124# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5202 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5203 a_12618_23470# a_11842_23762# a_12182_23755# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5204 a_6672_27227# sar9b_0.net58 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5205 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5206 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5207 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5208 a_6922_23534# sar9b_0.net54 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5209 a_8726_22954# a_8591_22855# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5210 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5211 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5212 a_9130_26198# sar9b_0.net41 a_9651_26138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5213 sar9b_0._15_ a_4467_24162# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.36323 ps=1.84 w=1.12 l=0.15
X5214 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5215 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5216 a_7188_22119# sar9b_0.net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5217 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5218 a_2847_26141# a_2706_26108# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5219 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5220 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5221 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5222 a_6058_18445# a_5844_18123# a_5394_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5223 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5224 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5225 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5226 VDPWR a_4332_23043# sar9b_0.clknet_0_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5227 VDPWR a_11466_23174# a_11718_23127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5228 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5229 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5230 VDPWR a_9760_22819# sar9b_0.net41 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5231 a_62748_16877# single_9b_cdac_1.SW[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5232 a_11430_24931# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5233 a_7978_22202# a_7188_22119# a_7470_22349# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5234 sar9b_0.net56 a_4771_18260# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5235 a_7602_16784# a_8057_17131# a_8006_17229# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5236 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5237 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5238 a_9372_23231# a_8202_23174# a_9162_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5239 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5240 single_9b_cdac_1.CF[1] a_12435_20806# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5241 a_12870_19603# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5242 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5243 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5244 sar9b_0.net59 a_3603_28156# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X5245 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5246 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5247 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5248 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5249 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5250 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5251 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5252 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5253 a_65367_15501# single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5254 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5255 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5256 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5257 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5258 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5259 a_3371_23106# a_3219_22860# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X5260 a_9414_23127# a_9162_23174# a_9552_23231# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5261 VDPWR sar9b_0.net8 a_11658_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5262 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5263 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5264 a_11178_27466# a_10218_27466# a_10742_27751# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5265 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5266 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5267 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5268 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X5269 VGND a_7284_20787# a_7289_21127# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X5270 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5271 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5272 a_3723_20140# a_2739_20140# a_3425_20244# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X5273 VGND a_10644_16791# a_10649_17131# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X5274 VGND sar9b_0.net47 a_5761_19487# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X5275 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5276 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5277 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5278 a_5846_26950# a_5711_26851# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5279 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5280 a_10025_24187# a_9546_24506# a_9935_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5281 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5282 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5283 a_9588_27045# sar9b_0.net45 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5284 a_40321_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5285 a_9449_20191# a_8970_20510# a_9359_20191# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5286 single_9b_cdac_0.SW[8] a_9323_27662# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5287 a_9472_23805# a_8874_23470# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5288 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5290 single_9b_cdac_1.SW[7] a_13011_19242# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5291 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5292 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5293 a_10644_16791# sar9b_0.net6 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5294 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5295 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5296 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5297 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5298 VGND sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X5299 VDPWR a_11008_17491# sar9b_0.net7 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5300 VDPWR a_4125_25958# a_4136_25584# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5301 a_8052_16791# sar9b_0.net5 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5302 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5303 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5304 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5305 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5306 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5307 VGND sar9b_0.net57 a_10218_24802# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5308 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5309 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5310 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5311 uo_out[5] a_7539_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5312 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5313 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5314 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5315 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5316 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5317 VGND a_9323_28371# single_9b_cdac_0.SW[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5318 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5319 VDPWR a_8874_19178# a_9126_19131# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5320 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5321 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5322 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5323 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5324 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5325 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5326 a_12246_18206# a_12182_18427# a_12168_18206# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5327 a_29134_16877# single_9b_cdac_1.SW[7] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5328 VGND a_5581_20992# sar9b_0._09_ VGND sky130_fd_pr__nfet_01v8_lvt ad=0.19322 pd=1.32 as=0.2109 ps=2.05 w=0.74 l=0.15
X5329 a_7498_21109# a_7289_21127# a_6834_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X5330 VDPWR a_8438_18958# a_8393_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5331 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5332 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5333 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5334 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5335 sar9b_0._02_ sar9b_0._12_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5336 VDPWR sar9b_0._04_ a_3027_21906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5337 VGND sar9b_0.net48 a_9261_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5338 a_10858_17113# a_10649_17131# a_10194_16784# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X5339 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5340 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5341 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5342 sar9b_0.clknet_1_1__leaf_CLK a_2508_23444# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5344 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5345 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5346 a_8726_22954# a_8591_22855# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5347 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5348 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5349 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5350 VGND a_4332_23043# sar9b_0.clknet_0_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5351 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5352 VGND a_8115_28566# uo_out[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5353 VDPWR a_11776_27801# sar9b_0.net25 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5354 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5355 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5356 a_10410_17846# a_9634_17478# a_9974_17626# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5357 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5358 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5359 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5360 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5361 a_12168_18206# a_11842_18434# a_12047_18525# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5362 a_30717_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5363 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5364 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5365 single_9b_cdac_1.SW[1] a_10803_19474# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5366 a_10502_18823# a_10239_19235# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5367 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5368 a_8393_18859# a_7914_19178# a_8303_18859# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5369 VDPWR sar9b_0.net56 a_5322_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5370 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5371 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5372 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5373 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5374 a_4698_25851# a_4125_25958# a_4365_25770# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.07875 ps=0.865 w=0.42 l=0.15
X5375 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5376 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5377 VGND a_2931_28566# uio_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5378 uo_out[7] a_5235_27466# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5380 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5381 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5382 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5383 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5384 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5385 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5386 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5387 a_3946_26198# sar9b_0.net59 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5388 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5389 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5390 a_33936_16877# single_9b_cdac_1.SW[6] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5391 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5392 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5393 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5394 a_60565_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5395 VDPWR sar9b_0._14_ a_2940_25096# VDPWR sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X5396 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5397 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5398 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5399 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5400 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5401 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5402 VGND ui_in[0] a_2451_27234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X5403 a_11339_27039# sar9b_0.net31 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X5404 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5405 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5406 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5407 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5408 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5409 a_36555_15501# single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5410 dw_12589_1395# a_10166_3438# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5411 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5412 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5413 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5414 VDPWR a_4018_24235# a_3926_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X5415 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5416 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5417 VDPWR sar9b_0.net42 a_13011_19242# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5418 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5419 VDPWR sar9b_0.net36 a_3946_27530# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5420 a_30012_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5421 VDPWR sar9b_0.net59 a_8031_26141# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5422 single_9b_cdac_1.SW[3] a_10803_18142# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5423 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5424 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5425 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5426 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5427 VDPWR a_12870_18271# a_12820_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X5428 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5429 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5430 VGND sar9b_0.net39 a_11859_17910# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5431 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5432 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5433 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5434 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.B VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X5435 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5436 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5437 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5438 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5439 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5440 a_57946_26999# single_9b_cdac_0.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5441 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5442 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5443 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5444 a_6534_27123# a_6282_27170# a_6672_27227# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5445 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5446 VGND a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5447 single_9b_cdac_1.CF[0] a_13011_20574# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5448 a_8874_19178# a_8098_18810# a_8438_18958# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5449 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5451 a_48343_26999# single_9b_cdac_0.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5453 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5454 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5455 a_4236_21738# sar9b_0._05_ VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5456 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5457 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5458 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5459 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5460 a_7914_27466# a_7138_27758# a_7478_27751# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5461 a_6484_26815# a_5506_26802# a_6282_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5462 sar9b_0.clknet_0_CLK a_4332_23043# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5463 sar9b_0.net46 a_6579_18832# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X5464 a_3206_22432# a_3027_22138# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5465 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5466 VDPWR sar9b_0.net11 a_11658_23470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5467 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5468 VGND a_13216_26469# sar9b_0.net33 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5469 a_5748_24381# sar9b_0.net13 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5470 VGND a_3922_20239# a_3880_20524# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X5471 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5472 VDPWR sar9b_0.net20 a_8115_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5473 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5474 VDPWR a_12618_19474# a_12870_19603# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5475 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5476 VGND sar9b_0.net53 a_10134_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5477 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5478 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5479 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5480 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5481 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5482 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5483 a_10758_24459# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5484 single_9b_cdac_1.SW[0] a_8595_17910# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5485 VGND a_8691_28566# uo_out[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5486 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5487 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5488 a_8334_17021# a_8057_17131# a_8664_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5489 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5490 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5491 VDPWR sar9b_0.clknet_0_CLK a_2508_20780# VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5492 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5493 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5494 a_3839_23194# sar9b_0.clk_div_0.COUNT\[2\] a_3725_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.1344 ps=1.06 w=0.64 l=0.15
X5495 sar9b_0.net6 a_7404_18116# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5496 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5497 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5498 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5499 VGND single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5500 VGND a_7539_28566# uo_out[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5501 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5502 VDPWR a_12684_20379# sar9b_0.net50 VDPWR sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5503 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5504 a_3454_22567# sar9b_0.net67 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X5505 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5506 VDPWR ui_in[0] a_2451_27234# VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5507 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5508 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5509 a_12246_22202# a_12182_22423# a_12168_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5510 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5511 a_9364_22819# a_8386_22806# a_9162_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5512 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5513 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5514 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5515 a_8664_16874# a_8266_17113# a_8586_16874# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5516 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5517 VDPWR sar9b_0.net56 a_9450_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5518 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5519 VDPWR sar9b_0.net37 a_4330_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5520 VDPWR a_3819_24136# a_4018_24235# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X5521 VGND a_11776_21141# sar9b_0.net8 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5522 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5523 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5524 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5525 single_9b_cdac_0.SW[4] a_11915_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5526 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5527 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5528 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5529 a_31753_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5530 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5531 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5532 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5533 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5534 a_12168_22202# a_11842_22430# a_12047_22521# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5535 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5536 a_6922_23534# a_6137_23791# a_6414_23681# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X5537 a_3273_20185# a_2918_20140# a_3166_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X5538 a_5622_18149# a_5394_18116# a_5535_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5539 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5540 VDPWR a_8940_24402# sar9b_0.net62 VDPWR sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5541 VGND a_6130_20239# a_6088_20524# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X5542 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5543 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5544 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5545 VDPWR a_11915_27039# single_9b_cdac_0.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5546 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5547 a_8586_16874# sar9b_0.net46 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X5548 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5549 sar9b_0._06_ a_12560_27128# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X5550 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5551 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5552 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5553 VGND a_8595_17910# single_9b_cdac_1.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5554 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5555 a_53154_16877# single_9b_cdac_1.SW[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5556 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5557 single_9b_cdac_0.cdac_sw_9b_0.S[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5558 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5559 a_10402_25094# a_10218_24802# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5560 VGND sar9b_0.net12 a_9546_24506# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5561 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5562 VGND a_5931_20140# a_6130_20239# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X5563 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5564 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5565 VGND sar9b_0.net55 a_5811_19178# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15198 pd=1.17 as=0.24915 ps=2.37 w=0.55 l=0.15
X5566 sar9b_0.clk_div_0.COUNT\[2\] a_4018_24235# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X5567 a_12137_18525# a_11658_18142# a_12047_18525# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5568 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y a_59529_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5569 VGND a_4749_27652# sar9b_0.net58 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X5570 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5571 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5572 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5573 sar9b_0.net48 a_10035_19474# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5574 a_3090_27163# a_3545_26914# a_3494_26815# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5575 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5576 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5577 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5578 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5579 a_12182_19759# a_12047_19857# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5580 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5581 VGND th_dif_sw_0.CKB a_21177_7457# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5582 a_3822_27060# a_3540_27045# a_4183_26851# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5583 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X5584 a_14897_9355# clk a_14871_9671# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5585 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5586 VDPWR sar9b_0.net54 a_5823_23477# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5587 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5588 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5589 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 a_57946_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5590 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5591 VDPWR sar9b_0.net74 a_11722_25838# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5592 a_11436_17742# sar9b_0.net2 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5593 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5594 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5595 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5596 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5597 VDPWR sar9b_0.net10 a_13011_23238# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5598 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5599 VGND a_12435_24802# single_9b_cdac_1.CF[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5600 a_6252_19074# sar9b_0.net15 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5601 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5602 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5603 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5604 a_4332_23043# clk VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X5605 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5606 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5607 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5608 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5609 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5610 a_4011_22488# a_3027_22138# a_3713_22522# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X5611 a_11338_19178# sar9b_0.net61 a_11859_19238# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5612 sar9b_0.net52 a_9165_24988# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.756 ps=3.59 w=1.12 l=0.15
X5613 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5614 a_5682_23444# a_6137_23791# a_6086_23889# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5615 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5616 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5617 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_26999# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5618 VDPWR sar9b_0.net52 a_11214_25728# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5619 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5620 uo_out[3] a_9939_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5621 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5622 a_9870_27060# a_9593_26914# a_10200_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5623 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5624 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5625 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5626 VGND a_8115_28566# uo_out[6] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5627 a_4183_26851# a_3754_26815# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X5628 sar9b_0.net57 a_5443_19074# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5629 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5630 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5631 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5632 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5633 a_9588_27045# sar9b_0.net45 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5634 a_12820_26553# a_11842_26426# a_12618_26134# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5635 a_16555_12412# tdc_0.phase_detector_0.pd_out_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5636 VGND single_9b_cdac_1.SW[1] a_58824_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5637 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5638 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5639 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5640 VDPWR sar9b_0.net68 a_3364_25120# VDPWR sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5641 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5642 a_10607_27849# a_10402_27758# a_9942_27470# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5643 sar9b_0.clknet_0_CLK a_4332_23043# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5644 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5645 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5646 VGND sar9b_0._07_ a_3795_19512# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14457 pd=1.15 as=0.15675 ps=1.67 w=0.55 l=0.15
X5647 VGND single_9b_cdac_1.SW[6] a_34814_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5648 a_7470_22349# a_7188_22119# a_7831_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5649 a_11859_19238# sar9b_0.net48 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5650 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5651 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5652 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5653 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5654 a_38738_26999# single_9b_cdac_0.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5655 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5656 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5657 VGND a_2931_28566# uio_out[1] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5658 VDPWR a_13011_25902# single_9b_cdac_1.CF[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5659 a_8334_17021# a_8052_16791# a_8695_17193# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X5660 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5661 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5662 VDPWR a_13011_20574# single_9b_cdac_1.CF[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5663 a_12047_19857# sar9b_0.net50 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5664 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5665 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5666 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5667 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5668 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5669 VDPWR sar9b_0.net46 a_5046_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X5670 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5671 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5672 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5673 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5674 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5675 VDPWR a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5676 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5677 a_6132_23451# sar9b_0.net57 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5678 a_6880_17491# a_6282_17846# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5679 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5680 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5681 VDPWR single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5682 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5683 a_5394_18116# a_5849_18463# a_5798_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5684 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5685 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5686 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5687 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5688 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5689 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5690 a_43540_26999# single_9b_cdac_0.SW[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5691 a_13216_26469# a_12618_26134# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5692 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5693 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5694 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5695 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5696 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5697 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5698 a_8695_17193# a_8266_17113# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X5699 single_9b_cdac_1.SW[5] a_13011_16810# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5700 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5701 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5702 single_9b_cdac_0.SW[7] a_10859_26330# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5703 a_64331_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5704 a_5133_17906# sar9b_0.net46 a_5046_17906# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5705 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5706 VGND single_9b_cdac_1.SW[0] a_63626_17740# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5707 a_63626_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5708 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5709 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5710 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5711 VDPWR a_10070_24286# a_10025_24187# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5712 VGND a_8019_17910# single_9b_cdac_1.SW[2] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5713 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5714 VGND sar9b_0.net57 a_9258_21842# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5716 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5717 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5718 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5719 uo_out[4] a_8691_28566# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5720 VGND a_3425_20244# a_3443_20547# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X5721 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5722 VGND sar9b_0.net19 a_5235_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5723 a_4812_21738# sar9b_0.clk_div_0.COUNT\[3\] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5724 th_dif_sw_0.th_sw_1.CK a_9132_7271# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5726 uio_out[0] a_4083_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5727 sar9b_0.net19 a_2892_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5728 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5729 VGND a_9363_20826# sar9b_0.net49 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5730 VGND sar9b_0.net40 a_13011_16810# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5731 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5732 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5733 single_9b_cdac_1.SW[4] a_11859_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5734 a_9132_7271# th_dif_sw_0.CK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5735 sar9b_0._16_ a_2893_24992# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X5736 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5737 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5738 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5739 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1764 ps=1.26 w=0.84 l=0.15
X5740 a_11434_16874# a_10644_16791# a_10926_17021# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5741 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5742 a_10607_25185# sar9b_0.net52 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5743 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5744 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5745 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5746 VGND a_13011_24802# single_9b_cdac_0.SW[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5747 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 a_29134_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5748 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5749 VDPWR sar9b_0.net46 a_7743_18149# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5750 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5751 VDPWR a_11915_27039# single_9b_cdac_0.SW[4] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5752 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5753 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5754 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5755 single_9b_cdac_1.CF[1] a_12435_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5756 VDPWR a_3425_20244# a_3380_20145# VDPWR sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X5757 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5758 VGND single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5759 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5760 a_9651_26138# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5761 a_7470_22349# a_7193_22459# a_7800_22202# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5762 sar9b_0.net37 a_9900_19047# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5763 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5764 a_9323_28371# sar9b_0.net32 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X5765 VDPWR a_13011_19242# single_9b_cdac_1.SW[7] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5766 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5767 a_10254_2858# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X5768 single_9b_cdac_1.CF[8] a_13011_25902# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5769 a_12137_22521# a_11658_22138# a_12047_22521# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5770 VGND sar9b_0.cyclic_flag_0.FINAL a_8883_27466# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5771 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5772 VGND a_13011_23238# single_9b_cdac_1.CF[5] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5773 VDPWR sar9b_0.net58 a_3822_27060# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5774 VGND sar9b_0.net48 a_5622_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X5775 a_7602_18116# a_8057_18463# a_8006_18561# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5776 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5777 a_7338_24802# a_6378_24802# a_6902_25087# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5778 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5779 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5780 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5781 a_12182_23755# a_12047_23853# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5782 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5783 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5784 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5785 VDPWR a_7284_20787# a_7289_21127# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5786 a_12870_18271# a_12618_18142# a_13008_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5787 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5788 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5789 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5790 ua[4] th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10166_3438# VGND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X5791 a_17125_9355# clk a_16331_9671# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5792 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5793 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5794 VDPWR VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5795 VGND a_11859_17910# single_9b_cdac_1.SW[4] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5796 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5797 VGND sar9b_0._17_ a_4922_20857# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X5798 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5799 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5800 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5801 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5802 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5803 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5804 VDPWR clk a_16331_9671# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X5805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5806 VDPWR a_8334_17021# a_8266_17113# VDPWR sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X5807 a_57946_16877# single_9b_cdac_1.SW[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5808 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5809 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5811 VDPWR a_8115_28566# uo_out[6] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5812 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5813 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5814 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5815 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5816 a_48343_16877# single_9b_cdac_1.SW[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5817 sar9b_0.net19 a_2892_27039# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5818 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 a_38738_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5819 VDPWR sar9b_0.net48 a_10239_19235# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X5820 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5821 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5822 VDPWR sar9b_0.net21 a_7539_28566# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5823 VGND sar9b_0.net65 a_3839_23194# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15182 pd=1.125 as=0.1152 ps=1 w=0.64 l=0.15
X5824 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5825 uo_out[3] a_9939_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5826 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5827 VDPWR sar9b_0.net47 a_7566_21017# VDPWR sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5828 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5829 a_8874_19178# a_7914_19178# a_8438_18958# VDPWR sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5830 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5831 VGND sar9b_0.net58 a_5910_27170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5832 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y a_45123_29917# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5833 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5834 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5835 VDPWR a_2931_28566# uio_out[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5836 sar9b_0.net37 a_9900_19047# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5837 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5838 VGND a_9132_7271# th_dif_sw_0.th_sw_1.CK VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5839 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5840 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5841 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5842 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5843 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X5844 VGND sar9b_0.clknet_1_1__leaf_CLK a_4755_22138# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X5845 th_dif_sw_0.CKB a_2603_17006# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X5846 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5847 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5848 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5849 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5850 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5851 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5852 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5853 a_7062_20813# a_6834_20780# a_6975_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5854 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5856 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5857 a_11568_27473# sar9b_0.net59 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5858 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1739 ps=1.21 w=0.74 l=0.15
X5859 a_12047_23853# sar9b_0.net53 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5860 sar9b_0.clk_div_0.COUNT\[3\] a_4210_22378# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X5861 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5862 VGND a_12870_18271# a_12828_18149# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5863 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5864 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5865 a_5010_28495# a_5460_28377# a_5412_28559# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X5866 VDPWR a_10995_28566# uo_out[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5867 a_4365_25770# a_4136_25584# a_4531_25875# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.0441 ps=0.63 w=0.42 l=0.15
X5868 VDPWR a_8019_17910# single_9b_cdac_1.SW[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5869 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5870 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5871 a_9472_18823# a_8874_19178# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5872 a_12047_18525# a_11658_18142# a_11382_18146# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5873 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5874 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5875 VDPWR sar9b_0.net44 a_5322_27170# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5876 VGND VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5877 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5878 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5879 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X5880 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5882 a_6834_20780# a_7284_20787# a_7236_20813# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X5883 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 a_43540_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5884 uo_out[6] a_8115_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5885 VDPWR sar9b_0.net19 a_5235_27466# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X5886 a_6678_27470# sar9b_0.net40 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5888 VGND a_11915_28371# uo_out[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X5889 single_9b_cdac_1.CF[3] a_13011_20806# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5890 a_38738_16877# single_9b_cdac_1.SW[5] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5891 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5892 VDPWR a_7914_27466# a_8166_27595# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5893 VGND sar9b_0.net54 a_8790_23174# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5894 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5895 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5896 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5897 single_9b_cdac_0.SW[4] a_11915_27039# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X5898 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5899 VGND a_12435_24802# single_9b_cdac_1.CF[7] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X5900 VGND sar9b_0.net49 a_10035_19474# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X5901 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5902 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5903 a_5412_28559# a_5151_28559# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X5904 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5905 sar9b_0.clknet_1_0__leaf_CLK a_2508_20780# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5906 a_12828_18149# a_11658_18142# a_12618_18142# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5907 VGND sar9b_0.net58 a_5133_27230# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5908 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5909 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5910 VDPWR sar9b_0.net5 a_8842_18206# VDPWR sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5911 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5912 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5913 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5914 a_11722_25838# a_10932_25713# a_11214_25728# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5915 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5916 a_5761_21100# sar9b_0._08_ VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2382 ps=1.555 w=1 l=0.15
X5917 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A a_35519_15495# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5918 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5919 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.S[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5920 VDPWR a_11339_27039# single_9b_cdac_0.SW[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5921 a_24332_26999# single_9b_cdac_0.SW[8] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5922 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5923 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5924 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5925 a_6086_23889# a_5823_23477# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5926 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5928 a_10710_25895# a_10482_25831# a_10623_25895# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X5929 a_4922_20857# sar9b_0.net65 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X5930 a_10528_20155# a_9930_20510# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5931 a_25915_15495# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5932 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5933 VDPWR sar9b_0.net11 a_8202_23174# VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5934 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5935 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5936 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5937 uo_out[1] a_12531_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5938 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5939 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5940 a_49221_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5941 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5942 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5943 a_13216_22473# a_12618_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5944 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5945 a_2508_23444# sar9b_0.clknet_0_CLK VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5946 a_3206_22432# a_3027_22138# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X5947 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5948 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5949 uo_out[2] a_10995_28566# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5950 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5951 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5952 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5953 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5954 single_9b_cdac_1.CF[6] a_13011_24570# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5955 a_6783_19481# a_6642_19448# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X5956 VDPWR a_6880_17491# sar9b_0.net5 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5957 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5958 VDPWR tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X5959 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5960 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5961 VDPWR a_13011_23238# single_9b_cdac_1.CF[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5963 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5964 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5965 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5966 VGND a_6579_18832# sar9b_0.net46 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5967 a_8266_18445# a_8052_18123# a_7602_18116# VDPWR sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5968 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5969 dw_17224_1400# a_21368_4076# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5970 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5971 VDPWR single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VDPWR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5972 VDPWR a_13216_19809# sar9b_0.net29 VDPWR sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5973 VGND sar9b_0.net54 a_8013_23234# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5974 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5975 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5976 a_3926_24136# a_3014_24136# a_3819_24136# VDPWR sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X5977 a_4292_19768# sar9b_0.net46 a_4072_19474# VDPWR sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.195 ps=1.39 w=1 l=0.15
X5978 a_7882_19538# sar9b_0.net62 a_8403_19478# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5979 single_9b_cdac_1.SW[2] a_8019_17910# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5980 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5981 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5982 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5983 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5984 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5985 VDPWR a_7539_28566# uo_out[5] VDPWR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5986 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5987 a_11104_24151# a_10506_24506# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5988 a_12870_22267# a_12618_22138# a_13008_22145# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5989 a_10612_17491# a_9634_17478# a_10410_17846# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5990 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5991 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5992 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# a_15265_9613# VDPWR sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X5993 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDPWR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5994 VGND sar9b_0.net60 a_3603_28156# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X5995 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5996 VGND a_6834_20780# a_6636_20780# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5997 a_5711_17527# a_5506_17478# a_5046_17906# VDPWR sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5998 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5999 a_10742_25087# a_10607_25185# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6000 a_5798_18561# a_5535_18149# VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X6001 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6002 a_11380_21225# a_10402_21098# a_11178_20806# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X6003 VDPWR sar9b_0.net48 a_10335_16817# VDPWR sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X6004 ua[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6005 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6006 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6007 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_53154_16877# VDPWR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6008 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6009 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6010 VGND single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6011 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6012 a_9737_21523# a_9258_21842# a_9647_21523# VDPWR sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X6013 VDPWR sar9b_0.net35 a_8595_17910# VDPWR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X6014 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6015 VGND single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6016 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6017 VGND a_4125_25958# a_4136_25584# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2553 ps=2.17 w=0.74 l=0.15
X6018 a_6282_17846# a_5506_17478# a_5846_17626# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X6019 th_dif_sw_0.VCP single_9b_cdac_1.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6020 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6021 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 single_9b_cdac_0.SW[6] uo_out[1] 0.04587f
C1 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.07579f
C2 sar9b_0._08_ sar9b_0._07_ 0.02717f
C3 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[8] 1.89002f
C4 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.36334f
C5 sar9b_0.net24 sar9b_0.net59 0.29571f
C6 a_7498_21109# sar9b_0.net10 0.03668f
C7 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.41793f
C8 sar9b_0.net49 a_9494_20290# 0.1204f
C9 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C10 sar9b_0.net72 a_4044_24776# 0.16551f
C11 VDPWR a_6880_26815# 0.20981f
C12 sar9b_0.net9 sar9b_0.net61 0.58982f
C13 sar9b_0.net13 sar9b_0.net53 0.0108f
C14 VDPWR sar9b_0.net30 0.61341f
C15 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C16 th_dif_sw_0.th_sw_1.CK ua[3] 0.42268f
C17 sar9b_0._13_ sar9b_0.net58 0.09533f
C18 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C19 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[8] 16.1938f
C20 sar9b_0.net38 a_10182_20463# 0.0163f
C21 single_9b_cdac_1.cdac_sw_9b_0.S[1] a_57946_16877# 0.59531f
C22 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[4] 0.26707f
C23 th_dif_sw_0.CK sar9b_0.net36 0.03321f
C24 a_4083_28566# sar9b_0.net59 0.10812f
C25 sar9b_0.net51 a_7443_21496# 0.28357f
C26 VDPWR a_10182_20463# 0.26691f
C27 VDPWR single_9b_cdac_1.SW[5] 2.51859f
C28 sar9b_0.net55 sar9b_0.net54 0.51028f
C29 sar9b_0.net56 sar9b_0.net57 0.1667f
C30 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.06503f
C31 a_9942_24806# sar9b_0.net38 0.01422f
C32 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C33 a_11382_19478# sar9b_0.net73 0.17436f
C34 a_10098_19171# sar9b_0.net48 0.29653f
C35 a_10548_19053# sar9b_0.net73 0.01967f
C36 VDPWR a_9942_24806# 0.28868f
C37 a_49926_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.01076f
C38 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22526f
C39 a_9939_28566# uo_out[3] 0.40366f
C40 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C41 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96978f
C42 a_7638_23474# sar9b_0.net62 0.01517f
C43 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] 1.15132f
C44 a_9900_19047# a_10098_19171# 0.06623f
C45 sar9b_0.net33 a_12618_26134# 0.07184f
C46 VDPWR a_7404_18116# 0.19099f
C47 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.12431f
C48 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[7] 0.06503f
C49 VDPWR a_10859_26330# 0.42645f
C50 a_9974_17626# a_10410_17846# 0.16939f
C51 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.62443f
C52 sar9b_0.net43 a_9935_24187# 0.09338f
C53 sar9b_0.net27 a_12870_26263# 0.0306f
C54 a_3161_26455# sar9b_0.net59 0.10291f
C55 a_8386_22806# a_9414_23127# 0.07826f
C56 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.81428f
C57 sar9b_0.net13 a_6562_25094# 0.12325f
C58 a_5682_23444# a_5823_23477# 0.27388f
C59 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.24288f
C60 a_5846_17626# a_6282_17846# 0.16939f
C61 VDPWR a_7890_26108# 0.33944f
C62 a_7404_17715# sar9b_0.net56 0.02799f
C63 a_7306_19777# sar9b_0.net35 0.01601f
C64 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[3] 0.02002f
C65 a_7602_18116# sar9b_0.net48 0.06506f
C66 sar9b_0.net7 sar9b_0.net9 0.36253f
C67 sar9b_0.net63 sar9b_0.net39 0.2717f
C68 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS ua[4] 0.93546f
C69 a_6879_22145# sar9b_0.net39 0.04509f
C70 sar9b_0.net26 a_12182_23755# 0.01551f
C71 VDPWR ua[0] 93.85329f
C72 sar9b_0.net44 a_3822_27060# 0.01345f
C73 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36044f
C74 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.02638f
C75 sar9b_0.net52 sar9b_0.net45 0.18401f
C76 a_6540_22112# sar9b_0._02_ 0.02465f
C77 sar9b_0.net7 sar9b_0.net61 0.28001f
C78 a_9546_24506# a_9730_24138# 0.43747f
C79 a_10402_21098# sar9b_0.net73 0.01426f
C80 a_11466_23174# a_12064_22819# 0.06623f
C81 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] 1.15113f
C82 sar9b_0.net35 clk 0.03859f
C83 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.62443f
C84 a_3946_27530# a_3156_27447# 0.1263f
C85 sar9b_0.net62 sar9b_0.net39 0.02577f
C86 a_11722_25838# sar9b_0.net31 0.01201f
C87 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[1] 1.81416f
C88 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.01152f
C89 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C90 VDPWR a_12047_26517# 0.26706f
C91 sar9b_0.net2 clk 0.03287f
C92 sar9b_0.net56 sar9b_0.net40 0.02195f
C93 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.12358f
C94 sar9b_0.net46 a_7914_19178# 0.07106f
C95 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0303f
C96 a_5083_21100# sar9b_0.net65 0.01754f
C97 a_2508_26108# a_2706_26108# 0.06623f
C98 a_8334_17021# sar9b_0.net5 0.01036f
C99 single_9b_cdac_1.SW[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.24456f
C100 a_5844_18123# a_5535_18149# 0.07766f
C101 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.10429f
C102 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.38397f
C103 a_7602_16784# a_7743_16817# 0.27388f
C104 a_8052_16791# a_8057_17131# 0.44098f
C105 a_5580_24776# sar9b_0._03_ 0.1431f
C106 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.81423f
C107 a_6678_27470# a_7138_27758# 0.26257f
C108 single_9b_cdac_1.SW[0] a_9174_17906# 0.04125f
C109 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[7] 0.21593f
C110 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.01175f
C111 a_21368_4076# th_dif_sw_0.CKB 0.01417f
C112 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[1] 0.22097f
C113 sar9b_0.net56 a_9174_17906# 0.04252f
C114 tdc_0.RDY tdc_0.OUTN 0.07358f
C115 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C116 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 1.71649f
C117 a_13011_20574# a_13216_19809# 0.01043f
C118 a_10607_25185# sar9b_0.net12 0.06942f
C119 a_3090_27163# a_3545_26914# 0.3578f
C120 uo_out[5] uo_out[6] 2.98352f
C121 a_8334_18353# sar9b_0.net5 0.06948f
C122 VDPWR a_10194_16784# 0.31773f
C123 sar9b_0.clknet_1_0__leaf_CLK a_3166_20145# 0.02652f
C124 a_11430_20935# a_11178_20806# 0.27388f
C125 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.10429f
C126 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.84061f
C127 a_11658_22138# a_12182_22423# 0.05022f
C128 a_8115_28566# uo_out[5] 0.03775f
C129 a_10932_25713# a_11214_25728# 0.06034f
C130 sar9b_0.net32 sar9b_0.net26 0.27199f
C131 sar9b_0.net32 single_9b_cdac_0.SW[7] 0.02288f
C132 VDPWR a_4496_20468# 0.33806f
C133 a_11382_19478# sar9b_0.net50 0.23074f
C134 a_10470_21795# a_10218_21842# 0.27388f
C135 a_10548_19053# sar9b_0.net50 0.02815f
C136 sar9b_0.net13 a_10932_25713# 0.23395f
C137 a_11146_25483# a_10937_25582# 0.24088f
C138 sar9b_0.net40 a_6902_25087# 0.0115f
C139 sar9b_0.net43 a_11859_20574# 0.20839f
C140 a_9126_23599# sar9b_0.net54 0.05162f
C141 sar9b_0.net15 a_5844_18123# 0.0119f
C142 a_7914_27466# a_8115_28566# 0.01021f
C143 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.38397f
C144 sar9b_0.net57 a_5394_18116# 0.02101f
C145 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C146 VDPWR a_2940_25096# 0.20267f
C147 ui_in[3] ui_in[2] 0.03102f
C148 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96835f
C149 sar9b_0.net26 sar9b_0.net51 0.02947f
C150 sar9b_0._07_ a_5523_21528# 0.18199f
C151 a_13011_19242# sar9b_0.net28 0.01241f
C152 single_9b_cdac_1.CF[0] single_9b_cdac_0.SW[0] 2.15297f
C153 sar9b_0.net5 single_9b_cdac_1.SW[2] 0.0302f
C154 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.363f
C155 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.62443f
C156 sar9b_0.net31 single_9b_cdac_1.CF[3] 0.01828f
C157 a_6540_22112# a_6879_22145# 0.07649f
C158 a_13011_24802# a_13011_24570# 0.02551f
C159 sar9b_0.net60 sar9b_0.net57 0.11607f
C160 sar9b_0.net48 a_7404_18116# 0.02507f
C161 sar9b_0.net49 sar9b_0.net2 0.02449f
C162 sar9b_0.net41 sar9b_0.net52 0.09293f
C163 sar9b_0.net60 a_5506_26802# 0.02734f
C164 VDPWR a_2547_28132# 0.36522f
C165 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.26942f
C166 a_13011_19242# single_9b_cdac_1.SW[7] 0.36033f
C167 VDPWR a_10410_17846# 0.32302f
C168 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.19147f
C169 sar9b_0.net43 sar9b_0.net51 0.39434f
C170 a_6130_20239# sar9b_0.net15 0.12036f
C171 sar9b_0._07_ sar9b_0._12_ 0.03077f
C172 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.24311f
C173 th_dif_sw_0.CK a_11382_18146# 0.05375f
C174 dw_12589_1395# th_dif_sw_0.CK 0.01665f
C175 sar9b_0.net38 a_9323_28371# 0.03711f
C176 a_8345_26455# a_8340_26115# 0.43491f
C177 VDPWR sar9b_0.net54 3.92712f
C178 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 1.71649f
C179 VDPWR a_9323_28371# 0.43901f
C180 sar9b_0.net12 a_11658_26134# 0.21062f
C181 sar9b_0._10_ a_5581_19664# 0.13526f
C182 a_8438_18958# sar9b_0.net61 0.0222f
C183 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C184 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[7] 0.01471f
C185 a_7882_19538# sar9b_0.net51 0.01799f
C186 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.01175f
C187 a_5322_27170# a_6534_27123# 0.07766f
C188 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.CF[3] 0.18985f
C189 VDPWR a_6834_20780# 0.32839f
C190 sar9b_0.net1 sar9b_0.net54 0.49885f
C191 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.71729f
C192 single_9b_cdac_1.SW[8] sar9b_0.net5 0.04994f
C193 a_58824_26990# single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22352f
C194 sar9b_0.net58 a_6534_27123# 0.17315f
C195 sar9b_0.net42 sar9b_0.net11 0.02571f
C196 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.CF[3] 0.105f
C197 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C198 a_7914_23470# clk 0.01168f
C199 VDPWR a_11776_21141# 0.20631f
C200 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[8] 1.08672f
C201 a_8386_22806# sar9b_0.net11 0.15667f
C202 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C203 a_8074_20870# sar9b_0.net62 0.01645f
C204 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[5] 0.0187f
C205 sar9b_0.net40 sar9b_0.net60 0.49844f
C206 a_21368_4076# th_dif_sw_0.th_sw_1.CKB 0.06647f
C207 sar9b_0._13_ a_4467_24162# 0.11876f
C208 sar9b_0.net53 sar9b_0.net62 0.14142f
C209 sar9b_0.net17 sar9b_0.net19 0.01908f
C210 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[2] 0.22184f
C211 sar9b_0._06_ clk 0.01579f
C212 a_11915_27039# sar9b_0.net30 0.22412f
C213 sar9b_0.net31 sar9b_0.net52 0.77905f
C214 sar9b_0.net26 sar9b_0.net12 0.02943f
C215 a_10553_18922# sar9b_0.net36 0.01892f
C216 sar9b_0.net41 a_9494_20290# 0.01451f
C217 sar9b_0.net8 a_11430_20935# 0.04729f
C218 a_15265_9613# th_dif_sw_0.VCP 0.10972f
C219 sar9b_0.net57 a_5443_19074# 0.25423f
C220 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.84082f
C221 a_5581_19664# sar9b_0.net4 0.01002f
C222 sar9b_0.net61 sar9b_0.net5 0.55611f
C223 a_10194_16784# sar9b_0.net48 0.24027f
C224 sar9b_0._11_ a_4947_20140# 0.14426f
C225 a_10230_23234# sar9b_0.net38 0.01802f
C226 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.22597f
C227 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C228 uo_out[5] uo_out[4] 2.90315f
C229 single_9b_cdac_0.cdac_sw_9b_0.S[4] th_dif_sw_0.VCN 13.5521f
C230 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[4] 0.12898f
C231 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.84426f
C232 VDPWR a_10230_23234# 0.30161f
C233 a_3713_22522# sar9b_0.clknet_1_1__leaf_CLK 0.04145f
C234 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.3196f
C235 a_6744_23238# sar9b_0.clk_div_0.COUNT\[1\] 0.02511f
C236 sar9b_0.net51 sar9b_0.net4 0.21881f
C237 VDPWR ui_in[0] 2.1737f
C238 a_8595_17910# sar9b_0.net35 0.20113f
C239 sar9b_0.net40 sar9b_0.net57 0.02758f
C240 VDPWR sar9b_0.net27 3.63493f
C241 a_38738_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.23864f
C242 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A a_59529_15495# 0.01076f
C243 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.22879f
C244 a_9363_20826# sar9b_0.net49 0.32854f
C245 sar9b_0.net43 sar9b_0.net12 0.38567f
C246 a_8334_17021# a_8842_16874# 0.19065f
C247 a_10762_18823# sar9b_0.net26 0.06684f
C248 VDPWR single_9b_cdac_0.SW[5] 2.59365f
C249 single_9b_cdac_1.cdac_sw_9b_0.S[7] ua[0] 1.97892f
C250 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.SW[4] 0.17175f
C251 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C252 single_9b_cdac_0.SW[3] ua[0] 0.16155f
C253 th_dif_sw_0.CKB clk 0.11297f
C254 a_10690_22806# sar9b_0.net31 0.01488f
C255 single_9b_cdac_0.SW[0] a_62748_26999# 0.28324f
C256 a_9930_20510# a_10182_20463# 0.27388f
C257 single_9b_cdac_0.cdac_sw_9b_0.S[7] th_dif_sw_0.VCN 1.61586f
C258 a_4947_20140# a_5374_20145# 0.04602f
C259 sar9b_0.net58 sar9b_0.net72 0.01694f
C260 a_4496_20468# sar9b_0.clknet_1_0__leaf_CLK 0.10004f
C261 sar9b_0.net1 sar9b_0.net27 0.07267f
C262 a_8970_20510# a_9154_20142# 0.43491f
C263 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.11216f
C264 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[8] 0.05215f
C265 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] 0.12898f
C266 sar9b_0.net36 a_10742_21091# 0.0132f
C267 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.81428f
C268 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.08121f
C269 sar9b_0.net21 uo_out[6] 0.34168f
C270 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02666f
C271 a_10742_25087# a_11178_24802# 0.16939f
C272 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.10984p
C273 a_10803_19474# sar9b_0.net73 0.03401f
C274 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.05472f
C275 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C276 sar9b_0.net48 a_10410_17846# 0.27687f
C277 a_8334_18353# a_8842_18206# 0.19065f
C278 single_9b_cdac_0.SW[1] a_58824_26990# 0.18991f
C279 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.11216f
C280 sar9b_0.net7 sar9b_0.net5 0.0215f
C281 th_dif_sw_0.th_sw_1.CKB a_10166_3438# 0.06536f
C282 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 3.10626f
C283 sar9b_0.net68 sar9b_0.clk_div_0.COUNT\[2\] 0.49269f
C284 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.12898f
C285 a_8019_17910# single_9b_cdac_1.SW[2] 0.35523f
C286 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.23864f
C287 sar9b_0.net60 uio_out[1] 0.27455f
C288 VDPWR a_3540_27045# 0.77744f
C289 a_5812_21028# sar9b_0._01_ 0.14953f
C290 a_6414_23681# sar9b_0.net11 0.02893f
C291 a_10402_27758# a_11430_27595# 0.07826f
C292 a_3540_27045# a_4330_27170# 0.1263f
C293 a_5682_23444# sar9b_0.net54 0.24995f
C294 a_8512_27801# sar9b_0.net45 0.03235f
C295 VDPWR a_13011_21906# 0.47029f
C296 single_9b_cdac_0.cdac_sw_9b_0.S[7] a_30012_26990# 0.22513f
C297 sar9b_0.net71 a_5196_19448# 0.14653f
C298 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.30106f
C299 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.net4 0.27294f
C300 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[2] 0.06503f
C301 sar9b_0.net69 sar9b_0.clk_div_0.COUNT\[1\] 0.04869f
C302 sar9b_0.net8 sar9b_0.net37 0.15963f
C303 sar9b_0.net65 a_4947_20140# 0.01364f
C304 sar9b_0.net10 a_7470_22349# 0.07606f
C305 single_9b_cdac_1.cdac_sw_9b_0.S[0] a_62748_16877# 0.59531f
C306 a_9935_24187# a_10070_24286# 0.35559f
C307 sar9b_0.net74 sar9b_0.net11 0.42192f
C308 sar9b_0.clk_div_0.COUNT\[2\] a_5580_24776# 0.02755f
C309 a_8622_26345# sar9b_0.cyclic_flag_0.FINAL 0.0786f
C310 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.12358f
C311 sar9b_0.net40 a_6861_22828# 0.01547f
C312 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C313 sar9b_0.net27 sar9b_0.net29 0.42418f
C314 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 1.55946f
C315 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[7] 0.42014f
C316 VDPWR a_11008_17491# 0.1898f
C317 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C318 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.26707f
C319 sar9b_0._18_ sar9b_0.clk_div_0.COUNT\[1\] 0.17343f
C320 sar9b_0.net36 sar9b_0.net38 0.92018f
C321 a_8202_23174# a_7926_23234# 0.1263f
C322 VDPWR sar9b_0.net36 1.87634f
C323 sar9b_0.net44 a_5711_26851# 0.06353f
C324 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] 3.10215f
C325 a_8052_16791# sar9b_0.net6 0.02602f
C326 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.969f
C327 a_7097_19795# a_7374_19685# 0.09983f
C328 sar9b_0.net40 a_12870_18271# 0.02062f
C329 a_59529_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.01076f
C330 sar9b_0.net48 sar9b_0.net27 0.34189f
C331 th_dif_sw_0.th_sw_1.CKB ua[3] 0.08416f
C332 single_9b_cdac_0.SW[1] th_dif_sw_0.VCN 0.09453f
C333 VDPWR single_9b_cdac_1.CF[4] 2.77384f
C334 th_dif_sw_0.th_sw_1.CKB clk 0.0198f
C335 a_7092_19455# a_7097_19795# 0.44098f
C336 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[2] 4.14971f
C337 a_6484_22845# sar9b_0._02_ 0.01922f
C338 single_9b_cdac_1.SW[8] a_12618_19474# 0.02801f
C339 VDPWR a_17125_9355# 0.01057f
C340 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C341 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.3601f
C342 sar9b_0.net20 a_5460_28377# 0.09259f
C343 a_5010_28495# a_5465_28246# 0.3578f
C344 sar9b_0.net1 sar9b_0.net36 0.01195f
C345 single_9b_cdac_1.CF[6] th_dif_sw_0.VCN 0.09453f
C346 sar9b_0.net35 a_7590_24931# 0.01235f
C347 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.19125f
C348 clk single_9b_cdac_1.SW[0] 0.21166f
C349 a_8019_17910# sar9b_0.net61 0.01405f
C350 a_11466_23174# sar9b_0.net53 0.28157f
C351 a_2892_23070# a_3219_22860# 0.09161f
C352 sar9b_0._18_ a_3371_23106# 0.05658f
C353 a_10690_22806# a_11718_23127# 0.07826f
C354 a_5846_17626# sar9b_0.net46 0.19277f
C355 a_8842_16874# sar9b_0.net61 0.2111f
C356 th_dif_sw_0.th_sw_1.CKB a_10254_2858# 0.42927f
C357 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.02618f
C358 sar9b_0.net41 sar9b_0.net2 0.36918f
C359 a_11030_22954# clk 0.01673f
C360 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[5] 1.26495f
C361 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[2] 17.4687f
C362 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.01175f
C363 a_10742_27751# a_10607_27849# 0.35559f
C364 ui_in[0] rst_n 0.03102f
C365 a_5322_27170# sar9b_0.net37 0.05304f
C366 a_7602_16784# sar9b_0.net27 0.05862f
C367 sar9b_0.net42 sar9b_0.net26 0.59576f
C368 sar9b_0.net42 single_9b_cdac_0.SW[7] 0.0472f
C369 sar9b_0.net55 sar9b_0.net51 0.50241f
C370 a_9279_27227# a_9593_26914# 0.07826f
C371 sar9b_0.net10 sar9b_0.clk_div_0.COUNT\[2\] 0.03438f
C372 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.36013f
C374 sar9b_0.net58 sar9b_0.net37 0.24097f
C375 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[4] 4.15153f
C376 a_8052_16791# sar9b_0.net46 0.1629f
C377 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.SW[4] 0.01837f
C378 a_48343_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.23864f
C379 VDPWR w_17430_1606# 0.44324f
C380 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.01003f
C381 VDPWR a_6534_17799# 0.26217f
C382 sar9b_0.net58 a_3438_27677# 0.2256f
C383 sar9b_0.net16 sar9b_0._00_ 0.01551f
C384 VDPWR a_3713_22522# 0.10433f
C385 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07517f
C386 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[8] 0.01285f
C387 sar9b_0.net43 sar9b_0.net42 0.4289f
C388 VDPWR a_3438_26345# 0.27271f
C389 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.17533f
C390 th_dif_sw_0.CK a_13216_18477# 0.04814f
C391 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.SW[7] 0.22983f
C392 VDPWR a_3922_20239# 0.38261f
C393 VDPWR a_9935_24187# 0.26083f
C394 sar9b_0.net64 a_6444_21738# 0.1416f
C395 sar9b_0.net23 a_8622_26345# 0.03011f
C396 a_14871_9671# a_15265_9613# 0.12812f
C397 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[4] 18.8692f
C398 sar9b_0.net45 sar9b_0._06_ 0.01013f
C399 sar9b_0.net40 a_6538_24506# 0.01312f
C400 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[8] 0.21771f
C401 a_8074_20870# a_7284_20787# 0.1263f
C402 single_9b_cdac_0.SW[6] uo_out[2] 0.04371f
C403 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.22609f
C404 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[3] 0.06162f
C405 sar9b_0.net36 a_8883_27466# 0.05427f
C406 sar9b_0.net24 sar9b_0.net36 0.37491f
C407 a_7638_23474# sar9b_0.net11 0.23589f
C408 VDPWR a_8057_18463# 0.24516f
C409 a_10858_17113# sar9b_0.net6 0.03245f
C410 a_12560_27128# VDPWR 0.33605f
C411 sar9b_0.net40 a_13011_17910# 0.02505f
C412 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_60565_15501# 0.01076f
C413 a_4332_23043# sar9b_0.clk_div_0.COUNT\[1\] 0.81462f
C414 VDPWR a_7478_27751# 0.20242f
C415 sar9b_0.net63 a_6484_22845# 0.05368f
C416 a_15151_10456# tdc_0.phase_detector_0.INP 0.10793f
C417 single_9b_cdac_0.cdac_sw_9b_0.S[0] a_62748_26999# 0.59531f
C418 sar9b_0.net19 a_5046_27230# 0.02764f
C419 sar9b_0.net56 sar9b_0.net49 0.45655f
C420 VDPWR a_12870_22267# 0.25924f
C421 a_6250_28502# a_5460_28377# 0.1263f
C422 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.03729f
C423 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[5] 1.06635f
C424 sar9b_0.net13 a_11430_24931# 0.03609f
C425 sar9b_0.net14 a_13164_28398# 0.14522f
C426 a_3027_22138# sar9b_0._05_ 0.07932f
C427 a_8057_18463# sar9b_0.net1 0.15171f
C428 VDPWR a_5151_28559# 0.26391f
C429 a_9323_27662# sar9b_0.net34 0.21484f
C430 single_9b_cdac_1.CF[4] sar9b_0.net29 0.03153f
C431 sar9b_0.net30 sar9b_0.net33 0.02513f
C432 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.12898f
C433 a_4467_24162# sar9b_0.net72 0.02699f
C434 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 1.71649f
C435 a_12870_19603# sar9b_0.net50 0.17286f
C436 sar9b_0.net54 a_6030_24396# 0.22581f
C437 sar9b_0.net61 single_9b_cdac_1.SW[1] 0.13622f
C438 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[2] 0.21948f
C439 sar9b_0.net31 a_12047_22521# 0.04699f
C440 sar9b_0.net36 sar9b_0.net48 0.17317f
C441 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26955f
C442 sar9b_0.net18 a_3946_27530# 0.02978f
C443 VDPWR a_12182_23755# 0.19519f
C444 sar9b_0.net42 a_11382_22142# 0.01996f
C445 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.03484f
C446 VDPWR a_3273_20185# 0.14496f
C447 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[0\] 0.01636f
C448 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.42784f
C449 sar9b_0.net11 sar9b_0.net39 0.01153f
C450 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 a_39616_17740# 0.14695f
C451 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_53154_16877# 0.04592f
C452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42784f
C453 a_10926_17021# sar9b_0.net27 0.03167f
C454 a_4211_19474# a_4072_19474# 0.02538f
C455 sar9b_0.net59 sar9b_0.net34 0.14932f
C456 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A a_25915_15495# 0.01076f
C457 a_10859_26330# sar9b_0.net33 0.22653f
C458 a_11382_23474# sar9b_0.net11 0.04486f
C459 a_8622_26345# a_9130_26198# 0.19065f
C460 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.31809f
C461 a_8303_23853# sar9b_0.net11 0.02489f
C462 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.04988f
C463 a_3219_22860# sar9b_0.clknet_1_1__leaf_CLK 0.01128f
C464 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.19266f
C465 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.3196f
C466 sar9b_0.net52 a_12182_26419# 0.14359f
C467 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C468 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] 1.14951f
C469 VDPWR a_11382_18146# 0.30035f
C470 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C471 sar9b_0.net46 a_4072_19474# 0.32046f
C472 VDPWR dw_12589_1395# 1.90366f
C473 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.01492f
C474 a_7638_23474# a_8098_23762# 0.26257f
C475 a_6954_27466# sar9b_0.net36 0.07226f
C476 sar9b_0.net60 clk 0.04516f
C477 VDPWR a_53154_16877# 1.81495f
C478 sar9b_0.net72 sar9b_0.clk_div_0.COUNT\[1\] 0.04678f
C479 sar9b_0.net71 sar9b_0.net46 0.29319f
C480 a_54737_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.01076f
C481 VDPWR single_9b_cdac_1.CF[8] 2.63907f
C482 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[8] 0.03384f
C483 sar9b_0.net59 sar9b_0.net58 0.82667f
C484 a_4947_20140# a_6130_20239# 0.0649f
C485 a_5126_20140# a_5931_20140# 0.29221f
C486 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[0] 0.02907f
C487 VDPWR a_11859_20574# 0.41872f
C488 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.10429f
C489 sar9b_0.net7 single_9b_cdac_1.SW[1] 0.70147f
C490 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C491 sar9b_0.net9 sar9b_0.net62 0.02856f
C492 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.02513f
C493 sar9b_0.net32 sar9b_0.net38 0.02088f
C494 VDPWR a_12588_16784# 0.22693f
C495 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C496 a_10553_18922# a_10762_18823# 0.24088f
C497 sar9b_0.net32 VDPWR 1.40875f
C498 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[7] 0.01285f
C499 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.05472f
C500 tdc_0.OUTN tdc_0.phase_detector_0.pd_out_0.A 0.11925f
C501 a_13011_25902# a_13011_24802# 0.0246f
C502 sar9b_0.net33 a_12047_26517# 0.04976f
C503 single_9b_cdac_1.CF[2] single_9b_cdac_0.SW[0] 0.35203f
C504 sar9b_0.net61 sar9b_0.net62 0.26134f
C505 sar9b_0.net57 clk 0.05645f
C506 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.1236f
C507 sar9b_0.net27 a_13216_26469# 0.01058f
C508 a_3370_26437# sar9b_0.net59 0.14542f
C509 a_6132_23451# a_6414_23681# 0.05462f
C510 a_5823_23477# a_6137_23791# 0.07826f
C511 a_8595_17910# single_9b_cdac_1.SW[0] 0.35058f
C512 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.08121f
C513 VDPWR a_5581_19664# 0.23366f
C514 sar9b_0.net43 a_8940_24402# 0.06556f
C515 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 2.81139f
C516 VDPWR a_8345_26455# 0.25217f
C517 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.0187f
C518 single_9b_cdac_1.cdac_sw_9b_0.S[8] th_dif_sw_0.VCP 0.85562f
C519 a_8595_17910# sar9b_0.net56 0.09371f
C520 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[3] 0.05403f
C521 sar9b_0.net38 sar9b_0.net51 0.1037f
C522 sar9b_0.net43 sar9b_0.net74 0.18429f
C523 a_5235_27466# uo_out[7] 0.39295f
C524 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.24399f
C525 a_16185_13034# tdc_0.RDY 0.06167f
C526 a_8057_18463# sar9b_0.net48 0.01239f
C527 VDPWR a_7402_22441# 0.20328f
C528 VDPWR sar9b_0.net51 1.04918f
C529 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C530 a_4755_22138# a_5938_22378# 0.0649f
C531 a_4934_22432# a_5289_22527# 0.18757f
C532 a_3161_26455# a_3438_26345# 0.09983f
C533 a_10402_27758# sar9b_0.net45 0.09798f
C534 sar9b_0.net26 a_12618_23470# 0.02755f
C535 a_41357_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C536 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[7] 0.31534f
C537 sar9b_0.net16 sar9b_0._10_ 0.06203f
C538 a_3922_20239# sar9b_0.clknet_1_0__leaf_CLK 0.09413f
C539 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.01664f
C540 a_8303_23853# a_8098_23762# 0.09983f
C541 a_9270_24566# a_9935_24187# 0.19065f
C542 a_8691_28566# a_9323_28371# 0.0245f
C543 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[4] 0.06951f
C544 sar9b_0.net1 sar9b_0.net51 0.16069f
C545 a_10995_28566# VDPWR 0.45062f
C546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.42509f
C547 a_3369_24181# a_3262_24141# 0.14439f
C548 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.06503f
C549 single_9b_cdac_1.CF[7] sar9b_0.net11 0.03981f
C550 a_7306_19777# sar9b_0.net40 0.02675f
C551 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.3545f
C552 single_9b_cdac_1.CF[1] th_dif_sw_0.VCN 0.09453f
C553 sar9b_0.net12 a_9165_24988# 0.01031f
C554 VDPWR a_13067_27662# 0.51166f
C555 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[5] 0.02149f
C556 a_2508_23444# sar9b_0.net69 0.06549f
C557 a_13011_23238# a_13216_22473# 0.01043f
C558 a_8019_17910# sar9b_0.net5 0.03181f
C559 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.01152f
C560 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.28523f
C561 a_7602_18116# a_7743_18149# 0.27388f
C562 a_8052_18123# a_8334_18353# 0.05462f
C563 sar9b_0.net43 a_10506_24506# 0.07702f
C564 a_3156_26115# a_2847_26141# 0.07766f
C565 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[7] 1.64863f
C566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.01003f
C567 a_8842_16874# sar9b_0.net5 0.04569f
C568 a_5394_18116# a_5849_18463# 0.3578f
C569 VDPWR a_5812_21028# 0.2311f
C570 a_7743_16817# a_8057_17131# 0.07826f
C571 sar9b_0.net40 clk 0.03834f
C572 sar9b_0._14_ sar9b_0.net68 0.7985f
C573 a_6954_27466# a_7478_27751# 0.05022f
C574 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.38397f
C575 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.69086f
C576 tdc_0.OUTN a_7404_16784# 0.05215f
C577 a_3545_26914# a_3754_26815# 0.24088f
C578 single_9b_cdac_1.CF[8] sar9b_0.net29 0.30185f
C579 sar9b_0.net49 sar9b_0.net57 0.18506f
C580 VDPWR a_10816_21487# 0.20703f
C581 a_8842_18206# sar9b_0.net5 0.21948f
C582 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.38397f
C583 VDPWR a_10649_17131# 0.21441f
C584 single_9b_cdac_1.CF[7] th_dif_sw_0.VCN 0.09453f
C585 sar9b_0.clknet_1_0__leaf_CLK a_3273_20185# 0.06919f
C586 a_11178_20806# a_11776_21141# 0.06623f
C587 th_dif_sw_0.CK tdc_0.OUTN 0.07179f
C588 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.75853f
C589 a_11842_22430# a_12182_22423# 0.24088f
C590 a_11658_22138# a_12618_22138# 0.03432f
C591 sar9b_0.net32 sar9b_0.net24 0.2487f
C592 a_2892_27039# a_3231_27227# 0.07649f
C593 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 1.55978f
C594 sar9b_0.net53 sar9b_0.net11 0.33023f
C595 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 2.82223f
C596 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] 3.10226f
C597 a_3521_24240# sar9b_0.clk_div_0.COUNT\[1\] 0.01149f
C598 sar9b_0.net31 a_11658_23470# 0.02378f
C599 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C600 a_10895_22855# sar9b_0.net11 0.04486f
C601 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C602 a_9258_21842# a_10218_21842# 0.03471f
C603 a_9442_21474# a_9782_21622# 0.24088f
C604 a_12531_28566# uo_out[0] 0.12656f
C605 sar9b_0.net32 sar9b_0.net29 0.02003f
C606 a_8340_26115# a_8940_27039# 0.0165f
C607 a_11915_28371# uo_out[0] 0.38176f
C608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.7611f
C609 a_6861_22828# clk 0.01643f
C610 a_2508_27440# a_2706_27440# 0.06623f
C611 a_3014_24136# a_3262_24141# 0.05308f
C612 sar9b_0.net12 sar9b_0.net38 0.02887f
C613 VDPWR sar9b_0.clk_div_0.COUNT\[0\] 0.52537f
C614 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.01003f
C615 a_8512_27801# sar9b_0.net22 0.27285f
C616 a_7289_21127# a_6975_20813# 0.07826f
C617 VDPWR sar9b_0.net12 1.09949f
C618 VDPWR a_5196_24776# 0.23838f
C619 a_6738_22112# a_7402_22441# 0.16939f
C620 sar9b_0.net56 a_10218_20806# 0.21365f
C621 sar9b_0.net13 sar9b_0.cyclic_flag_0.FINAL 0.03185f
C622 single_9b_cdac_1.cdac_sw_9b_0.S[0] th_dif_sw_0.VCP 0.21807p
C623 a_6636_20780# sar9b_0.net40 0.02169f
C624 sar9b_0.net1 sar9b_0.net12 0.03139f
C625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[6] 0.02149f
C626 VDPWR a_10762_18823# 0.20297f
C627 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01156f
C628 a_10607_25185# a_10402_25094# 0.09983f
C629 sar9b_0.net24 a_10995_28566# 0.21865f
C630 a_12560_27128# a_11915_27039# 0.02698f
C631 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[5] 0.01887f
C632 sar9b_0.net40 a_11658_19474# 0.07402f
C633 sar9b_0.net73 sar9b_0.net37 0.02388f
C634 a_8031_26141# sar9b_0.net59 0.20849f
C635 sar9b_0.net52 a_8438_23755# 0.13752f
C636 clk a_16331_9671# 0.37638f
C637 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[8] 0.36652f
C638 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C639 sar9b_0.net49 sar9b_0.net40 0.16393f
C640 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[0] 0.56248f
C641 VDPWR a_43540_26999# 1.81495f
C642 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.11216f
C643 a_7289_21127# a_7498_21109# 0.24088f
C644 sar9b_0.net29 a_13067_27662# 0.10621f
C645 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.01751f
C646 sar9b_0.net41 sar9b_0.net56 0.06968f
C647 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.69086f
C648 sar9b_0.net26 sar9b_0.net39 0.06931f
C649 a_5739_22488# sar9b_0.net39 0.01448f
C650 a_10553_18922# sar9b_0.net42 0.018f
C651 a_5812_21028# sar9b_0._17_ 0.04354f
C652 VDPWR a_3219_22860# 0.26196f
C653 a_6579_18832# a_5844_18123# 0.01182f
C654 VDPWR a_5289_22527# 0.14221f
C655 sar9b_0.net35 sar9b_0.net10 1.66696f
C656 sar9b_0.net16 a_3795_19512# 0.0476f
C657 a_10506_23174# a_10230_23234# 0.1263f
C658 sar9b_0.net43 a_5962_24151# 0.02064f
C659 a_7743_18149# a_7404_18116# 0.07649f
C660 a_5506_26802# a_5846_26950# 0.24088f
C661 sar9b_0.net30 a_11842_23762# 0.02126f
C662 a_5298_24499# a_5962_24151# 0.16939f
C663 sar9b_0.clknet_0_CLK a_4236_21738# 0.03044f
C664 a_10218_27466# sar9b_0.net38 0.01643f
C665 sar9b_0.net33 sar9b_0.net27 0.03715f
C666 sar9b_0.net2 sar9b_0.net10 0.02528f
C667 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.01879f
C668 a_10218_27466# VDPWR 0.8229f
C669 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[3] 0.01573f
C670 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C671 sar9b_0.net43 sar9b_0.net39 0.08882f
C672 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C673 sar9b_0.net6 sar9b_0.net37 0.05412f
C674 a_8726_22954# sar9b_0.net11 0.06796f
C675 sar9b_0._08_ a_5812_21028# 0.05999f
C676 a_24332_16877# single_9b_cdac_1.SW[8] 0.28324f
C677 a_7926_23234# sar9b_0.net54 0.22246f
C678 a_5298_24499# sar9b_0.net39 0.01755f
C679 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C680 VDPWR dw_17224_1400# 1.89831f
C681 a_3713_22522# sar9b_0._12_ 0.04441f
C682 sar9b_0.net68 sar9b_0._16_ 0.0172f
C683 a_4136_25584# a_4293_25852# 0.21226f
C684 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.26427f
C685 sar9b_0.net43 a_5439_24563# 0.02732f
C686 sar9b_0.net30 single_9b_cdac_0.SW[4] 0.11168f
C687 single_9b_cdac_1.CF[0] ua[0] 3.29077f
C688 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.19266f
C689 a_18214_3039# th_dif_sw_0.th_sw_1.CKB 0.42927f
C690 a_5298_24499# a_5439_24563# 0.27388f
C691 VDPWR a_7638_19238# 0.30428f
C692 sar9b_0.net60 sar9b_0.net45 1.09005f
C693 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.05472f
C694 a_7338_24802# a_6562_25094# 0.3578f
C695 sar9b_0.net32 single_9b_cdac_0.SW[3] 0.04904f
C696 a_6767_25185# a_6378_24802# 0.06034f
C697 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.47485f
C698 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36446f
C699 sar9b_0.net8 a_11776_21141# 0.3091f
C700 th_dif_sw_0.VCN th_dif_sw_0.VCP 0.69759f
C701 VDPWR a_6642_19448# 0.3497f
C702 a_6744_23238# sar9b_0.clk_div_0.COUNT\[2\] 0.03621f
C703 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.75899f
C704 single_9b_cdac_0.SW[2] th_dif_sw_0.VCN 0.09453f
C705 a_10649_17131# sar9b_0.net48 0.06775f
C706 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 0.19143f
C707 sar9b_0._11_ sar9b_0._10_ 0.03596f
C708 VDPWR a_7566_21017# 0.26799f
C709 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16331_9671# 0.18915f
C710 a_4210_22378# sar9b_0.clknet_1_1__leaf_CLK 0.09811f
C711 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C712 sar9b_0.clknet_0_CLK sar9b_0.clknet_1_1__leaf_CLK 0.04779f
C713 a_21368_4076# ua[3] 0.65763f
C714 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[1\] 1.08101f
C715 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22655f
C716 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] 0.17948f
C717 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.12431f
C718 uio_in[0] ui_in[7] 0.03102f
C719 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[1] 0.21792f
C720 single_9b_cdac_1.CF[1] sar9b_0.net26 0.05711f
C721 sar9b_0.net46 sar9b_0.net37 0.07123f
C722 a_10182_20463# a_10528_20155# 0.07649f
C723 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.02513f
C724 a_4125_25958# sar9b_0.net39 0.02409f
C725 a_5126_20140# a_5633_20244# 0.21226f
C726 a_7284_20787# sar9b_0.net61 0.01281f
C727 a_4947_20140# a_5481_20185# 0.35097f
C728 a_11382_22142# sar9b_0.net39 0.03507f
C729 VDPWR a_13216_18477# 0.21525f
C730 th_dif_sw_0.CK sar9b_0.net39 0.03714f
C731 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.SW[8] 0.22497f
C732 sar9b_0.net55 a_6414_23681# 0.0176f
C733 a_8970_20510# a_9494_20290# 0.04522f
C734 a_8694_20570# a_9359_20191# 0.19065f
C735 sar9b_0.net23 sar9b_0.cyclic_flag_0.FINAL 0.03316f
C736 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.19266f
C737 clk a_16527_10454# 0.20249f
C738 sar9b_0._09_ sar9b_0.net60 0.06706f
C739 single_9b_cdac_0.SW[4] ua[0] 0.17308f
C740 sar9b_0.net8 sar9b_0.net27 0.0426f
C741 a_10858_17113# tdc_0.OUTP 0.06033f
C742 a_4812_28371# sar9b_0.net60 0.02169f
C743 a_11430_24931# a_11776_25137# 0.07649f
C744 a_3371_23106# sar9b_0._07_ 0.18693f
C745 single_9b_cdac_1.CF[1] a_13011_20806# 0.06696f
C746 VDPWR a_9359_20191# 0.26316f
C747 a_13067_27662# single_9b_cdac_0.SW[3] 0.02544f
C748 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.26942f
C749 sar9b_0.net18 sar9b_0.net60 0.03658f
C750 a_10762_18823# sar9b_0.net48 0.14f
C751 tdc_0.phase_detector_0.pd_out_0.B a_15052_11404# 0.18949f
C752 a_9270_24566# sar9b_0.net12 0.04846f
C753 sar9b_0.net4 sar9b_0.net39 0.0209f
C754 a_9154_20142# sar9b_0.net37 0.02634f
C755 a_6975_20813# sar9b_0.net47 0.17348f
C756 a_5441_22522# a_5289_22527# 0.22517f
C757 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.SW[7] 0.03585f
C758 sar9b_0._11_ sar9b_0.net4 0.03423f
C759 sar9b_0._15_ sar9b_0.net39 0.09291f
C760 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C761 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C762 sar9b_0.net26 single_9b_cdac_1.CF[7] 0.18995f
C763 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.3545f
C764 single_9b_cdac_0.SW[7] single_9b_cdac_1.CF[7] 1.81115f
C765 a_10218_27466# sar9b_0.net24 0.03703f
C766 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C767 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.06503f
C768 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[8] 0.01791f
C769 a_5439_24563# sar9b_0._15_ 0.06796f
C770 a_9930_20510# sar9b_0.net51 0.07643f
C771 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A 0.74663f
C772 sar9b_0.net1 a_9359_20191# 0.01823f
C773 sar9b_0.net28 single_9b_cdac_0.SW[0] 0.1354f
C774 sar9b_0._09_ sar9b_0.net57 0.46567f
C775 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] 0.17948f
C776 sar9b_0._11_ sar9b_0._01_ 0.04965f
C777 sar9b_0.net52 a_12491_27662# 0.01099f
C778 a_10742_27751# a_11178_27466# 0.16939f
C779 a_6137_23791# sar9b_0.net54 0.06976f
C780 a_7890_26108# a_8031_26141# 0.27388f
C781 VDPWR a_2508_20780# 1.55529f
C782 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.19266f
C783 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.42509f
C784 a_7602_18116# sar9b_0.net73 0.08061f
C785 VDPWR w_12795_1601# 0.45037f
C786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.12431f
C787 VDPWR sar9b_0.net42 1.57366f
C788 sar9b_0.net40 sar9b_0.net45 0.05943f
C789 a_9942_27470# sar9b_0.net59 0.22307f
C790 single_9b_cdac_1.SW[3] a_49221_17740# 0.18991f
C791 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[4] 4.15222f
C792 sar9b_0.net10 a_7978_22202# 0.08861f
C793 VDPWR a_8386_22806# 0.24182f
C794 a_7498_21109# sar9b_0.net47 0.15768f
C795 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.SW[6] 0.03532f
C796 sar9b_0.net26 sar9b_0.net53 0.06847f
C797 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C798 a_7193_22459# a_7470_22349# 0.09983f
C799 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C800 sar9b_0._01_ a_5374_20145# 0.13551f
C801 a_9130_26198# sar9b_0.cyclic_flag_0.FINAL 0.05175f
C802 uio_in[4] uio_in[3] 0.03102f
C803 sar9b_0.net49 a_9647_21523# 0.22799f
C804 a_10166_3438# a_10254_2858# 0.99857f
C805 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[6] 0.09845f
C806 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[5] 0.0149f
C807 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.15428f
C808 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.62443f
C809 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C810 sar9b_0._18_ sar9b_0.clk_div_0.COUNT\[2\] 0.71169f
C811 a_7638_19238# sar9b_0.net48 0.22589f
C812 a_9323_28371# uo_out[3] 0.04123f
C813 a_16527_10454# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.09051f
C814 single_9b_cdac_0.cdac_sw_9b_0.S[7] VDPWR 4.1608f
C815 sar9b_0.net41 sar9b_0.net57 0.02983f
C816 VDPWR a_11859_17910# 0.40675f
C817 sar9b_0._07_ sar9b_0.net46 0.15475f
C818 single_9b_cdac_1.CF[3] single_9b_cdac_0.SW[0] 0.40374f
C819 a_8098_18810# a_9126_19131# 0.07826f
C820 sar9b_0.net43 sar9b_0.net53 0.57297f
C821 VDPWR a_4771_18260# 0.42657f
C822 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.42014f
C823 sar9b_0.net43 a_10895_22855# 0.02011f
C824 a_9450_17846# a_9634_17478# 0.43869f
C825 single_9b_cdac_1.SW[2] a_9634_17478# 0.01591f
C826 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C827 sar9b_0.net67 sar9b_0.clknet_0_CLK 0.0173f
C828 sar9b_0.net38 a_10482_25831# 0.01616f
C829 a_10926_17021# a_10649_17131# 0.09983f
C830 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[1] 4.15038f
C831 sar9b_0.net56 a_8874_19178# 0.01259f
C832 a_7743_16817# sar9b_0.net6 0.02026f
C833 VDPWR a_10482_25831# 0.34041f
C834 a_7097_19795# a_7882_19538# 0.26257f
C835 sar9b_0.net45 a_9588_27045# 0.25117f
C836 a_5506_17478# sar9b_0.net56 0.03523f
C837 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.01003f
C838 VDPWR a_21177_7457# 1.54446f
C839 sar9b_0.net20 a_5742_28392# 0.07038f
C840 a_5748_24381# a_5962_24151# 0.05022f
C841 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.19325f
C842 a_10070_24286# a_10506_24506# 0.16939f
C843 sar9b_0._18_ a_3695_23038# 0.02716f
C844 sar9b_0.net8 sar9b_0.net36 0.02461f
C845 a_10644_16791# sar9b_0.net61 0.02207f
C846 single_9b_cdac_0.SW[6] clk 0.22166f
C847 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.6919f
C848 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.42509f
C849 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C850 a_10859_26330# a_11382_26138# 0.04056f
C851 a_5439_24563# a_5748_24381# 0.07766f
C852 a_30012_17740# single_9b_cdac_1.SW[7] 0.18991f
C853 th_dif_sw_0.VCN single_9b_cdac_1.SW[2] 0.09468f
C854 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP a_38738_16877# 0.04592f
C855 sar9b_0.net27 single_9b_cdac_1.CF[0] 0.02972f
C856 a_5046_27230# sar9b_0.net37 0.04431f
C857 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.0313f
C858 a_8057_17131# sar9b_0.net27 0.01567f
C859 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.71729f
C860 sar9b_0.net41 sar9b_0.net40 0.06786f
C861 sar9b_0.net53 a_11382_22142# 0.2367f
C862 uo_out[0] uo_out[1] 3.57901f
C863 uo_out[3] ui_in[0] 0.06786f
C864 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[2] 0.01791f
C865 a_7602_18116# sar9b_0.net46 0.27602f
C866 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.6205f
C867 a_9588_27045# a_9870_27060# 0.06034f
C868 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C869 a_7743_16817# sar9b_0.net46 0.17057f
C870 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[2] 0.02195f
C871 sar9b_0.net73 a_7404_18116# 0.09233f
C872 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C873 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C874 sar9b_0.net58 a_3540_27045# 0.17959f
C875 sar9b_0.net39 sar9b_0.clknet_1_1__leaf_CLK 0.01422f
C876 VDPWR a_6414_23681# 0.26663f
C877 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.26707f
C878 VDPWR a_4210_22378# 0.37875f
C879 sar9b_0.net27 a_13011_20574# 0.04061f
C880 a_8052_18123# sar9b_0.net5 0.06414f
C881 VDPWR sar9b_0.clknet_0_CLK 2.46803f
C882 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0._12_ 0.30315f
C883 sar9b_0.net38 uo_out[5] 0.25815f
C884 VDPWR a_3946_26198# 0.30347f
C885 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.84424f
C886 a_2835_24136# sar9b_0.net69 0.01995f
C887 a_10378_27170# sar9b_0.net59 0.22839f
C888 a_10218_24802# a_9942_24806# 0.1263f
C889 sar9b_0.net42 sar9b_0.net48 0.07688f
C890 VDPWR uo_out[5] 0.89589f
C891 sar9b_0.net27 a_11842_23762# 0.01034f
C892 VDPWR sar9b_0.net16 1.35456f
C893 VDPWR a_12064_22819# 0.1986f
C894 sar9b_0.net23 a_9130_26198# 0.03663f
C895 a_14871_9671# th_dif_sw_0.VCN 0.11478f
C896 a_16331_9671# a_16357_9613# 0.12812f
C897 sar9b_0.net61 a_9634_17478# 0.16934f
C898 a_11382_26138# a_12047_26517# 0.19065f
C899 a_4332_23043# sar9b_0.clk_div_0.COUNT\[2\] 0.1269f
C900 VDPWR a_8940_24402# 0.29362f
C901 sar9b_0.net74 sar9b_0.net38 0.03312f
C902 sar9b_0.net36 sar9b_0.net34 0.04627f
C903 a_10194_16784# a_10335_16817# 0.27388f
C904 single_9b_cdac_1.SW[8] th_dif_sw_0.VCN 0.09453f
C905 a_2508_20780# sar9b_0.clknet_1_0__leaf_CLK 1.89917f
C906 sar9b_0.net55 sar9b_0.net39 0.04945f
C907 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C908 VDPWR sar9b_0.net74 1.07986f
C909 a_6922_23534# sar9b_0.net11 0.05827f
C910 sar9b_0.net56 a_5322_17846# 0.23955f
C911 single_9b_cdac_0.SW[1] VDPWR 2.63243f
C912 VDPWR a_7914_27466# 0.35464f
C913 sar9b_0._04_ a_3027_21906# 0.24347f
C914 sar9b_0.net63 sar9b_0._02_ 0.07961f
C915 a_7188_22119# sar9b_0.net10 0.01911f
C916 sar9b_0.net18 uio_out[1] 0.0124f
C917 VDPWR a_2893_24992# 0.23635f
C918 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.76578f
C919 VDPWR tdc_0.OUTN 0.62093f
C920 sar9b_0.net6 a_7404_18116# 0.28739f
C921 single_9b_cdac_0.SW[4] sar9b_0.net27 0.05602f
C922 VDPWR single_9b_cdac_1.CF[6] 2.73682f
C923 sar9b_0.net65 a_4236_21738# 0.08898f
C924 a_6250_28502# a_5742_28392# 0.19065f
C925 VDPWR a_13216_22473# 0.20771f
C926 sar9b_0.net13 a_11776_25137# 0.29958f
C927 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[4] 10.4962f
C928 sar9b_0._04_ sar9b_0._05_ 0.2432f
C929 sar9b_0.net4 a_6562_25094# 0.01993f
C930 VDPWR a_5465_28246# 0.21298f
C931 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.27713f
C932 sar9b_0.net60 uo_out[7] 0.02565f
C933 a_21368_4076# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.16499f
C934 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.6919f
C935 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[6] 4.16106f
C936 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.81428f
C937 clk tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.09743f
C938 sar9b_0.net58 sar9b_0.net36 0.27889f
C939 sar9b_0.net1 tdc_0.OUTN 0.04134f
C940 a_4934_22432# sar9b_0.net39 0.0126f
C941 a_9162_23174# clk 0.02449f
C942 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 2.71729f
C943 VDPWR a_12618_23470# 0.32668f
C944 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C945 th_dif_sw_0.CK th_dif_sw_0.VCP 0.0144f
C946 a_5289_22527# sar9b_0._12_ 0.0393f
C947 VDPWR a_3723_20140# 0.08905f
C948 sar9b_0.net38 a_10506_24506# 0.02782f
C949 VDPWR a_62748_16877# 1.81495f
C950 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C951 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.A 0.02054f
C952 VDPWR a_10506_24506# 0.34709f
C953 sar9b_0.net32 sar9b_0.net33 0.02518f
C954 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[2] 54.8348f
C955 a_6052_19792# a_5581_19664# 0.01114f
C956 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.7611f
C957 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.08121f
C958 sar9b_0.net60 a_5484_23444# 0.01027f
C959 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[3] 0.08999f
C960 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_53154_26999# 0.04592f
C961 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02632f
C962 sar9b_0.net60 a_5126_20140# 0.02835f
C963 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C964 a_4922_20857# sar9b_0._18_ 0.14576f
C965 VDPWR a_8940_27039# 0.24411f
C966 a_16222_11316# tdc_0.phase_detector_0.INN 0.02415f
C967 sar9b_0.net72 sar9b_0.clk_div_0.COUNT\[2\] 0.29657f
C968 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[1] 0.21746f
C969 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.45521f
C970 sar9b_0.net65 sar9b_0.clknet_1_1__leaf_CLK 0.19718f
C971 sar9b_0.net52 a_12618_26134# 0.26209f
C972 a_5581_20992# sar9b_0._01_ 0.01832f
C973 a_10182_20463# a_9154_20142# 0.07826f
C974 a_7914_23470# a_8438_23755# 0.05022f
C975 a_7138_27758# sar9b_0.net36 0.13653f
C976 a_5235_27466# sar9b_0.net19 0.19875f
C977 sar9b_0.net59 a_5046_27230# 0.01797f
C978 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07579f
C979 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[8] 0.2453f
C980 a_13011_19242# sar9b_0.net40 0.03f
C981 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[0] 0.03109f
C982 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.75853f
C983 sar9b_0.net57 a_5484_23444# 0.04904f
C984 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C985 sar9b_0.net57 a_5126_20140# 0.01075f
C986 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.17533f
C987 a_10194_16784# sar9b_0.net6 0.07207f
C988 a_3369_24181# sar9b_0.clknet_1_1__leaf_CLK 0.06961f
C989 sar9b_0.net18 a_3156_27447# 0.02909f
C990 single_9b_cdac_1.SW[3] ua[0] 0.14032f
C991 a_10548_19053# a_11338_19178# 0.1263f
C992 a_2547_28132# sar9b_0.net17 0.0815f
C993 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.12431f
C994 sar9b_0.net70 a_3027_21906# 0.15443f
C995 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.94957f
C996 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[7] 0.02149f
C997 sar9b_0._08_ sar9b_0.net16 0.13446f
C998 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.CF[5] 0.03484f
C999 sar9b_0.net41 a_13011_17910# 0.2244f
C1000 single_9b_cdac_0.SW[1] sar9b_0.net29 0.30909f
C1001 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.01003f
C1002 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 ua[0] 0.12076f
C1003 sar9b_0.net70 sar9b_0._05_ 0.12818f
C1004 sar9b_0.net60 a_6102_24806# 0.02205f
C1005 a_6282_17846# a_6534_17799# 0.27388f
C1006 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.10429f
C1007 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 3.04383f
C1008 sar9b_0.net8 a_11859_20574# 0.0265f
C1009 single_9b_cdac_1.CF[6] sar9b_0.net29 0.19274f
C1010 sar9b_0.net29 a_13216_22473# 0.01568f
C1011 VDPWR a_7638_23474# 0.28218f
C1012 sar9b_0.net2 a_10803_19474# 0.02668f
C1013 single_9b_cdac_0.SW[0] a_63626_26990# 0.18991f
C1014 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 ua[0] 0.12069f
C1015 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.42509f
C1016 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C1017 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.SW[6] 0.17155f
C1018 sar9b_0.clknet_1_0__leaf_CLK sar9b_0.clknet_0_CLK 0.03854f
C1019 VDPWR a_3372_25734# 0.23391f
C1020 a_8303_18859# a_7914_19178# 0.05462f
C1021 a_3161_26455# a_3946_26198# 0.26257f
C1022 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.24443f
C1023 a_3370_26437# a_3438_26345# 0.35559f
C1024 sar9b_0._13_ sar9b_0._14_ 0.15271f
C1025 sar9b_0.net41 a_9647_21523# 0.0288f
C1026 a_34814_17740# single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.22352f
C1027 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0313f
C1028 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[7] 0.06503f
C1029 sar9b_0.net16 sar9b_0.clknet_1_0__leaf_CLK 0.0448f
C1030 a_6130_20239# sar9b_0.net4 0.03123f
C1031 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36322f
C1032 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 1.71649f
C1033 a_3855_25792# a_4136_25584# 0.29207f
C1034 a_9472_23805# a_8874_23470# 0.06623f
C1035 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[4] 1.90123f
C1036 a_10335_16817# sar9b_0.net27 0.02939f
C1037 sar9b_0.net58 a_5151_28559# 0.19397f
C1038 a_9730_24138# a_9935_24187# 0.09983f
C1039 VDPWR a_13164_28398# 0.25851f
C1040 VDPWR a_7343_27849# 0.26147f
C1041 a_13011_16810# single_9b_cdac_1.SW[4] 0.01587f
C1042 sar9b_0.net44 a_3161_27787# 0.02151f
C1043 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1044 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.05472f
C1045 a_8266_17113# a_8052_16791# 0.04522f
C1046 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.81428f
C1047 a_8940_24402# a_9270_24566# 0.04271f
C1048 sar9b_0.net2 a_9546_24506# 0.05795f
C1049 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1050 VDPWR a_5962_24151# 0.19439f
C1051 sar9b_0.net38 sar9b_0.net21 0.04603f
C1052 a_3014_24136# sar9b_0.clknet_1_1__leaf_CLK 0.09139f
C1053 sar9b_0.net8 sar9b_0.net51 0.28615f
C1054 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.SW[7] 0.14951f
C1055 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.0303f
C1056 VDPWR sar9b_0.net21 0.42201f
C1057 sar9b_0.net24 a_8940_27039# 0.28492f
C1058 sar9b_0.net36 a_10528_20155# 0.0105f
C1059 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.19266f
C1060 sar9b_0.net33 sar9b_0.net12 0.05295f
C1061 sar9b_0.net38 sar9b_0.net39 0.02578f
C1062 a_7743_18149# a_8057_18463# 0.07826f
C1063 a_8052_18123# a_8842_18206# 0.1263f
C1064 sar9b_0.net43 a_11104_24151# 0.02813f
C1065 VDPWR sar9b_0.net39 1.30812f
C1066 a_6834_20780# a_6975_20813# 0.27388f
C1067 single_9b_cdac_0.cdac_sw_9b_0.S[3] ua[0] 1.59042f
C1068 a_5394_18116# a_6058_18445# 0.16939f
C1069 a_5844_18123# a_6126_18353# 0.05462f
C1070 a_21368_4076# a_18214_3039# 0.99857f
C1071 VDPWR sar9b_0._11_ 0.2748f
C1072 a_7138_27758# a_7478_27751# 0.24088f
C1073 a_6954_27466# a_7914_27466# 0.03432f
C1074 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.22875f
C1075 single_9b_cdac_1.SW[0] a_9839_17527# 0.03009f
C1076 VDPWR a_5439_24563# 0.25892f
C1077 single_9b_cdac_1.CF[2] ua[0] 3.58697f
C1078 VDPWR a_2603_17006# 0.51948f
C1079 tdc_0.OUTN a_7602_16784# 0.07198f
C1080 VDPWR a_11382_23474# 0.29464f
C1081 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.62443f
C1082 sar9b_0.net26 single_9b_cdac_1.SW[8] 0.03854f
C1083 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS ua[3] 0.93526f
C1084 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.59531f
C1085 sar9b_0.net1 sar9b_0.net39 0.02611f
C1086 sar9b_0._14_ sar9b_0.net69 0.03025f
C1087 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 3.10626f
C1088 VDPWR a_8982_21902# 0.33673f
C1089 a_3090_27163# a_3754_26815# 0.16939f
C1090 VDPWR a_8303_23853# 0.26302f
C1091 sar9b_0.net67 sar9b_0.net65 0.11461f
C1092 sar9b_0.net17 ui_in[0] 0.02606f
C1093 sar9b_0.clknet_1_0__leaf_CLK a_3723_20140# 0.07189f
C1094 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.3196f
C1095 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.71729f
C1096 a_9258_21842# sar9b_0.net37 0.02924f
C1097 a_11842_22430# a_12618_22138# 0.3578f
C1098 a_11658_22138# a_12047_22521# 0.06034f
C1099 VDPWR a_15400_11316# 0.52162f
C1100 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP a_57946_16877# 0.04592f
C1101 VDPWR a_5374_20145# 0.01375f
C1102 a_9546_24506# a_10758_24459# 0.07766f
C1103 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[7] 0.02552f
C1104 sar9b_0._06_ uo_out[0] 0.19708f
C1105 a_8982_21902# sar9b_0.net1 0.01917f
C1106 sar9b_0.net53 a_10070_24286# 0.1338f
C1107 a_3156_27447# a_2847_27473# 0.07766f
C1108 sar9b_0.net9 sar9b_0.net26 0.02943f
C1109 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[3] 0.02468f
C1110 sar9b_0.net47 a_6444_19448# 0.06747f
C1111 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C1112 sar9b_0.net40 a_6102_24806# 0.01823f
C1113 a_10548_19053# a_10803_18142# 0.04032f
C1114 single_9b_cdac_0.SW[5] a_39616_26990# 0.18991f
C1115 a_7498_21109# a_6834_20780# 0.16939f
C1116 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.83441f
C1117 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[3] 0.02012f
C1118 th_dif_sw_0.CK single_9b_cdac_1.SW[2] 0.04691f
C1119 sar9b_0.net26 sar9b_0.net61 0.01357f
C1120 sar9b_0.net47 a_7470_22349# 0.22357f
C1121 sar9b_0.net56 a_10402_21098# 0.01558f
C1122 a_12560_27128# single_9b_cdac_0.SW[4] 0.03746f
C1123 sar9b_0.net57 sar9b_0.net10 0.09558f
C1124 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[7] 14.2348f
C1125 sar9b_0.net43 sar9b_0.net9 0.0248f
C1126 sar9b_0.net25 a_12531_28566# 0.21118f
C1127 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C1128 sar9b_0.net27 sar9b_0.net6 1.39158f
C1129 a_11915_28371# sar9b_0.net25 0.11385f
C1130 a_11842_23762# a_12182_23755# 0.24088f
C1131 sar9b_0.net19 a_3545_26914# 0.17405f
C1132 sar9b_0.net49 a_10227_18142# 0.20483f
C1133 sar9b_0.net40 a_11842_19766# 0.1379f
C1134 sar9b_0.net54 a_6378_24802# 0.1648f
C1135 single_9b_cdac_1.CF[5] sar9b_0.net28 0.03576f
C1136 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C1137 clk a_16357_9613# 0.01204f
C1138 sar9b_0.net52 a_8874_23470# 0.26484f
C1139 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[0] 0.01464f
C1140 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 1.71649f
C1141 VDPWR single_9b_cdac_1.CF[1] 2.73909f
C1142 a_3425_20244# a_3273_20185# 0.22338f
C1143 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[6] 0.26707f
C1144 sar9b_0._06_ a_12491_27662# 0.04301f
C1145 th_dif_sw_0.CK a_12182_18427# 0.06686f
C1146 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.38397f
C1147 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C1148 a_8622_26345# a_8340_26115# 0.05462f
C1149 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.15052f
C1150 a_10335_16817# sar9b_0.net36 0.02026f
C1151 a_10402_25094# sar9b_0.net38 0.0296f
C1152 sar9b_0._17_ sar9b_0.net39 0.02501f
C1153 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24495f
C1154 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.36006f
C1155 a_6738_22112# sar9b_0.net39 0.05411f
C1156 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C1157 VDPWR sar9b_0.net65 0.94256f
C1158 a_9165_24988# sar9b_0.net53 0.20816f
C1159 sar9b_0._11_ sar9b_0._17_ 0.45057f
C1160 a_6922_23534# a_6132_23451# 0.1263f
C1161 VDPWR a_10402_25094# 0.21159f
C1162 VDPWR a_6540_22112# 0.20318f
C1163 a_7882_19538# sar9b_0.net61 0.01172f
C1164 sar9b_0.net63 a_4811_23656# 0.08526f
C1165 a_5441_22522# sar9b_0.net39 0.01163f
C1166 sar9b_0.net32 uo_out[3] 0.13894f
C1167 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VDPWR 2.81428f
C1168 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[2] 0.0313f
C1169 sar9b_0.net35 a_7193_22459# 0.01725f
C1170 sar9b_0.net41 clk 0.05496f
C1171 VDPWR single_9b_cdac_1.CF[7] 2.59279f
C1172 single_9b_cdac_0.SW[1] a_57946_26999# 0.28324f
C1173 sar9b_0.net7 sar9b_0.net26 0.07618f
C1174 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.26707f
C1175 single_9b_cdac_1.SW[5] a_38738_16877# 0.28324f
C1176 sar9b_0.net31 a_11178_24802# 0.01626f
C1177 sar9b_0._08_ sar9b_0._11_ 0.26992f
C1178 sar9b_0.net27 sar9b_0.net46 0.77693f
C1179 sar9b_0.net27 sar9b_0.net50 0.03263f
C1180 a_4210_22378# sar9b_0._12_ 0.04138f
C1181 VDPWR a_3369_24181# 0.15274f
C1182 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.11216f
C1183 sar9b_0.net48 sar9b_0.net39 0.0236f
C1184 sar9b_0.net52 sar9b_0.net37 0.74767f
C1185 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[3] 0.02744f
C1186 single_9b_cdac_1.SW[3] sar9b_0.net27 0.02529f
C1187 sar9b_0.net40 sar9b_0.net10 0.35246f
C1188 sar9b_0.clknet_0_CLK sar9b_0._12_ 0.02864f
C1189 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.42784f
C1190 a_7092_19455# sar9b_0.net62 0.03046f
C1191 sar9b_0.net27 a_12618_18142# 0.02447f
C1192 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[4] 0.0154f
C1193 sar9b_0.net15 a_6579_18832# 0.01202f
C1194 sar9b_0.net43 sar9b_0.net7 0.59584f
C1195 VDPWR a_8098_18810# 0.26718f
C1196 sar9b_0.net36 sar9b_0.net73 0.03096f
C1197 th_dif_sw_0.CK sar9b_0.net61 0.02316f
C1198 a_4365_25770# a_4698_25851# 0.14439f
C1199 sar9b_0._16_ sar9b_0.net69 0.04762f
C1200 VDPWR a_7097_19795# 0.22516f
C1201 sar9b_0.net49 a_10218_20806# 0.2026f
C1202 a_6954_27466# a_7343_27849# 0.06034f
C1203 sar9b_0.net53 sar9b_0.net38 0.33144f
C1204 a_12182_19759# single_9b_cdac_1.SW[8] 0.01333f
C1205 VDPWR a_8074_20870# 0.30584f
C1206 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[2\] 0.04613f
C1207 a_3521_24240# a_2835_24136# 0.27693f
C1208 a_13011_20574# sar9b_0.net51 0.0305f
C1209 sar9b_0._11_ sar9b_0.clknet_1_0__leaf_CLK 0.08207f
C1210 a_4755_22138# sar9b_0.net60 0.01468f
C1211 a_10166_3438# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.16499f
C1212 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] 3.10214f
C1213 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_16357_9613# 0.16728f
C1214 VDPWR sar9b_0.net53 3.3527f
C1215 VDPWR a_10895_22855# 0.26689f
C1216 sar9b_0.net32 single_9b_cdac_0.SW[4] 0.02994f
C1217 single_9b_cdac_0.SW[1] a_13216_26469# 0.02143f
C1218 a_6954_27466# sar9b_0.net21 0.03499f
C1219 a_18214_3039# ua[3] 0.12559f
C1220 single_9b_cdac_0.cdac_sw_9b_0.S[0] a_63626_26990# 0.22513f
C1221 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.12358f
C1222 sar9b_0.net1 sar9b_0.net53 0.19803f
C1223 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C1224 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.71729f
C1225 single_9b_cdac_1.SW[4] th_dif_sw_0.VCN 0.09453f
C1226 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.84423f
C1227 single_9b_cdac_1.CF[1] sar9b_0.net29 0.04096f
C1228 sar9b_0.net31 clk 0.0477f
C1229 a_4755_22138# sar9b_0.net57 0.01782f
C1230 VDPWR a_3014_24136# 0.9015f
C1231 sar9b_0.net42 sar9b_0.net33 0.01652f
C1232 sar9b_0.net41 sar9b_0.net49 0.52224f
C1233 sar9b_0.net36 sar9b_0.net6 0.05014f
C1234 clk tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.09625f
C1235 sar9b_0.net41 a_9162_23174# 0.01093f
C1236 sar9b_0.net65 sar9b_0._17_ 0.17308f
C1237 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.31534f
C1238 sar9b_0.net20 sar9b_0.net60 0.0552f
C1239 VDPWR a_6562_25094# 0.22221f
C1240 a_6540_22112# a_6738_22112# 0.06623f
C1241 a_3695_23038# sar9b_0._07_ 0.02799f
C1242 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.01003f
C1243 sar9b_0.net7 th_dif_sw_0.CK 0.17128f
C1244 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INN 0.0434f
C1245 a_9730_24138# sar9b_0.net12 0.06386f
C1246 a_11722_25838# sar9b_0.net30 0.01802f
C1247 a_7284_20787# sar9b_0.net62 0.023f
C1248 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 ua[0] 0.12378f
C1249 sar9b_0.net3 a_2508_27440# 0.02829f
C1250 a_10218_27466# sar9b_0.net34 0.05477f
C1251 sar9b_0.net27 single_9b_cdac_1.CF[2] 0.07174f
C1252 a_10742_27751# single_9b_cdac_0.SW[7] 0.02243f
C1253 a_10528_20155# sar9b_0.net51 0.04328f
C1254 single_9b_cdac_1.CF[7] sar9b_0.net29 0.04004f
C1255 single_9b_cdac_0.SW[4] a_13067_27662# 0.0479f
C1256 a_11436_17742# sar9b_0.net27 0.04295f
C1257 a_11430_27595# a_11776_27801# 0.07649f
C1258 a_6346_23773# sar9b_0.net54 0.1286f
C1259 a_62748_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.23864f
C1260 VDPWR a_5581_20992# 0.1971f
C1261 a_8031_26141# a_8345_26455# 0.07826f
C1262 sar9b_0.net72 sar9b_0._14_ 1.15565f
C1263 a_10830_19068# sar9b_0.net2 0.018f
C1264 a_8057_18463# sar9b_0.net73 0.07314f
C1265 VDPWR th_dif_sw_0.VCP 6.87158f
C1266 VDPWR single_9b_cdac_0.SW[2] 2.53031f
C1267 sar9b_0.net13 a_7338_24802# 0.07649f
C1268 a_6783_19481# sar9b_0.net47 0.24046f
C1269 sar9b_0.net65 sar9b_0.clknet_1_0__leaf_CLK 0.03848f
C1270 single_9b_cdac_1.SW[5] sar9b_0.net28 0.01641f
C1271 VDPWR a_8726_22954# 0.22795f
C1272 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02513f
C1273 single_9b_cdac_1.SW[3] sar9b_0.net36 0.01142f
C1274 sar9b_0.net40 a_11382_19478# 0.06135f
C1275 a_8591_22855# sar9b_0.net37 0.01032f
C1276 a_7347_24160# sar9b_0.net54 0.37926f
C1277 a_7193_22459# a_7978_22202# 0.26257f
C1278 sar9b_0._01_ a_5481_20185# 0.0279f
C1279 sar9b_0.net55 a_6484_22845# 0.01609f
C1280 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02589f
C1281 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[4] 0.0149f
C1282 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_10254_2858# 1.3306f
C1283 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[7] 0.06961f
C1284 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96985f
C1285 sar9b_0.net8 sar9b_0.net42 0.01991f
C1286 a_8098_18810# sar9b_0.net48 0.09937f
C1287 sar9b_0._04_ sar9b_0.net69 0.13306f
C1288 sar9b_0.net13 a_10607_25185# 0.06161f
C1289 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.42014f
C1290 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.12898f
C1291 VDPWR a_2508_26108# 0.21993f
C1292 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 2.71729f
C1293 sar9b_0.net57 a_8438_23755# 0.02145f
C1294 a_13011_21906# single_9b_cdac_1.CF[2] 0.08337f
C1295 VDPWR a_5844_18123# 0.83758f
C1296 a_9174_17906# a_9839_17527# 0.19065f
C1297 a_9450_17846# a_9974_17626# 0.04522f
C1298 a_58824_17740# single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22352f
C1299 a_7926_23234# a_8386_22806# 0.26257f
C1300 a_8202_23174# a_8591_22855# 0.05462f
C1301 single_9b_cdac_1.SW[2] a_9974_17626# 0.02309f
C1302 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 2.82231f
C1303 tdc_0.OUTP a_10194_16784# 0.02444f
C1304 a_11434_16874# a_10649_17131# 0.26257f
C1305 uo_out[2] uo_out[0] 0.01052f
C1306 sar9b_0.net44 a_6282_27170# 0.02958f
C1307 sar9b_0.net60 a_6250_28502# 0.06687f
C1308 VDPWR a_10932_25713# 0.81346f
C1309 sar9b_0.net26 sar9b_0.net5 0.02305f
C1310 a_5846_17626# sar9b_0.net56 0.02562f
C1311 VDPWR a_2931_28566# 0.47184f
C1312 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1313 a_7092_19455# a_7374_19685# 0.05462f
C1314 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26955f
C1315 a_7289_21127# sar9b_0.net35 0.02113f
C1316 a_5010_28495# a_5674_28147# 0.16939f
C1317 a_6030_24396# a_5962_24151# 0.35559f
C1318 ua[0] single_9b_cdac_1.SW[7] 0.13071f
C1319 a_11382_18146# sar9b_0.net73 0.16947f
C1320 single_9b_cdac_0.SW[7] a_10607_27849# 0.02998f
C1321 a_10378_27170# sar9b_0.net36 0.05314f
C1322 a_9270_24566# sar9b_0.net53 0.22967f
C1323 a_6534_17799# sar9b_0.net46 0.2223f
C1324 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.03729f
C1325 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[6] 0.01887f
C1326 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.37833f
C1327 VDPWR a_6130_20239# 0.38534f
C1328 single_9b_cdac_0.SW[4] a_43540_26999# 0.28324f
C1329 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[3] 0.02029f
C1330 sar9b_0._12_ sar9b_0.net39 0.48411f
C1331 a_11718_23127# clk 0.01747f
C1332 sar9b_0.net41 a_10227_18142# 0.01117f
C1333 a_5581_20992# sar9b_0._17_ 0.04255f
C1334 a_10506_23174# sar9b_0.net74 0.05564f
C1335 a_3206_22432# sar9b_0.clknet_1_1__leaf_CLK 0.06142f
C1336 a_11008_17491# a_11436_17742# 0.01819f
C1337 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A a_30717_15495# 0.01076f
C1338 sar9b_0.net33 sar9b_0.net74 0.12313f
C1339 single_9b_cdac_0.SW[1] sar9b_0.net33 0.06514f
C1340 VDPWR a_16185_13034# 0.19332f
C1341 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.01514f
C1342 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.69086f
C1343 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] 1.15121f
C1344 a_8057_18463# sar9b_0.net46 0.10239f
C1345 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.11216f
C1346 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[2] 0.07133f
C1347 a_5331_16810# sar9b_0.net27 0.05702f
C1348 single_9b_cdac_0.SW[2] sar9b_0.net29 0.33939f
C1349 single_9b_cdac_1.CF[3] ua[0] 3.58897f
C1350 sar9b_0.net27 a_12618_22138# 0.02584f
C1351 a_5581_20992# sar9b_0._08_ 0.16775f
C1352 sar9b_0.net72 sar9b_0._16_ 0.06363f
C1353 VDPWR a_8334_17021# 0.2535f
C1354 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP a_62748_16877# 0.04592f
C1355 sar9b_0.net30 sar9b_0.net52 0.05789f
C1356 single_9b_cdac_1.SW[1] th_dif_sw_0.VCN 0.0955f
C1357 sar9b_0.net51 sar9b_0.net73 0.03243f
C1358 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07579f
C1359 sar9b_0.net70 sar9b_0.net69 0.12146f
C1360 sar9b_0.net35 sar9b_0.net37 0.35869f
C1361 sar9b_0.net27 a_12870_23599# 0.02852f
C1362 sar9b_0.net25 uo_out[1] 0.06669f
C1363 sar9b_0.net61 a_9974_17626# 0.04925f
C1364 a_10470_21795# a_10816_21487# 0.07649f
C1365 sar9b_0.net6 a_11859_20574# 0.01121f
C1366 a_10335_16817# a_10649_17131# 0.07826f
C1367 VDPWR a_8334_18353# 0.25378f
C1368 a_25915_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.01076f
C1369 sar9b_0.net2 sar9b_0.net37 0.03346f
C1370 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C1371 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[0] 0.06503f
C1372 ui_in[2] ui_in[1] 0.03102f
C1373 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[3] 0.26707f
C1374 sar9b_0.net63 sar9b_0.net11 0.60944f
C1375 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 ua[0] 0.12358f
C1376 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.SW[2] 0.17199f
C1377 sar9b_0.net52 a_9942_24806# 0.20968f
C1378 VDPWR a_6307_27584# 0.36193f
C1379 a_7188_22119# a_7193_22459# 0.43491f
C1380 a_8334_18353# sar9b_0.net1 0.01172f
C1381 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.11216f
C1382 sar9b_0.net70 sar9b_0._18_ 0.03792f
C1383 sar9b_0.net23 single_9b_cdac_0.SW[8] 0.02815f
C1384 sar9b_0.net48 a_5844_18123# 0.18591f
C1385 a_18214_3039# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.33121f
C1386 sar9b_0.net11 sar9b_0.net62 0.20455f
C1387 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46159_29911# 0.01076f
C1388 a_9760_22819# clk 0.01624f
C1389 a_11382_18146# sar9b_0.net50 0.23307f
C1390 sar9b_0.net6 sar9b_0.net51 0.0241f
C1391 a_8115_28566# uo_out[6] 0.42188f
C1392 VDPWR a_9450_17846# 0.85429f
C1393 VDPWR a_12047_23853# 0.26429f
C1394 single_9b_cdac_1.SW[3] a_11382_18146# 0.03693f
C1395 sar9b_0.net31 sar9b_0.net45 0.06702f
C1396 sar9b_0.net65 sar9b_0._12_ 0.02841f
C1397 VDPWR single_9b_cdac_1.SW[2] 2.86879f
C1398 sar9b_0.net43 sar9b_0.net13 0.02924f
C1399 VDPWR a_6484_22845# 0.26318f
C1400 a_10553_18922# sar9b_0.net7 0.06335f
C1401 VDPWR a_11104_24151# 0.19368f
C1402 a_11382_26138# sar9b_0.net12 0.03109f
C1403 sar9b_0.net50 a_11859_20574# 0.05205f
C1404 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.10429f
C1405 a_7306_19777# sar9b_0.net10 0.04467f
C1406 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[3] 0.06019f
C1407 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_26951_15501# 0.01076f
C1408 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.03484f
C1409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] 3.1021f
C1410 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.clk_div_0.COUNT\[1\] 0.46155f
C1411 a_12588_16784# single_9b_cdac_1.SW[3] 0.02701f
C1412 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[4] 0.36316f
C1413 single_9b_cdac_1.cdac_sw_9b_0.S[7] th_dif_sw_0.VCP 1.61586f
C1414 a_16527_10454# tdc_0.phase_detector_0.INN 0.10585f
C1415 VDPWR a_9279_27227# 0.27846f
C1416 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.6205f
C1417 a_9472_23805# sar9b_0.net54 0.08291f
C1418 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[3] 14.7461f
C1419 sar9b_0.net52 a_12047_26517# 0.22373f
C1420 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[8] 0.01887f
C1421 a_3206_22432# sar9b_0.net67 0.25532f
C1422 a_9138_27163# sar9b_0.net37 0.04632f
C1423 VDPWR a_12182_18427# 0.20217f
C1424 a_25210_17740# single_9b_cdac_1.SW[8] 0.18991f
C1425 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 3.27833f
C1426 single_9b_cdac_1.SW[6] th_dif_sw_0.VCN 0.09453f
C1427 single_9b_cdac_1.SW[4] th_dif_sw_0.CK 0.04291f
C1428 sar9b_0.net10 clk 0.1264f
C1429 a_11178_20806# sar9b_0.net39 0.01531f
C1430 a_7914_23470# a_8874_23470# 0.03432f
C1431 a_8340_26115# sar9b_0.cyclic_flag_0.FINAL 0.2316f
C1432 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN ua[0] 3.10229f
C1433 a_8166_27595# sar9b_0.net36 0.06865f
C1434 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP 0.04344f
C1435 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C1436 sar9b_0.net47 sar9b_0.net35 0.11331f
C1437 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.12898f
C1438 VDPWR a_14871_9671# 0.67026f
C1439 a_6678_27470# sar9b_0.net60 0.21743f
C1440 a_11658_19474# a_11842_19766# 0.44532f
C1441 sar9b_0.net46 sar9b_0.net51 0.64278f
C1442 VDPWR single_9b_cdac_1.SW[8] 2.60138f
C1443 single_9b_cdac_1.cdac_sw_9b_0.S[8] a_24332_16877# 0.59531f
C1444 sar9b_0.net50 sar9b_0.net51 0.03079f
C1445 a_9802_26815# a_9138_27163# 0.16939f
C1446 sar9b_0.net7 a_10742_21091# 0.06412f
C1447 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP a_29134_26999# 0.04592f
C1448 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.22983f
C1449 a_10649_17131# sar9b_0.net6 0.09326f
C1450 a_3819_24136# sar9b_0.clknet_1_1__leaf_CLK 0.01525f
C1451 sar9b_0.net18 a_2847_27473# 0.03049f
C1452 sar9b_0.net4 a_5535_18149# 0.03052f
C1453 sar9b_0.net26 a_12618_19474# 0.03006f
C1454 a_10830_19068# a_11338_19178# 0.19065f
C1455 single_9b_cdac_0.SW[5] a_12531_28566# 0.03035f
C1456 a_9363_20826# sar9b_0.net37 0.01328f
C1457 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.17533f
C1458 a_10218_24802# sar9b_0.net12 0.06895f
C1459 a_8098_23762# sar9b_0.net62 0.02357f
C1460 a_11915_28371# single_9b_cdac_0.SW[5] 0.0323f
C1461 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.CF[4] 0.12358f
C1462 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.71729f
C1463 sar9b_0.net40 a_6744_23238# 0.02487f
C1464 sar9b_0.net9 sar9b_0.net38 0.32278f
C1465 sar9b_0.net35 sar9b_0.net59 0.93479f
C1466 sar9b_0.net27 sar9b_0.net28 0.01665f
C1467 a_9162_23174# a_9760_22819# 0.06623f
C1468 VDPWR sar9b_0.net9 1.21348f
C1469 sar9b_0.net61 a_8694_20570# 0.18235f
C1470 a_9154_20142# sar9b_0.net51 0.06402f
C1471 a_6137_23791# a_6414_23681# 0.09983f
C1472 a_6534_17799# a_6880_17491# 0.07649f
C1473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[8] 1.50844f
C1474 VDPWR a_8622_26345# 0.28256f
C1475 a_3219_22860# sar9b_0.clk_div_0.COUNT\[1\] 0.21033f
C1476 sar9b_0.net13 sar9b_0.net4 0.20455f
C1477 a_3713_22522# a_3561_22527# 0.22517f
C1478 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[2] 0.01481f
C1479 sar9b_0.net13 sar9b_0._15_ 0.03815f
C1480 sar9b_0._18_ sar9b_0.net60 0.06258f
C1481 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C1482 VDPWR a_6922_23534# 0.2895f
C1483 VDPWR sar9b_0.net61 2.29778f
C1484 a_8334_18353# sar9b_0.net48 0.04696f
C1485 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.05472f
C1486 a_4934_22432# a_5182_22567# 0.05308f
C1487 VDPWR sar9b_0.net44 0.51556f
C1488 sar9b_0.net45 uo_out[7] 0.02028f
C1489 sar9b_0.net9 sar9b_0.net1 0.02842f
C1490 a_6636_20780# sar9b_0.net10 0.29165f
C1491 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C1492 sar9b_0.net44 a_4330_27170# 0.07062f
C1493 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.42784f
C1494 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.03729f
C1495 sar9b_0.net15 sar9b_0.net4 0.47161f
C1496 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[2] 4.15039f
C1497 a_5235_27466# sar9b_0.net59 0.05706f
C1498 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[5] 0.31534f
C1499 sar9b_0.net40 a_10803_19474# 0.07638f
C1500 a_6861_22828# a_6744_23238# 0.3009f
C1501 a_6484_22845# sar9b_0._17_ 0.03367f
C1502 a_3855_25792# a_4293_25852# 0.02614f
C1503 a_4125_25958# a_4365_25770# 0.35097f
C1504 sar9b_0.net58 a_5465_28246# 0.07923f
C1505 sar9b_0.net1 sar9b_0.net61 0.02364f
C1506 VDPWR a_3206_22432# 0.86795f
C1507 a_3946_27530# a_3438_27677# 0.19065f
C1508 a_2739_20140# sar9b_0._00_ 0.0764f
C1509 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.02638f
C1510 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.SW[7] 0.15499f
C1511 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.84426f
C1512 a_3371_23106# a_3219_22860# 0.24998f
C1513 sar9b_0._18_ sar9b_0.net57 0.25105f
C1514 sar9b_0.net24 a_9279_27227# 0.03138f
C1515 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0313f
C1516 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.36013f
C1517 sar9b_0.net48 a_9450_17846# 0.17495f
C1518 a_7638_19238# sar9b_0.net73 0.17598f
C1519 sar9b_0.net27 single_9b_cdac_1.CF[3] 0.12277f
C1520 a_7602_18116# a_8266_18445# 0.16939f
C1521 sar9b_0.net43 sar9b_0.net23 0.30643f
C1522 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31753_15501# 0.01076f
C1523 sar9b_0.net48 single_9b_cdac_1.SW[2] 0.7306f
C1524 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.17533f
C1525 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR 0.62553f
C1526 sar9b_0.net52 sar9b_0.net54 0.82593f
C1527 a_5849_18463# a_6058_18445# 0.24088f
C1528 a_5844_18123# a_6634_18206# 0.1263f
C1529 sar9b_0.net26 single_9b_cdac_1.SW[1] 0.02116f
C1530 a_7138_27758# a_7914_27466# 0.3578f
C1531 VDPWR a_3822_27060# 0.26946f
C1532 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[0] 0.02666f
C1533 tdc_0.OUTN a_8057_17131# 0.03327f
C1534 sar9b_0.net7 sar9b_0.net38 0.02694f
C1535 a_3822_27060# a_4330_27170# 0.19065f
C1536 VDPWR a_2892_27039# 0.25024f
C1537 sar9b_0.net40 a_6678_27470# 0.17609f
C1538 a_9442_21474# sar9b_0.net38 0.01689f
C1539 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.11216f
C1540 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 0.19147f
C1541 a_4812_28371# uo_out[7] 0.0141f
C1542 sar9b_0.net43 a_9593_26914# 0.01648f
C1543 VDPWR sar9b_0.net7 1.0007f
C1544 sar9b_0.net23 a_8340_26115# 0.02021f
C1545 a_11859_21906# sar9b_0.net39 0.01794f
C1546 VDPWR a_9442_21474# 0.23612f
C1547 a_9942_27470# a_10218_27466# 0.1263f
C1548 VDPWR a_2508_27440# 0.21708f
C1549 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.7611f
C1550 sar9b_0.net59 a_9138_27163# 0.3052f
C1551 sar9b_0.net29 single_9b_cdac_1.SW[8] 0.04274f
C1552 a_12870_22267# a_12618_22138# 0.27388f
C1553 a_11842_22430# a_12047_22521# 0.09983f
C1554 sar9b_0.net4 a_5811_19178# 0.07105f
C1555 VDPWR a_15151_10456# 0.3789f
C1556 sar9b_0.net8 sar9b_0.net39 0.1827f
C1557 single_9b_cdac_1.cdac_sw_9b_0.S[3] a_49221_17740# 0.22497f
C1558 single_9b_cdac_0.SW[3] a_49221_26990# 0.18991f
C1559 VDPWR a_5481_20185# 0.14537f
C1560 a_11466_23174# sar9b_0.net11 0.0513f
C1561 a_9730_24138# a_10506_24506# 0.3578f
C1562 a_5151_28559# a_5460_28377# 0.07766f
C1563 clk tdc_0.phase_detector_0.INN 0.04168f
C1564 a_9442_21474# sar9b_0.net1 0.02634f
C1565 a_2706_27440# a_3161_27787# 0.3578f
C1566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02813f
C1567 sar9b_0.net27 a_13011_24570# 0.04167f
C1568 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1569 sar9b_0.net8 a_8982_21902# 0.17036f
C1570 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.3196f
C1571 sar9b_0._09_ a_5126_20140# 0.01059f
C1572 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_50962_29911# 0.01076f
C1573 sar9b_0.net47 a_7978_22202# 0.20624f
C1574 sar9b_0.net41 a_10662_17799# 0.06166f
C1575 sar9b_0.net22 sar9b_0.net45 0.14216f
C1576 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1577 sar9b_0.net60 uio_out[0] 0.09917f
C1578 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[4] 0.05054f
C1579 sar9b_0.net60 a_5753_24250# 0.01748f
C1580 sar9b_0.net60 a_4332_23043# 0.05573f
C1581 a_13011_21906# single_9b_cdac_1.CF[3] 0.02875f
C1582 a_12182_19759# a_12618_19474# 0.16939f
C1583 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[5] 0.17948f
C1584 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C1585 VDPWR a_4749_27652# 0.4017f
C1586 sar9b_0.net13 a_5748_24381# 0.24967f
C1587 sar9b_0.net60 a_6534_27123# 0.01098f
C1588 a_11842_23762# a_12618_23470# 0.3578f
C1589 single_9b_cdac_1.CF[4] sar9b_0.net28 0.36381f
C1590 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[4] 0.02008f
C1591 sar9b_0.net40 a_12870_19603# 0.07154f
C1592 a_8554_26437# sar9b_0.net59 0.1439f
C1593 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.84059f
C1594 sar9b_0.net52 sar9b_0.net27 0.01796f
C1595 sar9b_0._02_ sar9b_0.net4 0.02372f
C1596 a_3090_27163# sar9b_0.net19 0.05411f
C1597 sar9b_0.net52 single_9b_cdac_0.SW[5] 0.12211f
C1598 a_3425_20244# a_3723_20140# 0.02614f
C1599 single_9b_cdac_1.SW[8] a_12047_19857# 0.03035f
C1600 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1601 sar9b_0.net43 sar9b_0.net63 0.0282f
C1602 a_10707_23470# sar9b_0.net36 0.02924f
C1603 sar9b_0.net61 sar9b_0.net48 0.8171f
C1604 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.11216f
C1605 sar9b_0.net35 a_7404_18116# 0.01538f
C1606 th_dif_sw_0.CK single_9b_cdac_1.SW[1] 0.06557f
C1607 a_9130_26198# a_8340_26115# 0.1263f
C1608 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.17533f
C1609 a_7289_21127# sar9b_0.net56 0.01572f
C1610 a_7498_21109# a_7566_21017# 0.35559f
C1611 a_11382_19478# a_11658_19474# 0.1263f
C1612 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.23119f
C1613 sar9b_0.net57 a_4332_23043# 0.0332f
C1614 sar9b_0.net42 sar9b_0.net73 1.30182f
C1615 a_7638_19238# sar9b_0.net46 0.03287f
C1616 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1617 VDPWR a_11430_24931# 0.26219f
C1618 VDPWR a_5182_22567# 0.0129f
C1619 a_10506_23174# sar9b_0.net53 0.17591f
C1620 sar9b_0.net16 a_5196_19448# 0.27599f
C1621 a_10230_23234# a_10690_22806# 0.26257f
C1622 a_10506_23174# a_10895_22855# 0.05462f
C1623 sar9b_0.net43 sar9b_0.net62 0.65145f
C1624 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[0] 0.06019f
C1625 a_5506_26802# a_6534_27123# 0.07826f
C1626 sar9b_0.net8 single_9b_cdac_1.CF[1] 0.12551f
C1627 single_9b_cdac_0.cdac_sw_9b_0.S[8] th_dif_sw_0.VCN 0.85562f
C1628 a_3161_26455# sar9b_0.net44 0.01837f
C1629 sar9b_0.net20 a_7539_28566# 0.08083f
C1630 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0._05_ 0.02778f
C1631 a_5322_27170# sar9b_0.net39 0.02945f
C1632 single_9b_cdac_0.SW[6] a_33936_26999# 0.28324f
C1633 a_10742_27751# VDPWR 0.20368f
C1634 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38715f
C1635 a_9414_23127# sar9b_0.net11 0.06993f
C1636 sar9b_0.net58 sar9b_0.net39 0.55587f
C1637 a_8591_22855# sar9b_0.net54 0.22373f
C1638 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C1639 a_7882_19538# sar9b_0.net62 0.20424f
C1640 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[3] 12.1694f
C1641 a_3206_22432# sar9b_0.clknet_1_0__leaf_CLK 0.05926f
C1642 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1643 VDPWR a_3819_24136# 0.09178f
C1644 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.03729f
C1645 dw_12589_1395# ua[4] 1.41177f
C1646 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.01472f
C1647 sar9b_0._07_ a_5633_20244# 0.0155f
C1648 a_6954_27466# sar9b_0.net44 0.22029f
C1649 sar9b_0.net32 a_12870_23599# 0.0306f
C1650 a_10926_17021# single_9b_cdac_1.SW[2] 0.01526f
C1651 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.62443f
C1652 VDPWR a_8438_18958# 0.21428f
C1653 a_6767_25185# a_6902_25087# 0.35559f
C1654 a_11382_18146# a_11658_18142# 0.1263f
C1655 a_4365_25770# sar9b_0.clknet_1_1__leaf_CLK 0.06633f
C1656 sar9b_0.net42 sar9b_0.net6 0.02813f
C1657 sar9b_0.net7 sar9b_0.net48 0.22803f
C1658 single_9b_cdac_1.SW[0] sar9b_0.net37 0.06363f
C1659 sar9b_0.net55 sar9b_0.net15 0.43777f
C1660 sar9b_0.net49 a_10402_21098# 0.10002f
C1661 a_7138_27758# a_7343_27849# 0.09983f
C1662 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C1663 a_53154_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.23864f
C1664 a_12618_18142# a_13216_18477# 0.06623f
C1665 sar9b_0.net64 sar9b_0.net60 0.08504f
C1666 sar9b_0.net56 sar9b_0.net37 1.42615f
C1667 sar9b_0.net40 a_5753_24250# 0.01091f
C1668 a_7138_27758# sar9b_0.net21 0.0211f
C1669 sar9b_0.net63 sar9b_0.net4 0.04374f
C1670 sar9b_0.net63 sar9b_0._15_ 0.04597f
C1671 sar9b_0.net40 a_6534_27123# 0.03801f
C1672 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.26707f
C1673 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.84426f
C1674 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.SW[8] 0.22497f
C1675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 a_63626_26990# 0.14695f
C1676 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 ua[0] 0.11944f
C1677 a_11718_23127# sar9b_0.net31 0.01022f
C1678 a_10218_24802# a_10482_25831# 0.02278f
C1679 single_9b_cdac_1.SW[6] th_dif_sw_0.CK 0.11297f
C1680 sar9b_0.net64 sar9b_0.net57 0.02277f
C1681 a_10227_23490# clk 0.01166f
C1682 a_7284_20787# a_7443_21496# 0.02666f
C1683 a_9154_20142# a_9359_20191# 0.09983f
C1684 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.04988f
C1685 sar9b_0.net38 sar9b_0.net5 0.08475f
C1686 a_5196_24776# sar9b_0._03_ 0.10899f
C1687 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C1688 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.6919f
C1689 sar9b_0.net41 a_9760_22819# 0.28794f
C1690 VDPWR sar9b_0.net5 1.99906f
C1691 a_12588_16784# tdc_0.OUTP 0.28954f
C1692 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.06503f
C1693 sar9b_0.net52 sar9b_0.net36 0.10328f
C1694 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62573f
C1695 a_7188_22119# sar9b_0.net47 0.17293f
C1696 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.58106f
C1697 sar9b_0.net42 sar9b_0.net50 0.03413f
C1698 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.0303f
C1699 single_9b_cdac_0.SW[4] a_13164_28398# 0.01356f
C1700 sar9b_0.net55 a_5811_19178# 0.26511f
C1701 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.01173f
C1702 sar9b_0.net1 sar9b_0.net5 0.83129f
C1703 VDPWR a_10607_27849# 0.26664f
C1704 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[1\] 0.17923f
C1705 single_9b_cdac_0.SW[6] uo_out[0] 0.04513f
C1706 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDPWR 0.62555f
C1707 sar9b_0.net74 a_11382_26138# 0.17525f
C1708 sar9b_0.clk_div_0.COUNT\[3\] a_4755_22138# 0.02068f
C1709 a_11382_23474# a_11842_23762# 0.26257f
C1710 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[0] 0.31534f
C1711 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.07579f
C1712 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.03482f
C1713 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.28813f
C1714 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 2.82223f
C1715 uo_out[1] ui_in[0] 0.06797f
C1716 uo_out[0] clk 0.48415f
C1717 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[0] 0.22459f
C1718 sar9b_0._14_ a_2940_25096# 0.01562f
C1719 a_2893_24992# a_3364_25120# 0.01114f
C1720 a_10690_22806# sar9b_0.net36 0.01892f
C1721 sar9b_0.net27 a_5196_18116# 0.2837f
C1722 sar9b_0.net49 a_8970_20510# 0.17751f
C1723 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.02149f
C1724 a_7890_26108# a_8554_26437# 0.16939f
C1725 single_9b_cdac_0.SW[5] uo_out[1] 0.07247f
C1726 a_3713_22522# a_3027_22138# 0.27693f
C1727 sar9b_0.net41 sar9b_0.net10 0.02787f
C1728 single_9b_cdac_1.CF[8] sar9b_0.net28 0.04086f
C1729 a_11859_17910# single_9b_cdac_1.SW[3] 0.01458f
C1730 sar9b_0.net46 a_4771_18260# 0.03699f
C1731 sar9b_0.net35 sar9b_0.net54 0.19733f
C1732 sar9b_0.net13 a_9165_24988# 0.11202f
C1733 sar9b_0.net32 a_12531_28566# 0.02777f
C1734 a_10402_27758# sar9b_0.net59 0.08863f
C1735 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[0] 18.6433f
C1736 sar9b_0.net32 a_11915_28371# 0.04795f
C1737 sar9b_0.net56 sar9b_0.net47 0.18012f
C1738 uio_out[1] uio_out[0] 2.82713f
C1739 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C1740 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.04988f
C1741 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A a_45123_15495# 0.01076f
C1742 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.7611f
C1743 a_7402_22441# a_7470_22349# 0.35559f
C1744 a_6834_20780# sar9b_0.net35 0.03194f
C1745 sar9b_0.net55 sar9b_0._02_ 0.49529f
C1746 a_6744_23238# clk 0.01136f
C1747 sar9b_0.net49 a_10218_21842# 0.2811f
C1748 single_9b_cdac_1.cdac_sw_9b_0.S[3] ua[0] 1.59889f
C1749 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] 3.11836f
C1750 a_10378_27170# sar9b_0.net42 0.16789f
C1751 a_8438_18958# sar9b_0.net48 0.14544f
C1752 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95338f
C1753 VDPWR single_9b_cdac_1.SW[4] 2.6945f
C1754 single_9b_cdac_1.CF[1] a_13011_20574# 0.01474f
C1755 VDPWR a_2706_26108# 0.40591f
C1756 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.SW[8] 0.17661f
C1757 VDPWR a_5535_18149# 0.2712f
C1758 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[0] 0.02356f
C1759 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.19147f
C1760 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[3] 14.7603f
C1761 sar9b_0.net70 sar9b_0._07_ 0.01892f
C1762 tdc_0.OUTP a_10649_17131# 0.06549f
C1763 VDPWR a_11214_25728# 0.25894f
C1764 a_7374_19685# a_7882_19538# 0.19065f
C1765 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[3] 0.01497f
C1766 sar9b_0.net13 sar9b_0.net38 0.02597f
C1767 a_12560_27128# sar9b_0.net52 0.08336f
C1768 a_3206_22432# sar9b_0._12_ 0.04817f
C1769 sar9b_0.net60 sar9b_0.net37 0.02643f
C1770 a_7092_19455# a_7882_19538# 0.1263f
C1771 a_4947_20140# sar9b_0._10_ 0.0624f
C1772 VDPWR sar9b_0.net13 2.18619f
C1773 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.37833f
C1774 sar9b_0.net20 sar9b_0.net45 0.05044f
C1775 a_5753_24250# a_6538_24506# 0.26257f
C1776 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36041f
C1777 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.51772f
C1778 sar9b_0.net31 sar9b_0.net10 0.16278f
C1779 VDPWR a_29134_16877# 1.81495f
C1780 a_9730_24138# sar9b_0.net53 0.08408f
C1781 th_dif_sw_0.CKB ua[0] 0.02532f
C1782 a_8266_17113# sar9b_0.net27 0.02296f
C1783 sar9b_0.net63 sar9b_0.clknet_1_1__leaf_CLK 0.02378f
C1784 VDPWR sar9b_0.cyclic_flag_0.FINAL 0.90593f
C1785 sar9b_0.net35 sar9b_0.net27 0.08696f
C1786 single_9b_cdac_0.SW[8] uo_out[4] 0.18749f
C1787 a_35519_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A 0.01076f
C1788 VDPWR sar9b_0.net15 0.41783f
C1789 a_13067_27662# sar9b_0.net28 0.22031f
C1790 sar9b_0.net48 sar9b_0.net5 0.3854f
C1791 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.93403f
C1792 single_9b_cdac_0.cdac_sw_9b_0.S[1] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.31809f
C1793 sar9b_0.net16 sar9b_0.net46 0.16498f
C1794 sar9b_0.net2 sar9b_0.net27 0.34591f
C1795 a_11436_17742# a_11859_17910# 0.05125f
C1796 VDPWR a_5711_26851# 0.26739f
C1797 sar9b_0.net57 sar9b_0.net37 0.18597f
C1798 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.02513f
C1799 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.01515f
C1800 a_5506_26802# sar9b_0.net37 0.11789f
C1801 sar9b_0.net40 a_6767_25185# 0.02519f
C1802 sar9b_0.net53 a_12182_22423# 0.14409f
C1803 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C1804 sar9b_0.net27 a_13011_27234# 0.22439f
C1805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.03729f
C1806 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[4] 0.02019f
C1807 VDPWR a_4365_25770# 0.1412f
C1808 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.84061f
C1809 sar9b_0.net63 sar9b_0.net55 0.27808f
C1810 a_11722_25838# sar9b_0.net12 0.01432f
C1811 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36555_29911# 0.01076f
C1812 tdc_0.OUTN sar9b_0.net46 0.09655f
C1813 a_2940_25096# sar9b_0._16_ 0.11593f
C1814 VDPWR a_8019_17910# 0.39892f
C1815 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.75849f
C1816 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.81423f
C1817 a_4812_28371# sar9b_0.net20 0.3101f
C1818 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[6] 0.0149f
C1819 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.03729f
C1820 sar9b_0.net53 a_11842_23762# 0.09947f
C1821 sar9b_0.net57 a_8202_23174# 0.01828f
C1822 th_dif_sw_0.CK tdc_0.RDY 0.05459f
C1823 sar9b_0.net41 a_9839_17527# 0.06481f
C1824 VDPWR a_8842_16874# 0.29337f
C1825 sar9b_0.net36 a_10623_25895# 0.01701f
C1826 a_3747_25724# a_4125_25958# 0.0649f
C1827 a_3372_25734# sar9b_0.clk_div_0.COUNT\[1\] 0.12822f
C1828 a_10218_20806# a_10402_21098# 0.44532f
C1829 VDPWR tdc_0.phase_detector_0.INP 0.59622f
C1830 sar9b_0.net49 a_10607_21189# 0.22001f
C1831 sar9b_0.net55 sar9b_0.net62 0.19573f
C1832 a_10284_25707# a_10482_25831# 0.06623f
C1833 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.02666f
C1834 sar9b_0.net27 a_13216_23805# 0.01206f
C1835 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 1.71649f
C1836 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1837 a_8019_17910# sar9b_0.net1 0.01265f
C1838 sar9b_0._01_ a_4947_20140# 0.16646f
C1839 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.81434f
C1840 VDPWR a_5811_19178# 0.21566f
C1841 a_5506_17478# a_5322_17846# 0.43491f
C1842 a_11658_26134# a_11842_26426# 0.44532f
C1843 a_8098_23762# sar9b_0.net11 0.05862f
C1844 VDPWR a_8842_18206# 0.30615f
C1845 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VDPWR 0.75853f
C1846 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 3.10626f
C1847 a_7914_23470# sar9b_0.net54 0.03451f
C1848 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[2] 0.42016f
C1849 VDPWR a_12618_19474# 0.35538f
C1850 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.22879f
C1851 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.SW[0] 0.14962f
C1852 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[7] 0.12898f
C1853 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0313f
C1854 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.95338f
C1855 sar9b_0.net32 sar9b_0.net52 0.06191f
C1856 sar9b_0._07_ sar9b_0.net60 0.56326f
C1857 a_6250_28502# sar9b_0.net45 0.03629f
C1858 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.12431f
C1859 clk single_9b_cdac_0.SW[0] 0.23595f
C1860 sar9b_0.net40 sar9b_0.net37 0.05789f
C1861 a_8842_18206# sar9b_0.net1 0.03616f
C1862 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.75853f
C1863 VDPWR a_5674_28147# 0.19864f
C1864 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.SW[7] 0.05167f
C1865 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[0] 0.02181f
C1866 sar9b_0.clk_div_0.COUNT\[1\] sar9b_0.net39 0.0203f
C1867 a_11842_18434# sar9b_0.net27 0.01125f
C1868 single_9b_cdac_1.cdac_sw_9b_0.S[0] a_63626_17740# 0.22513f
C1869 sar9b_0.net59 a_3156_26115# 0.17719f
C1870 a_9472_23805# sar9b_0.net12 0.27258f
C1871 sar9b_0.net48 a_5535_18149# 0.17429f
C1872 sar9b_0.net73 sar9b_0.net39 0.09841f
C1873 sar9b_0.cyclic_flag_0.FINAL a_8883_27466# 0.28976f
C1874 sar9b_0.net24 sar9b_0.cyclic_flag_0.FINAL 0.01327f
C1875 a_5580_24776# a_6102_24806# 0.01519f
C1876 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.17461f
C1877 a_5182_22567# sar9b_0._12_ 0.01992f
C1878 a_9174_17906# sar9b_0.net37 0.03941f
C1879 sar9b_0.net23 sar9b_0.net38 0.02577f
C1880 sar9b_0.net59 sar9b_0.net60 0.37207f
C1881 a_11382_18146# a_12047_18525# 0.19065f
C1882 sar9b_0.net47 sar9b_0.net57 0.03056f
C1883 sar9b_0._07_ sar9b_0.net57 1.15961f
C1884 a_3161_26455# a_2706_26108# 0.3578f
C1885 VDPWR sar9b_0._02_ 0.67644f
C1886 sar9b_0.net23 VDPWR 1.79675f
C1887 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[2] 0.03797f
C1888 a_6642_19448# a_6444_19448# 0.06623f
C1889 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.clk_div_0.COUNT\[2\] 0.31022f
C1890 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 2.82223f
C1891 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.SW[3] 0.019f
C1892 sar9b_0.net60 a_5823_23477# 0.03124f
C1893 a_11008_17491# sar9b_0.net2 0.03502f
C1894 single_9b_cdac_0.SW[8] th_dif_sw_0.VCN 0.15316f
C1895 a_7590_24931# a_7936_25137# 0.07649f
C1896 sar9b_0.net9 a_10506_23174# 0.21399f
C1897 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[2] 0.02038f
C1898 sar9b_0.net38 a_9593_26914# 0.0231f
C1899 a_5196_24776# sar9b_0.clk_div_0.COUNT\[2\] 0.28871f
C1900 a_13011_16810# th_dif_sw_0.CK 0.0156f
C1901 single_9b_cdac_1.SW[0] ua[0] 1.99402f
C1902 a_11718_23127# sar9b_0.net10 0.07252f
C1903 VDPWR a_9593_26914# 0.22537f
C1904 sar9b_0.net2 sar9b_0.net36 1.60268f
C1905 VDPWR a_5083_21100# 0.18914f
C1906 a_9930_20510# sar9b_0.net5 0.07266f
C1907 sar9b_0.net6 sar9b_0.net39 0.02562f
C1908 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.31534f
C1909 VDPWR single_9b_cdac_1.SW[1] 2.46863f
C1910 a_8512_27801# sar9b_0.net36 0.04404f
C1911 VDPWR a_3603_28156# 0.4289f
C1912 ua[4] w_12795_1601# 0.89427f
C1913 VDPWR a_15265_9613# 0.18873f
C1914 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.26942f
C1915 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.11216f
C1916 a_5235_27466# sar9b_0.net36 0.073f
C1917 a_13011_25902# sar9b_0.net27 0.0399f
C1918 sar9b_0.net57 a_5823_23477# 0.0298f
C1919 a_11658_19474# a_12870_19603# 0.07766f
C1920 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46159_15501# 0.01076f
C1921 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[4] 0.20642f
C1922 a_9802_26815# a_9588_27045# 0.05022f
C1923 sar9b_0.net7 a_11178_20806# 0.04419f
C1924 sar9b_0._07_ a_5443_19074# 0.02952f
C1925 a_10218_21842# a_10218_20806# 0.01915f
C1926 a_3695_23038# sar9b_0.clk_div_0.COUNT\[0\] 0.14551f
C1927 sar9b_0.net27 sar9b_0._06_ 0.01706f
C1928 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1929 a_5938_22378# sar9b_0.clk_div_0.COUNT\[0\] 0.11986f
C1930 single_9b_cdac_0.SW[5] sar9b_0._06_ 0.01662f
C1931 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C1932 a_4332_23043# clk 0.4678f
C1933 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.SW[2] 0.15027f
C1934 sar9b_0.net47 sar9b_0.net40 0.3867f
C1935 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.7611f
C1936 a_6346_23773# a_6414_23681# 0.35559f
C1937 a_9494_20290# sar9b_0.net51 0.05999f
C1938 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C1939 VDPWR a_9130_26198# 0.30205f
C1940 sar9b_0.net8 single_9b_cdac_1.SW[8] 0.05906f
C1941 sar9b_0.net36 a_10758_24459# 0.02391f
C1942 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[1\] 0.02971f
C1943 a_10194_16784# single_9b_cdac_1.SW[0] 0.02286f
C1944 ui_in[7] ui_in[6] 0.03102f
C1945 sar9b_0.net52 sar9b_0.net12 0.59278f
C1946 a_10239_19235# sar9b_0.net26 0.06761f
C1947 a_8842_18206# sar9b_0.net48 0.06788f
C1948 sar9b_0.net28 a_13216_18477# 0.28248f
C1949 a_2508_23444# sar9b_0.clknet_0_CLK 0.46608f
C1950 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C1951 a_8874_19178# a_7914_19178# 0.03471f
C1952 a_11859_21906# sar9b_0.net9 0.06677f
C1953 sar9b_0.net50 sar9b_0.net39 0.78191f
C1954 VDPWR sar9b_0.net63 1.51034f
C1955 a_2451_27234# ui_in[0] 0.24933f
C1956 VDPWR a_6879_22145# 0.27369f
C1957 single_9b_cdac_1.SW[3] sar9b_0.net39 0.0537f
C1958 a_43540_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.23864f
C1959 tdc_0.phase_detector_0.pd_out_0.A a_16970_11404# 0.18949f
C1960 single_9b_cdac_1.cdac_sw_9b_0.S[7] a_29134_16877# 0.59531f
C1961 sar9b_0.net36 a_9138_27163# 0.04377f
C1962 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.27833f
C1963 sar9b_0.net23 sar9b_0.net24 0.18313f
C1964 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.19143f
C1965 sar9b_0.net40 sar9b_0.net59 0.03006f
C1966 sar9b_0._02_ sar9b_0._17_ 0.15132f
C1967 sar9b_0.net9 sar9b_0.net8 0.25322f
C1968 sar9b_0.net26 sar9b_0.net11 0.03443f
C1969 a_8595_17910# a_8052_16791# 0.03549f
C1970 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C1971 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.11216f
C1972 a_7188_22119# sar9b_0.net54 0.01061f
C1973 m2_23774_26966# single_9b_cdac_0.SW[8] 0.02037f
C1974 a_3369_24181# sar9b_0.clk_div_0.COUNT\[1\] 0.0204f
C1975 a_8334_17021# a_8057_17131# 0.09983f
C1976 sar9b_0.net2 a_9935_24187# 0.06094f
C1977 sar9b_0.net7 a_9942_20810# 0.21228f
C1978 VDPWR sar9b_0.net62 2.17291f
C1979 a_4125_25958# a_4698_25851# 0.04602f
C1980 a_3747_25724# sar9b_0.clknet_1_1__leaf_CLK 0.10609f
C1981 a_3371_23106# sar9b_0.net65 0.03052f
C1982 a_3219_22860# a_3695_23038# 0.08279f
C1983 single_9b_cdac_1.CF[1] sar9b_0.net6 0.01228f
C1984 sar9b_0.net8 sar9b_0.net61 0.19337f
C1985 a_10218_24802# a_10402_25094# 0.44532f
C1986 VDPWR a_2739_20140# 0.47557f
C1987 sar9b_0.net24 a_9593_26914# 0.11222f
C1988 VDPWR single_9b_cdac_1.SW[6] 2.4631f
C1989 a_5083_21100# sar9b_0._17_ 0.01853f
C1990 sar9b_0.net32 uo_out[1] 0.22658f
C1991 a_8057_18463# a_8266_18445# 0.24088f
C1992 sar9b_0.net43 sar9b_0.net11 0.02461f
C1993 a_14897_9355# a_14871_9671# 0.06748f
C1994 a_21684_3438# VDPWR 0.07087f
C1995 a_8166_27595# a_7914_27466# 0.27388f
C1996 single_9b_cdac_1.SW[0] a_10410_17846# 0.04572f
C1997 single_9b_cdac_0.SW[7] th_dif_sw_0.VCN 0.0955f
C1998 sar9b_0.net53 sar9b_0.net73 0.13314f
C1999 VDPWR a_3231_27227# 0.28136f
C2000 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.36301f
C2001 a_10859_26330# a_10937_25582# 0.01019f
C2002 sar9b_0.net20 uo_out[7] 0.0338f
C2003 a_6132_23451# sar9b_0.net11 0.06939f
C2004 VDPWR a_9782_21622# 0.20774f
C2005 a_3540_27045# a_3545_26914# 0.44532f
C2006 VDPWR a_11339_27039# 0.48115f
C2007 a_6678_27470# sar9b_0.net45 0.08442f
C2008 VDPWR a_2706_27440# 0.37404f
C2009 sar9b_0.net59 a_9588_27045# 0.18035f
C2010 a_12618_22138# a_13216_22473# 0.06623f
C2011 a_10218_20806# a_10607_21189# 0.06034f
C2012 sar9b_0.net42 single_9b_cdac_1.SW[7] 0.01299f
C2013 a_3946_27530# sar9b_0.net36 0.17818f
C2014 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 2.82171f
C2015 sar9b_0.net48 single_9b_cdac_1.SW[1] 0.05838f
C2016 a_5460_28377# a_5465_28246# 0.44532f
C2017 single_9b_cdac_0.SW[4] a_44418_26990# 0.18991f
C2018 sar9b_0.net7 a_11859_21906# 0.21737f
C2019 a_3603_28156# a_4083_28566# 0.03385f
C2020 a_3014_24136# sar9b_0.clk_div_0.COUNT\[1\] 0.0121f
C2021 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[2] 0.34042f
C2022 single_9b_cdac_0.cdac_sw_9b_0.S[5] th_dif_sw_0.VCN 6.58553f
C2023 a_2706_27440# a_3370_27769# 0.16939f
C2024 a_3156_27447# a_3438_27677# 0.05462f
C2025 uio_in[3] uio_in[2] 0.03102f
C2026 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.CF[4] 0.01514f
C2027 sar9b_0.net57 a_9942_24806# 0.04118f
C2028 sar9b_0.net7 sar9b_0.net8 0.39284f
C2029 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[2] 16.7662f
C2030 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01175f
C2031 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.84427f
C2032 a_38738_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.23864f
C2033 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.17533f
C2034 sar9b_0._05_ a_3027_21906# 0.07466f
C2035 sar9b_0.net63 sar9b_0._17_ 0.1985f
C2036 a_11436_17742# sar9b_0.net39 0.01601f
C2037 single_9b_cdac_0.cdac_sw_9b_0.S[0] clk 0.03331f
C2038 a_6738_22112# a_6879_22145# 0.27388f
C2039 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[0] 0.17948f
C2040 single_9b_cdac_0.SW[7] a_30012_26990# 0.18991f
C2041 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] 1.20704f
C2042 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.42016f
C2043 a_12870_23599# a_12618_23470# 0.27388f
C2044 a_11842_23762# a_12047_23853# 0.09983f
C2045 sar9b_0.net19 a_3754_26815# 0.0389f
C2046 a_10402_27758# single_9b_cdac_0.SW[5] 0.013f
C2047 sar9b_0.net54 a_6902_25087# 0.12912f
C2048 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.95338f
C2049 sar9b_0.net40 a_6880_26815# 0.01367f
C2050 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[7] 0.0149f
C2051 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[8] 4.67496f
C2052 sar9b_0.net44 a_5322_27170# 0.25565f
C2053 VDPWR a_10482_3438# 0.07094f
C2054 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.19266f
C2055 sar9b_0.net11 sar9b_0.net4 0.02493f
C2056 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.3196f
C2057 a_6642_19448# a_6783_19481# 0.27388f
C2058 sar9b_0.net58 sar9b_0.net44 1.08603f
C2059 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.03729f
C2060 single_9b_cdac_1.SW[8] single_9b_cdac_1.CF[0] 3.87975f
C2061 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[3] 14.7603f
C2062 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.31534f
C2063 a_12588_16784# sar9b_0.net2 0.14533f
C2064 a_11382_19478# a_11842_19766# 0.26257f
C2065 a_2892_23070# sar9b_0.net66 0.14576f
C2066 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C2067 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C2068 sar9b_0.net27 single_9b_cdac_1.SW[0] 0.02138f
C2069 a_8098_18810# sar9b_0.net46 0.03666f
C2070 a_6922_23534# a_6137_23791# 0.26257f
C2071 VDPWR a_11776_25137# 0.19971f
C2072 single_9b_cdac_1.SW[5] sar9b_0.net40 0.09333f
C2073 a_34814_17740# single_9b_cdac_1.SW[6] 0.18991f
C2074 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C2075 sar9b_0.net41 a_9546_24506# 0.01299f
C2076 sar9b_0.clk_div_0.COUNT\[3\] a_4812_21738# 0.29499f
C2077 sar9b_0.net56 sar9b_0.net27 0.19838f
C2078 sar9b_0.net63 a_5682_23444# 0.04284f
C2079 a_11842_26426# a_12870_26263# 0.07826f
C2080 tdc_0.OUTP tdc_0.OUTN 1.54073f
C2081 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.02632f
C2082 sar9b_0.net35 a_7402_22441# 0.01975f
C2083 sar9b_0.net35 sar9b_0.net51 0.08262f
C2084 sar9b_0.net60 a_4496_20468# 0.09564f
C2085 single_9b_cdac_1.SW[8] a_13011_20574# 0.01361f
C2086 sar9b_0._09_ sar9b_0._18_ 0.1776f
C2087 a_11178_27466# VDPWR 0.35818f
C2088 a_5046_27230# sar9b_0.net39 0.19915f
C2089 a_8874_23470# clk 0.01286f
C2090 sar9b_0.net2 sar9b_0.net51 0.02425f
C2091 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36044f
C2092 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[2] 16.4998f
C2093 sar9b_0.net61 a_8057_17131# 0.03749f
C2094 a_7138_27758# sar9b_0.net44 0.0155f
C2095 sar9b_0.net58 a_3822_27060# 0.22673f
C2096 a_11722_25838# sar9b_0.net74 0.21463f
C2097 sar9b_0.net32 a_13216_23805# 0.28438f
C2098 sar9b_0.net17 a_2508_26108# 0.28355f
C2099 sar9b_0.net39 sar9b_0._03_ 0.13967f
C2100 a_9270_24566# sar9b_0.net62 0.16799f
C2101 sar9b_0.clknet_1_0__leaf_CLK a_2739_20140# 0.35818f
C2102 a_11382_18146# a_11842_18434# 0.26257f
C2103 VDPWR a_4811_23656# 0.24092f
C2104 sar9b_0.net27 a_12684_20379# 0.01643f
C2105 VDPWR a_7374_19685# 0.26931f
C2106 a_12560_27128# sar9b_0._06_ 0.0956f
C2107 sar9b_0.net49 a_11430_20935# 0.17358f
C2108 sar9b_0.net42 sar9b_0.net52 0.15052f
C2109 VDPWR a_4947_20140# 0.39022f
C2110 sar9b_0.net17 a_2931_28566# 0.22067f
C2111 a_2547_28132# sar9b_0.net60 0.23163f
C2112 a_4698_25851# sar9b_0.clknet_1_1__leaf_CLK 0.02594f
C2113 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 a_39616_26990# 0.14695f
C2114 VDPWR a_7092_19455# 0.85935f
C2115 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[2] 0.02011f
C2116 VDPWR a_11466_23174# 0.34557f
C2117 single_9b_cdac_0.SW[1] sar9b_0.net28 0.04119f
C2118 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 ua[0] 0.11907f
C2119 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 2.71729f
C2120 a_13011_27234# a_13067_27662# 0.01136f
C2121 VDPWR a_8052_18123# 0.76662f
C2122 single_9b_cdac_1.CF[6] sar9b_0.net28 0.04016f
C2123 sar9b_0.net60 sar9b_0.net54 0.10669f
C2124 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C2125 a_10926_17021# single_9b_cdac_1.SW[1] 0.02544f
C2126 a_10742_25087# sar9b_0.net36 0.01344f
C2127 clk sar9b_0.net37 0.04254f
C2128 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.31534f
C2129 uo_out[2] ui_in[0] 0.0679f
C2130 a_65367_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C2131 a_10218_24802# a_10932_25713# 0.04762f
C2132 VDPWR tdc_0.RDY 0.57898f
C2133 sar9b_0.net19 uo_out[7] 0.03323f
C2134 single_9b_cdac_0.SW[5] uo_out[2] 0.04146f
C2135 a_6378_24802# a_6562_25094# 0.44532f
C2136 VDPWR a_3747_25724# 0.37697f
C2137 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.26684f
C2138 sar9b_0.net6 a_5844_18123# 0.23512f
C2139 a_10707_23470# sar9b_0.net74 0.16592f
C2140 a_10690_22806# sar9b_0.net42 0.01178f
C2141 sar9b_0._09_ a_4072_19474# 0.06295f
C2142 a_9359_20191# a_9494_20290# 0.35559f
C2143 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] 1.15121f
C2144 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.45521f
C2145 sar9b_0._09_ sar9b_0.net71 0.06932f
C2146 a_8052_18123# sar9b_0.net1 0.02679f
C2147 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 2.82181f
C2148 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.08121f
C2149 sar9b_0.net58 a_4749_27652# 0.34567f
C2150 sar9b_0._12_ sar9b_0._02_ 0.12883f
C2151 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[8] 4.16613f
C2152 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.12431f
C2153 sar9b_0.net38 uo_out[6] 0.72968f
C2154 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01152f
C2155 sar9b_0.net52 a_10482_25831# 0.33514f
C2156 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[2\] 1.2616f
C2157 a_8202_23174# clk 0.02077f
C2158 sar9b_0.net57 sar9b_0.net54 1.01482f
C2159 sar9b_0.net31 a_11658_22138# 0.02838f
C2160 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.45521f
C2161 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.28523f
C2162 a_13011_24802# single_9b_cdac_0.SW[0] 0.35451f
C2163 VDPWR uo_out[6] 0.80816f
C2164 sar9b_0.net55 a_6579_18832# 0.01696f
C2165 VDPWR a_24332_16877# 1.81495f
C2166 sar9b_0.net38 a_8115_28566# 0.08106f
C2167 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 1.71649f
C2168 a_3262_24141# sar9b_0.clknet_1_1__leaf_CLK 0.01978f
C2169 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.12358f
C2170 single_9b_cdac_1.CF[8] a_13011_25902# 0.35919f
C2171 sar9b_0.net2 sar9b_0.net12 0.20768f
C2172 VDPWR a_8115_28566# 0.46684f
C2173 sar9b_0.net36 single_9b_cdac_1.SW[0] 0.14f
C2174 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[3] 0.01995f
C2175 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.12898f
C2176 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.69086f
C2177 a_11658_23470# a_12182_23755# 0.05022f
C2178 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.net64 0.02988f
C2179 sar9b_0.net8 sar9b_0.net5 0.02967f
C2180 a_9363_20826# sar9b_0.net51 0.24159f
C2181 a_11434_16874# sar9b_0.net61 0.25057f
C2182 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[0] 0.22459f
C2183 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[3] 0.02091f
C2184 VDPWR a_7284_20787# 0.86664f
C2185 sar9b_0.net18 uio_out[0] 0.11108f
C2186 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.02778f
C2187 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.26942f
C2188 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07517f
C2189 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.07579f
C2190 a_8345_26455# a_8554_26437# 0.24088f
C2191 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[6] 0.363f
C2192 a_4210_22378# a_3027_22138# 0.0649f
C2193 a_13011_19242# a_13216_19809# 0.01179f
C2194 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.42509f
C2195 a_10762_18823# sar9b_0.net2 0.01126f
C2196 a_8334_18353# sar9b_0.net73 0.02504f
C2197 a_11658_18142# sar9b_0.net39 0.02313f
C2198 a_3561_22527# sar9b_0.net65 0.0125f
C2199 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C2200 a_7306_19777# sar9b_0.net47 0.19638f
C2201 a_11430_27595# sar9b_0.net59 0.17391f
C2202 sar9b_0.net32 sar9b_0._06_ 0.10957f
C2203 a_11008_17491# a_10803_18142# 0.01179f
C2204 a_3695_23038# sar9b_0.clknet_0_CLK 0.01593f
C2205 VDPWR a_9414_23127# 0.27453f
C2206 sar9b_0.net43 a_5298_24499# 0.06128f
C2207 single_9b_cdac_1.cdac_sw_9b_0.S[8] a_25210_17740# 0.22352f
C2208 sar9b_0.net49 sar9b_0.net37 0.07403f
C2209 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.45521f
C2210 single_9b_cdac_1.SW[5] a_13011_17910# 0.02888f
C2211 single_9b_cdac_1.CF[5] clk 0.48018f
C2212 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38702f
C2213 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C2214 a_9162_23174# sar9b_0.net37 0.02849f
C2215 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.84424f
C2216 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02632f
C2217 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.03729f
C2218 a_10803_18142# sar9b_0.net36 0.02932f
C2219 sar9b_0.net55 sar9b_0.net11 0.02067f
C2220 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.11216f
C2221 VDPWR a_13011_16810# 0.4276f
C2222 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.42784f
C2223 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.42509f
C2224 a_8334_17021# sar9b_0.net6 0.03019f
C2225 sar9b_0.net1 a_9414_23127# 0.02489f
C2226 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[8] 4.16545f
C2227 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.7611f
C2228 sar9b_0.net40 sar9b_0.net54 0.09214f
C2229 a_10239_19235# a_10553_18922# 0.07826f
C2230 single_9b_cdac_1.CF[6] a_13011_24570# 0.35426f
C2231 a_8874_19178# a_9472_18823# 0.06623f
C2232 sar9b_0.net57 sar9b_0.net27 0.10308f
C2233 a_6484_22845# sar9b_0.clk_div_0.COUNT\[1\] 0.04883f
C2234 a_3180_19448# sar9b_0._00_ 0.1679f
C2235 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.17533f
C2236 a_9634_17478# a_9974_17626# 0.24088f
C2237 a_8386_22806# a_8591_22855# 0.09983f
C2238 a_8202_23174# a_9162_23174# 0.03529f
C2239 sar9b_0.net63 sar9b_0._12_ 0.07563f
C2240 a_5506_17478# a_5846_17626# 0.24088f
C2241 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[2] 2.01677f
C2242 a_6834_20780# sar9b_0.net40 0.01162f
C2243 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 1.56012f
C2244 a_3540_27045# a_3156_26115# 0.15019f
C2245 a_12531_28566# a_13164_28398# 0.02384f
C2246 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.22497f
C2247 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.22879f
C2248 a_6534_17799# sar9b_0.net56 0.02731f
C2249 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.10626f
C2250 sar9b_0.net52 sar9b_0.net74 0.7241f
C2251 a_7470_22349# sar9b_0.net39 0.03069f
C2252 a_6642_19448# sar9b_0.net35 0.01573f
C2253 a_8052_18123# sar9b_0.net48 0.02566f
C2254 a_10470_21795# sar9b_0.net9 0.03298f
C2255 a_57946_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.23864f
C2256 a_4947_20140# sar9b_0.clknet_1_0__leaf_CLK 0.21937f
C2257 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 3.27803f
C2258 sar9b_0._06_ a_13067_27662# 0.01122f
C2259 a_21368_4076# ua[0] 0.17332f
C2260 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.95338f
C2261 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C2262 sar9b_0.net56 a_8057_18463# 0.01557f
C2263 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.SW[6] 0.14966f
C2264 a_8334_17021# sar9b_0.net46 0.19846f
C2265 sar9b_0.net6 single_9b_cdac_1.SW[2] 0.15073f
C2266 sar9b_0.net43 sar9b_0.net4 0.0207f
C2267 a_10690_22806# sar9b_0.net74 0.04092f
C2268 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.7611f
C2269 VDPWR a_11842_26426# 0.23378f
C2270 sar9b_0.net43 sar9b_0._15_ 0.16183f
C2271 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.CF[2] 0.03547f
C2272 a_5298_24499# sar9b_0._15_ 0.079f
C2273 a_5846_26950# sar9b_0.net37 0.0568f
C2274 a_3014_24136# a_2508_23444# 0.01366f
C2275 sar9b_0.net38 uo_out[4] 0.07167f
C2276 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 a_44418_26990# 0.14695f
C2277 sar9b_0.net53 a_12618_22138# 0.26166f
C2278 a_8334_18353# sar9b_0.net46 0.22365f
C2279 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.38397f
C2280 VDPWR uo_out[4] 0.83671f
C2281 a_2547_28132# uio_out[1] 0.03336f
C2282 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.75853f
C2283 sar9b_0.net40 sar9b_0.net27 0.81488f
C2284 a_6252_20780# sar9b_0._11_ 0.27844f
C2285 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 2.82172f
C2286 a_5711_17527# sar9b_0.net4 0.01409f
C2287 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[8] 0.31534f
C2288 sar9b_0.net9 sar9b_0.net73 0.02088f
C2289 VDPWR a_4698_25851# 0.01249f
C2290 sar9b_0.net63 a_4044_24776# 0.04322f
C2291 a_12182_18427# sar9b_0.net6 0.02363f
C2292 a_8595_17910# sar9b_0.net37 0.04816f
C2293 sar9b_0.net53 a_12870_23599# 0.17313f
C2294 a_7743_18149# sar9b_0.net5 0.0249f
C2295 VDPWR a_10644_16791# 0.84151f
C2296 sar9b_0.net5 single_9b_cdac_1.CF[0] 0.02589f
C2297 sar9b_0.net36 a_10937_25582# 0.02011f
C2298 a_10218_20806# a_11430_20935# 0.07766f
C2299 a_8057_17131# sar9b_0.net5 0.05766f
C2300 sar9b_0.net61 sar9b_0.net73 0.22051f
C2301 sar9b_0.net60 sar9b_0.net36 0.25636f
C2302 a_10482_25831# a_10623_25895# 0.27388f
C2303 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 a_49221_26990# 0.14695f
C2304 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.28813f
C2305 sar9b_0._01_ sar9b_0._10_ 0.03463f
C2306 a_10470_21795# a_9442_21474# 0.07826f
C2307 sar9b_0.net6 single_9b_cdac_1.SW[8] 0.1227f
C2308 VDPWR a_6579_18832# 0.41927f
C2309 a_9258_21842# a_8982_21902# 0.1263f
C2310 a_5846_17626# a_5322_17846# 0.04522f
C2311 a_5711_17527# a_5046_17906# 0.19065f
C2312 dw_12589_1395# th_dif_sw_0.th_sw_1.CKB 0.24188f
C2313 a_11658_26134# a_12870_26263# 0.07766f
C2314 sar9b_0.net46 single_9b_cdac_1.SW[2] 0.02228f
C2315 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.0303f
C2316 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[0] 4.15031f
C2317 sar9b_0.net49 a_10098_19171# 0.02393f
C2318 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[2] 15.0435f
C2319 sar9b_0.net5 a_13011_20574# 0.2669f
C2320 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[0] 0.22444f
C2321 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net39 0.06168f
C2322 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.3196f
C2323 a_7188_22119# a_7402_22441# 0.04522f
C2324 sar9b_0.net42 sar9b_0.net2 0.15479f
C2325 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP ua[0] 1.15122f
C2326 a_12870_18271# sar9b_0.net27 0.02288f
C2327 sar9b_0.net59 a_2847_26141# 0.17414f
C2328 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.03729f
C2329 single_9b_cdac_1.CF[1] sar9b_0.net28 0.04257f
C2330 sar9b_0.net30 clk 0.0304f
C2331 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.84061f
C2332 VDPWR a_3262_24141# 0.01376f
C2333 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C2334 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38733f
C2335 sar9b_0.net54 a_6538_24506# 0.22653f
C2336 VDPWR a_10239_19235# 0.26788f
C2337 a_49221_26990# single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.22497f
C2338 sar9b_0.net61 sar9b_0.net6 0.4224f
C2339 a_12182_18427# sar9b_0.net50 0.14036f
C2340 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN ua[0] 3.10218f
C2341 sar9b_0.net52 a_7638_23474# 0.19487f
C2342 VDPWR a_9634_17478# 0.21868f
C2343 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.07579f
C2344 a_12182_18427# a_12618_18142# 0.16939f
C2345 VDPWR sar9b_0.net14 0.26926f
C2346 sar9b_0.net38 sar9b_0.net11 0.02613f
C2347 sar9b_0.net17 a_2892_27039# 0.01295f
C2348 single_9b_cdac_1.SW[5] clk 0.08628f
C2349 sar9b_0.net7 sar9b_0.net73 1.54797f
C2350 a_3370_26437# a_2706_26108# 0.16939f
C2351 a_3438_26345# a_3156_26115# 0.05462f
C2352 sar9b_0._01_ sar9b_0.net4 0.03109f
C2353 VDPWR sar9b_0.net11 1.08113f
C2354 VDPWR sar9b_0.net66 0.70022f
C2355 sar9b_0.net17 a_2508_27440# 0.01561f
C2356 uio_out[0] uo_out[7] 2.91188f
C2357 uio_out[1] ui_in[0] 1.11045f
C2358 sar9b_0.net50 single_9b_cdac_1.SW[8] 0.1731f
C2359 a_11859_17910# sar9b_0.net2 0.11023f
C2360 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[8] 0.06897f
C2361 a_5046_17906# sar9b_0.net4 0.01394f
C2362 a_5938_22378# sar9b_0.net39 0.0251f
C2363 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.01152f
C2364 single_9b_cdac_1.CF[7] sar9b_0.net28 0.03957f
C2365 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[0] 0.45278f
C2366 sar9b_0.net43 a_5748_24381# 0.02206f
C2367 a_5322_27170# a_5711_26851# 0.05462f
C2368 sar9b_0.net1 sar9b_0.net11 0.03134f
C2369 a_5298_24499# a_5748_24381# 0.03432f
C2370 sar9b_0.net56 sar9b_0.net51 0.81695f
C2371 sar9b_0.net60 a_3922_20239# 0.01343f
C2372 a_10528_20155# sar9b_0.net5 0.02721f
C2373 sar9b_0.net20 a_6250_28502# 0.0646f
C2374 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[7] 2.07035f
C2375 single_9b_cdac_0.SW[6] ua[0] 0.22043f
C2376 sar9b_0.net42 a_10758_24459# 0.01335f
C2377 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.71729f
C2378 sar9b_0.net58 a_5711_26851# 0.21873f
C2379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.SW[4] 0.1516f
C2380 VDPWR a_5010_28495# 0.34506f
C2381 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C2382 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.06503f
C2383 a_8098_23762# a_9126_23599# 0.07826f
C2384 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] 3.10048f
C2385 ua[4] th_dif_sw_0.VCP 3.30291f
C2386 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[3] 0.05125f
C2387 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.01003f
C2388 VDPWR th_dif_sw_0.VCN 1.99513f
C2389 a_6132_23451# a_5748_24381# 0.15019f
C2390 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.03729f
C2391 sar9b_0.net40 sar9b_0.net36 0.14787f
C2392 a_7478_27751# sar9b_0.net60 0.13192f
C2393 sar9b_0.net58 a_4365_25770# 0.01101f
C2394 a_11842_19766# a_12870_19603# 0.07826f
C2395 single_9b_cdac_1.CF[2] single_9b_cdac_1.SW[2] 1.79549f
C2396 sar9b_0.net61 sar9b_0.net46 0.5339f
C2397 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.84425f
C2398 sar9b_0.net61 sar9b_0.net50 0.03896f
C2399 sar9b_0.net10 a_11658_22138# 0.24856f
C2400 a_9802_26815# a_9870_27060# 0.35559f
C2401 single_9b_cdac_1.SW[3] sar9b_0.net61 0.02878f
C2402 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[7] 16.1938f
C2403 th_dif_sw_0.CKB dw_17224_1400# 0.01749f
C2404 sar9b_0.net18 a_3438_27677# 0.04725f
C2405 sar9b_0.net60 a_5151_28559# 0.02736f
C2406 sar9b_0.net52 a_8303_23853# 0.19552f
C2407 a_10742_25087# sar9b_0.net12 0.06525f
C2408 single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.10499f
C2409 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[2\] 0.26122f
C2410 a_12684_20379# sar9b_0.net51 0.25465f
C2411 a_10644_16791# sar9b_0.net48 0.15925f
C2412 sar9b_0.net45 a_9323_27662# 0.10552f
C2413 single_9b_cdac_1.CF[7] single_9b_cdac_1.CF[3] 0.02038f
C2414 sar9b_0.net32 uo_out[2] 0.09101f
C2415 VDPWR a_7338_24802# 0.35888f
C2416 a_13011_17910# sar9b_0.net27 0.03831f
C2417 a_10649_17131# single_9b_cdac_1.SW[0] 0.02173f
C2418 sar9b_0.net49 a_10182_20463# 0.2021f
C2419 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[7] 0.0313f
C2420 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.26427f
C2421 a_3713_22522# a_4011_22488# 0.02614f
C2422 sar9b_0.net41 sar9b_0.net37 0.12296f
C2423 VDPWR a_8098_23762# 0.25671f
C2424 sar9b_0.net43 sar9b_0.net55 0.27955f
C2425 a_10707_23470# sar9b_0.net53 0.05847f
C2426 a_10553_18922# sar9b_0.net26 0.13039f
C2427 a_4934_22432# a_5739_22488# 0.29207f
C2428 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C2429 a_16159_13315# tdc_0.OUTN 0.01845f
C2430 VDPWR a_7443_21496# 0.44805f
C2431 a_3946_26198# sar9b_0.net35 0.17078f
C2432 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.69086f
C2433 a_9472_23805# sar9b_0.net53 0.01787f
C2434 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.07517f
C2435 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.10499f
C2436 sar9b_0.net36 a_9588_27045# 0.07056f
C2437 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.62443f
C2438 sar9b_0.net23 sar9b_0.net34 0.07163f
C2439 a_10607_25185# sar9b_0.net38 0.01125f
C2440 sar9b_0.net38 single_9b_cdac_0.SW[8] 0.02501f
C2441 sar9b_0.net58 a_5674_28147# 0.12675f
C2442 sar9b_0.net65 a_3027_22138# 0.01967f
C2443 VDPWR a_10607_25185# 0.25735f
C2444 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C2445 sar9b_0.net59 sar9b_0.net45 0.55332f
C2446 VDPWR single_9b_cdac_0.SW[8] 2.48304f
C2447 sar9b_0.net7 sar9b_0.net50 0.20371f
C2448 a_8842_16874# a_8057_17131# 0.26257f
C2449 sar9b_0.net7 single_9b_cdac_1.SW[3] 0.03478f
C2450 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 1.55942f
C2451 a_4125_25958# sar9b_0.clknet_1_1__leaf_CLK 0.31513f
C2452 a_3695_23038# sar9b_0.net65 0.11374f
C2453 a_10218_24802# a_11430_24931# 0.07766f
C2454 a_5938_22378# a_6540_22112# 0.01219f
C2455 a_8940_24402# sar9b_0.net2 0.24809f
C2456 single_9b_cdac_1.CF[7] a_13011_24570# 0.03372f
C2457 sar9b_0.net9 single_9b_cdac_1.CF[2] 0.25447f
C2458 a_10239_19235# sar9b_0.net48 0.22117f
C2459 sar9b_0.net34 a_9593_26914# 0.02203f
C2460 VDPWR sar9b_0._00_ 0.73774f
C2461 sar9b_0.net35 tdc_0.OUTN 0.05242f
C2462 a_10995_28566# uo_out[2] 0.42572f
C2463 sar9b_0.net48 a_9634_17478# 0.1085f
C2464 sar9b_0.net2 sar9b_0.net74 0.26355f
C2465 a_10239_19235# a_9900_19047# 0.07649f
C2466 a_17125_9355# a_16331_9671# 0.06748f
C2467 sar9b_0._09_ sar9b_0._07_ 0.58193f
C2468 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.23864f
C2469 m2_23774_26966# VDPWR 0.19016f
C2470 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[6] 0.06019f
C2471 sar9b_0.net43 a_10070_24286# 0.04223f
C2472 single_9b_cdac_0.SW[1] a_13011_27234# 0.35197f
C2473 a_7914_27466# a_8512_27801# 0.06623f
C2474 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.S[3] 16.7662f
C2475 sar9b_0.net52 a_10402_25094# 0.0792f
C2476 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.10499f
C2477 a_2893_24992# sar9b_0._14_ 0.34774f
C2478 sar9b_0.net72 sar9b_0.net68 0.02728f
C2479 a_11436_17742# sar9b_0.net61 0.18223f
C2480 single_9b_cdac_0.SW[2] sar9b_0.net28 0.04952f
C2481 a_7926_23234# sar9b_0.net62 0.21091f
C2482 a_5682_23444# sar9b_0.net11 0.04944f
C2483 a_10218_27466# a_10402_27758# 0.44532f
C2484 VDPWR a_3161_27787# 0.24214f
C2485 a_4922_20857# sar9b_0._11_ 0.07006f
C2486 a_3180_19448# a_3795_19512# 0.02106f
C2487 sar9b_0.net59 a_9870_27060# 0.26796f
C2488 a_10402_21098# a_10607_21189# 0.09983f
C2489 a_3090_27163# a_3540_27045# 0.03432f
C2490 a_6307_27584# a_5460_28377# 0.01439f
C2491 sar9b_0.net66 sar9b_0.clknet_1_0__leaf_CLK 0.08897f
C2492 single_9b_cdac_0.SW[6] a_9323_28371# 0.38985f
C2493 sar9b_0.net59 a_4812_28371# 0.01553f
C2494 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.42509f
C2495 a_5465_28246# a_5742_28392# 0.09983f
C2496 sar9b_0.net55 sar9b_0.net4 0.82102f
C2497 sar9b_0.net10 a_7193_22459# 0.01351f
C2498 sar9b_0.net18 sar9b_0.net59 0.09486f
C2499 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.27554f
C2500 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.42509f
C2501 a_3161_27787# a_3370_27769# 0.24088f
C2502 a_11722_25838# a_10932_25713# 0.1263f
C2503 sar9b_0.net2 a_10506_24506# 0.076f
C2504 sar9b_0.net54 clk 0.11407f
C2505 th_dif_sw_0.th_sw_1.CKB dw_17224_1400# 0.24436f
C2506 a_8031_26141# sar9b_0.cyclic_flag_0.FINAL 0.03467f
C2507 sar9b_0.net5 sar9b_0.net73 1.10057f
C2508 VDPWR a_11658_26134# 0.83989f
C2509 sar9b_0.net23 uo_out[3] 0.10721f
C2510 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.17533f
C2511 sar9b_0._05_ a_4812_21738# 0.01191f
C2512 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C2513 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C2514 a_7638_19238# a_8303_18859# 0.19065f
C2515 sar9b_0.net52 sar9b_0.net53 0.37319f
C2516 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.SW[5] 0.03636f
C2517 a_12618_23470# a_13216_23805# 0.06623f
C2518 sar9b_0.net70 a_3219_22860# 0.03435f
C2519 a_8883_27466# single_9b_cdac_0.SW[8] 0.0266f
C2520 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[3] 0.04427f
C2521 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.22549f
C2522 a_11430_27595# single_9b_cdac_0.SW[5] 0.03357f
C2523 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[0] 0.30922f
C2524 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 3.27795f
C2525 sar9b_0.net41 sar9b_0.net59 0.1373f
C2526 a_10926_17021# a_10644_16791# 0.05462f
C2527 a_4755_22138# sar9b_0._18_ 0.01306f
C2528 sar9b_0.net44 a_5046_27230# 0.06448f
C2529 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 1.71649f
C2530 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.3196f
C2531 a_6783_19481# a_7097_19795# 0.07826f
C2532 a_5812_21028# sar9b_0.net60 0.24213f
C2533 a_62748_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.23864f
C2534 a_8691_28566# uo_out[6] 0.03562f
C2535 sar9b_0.net63 sar9b_0.net58 0.25917f
C2536 sar9b_0.net30 sar9b_0.net45 0.11616f
C2537 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.01152f
C2538 a_10506_24506# a_10758_24459# 0.27388f
C2539 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 3.10626f
C2540 sar9b_0.net26 sar9b_0.net38 0.02477f
C2541 single_9b_cdac_0.SW[7] sar9b_0.net38 0.18897f
C2542 a_11338_19178# sar9b_0.net42 0.02024f
C2543 VDPWR tdc_0.phase_detector_0.pd_out_0.A 1.77491f
C2544 a_21177_7457# th_dif_sw_0.CKB 0.6816f
C2545 sar9b_0.net6 sar9b_0.net5 0.134f
C2546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02519f
C2547 VDPWR sar9b_0.net26 0.97073f
C2548 VDPWR a_5739_22488# 0.09539f
C2549 a_10690_22806# sar9b_0.net53 0.11211f
C2550 a_3369_24181# a_2835_24136# 0.35097f
C2551 VDPWR single_9b_cdac_0.SW[7] 2.68913f
C2552 a_10690_22806# a_10895_22855# 0.09983f
C2553 a_10506_23174# a_11466_23174# 0.03471f
C2554 sar9b_0.net63 a_6137_23791# 0.04828f
C2555 a_12182_26419# a_12618_26134# 0.16939f
C2556 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[5] 8.69008f
C2557 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[7] 0.06019f
C2558 a_10230_23234# clk 0.01685f
C2559 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.12077f
C2560 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C2561 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[2] 0.3633f
C2562 a_9942_27470# a_10607_27849# 0.19065f
C2563 single_9b_cdac_1.cdac_sw_9b_0.S[5] ua[0] 1.57219f
C2564 ui_in[0] clk 0.23226f
C2565 a_4922_20857# sar9b_0.net65 0.08585f
C2566 sar9b_0.net26 sar9b_0.net1 0.04547f
C2567 sar9b_0.net27 clk 0.04404f
C2568 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.3196f
C2569 a_6636_20780# a_6834_20780# 0.06623f
C2570 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 ua[0] 0.14027f
C2571 sar9b_0.net43 sar9b_0.net38 0.17602f
C2572 single_9b_cdac_0.SW[3] th_dif_sw_0.VCN 0.09453f
C2573 VDPWR a_13011_20806# 0.49978f
C2574 single_9b_cdac_0.SW[5] clk 0.153f
C2575 a_3206_22432# a_3561_22527# 0.18757f
C2576 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[0\] 0.03041f
C2577 sar9b_0.net12 a_10937_25582# 0.02312f
C2578 sar9b_0.net43 VDPWR 3.08648f
C2579 a_9162_23174# sar9b_0.net54 0.27476f
C2580 sar9b_0.net42 a_10742_25087# 0.02075f
C2581 VDPWR a_5298_24499# 0.32802f
C2582 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[5] 4.15421f
C2583 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02552f
C2584 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.12898f
C2585 a_8940_27039# a_9138_27163# 0.06623f
C2586 VDPWR a_10035_19474# 0.46118f
C2587 sar9b_0.net17 a_2706_26108# 0.01317f
C2588 tdc_0.OUTP single_9b_cdac_1.SW[2] 0.36499f
C2589 a_2893_24992# sar9b_0._16_ 0.18199f
C2590 sar9b_0.net56 a_9359_20191# 0.01326f
C2591 sar9b_0.net40 sar9b_0.net51 0.02551f
C2592 sar9b_0.net58 a_3231_27227# 0.17354f
C2593 VDPWR a_9126_19131# 0.28669f
C2594 a_11658_18142# a_12182_18427# 0.05022f
C2595 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._00_ 0.1706f
C2596 VDPWR a_6132_23451# 0.78916f
C2597 VDPWR a_5711_17527# 0.25721f
C2598 a_8874_19178# sar9b_0.net37 0.03852f
C2599 VDPWR a_8340_26115# 0.87266f
C2600 sar9b_0.net58 a_2706_27440# 0.26179f
C2601 VDPWR a_7882_19538# 0.30688f
C2602 a_6767_25185# a_6102_24806# 0.19065f
C2603 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.07579f
C2604 sar9b_0.net35 sar9b_0.net39 0.0534f
C2605 VDPWR sar9b_0._10_ 0.48054f
C2606 sar9b_0.net46 sar9b_0.net5 1.36216f
C2607 VDPWR a_13011_23238# 0.48316f
C2608 sar9b_0.net55 a_5748_24381# 0.0128f
C2609 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[0\] 0.01565f
C2610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.0303f
C2611 sar9b_0.net50 sar9b_0.net5 0.49397f
C2612 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.76578f
C2613 sar9b_0.net57 sar9b_0.net12 0.27108f
C2614 a_2835_24136# a_3014_24136# 0.54426f
C2615 sar9b_0.net23 a_8031_26141# 0.02315f
C2616 a_44418_17740# single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.22513f
C2617 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[0] 0.74373f
C2618 sar9b_0.net2 sar9b_0.net39 0.23235f
C2619 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.02638f
C2620 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.42509f
C2621 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.01427f
C2622 a_9996_16784# a_10194_16784# 0.06623f
C2623 sar9b_0._02_ a_6444_21738# 0.25486f
C2624 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.06503f
C2625 VDPWR a_7404_16784# 0.19127f
C2626 single_9b_cdac_1.SW[4] sar9b_0.net6 0.02588f
C2627 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.81428f
C2628 a_9546_24506# a_10227_23490# 0.02456f
C2629 sar9b_0.net5 a_9154_20142# 0.01312f
C2630 th_dif_sw_0.CK sar9b_0.net38 0.21539f
C2631 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.83441f
C2632 VDPWR a_4125_25958# 0.4305f
C2633 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.1507f
C2634 a_11030_22954# sar9b_0.net42 0.0141f
C2635 VDPWR a_11382_22142# 0.28804f
C2636 sar9b_0.net13 a_10218_24802# 0.02005f
C2637 VDPWR th_dif_sw_0.CK 1.56597f
C2638 single_9b_cdac_0.SW[8] single_9b_cdac_0.SW[3] 0.026f
C2639 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.01175f
C2640 th_dif_sw_0.CKB tdc_0.OUTN 2.99096f
C2641 VDPWR sar9b_0.net3 0.45768f
C2642 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.02632f
C2643 sar9b_0.net24 single_9b_cdac_0.SW[7] 0.05134f
C2644 a_11658_18142# sar9b_0.net61 0.01086f
C2645 a_2918_20140# a_3166_20145# 0.05308f
C2646 a_2739_20140# a_3425_20244# 0.27693f
C2647 sar9b_0.net66 sar9b_0._12_ 0.16928f
C2648 sar9b_0.net52 a_10932_25713# 0.17701f
C2649 sar9b_0.net31 a_11842_22430# 0.01313f
C2650 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.17533f
C2651 VDPWR sar9b_0.net4 1.04258f
C2652 a_5441_22522# a_5739_22488# 0.02614f
C2653 a_11776_27801# sar9b_0.net25 0.26874f
C2654 VDPWR sar9b_0._15_ 0.37538f
C2655 single_9b_cdac_1.SW[2] single_9b_cdac_1.SW[7] 0.2192f
C2656 sar9b_0.net56 a_4771_18260# 0.23559f
C2657 VDPWR a_2892_23070# 0.30728f
C2658 a_11658_23470# a_12618_23470# 0.03432f
C2659 sar9b_0.net43 sar9b_0.net24 0.02255f
C2660 a_21177_7457# th_dif_sw_0.th_sw_1.CKB 2.27999f
C2661 a_8691_28566# uo_out[4] 0.37881f
C2662 sar9b_0.net67 a_4236_21738# 0.14162f
C2663 sar9b_0.net20 uio_out[0] 0.01201f
C2664 sar9b_0.net1 sar9b_0.net4 0.01778f
C2665 tdc_0.OUTP sar9b_0.net61 0.10662f
C2666 VDPWR sar9b_0._01_ 0.28816f
C2667 sar9b_0.net29 a_13011_20806# 0.01682f
C2668 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02784f
C2669 sar9b_0.net26 sar9b_0.net48 0.4034f
C2670 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.01003f
C2671 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.95338f
C2672 a_7289_21127# sar9b_0.net10 0.01176f
C2673 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP a_33936_26999# 0.04592f
C2674 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.05472f
C2675 VDPWR a_12182_19759# 0.20727f
C2676 VDPWR a_5046_17906# 0.28567f
C2677 a_8842_18206# sar9b_0.net73 0.04312f
C2678 a_9900_19047# sar9b_0.net26 0.04584f
C2679 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[3] 12.6046f
C2680 sar9b_0.net36 clk 0.03715f
C2681 single_9b_cdac_1.cdac_sw_9b_0.S[1] ua[0] 1.19426f
C2682 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C2683 sar9b_0.net59 uo_out[7] 0.02838f
C2684 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C2685 a_7638_23474# a_7914_23470# 0.1263f
C2686 sar9b_0.net28 single_9b_cdac_1.SW[8] 0.04546f
C2687 single_9b_cdac_1.CF[4] clk 0.14003f
C2688 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.45521f
C2689 a_11339_27039# single_9b_cdac_0.SW[4] 0.03465f
C2690 a_4922_20857# a_5581_20992# 0.01403f
C2691 sar9b_0._07_ a_5126_20140# 0.02529f
C2692 single_9b_cdac_1.CF[3] single_9b_cdac_1.SW[2] 0.01297f
C2693 a_17125_9355# clk 0.02939f
C2694 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.02784f
C2695 sar9b_0.net7 a_11658_18142# 0.21927f
C2696 a_13011_23238# sar9b_0.net29 0.02021f
C2697 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.03729f
C2698 a_3372_25734# sar9b_0._16_ 0.26724f
C2699 a_10035_19474# sar9b_0.net48 0.35551f
C2700 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 1.71649f
C2701 sar9b_0.net31 sar9b_0.net30 0.08627f
C2702 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[7] 3.98346f
C2703 a_8842_16874# sar9b_0.net6 0.05357f
C2704 a_6484_22845# sar9b_0.clk_div_0.COUNT\[2\] 0.0424f
C2705 a_9126_19131# sar9b_0.net48 0.21244f
C2706 sar9b_0._08_ sar9b_0._10_ 0.25501f
C2707 a_10548_19053# a_10830_19068# 0.06034f
C2708 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.95338f
C2709 a_7692_26108# sar9b_0.net59 0.04276f
C2710 a_4755_22138# sar9b_0.net64 0.07292f
C2711 single_9b_cdac_1.cdac_sw_9b_0.S[2] a_54032_17740# 0.22367f
C2712 sar9b_0.net33 a_11842_26426# 0.13675f
C2713 sar9b_0._02_ sar9b_0.clk_div_0.COUNT\[1\] 0.01796f
C2714 VDPWR a_6126_18353# 0.26525f
C2715 sar9b_0.net43 a_9270_24566# 0.05226f
C2716 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.07517f
C2717 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] 1.15122f
C2718 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 3.10626f
C2719 a_8591_22855# a_8726_22954# 0.35559f
C2720 sar9b_0.net13 a_6378_24802# 0.08313f
C2721 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C2722 a_5484_23444# a_5823_23477# 0.07649f
C2723 a_6132_23451# a_5682_23444# 0.03529f
C2724 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26427f
C2725 VDPWR a_3795_19512# 0.60141f
C2726 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[5] 0.12898f
C2727 a_13164_28398# sar9b_0._06_ 0.28405f
C2728 VDPWR a_3180_19448# 0.26779f
C2729 a_11915_27039# a_11658_26134# 0.04032f
C2730 a_7978_22202# sar9b_0.net39 0.04787f
C2731 sar9b_0.net10 sar9b_0.net37 0.02841f
C2732 a_7097_19795# sar9b_0.net35 0.01811f
C2733 w_17430_1606# ua[3] 0.88896f
C2734 VDPWR a_4236_21738# 0.23821f
C2735 sar9b_0._17_ sar9b_0.net4 0.77945f
C2736 sar9b_0._10_ sar9b_0.clknet_1_0__leaf_CLK 0.20402f
C2737 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[3] 0.026f
C2738 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP a_43540_26999# 0.04592f
C2739 a_8019_17910# sar9b_0.net46 0.05518f
C2740 single_9b_cdac_1.SW[1] sar9b_0.net73 0.05555f
C2741 a_9996_16784# sar9b_0.net27 0.02177f
C2742 a_8303_23853# a_7914_23470# 0.06034f
C2743 th_dif_sw_0.CK sar9b_0.net48 0.03264f
C2744 sar9b_0.net49 sar9b_0.net36 0.04379f
C2745 sar9b_0.net42 a_10937_25582# 0.02311f
C2746 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.02149f
C2747 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 1.55982f
C2748 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.01402f
C2749 sar9b_0.net2 sar9b_0.net53 0.39622f
C2750 a_8842_16874# sar9b_0.net46 0.19416f
C2751 sar9b_0._01_ sar9b_0._17_ 0.03752f
C2752 a_10895_22855# sar9b_0.net2 0.01734f
C2753 dw_12589_1395# a_10166_3438# 26.7601f
C2754 tdc_0.OUTN single_9b_cdac_1.SW[0] 0.44367f
C2755 VDPWR a_5748_24381# 0.75977f
C2756 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCP 1.0224f
C2757 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[0] 0.22459f
C2758 a_11146_25483# sar9b_0.net42 0.01506f
C2759 a_6642_19448# sar9b_0.net40 0.06124f
C2760 a_11030_22954# sar9b_0.net74 0.01098f
C2761 VDPWR a_12870_26263# 0.2717f
C2762 VDPWR a_6282_27170# 0.35695f
C2763 a_9942_27470# sar9b_0.net23 0.02292f
C2764 sar9b_0.net58 uo_out[6] 0.11715f
C2765 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.02778f
C2766 sar9b_0.net48 sar9b_0.net4 0.02286f
C2767 a_6880_17491# sar9b_0.net5 0.27459f
C2768 a_8052_18123# a_7743_18149# 0.07766f
C2769 sar9b_0.net53 a_12047_22521# 0.22562f
C2770 a_8842_18206# sar9b_0.net46 0.221f
C2771 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C2772 a_7404_16784# a_7602_16784# 0.06623f
C2773 sar9b_0._08_ sar9b_0._01_ 0.05213f
C2774 sar9b_0.net50 a_12618_19474# 0.26154f
C2775 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C2776 sar9b_0.net35 a_6562_25094# 0.02907f
C2777 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.CF[8] 0.19143f
C2778 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07517f
C2779 a_10218_27466# a_9588_27045# 0.01007f
C2780 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.01472f
C2781 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 2.7611f
C2782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C2783 VDPWR sar9b_0.clknet_1_1__leaf_CLK 3.19348f
C2784 a_62748_16877# single_9b_cdac_1.SW[0] 0.28324f
C2785 sar9b_0.net45 single_9b_cdac_0.SW[5] 0.0907f
C2786 a_2603_17006# th_dif_sw_0.CKB 0.35268f
C2787 sar9b_0.net57 a_8386_22806# 0.03019f
C2788 sar9b_0.net41 a_10410_17846# 0.06272f
C2789 single_9b_cdac_1.SW[1] sar9b_0.net6 0.04631f
C2790 sar9b_0.net40 a_13216_18477# 0.01664f
C2791 a_10402_21098# a_11430_20935# 0.07826f
C2792 a_11382_23474# a_11658_23470# 0.1263f
C2793 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[1\] 0.89565f
C2794 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP ua[0] 1.15133f
C2795 a_10482_25831# a_10937_25582# 0.3578f
C2796 a_10623_25895# a_10932_25713# 0.07766f
C2797 sar9b_0.net53 a_10758_24459# 0.16837f
C2798 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP ua[0] 1.15113f
C2799 a_10506_23174# sar9b_0.net11 0.06113f
C2800 a_7590_24931# sar9b_0.net54 0.20557f
C2801 sar9b_0.net7 a_9258_21842# 0.01005f
C2802 sar9b_0.net41 sar9b_0.net54 0.04048f
C2803 a_9258_21842# a_9442_21474# 0.44098f
C2804 a_11146_25483# a_10482_25831# 0.16939f
C2805 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.95338f
C2806 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.24288f
C2807 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C2808 VDPWR sar9b_0.net55 0.724f
C2809 sar9b_0.net47 sar9b_0.net10 1.99512f
C2810 sar9b_0.net57 a_4771_18260# 0.29258f
C2811 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.12431f
C2812 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.36041f
C2813 a_12182_19759# a_12047_19857# 0.35559f
C2814 a_12870_19603# a_13216_19809# 0.07649f
C2815 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.38397f
C2816 a_3206_22432# a_3027_22138# 0.54361f
C2817 sar9b_0.net48 a_6126_18353# 0.22812f
C2818 a_10553_18922# sar9b_0.net38 0.02338f
C2819 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.28813f
C2820 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.22875f
C2821 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.75853f
C2822 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.42784f
C2823 VDPWR a_10553_18922# 0.21937f
C2824 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.0303f
C2825 single_9b_cdac_1.CF[8] clk 0.12991f
C2826 VDPWR a_4934_22432# 0.89137f
C2827 single_9b_cdac_0.SW[2] a_13011_27234# 0.04188f
C2828 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 1.71649f
C2829 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.3196f
C2830 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.04988f
C2831 VDPWR a_9974_17626# 0.19746f
C2832 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96841f
C2833 sar9b_0.net40 sar9b_0.net42 0.0514f
C2834 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.26709f
C2835 a_5739_22488# sar9b_0._12_ 0.0684f
C2836 sar9b_0.net32 single_9b_cdac_0.SW[6] 0.05164f
C2837 a_12870_18271# a_13216_18477# 0.07649f
C2838 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[1] 0.26555f
C2839 a_12182_18427# a_12047_18525# 0.35559f
C2840 a_5931_20140# a_6130_20239# 0.29821f
C2841 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.11216f
C2842 a_3946_26198# a_3156_26115# 0.1263f
C2843 dw_12589_1395# a_10254_2858# 1.98316f
C2844 a_7890_26108# a_7692_26108# 0.06623f
C2845 sar9b_0.net38 a_10070_24286# 0.01531f
C2846 sar9b_0.net17 a_2706_27440# 0.02173f
C2847 a_9996_16784# sar9b_0.net36 0.27514f
C2848 VDPWR a_10070_24286# 0.20147f
C2849 a_7188_22119# sar9b_0.net39 0.05015f
C2850 sar9b_0.net9 a_10690_22806# 0.03973f
C2851 sar9b_0.net60 sar9b_0.clknet_0_CLK 0.01871f
C2852 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.22875f
C2853 sar9b_0.net43 a_6030_24396# 0.04681f
C2854 a_5046_27230# a_5711_26851# 0.19065f
C2855 sar9b_0.net60 sar9b_0.net16 0.01459f
C2856 sar9b_0.net41 sar9b_0.net27 0.03867f
C2857 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.24495f
C2858 a_16159_13315# a_16185_13034# 0.19021f
C2859 a_8438_23755# a_8874_23470# 0.16939f
C2860 VDPWR a_10742_21091# 0.20336f
C2861 sar9b_0.net74 a_10937_25582# 0.05953f
C2862 a_6286_22804# sar9b_0._02_ 0.01706f
C2863 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C2864 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.SW[4] 0.1498f
C2865 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C2866 a_7926_23234# sar9b_0.net11 0.05391f
C2867 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.84425f
C2868 a_7914_27466# sar9b_0.net60 0.24386f
C2869 sar9b_0.net57 a_6414_23681# 0.05577f
C2870 a_21368_4076# dw_17224_1400# 26.7601f
C2871 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.55985f
C2872 single_9b_cdac_0.SW[6] a_10995_28566# 0.01025f
C2873 a_11146_25483# sar9b_0.net74 0.0492f
C2874 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.42784f
C2875 sar9b_0.net36 sar9b_0.net45 0.56715f
C2876 sar9b_0.net10 a_11842_22430# 0.03989f
C2877 a_10378_27170# a_9593_26914# 0.26257f
C2878 sar9b_0.net57 sar9b_0.clknet_0_CLK 0.03539f
C2879 VDPWR sar9b_0.net67 0.30253f
C2880 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.6919f
C2881 a_13011_24802# sar9b_0.net27 0.04101f
C2882 sar9b_0.net55 sar9b_0._17_ 0.77591f
C2883 sar9b_0.net60 a_5465_28246# 0.02116f
C2884 sar9b_0.net57 sar9b_0.net16 0.01547f
C2885 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C2886 a_11178_24802# sar9b_0.net12 0.08132f
C2887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN ua[0] 3.14416f
C2888 a_26951_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C2889 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.07517f
C2890 a_11658_19474# a_11859_20574# 0.03761f
C2891 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[5] 18.8692f
C2892 VDPWR a_9165_24988# 0.44778f
C2893 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A a_35519_15495# 0.01076f
C2894 uo_out[0] uio_in[7] 0.03102f
C2895 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[2] 0.22161f
C2896 sar9b_0.clknet_1_0__leaf_CLK sar9b_0.clknet_1_1__leaf_CLK 0.01438f
C2897 a_4210_22378# a_4011_22488# 0.29821f
C2898 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C2899 VDPWR a_9126_23599# 0.28311f
C2900 a_11658_23470# sar9b_0.net53 0.18176f
C2901 a_4011_22488# sar9b_0.clknet_0_CLK 0.01809f
C2902 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 ua[0] 0.15943f
C2903 a_8266_17113# a_8334_17021# 0.35559f
C2904 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[3] 0.06971f
C2905 tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTN 0.19342f
C2906 a_4755_22138# sar9b_0._07_ 0.01014f
C2907 sar9b_0._18_ a_4812_21738# 0.01257f
C2908 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.12358f
C2909 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A 0.38397f
C2910 a_13011_17910# a_13216_18477# 0.01179f
C2911 uo_out[4] uo_out[3] 2.93276f
C2912 a_2540_22432# sar9b_0._04_ 0.0164f
C2913 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.81428f
C2914 a_3819_24136# sar9b_0.clk_div_0.COUNT\[2\] 0.01683f
C2915 a_4934_22432# a_5441_22522# 0.21226f
C2916 sar9b_0.net36 a_9870_27060# 0.04885f
C2917 sar9b_0._13_ sar9b_0.net72 0.1941f
C2918 sar9b_0.net31 sar9b_0.net27 0.03712f
C2919 sar9b_0._12_ sar9b_0.net4 0.24818f
C2920 sar9b_0.net4 a_6030_24396# 0.01963f
C2921 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 3.27824f
C2922 a_10662_17799# a_10410_17846# 0.27388f
C2923 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C2924 sar9b_0.net31 single_9b_cdac_0.SW[5] 0.01126f
C2925 sar9b_0.net30 sar9b_0.net10 0.07137f
C2926 sar9b_0.net40 a_6414_23681# 0.0209f
C2927 single_9b_cdac_1.cdac_sw_9b_0.S[3] th_dif_sw_0.VCP 27.3302f
C2928 a_10402_25094# a_10742_25087# 0.24088f
C2929 sar9b_0._18_ a_4332_23043# 0.03742f
C2930 VDPWR a_8694_20570# 0.32519f
C2931 sar9b_0.net49 sar9b_0.net51 0.50265f
C2932 a_10553_18922# sar9b_0.net48 0.08167f
C2933 a_16159_13315# a_16185_12837# 0.01114f
C2934 w_17430_1606# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.3776f
C2935 a_8970_20510# sar9b_0.net37 0.02159f
C2936 sar9b_0.net48 a_9974_17626# 0.13813f
C2937 sar9b_0.clk_div_0.COUNT\[0\] clk 0.21954f
C2938 a_8266_18445# a_8334_18353# 0.35559f
C2939 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.SW[3] 0.14997f
C2940 VDPWR sar9b_0.net38 3.13581f
C2941 a_10548_19053# a_10098_19171# 0.03432f
C2942 sar9b_0.net33 a_11658_26134# 0.07465f
C2943 a_14897_9355# th_dif_sw_0.VCN 0.05461f
C2944 a_6126_18353# a_6634_18206# 0.19065f
C2945 single_9b_cdac_0.SW[2] sar9b_0._06_ 0.01711f
C2946 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C2947 sar9b_0.net41 a_11008_17491# 0.03875f
C2948 a_39616_17740# single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.22512f
C2949 VDPWR a_4330_27170# 0.29064f
C2950 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[0] 0.23282f
C2951 sar9b_0.net68 a_2940_25096# 0.01396f
C2952 sar9b_0.net52 a_11430_24931# 0.16913f
C2953 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.27794f
C2954 sar9b_0.net1 sar9b_0.net38 0.03587f
C2955 a_6137_23791# sar9b_0.net11 0.11829f
C2956 sar9b_0.net41 sar9b_0.net36 0.03019f
C2957 a_12560_27128# sar9b_0.net45 0.20749f
C2958 sar9b_0.net35 single_9b_cdac_1.SW[2] 0.05528f
C2959 a_3795_19512# a_3991_19768# 0.0388f
C2960 a_10218_27466# a_11430_27595# 0.07766f
C2961 a_3540_27045# a_3754_26815# 0.05022f
C2962 VDPWR sar9b_0.net1 1.19391f
C2963 a_7478_27751# sar9b_0.net45 0.02536f
C2964 VDPWR a_3370_27769# 0.20008f
C2965 a_13011_19242# sar9b_0.net27 0.02433f
C2966 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.S[1] 16.8012f
C2967 sar9b_0.net71 a_4072_19474# 0.10694f
C2968 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C2969 a_8052_18123# sar9b_0.net73 0.05137f
C2970 sar9b_0.net72 sar9b_0.net69 0.04519f
C2971 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 2.71729f
C2972 a_5010_28495# sar9b_0.net58 0.2625f
C2973 sar9b_0.net43 a_11178_20806# 0.01951f
C2974 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C2975 sar9b_0.net59 sar9b_0.net20 0.0752f
C2976 a_3747_25724# sar9b_0.clk_div_0.COUNT\[1\] 0.11932f
C2977 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.05472f
C2978 th_dif_sw_0.CKB th_dif_sw_0.VCP 0.21902f
C2979 a_5460_28377# a_5674_28147# 0.05022f
C2980 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.05472f
C2981 a_11722_25838# a_11214_25728# 0.19065f
C2982 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[0] 0.22459f
C2983 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07517f
C2984 single_9b_cdac_0.SW[7] sar9b_0.net33 0.01742f
C2985 sar9b_0.net13 a_11722_25838# 0.05888f
C2986 tdc_0.OUTN a_16555_12412# 0.01287f
C2987 a_6444_19448# sar9b_0.net15 0.01357f
C2988 a_12435_24802# sar9b_0.net27 0.01432f
C2989 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C2990 sar9b_0.net60 a_7343_27849# 0.20041f
C2991 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[7] 0.05361f
C2992 sar9b_0.net60 a_5962_24151# 0.02401f
C2993 uo_out[7] ui_in[0] 0.06786f
C2994 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.42014f
C2995 a_8098_18810# a_8303_18859# 0.09983f
C2996 sar9b_0.net57 a_7638_23474# 0.06419f
C2997 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.3186f
C2998 sar9b_0.net60 sar9b_0.net21 0.08339f
C2999 sar9b_0.net34 single_9b_cdac_0.SW[8] 0.01408f
C3000 sar9b_0.net19 sar9b_0.net37 0.21509f
C3001 a_11776_27801# single_9b_cdac_0.SW[5] 0.01854f
C3002 sar9b_0.net27 a_12435_20806# 0.01148f
C3003 sar9b_0.net67 sar9b_0.clknet_1_0__leaf_CLK 0.18709f
C3004 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.42014f
C3005 a_11434_16874# a_10644_16791# 0.1263f
C3006 sar9b_0.net64 sar9b_0._18_ 0.2077f
C3007 ua[3] dw_17224_1400# 1.4136f
C3008 single_9b_cdac_1.CF[0] th_dif_sw_0.VCN 0.09453f
C3009 a_6642_19448# a_7306_19777# 0.16939f
C3010 sar9b_0.net60 sar9b_0.net39 0.1395f
C3011 a_11842_23762# sar9b_0.net11 0.05371f
C3012 sar9b_0.net54 a_6102_24806# 0.21862f
C3013 sar9b_0._11_ sar9b_0.net60 0.60917f
C3014 a_3695_23038# a_3725_23194# 0.0101f
C3015 a_8074_20870# sar9b_0.net56 0.0467f
C3016 a_4812_28371# a_5151_28559# 0.07649f
C3017 a_5748_24381# a_6030_24396# 0.06034f
C3018 a_10758_24459# a_11104_24151# 0.07649f
C3019 sar9b_0.net24 sar9b_0.net38 0.18f
C3020 VDPWR a_8883_27466# 0.46906f
C3021 sar9b_0.net24 VDPWR 0.56782f
C3022 VDPWR sar9b_0._17_ 1.32705f
C3023 VDPWR a_6738_22112# 0.36714f
C3024 a_11030_22954# sar9b_0.net53 0.14085f
C3025 a_3819_24136# a_2835_24136# 0.08669f
C3026 a_3369_24181# sar9b_0.net70 0.01723f
C3027 a_29134_16877# single_9b_cdac_1.SW[7] 0.28324f
C3028 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.22875f
C3029 a_10895_22855# a_11030_22954# 0.35559f
C3030 sar9b_0.net63 a_6346_23773# 0.03952f
C3031 a_12870_26263# a_13216_26469# 0.07649f
C3032 a_12182_26419# a_12047_26517# 0.35559f
C3033 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36037f
C3034 a_33936_26999# single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.59531f
C3035 a_8266_17113# sar9b_0.net61 0.04067f
C3036 sar9b_0.net9 sar9b_0.net2 0.0459f
C3037 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.26942f
C3038 VDPWR a_5441_22522# 0.10419f
C3039 sar9b_0.net35 a_6922_23534# 0.02301f
C3040 sar9b_0.net35 sar9b_0.net61 0.03955f
C3041 VDPWR sar9b_0.net29 1.26137f
C3042 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C3043 sar9b_0.net35 sar9b_0.net44 0.01492f
C3044 sar9b_0.net57 sar9b_0.net39 0.68049f
C3045 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3046 sar9b_0._11_ sar9b_0.net57 0.0163f
C3047 sar9b_0.net32 sar9b_0.net45 0.02882f
C3048 a_11859_21906# sar9b_0.net26 0.01146f
C3049 a_7284_20787# a_6975_20813# 0.07766f
C3050 sar9b_0.net51 a_6252_19074# 0.05727f
C3051 sar9b_0.net2 sar9b_0.net61 0.18227f
C3052 VDPWR sar9b_0._08_ 0.41847f
C3053 a_3206_22432# a_3454_22567# 0.05308f
C3054 sar9b_0._12_ sar9b_0.clknet_1_1__leaf_CLK 0.30353f
C3055 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.SW[0] 0.22983f
C3056 a_8266_18445# sar9b_0.net61 0.01651f
C3057 sar9b_0.net42 a_11178_24802# 0.01588f
C3058 a_6867_16810# sar9b_0.net27 0.04386f
C3059 sar9b_0.net48 sar9b_0.net38 0.55083f
C3060 sar9b_0.net8 sar9b_0.net26 0.0267f
C3061 a_8052_18123# sar9b_0.net46 0.16885f
C3062 a_9138_27163# a_9279_27227# 0.27388f
C3063 VDPWR a_4083_28566# 0.47299f
C3064 a_8982_21902# sar9b_0.net57 0.05351f
C3065 VDPWR sar9b_0.net48 5.69977f
C3066 sar9b_0.net57 a_8303_23853# 0.04177f
C3067 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP a_29134_16877# 0.04592f
C3068 tdc_0.OUTP a_16555_12124# 0.01017f
C3069 a_18214_3039# w_17430_1606# 0.14276f
C3070 VDPWR a_9900_19047# 0.20374f
C3071 a_11842_18434# a_12182_18427# 0.24088f
C3072 single_9b_cdac_0.SW[4] th_dif_sw_0.VCN 0.09453f
C3073 VDPWR a_5682_23444# 0.35048f
C3074 a_9472_18823# sar9b_0.net37 0.03442f
C3075 sar9b_0.net57 a_5374_20145# 0.01527f
C3076 sar9b_0.net58 a_3161_27787# 0.10647f
C3077 a_7347_24160# sar9b_0.net62 0.09083f
C3078 a_3922_20239# a_2918_20140# 0.06302f
C3079 tdc_0.phase_detector_0.pd_out_0.B a_15400_11316# 0.48689f
C3080 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.45521f
C3081 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C3082 sar9b_0.net8 a_13011_20806# 0.22594f
C3083 sar9b_0.net1 sar9b_0.net48 0.20331f
C3084 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.02624f
C3085 sar9b_0.net43 sar9b_0.net8 0.04888f
C3086 VDPWR sar9b_0.clknet_1_0__leaf_CLK 2.99385f
C3087 VDPWR a_3161_26455# 0.25277f
C3088 single_9b_cdac_0.SW[8] uo_out[3] 0.28955f
C3089 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.19129f
C3090 sar9b_0.net25 uo_out[0] 0.27942f
C3091 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[7] 1.56115f
C3092 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.VCP 0.31462f
C3093 VDPWR a_9270_24566# 0.29709f
C3094 a_3014_24136# sar9b_0.net70 0.26822f
C3095 a_11382_26138# a_11842_26426# 0.26257f
C3096 a_7498_21109# a_7284_20787# 0.04522f
C3097 VDPWR a_12047_19857# 0.26705f
C3098 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36555_15501# 0.01076f
C3099 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.05472f
C3100 sar9b_0.net10 sar9b_0.net54 0.15482f
C3101 a_10644_16791# a_10335_16817# 0.07766f
C3102 sar9b_0.net40 sar9b_0.net21 0.06941f
C3103 a_10662_17799# a_11008_17491# 0.07649f
C3104 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C3105 tdc_0.OUTP single_9b_cdac_1.SW[1] 0.10358f
C3106 VDPWR a_7602_16784# 0.3319f
C3107 VDPWR a_6954_27466# 0.83781f
C3108 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C3109 sar9b_0.net5 a_9494_20290# 0.0262f
C3110 sar9b_0.net40 sar9b_0.net39 0.04664f
C3111 a_6562_25094# a_6902_25087# 0.24088f
C3112 sar9b_0.net7 sar9b_0.net2 0.26633f
C3113 a_4934_22432# sar9b_0._12_ 0.06662f
C3114 a_6834_20780# sar9b_0.net10 0.0738f
C3115 a_10662_17799# sar9b_0.net36 0.03369f
C3116 sar9b_0.net27 a_5322_17846# 0.0316f
C3117 sar9b_0.net36 uo_out[7] 0.10138f
C3118 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[6] 0.01887f
C3119 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.26707f
C3120 sar9b_0.net42 clk 0.03904f
C3121 sar9b_0.net59 sar9b_0.net19 0.15362f
C3122 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.3196f
C3123 a_2918_20140# a_3273_20185# 0.18752f
C3124 a_8386_22806# clk 0.03185f
C3125 sar9b_0.net52 a_11214_25728# 0.27195f
C3126 sar9b_0.net31 a_12870_22267# 0.03044f
C3127 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.28523f
C3128 single_9b_cdac_0.SW[4] single_9b_cdac_0.SW[8] 0.03894f
C3129 a_10254_2858# w_12795_1601# 0.14391f
C3130 sar9b_0.net13 sar9b_0.net52 1.35209f
C3131 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[7] 4.16011f
C3132 sar9b_0.net57 a_10402_25094# 0.01621f
C3133 VDPWR single_9b_cdac_0.SW[3] 2.47465f
C3134 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.69086f
C3135 sar9b_0._08_ sar9b_0._17_ 0.25385f
C3136 sar9b_0.net43 sar9b_0.net34 0.26137f
C3137 a_11658_23470# a_12047_23853# 0.06034f
C3138 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[3] 0.02149f
C3139 single_9b_cdac_1.CF[8] a_13011_24802# 0.02059f
C3140 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.02624f
C3141 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.SW[3] 0.17268f
C3142 single_9b_cdac_1.SW[1] a_57946_16877# 0.28324f
C3143 a_13011_16810# single_9b_cdac_1.SW[3] 0.03223f
C3144 sar9b_0.net49 a_9359_20191# 0.18621f
C3145 a_8554_26437# a_8622_26345# 0.35559f
C3146 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.62443f
C3147 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.02618f
C3148 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 a_44418_17740# 0.14695f
C3149 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.17533f
C3150 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.03543f
C3151 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.38037f
C3152 sar9b_0.net9 a_7978_22202# 0.04916f
C3153 clk single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.02119f
C3154 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.81428f
C3155 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.CF[0] 0.10499f
C3156 VDPWR a_11915_27039# 0.44729f
C3157 sar9b_0.net10 sar9b_0.net27 0.03534f
C3158 a_4011_22488# sar9b_0.net65 0.01096f
C3159 sar9b_0.net41 sar9b_0.net51 0.02663f
C3160 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.11216f
C3161 a_10182_20463# a_8970_20510# 0.07766f
C3162 sar9b_0.net67 sar9b_0._12_ 0.06679f
C3163 a_5235_27466# a_4749_27652# 0.13237f
C3164 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[7] 0.21737f
C3165 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.42014f
C3166 a_7978_22202# sar9b_0.net61 0.17441f
C3167 sar9b_0.net38 a_9930_20510# 0.02335f
C3168 sar9b_0.net7 a_11842_18434# 0.01552f
C3169 a_3946_27530# sar9b_0.net44 0.05385f
C3170 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.10429f
C3171 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C3172 VDPWR a_9930_20510# 0.34995f
C3173 a_10816_21487# a_10218_20806# 0.0165f
C3174 sar9b_0._02_ sar9b_0.clk_div_0.COUNT\[2\] 0.09854f
C3175 a_10644_16791# sar9b_0.net6 0.22613f
C3176 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.69086f
C3177 a_9900_19047# sar9b_0.net48 0.04064f
C3178 sar9b_0.net57 sar9b_0.net53 0.08138f
C3179 VDPWR a_10926_17021# 0.26037f
C3180 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.12431f
C3181 a_11178_24802# sar9b_0.net74 0.03041f
C3182 sar9b_0.net49 sar9b_0.net42 0.02948f
C3183 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[7] 0.01887f
C3184 single_9b_cdac_0.SW[7] uo_out[3] 0.06777f
C3185 sar9b_0.net33 a_12870_26263# 0.07013f
C3186 VDPWR a_6634_18206# 0.28909f
C3187 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.04988f
C3188 a_6540_22112# sar9b_0.net40 0.01639f
C3189 sar9b_0.net43 a_9730_24138# 0.06642f
C3190 sar9b_0.net26 a_12182_22423# 0.0187f
C3191 sar9b_0.net7 a_9363_20826# 0.03016f
C3192 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.17533f
C3193 VDPWR a_57946_26999# 1.81495f
C3194 a_8386_22806# a_9162_23174# 0.3578f
C3195 sar9b_0.net36 sar9b_0.net22 0.02611f
C3196 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.22875f
C3197 a_6132_23451# a_6137_23791# 0.43491f
C3198 a_5506_17478# a_6534_17799# 0.07826f
C3199 ui_in[6] ui_in[5] 0.03102f
C3200 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[0] 0.12898f
C3201 single_9b_cdac_1.SW[1] single_9b_cdac_1.CF[3] 0.22098f
C3202 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.12358f
C3203 VDPWR a_5523_21528# 0.22726f
C3204 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.01134f
C3205 a_5151_28559# uo_out[7] 0.02535f
C3206 a_10218_27466# sar9b_0.net45 0.24807f
C3207 sar9b_0.net26 a_11842_23762# 0.0241f
C3208 sar9b_0.net44 a_3545_26914# 0.05842f
C3209 single_9b_cdac_1.cdac_sw_9b_0.S[4] a_43540_16877# 0.59531f
C3210 sar9b_0.net58 a_4125_25958# 0.03759f
C3211 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.75853f
C3212 a_5581_20992# sar9b_0.net60 0.06229f
C3213 sar9b_0._18_ sar9b_0._07_ 0.02201f
C3214 a_13011_20806# a_13011_20574# 0.02551f
C3215 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.69086f
C3216 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.22875f
C3217 sar9b_0.net29 single_9b_cdac_0.SW[3] 0.06969f
C3218 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[0] 0.584f
C3219 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS dw_17224_1400# 1.26208f
C3220 dw_12589_1395# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.26214f
C3221 single_9b_cdac_1.SW[6] sar9b_0.net28 0.14409f
C3222 VDPWR a_6030_24396# 0.2481f
C3223 VDPWR sar9b_0._12_ 1.04527f
C3224 a_12064_22819# clk 0.01615f
C3225 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[1] 0.01285f
C3226 a_7097_19795# sar9b_0.net40 0.16334f
C3227 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 2.82172f
C3228 VDPWR a_13216_26469# 0.21606f
C3229 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[4] 0.03897f
C3230 sar9b_0.net41 sar9b_0.net12 0.51525f
C3231 sar9b_0.net58 sar9b_0._15_ 0.04426f
C3232 single_9b_cdac_0.SW[6] single_9b_cdac_1.CF[6] 1.79589f
C3233 sar9b_0.net46 a_6579_18832# 0.31908f
C3234 a_6534_27123# sar9b_0.net37 0.0697f
C3235 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[7] 6.17399f
C3236 sar9b_0.net74 clk 0.07221f
C3237 single_9b_cdac_0.SW[1] clk 0.13072f
C3238 a_5844_18123# a_5394_18116# 0.03471f
C3239 a_5196_18116# a_5535_18149# 0.07649f
C3240 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.02666f
C3241 sar9b_0.net35 sar9b_0.net5 0.0951f
C3242 a_8052_16791# a_7743_16817# 0.07766f
C3243 VDPWR a_48343_16877# 1.81495f
C3244 a_6137_23791# sar9b_0.net4 0.01198f
C3245 single_9b_cdac_1.CF[6] clk 0.13098f
C3246 single_9b_cdac_1.SW[0] a_9450_17846# 0.02044f
C3247 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[0] 0.31534f
C3248 single_9b_cdac_1.SW[2] single_9b_cdac_1.SW[0] 0.98657f
C3249 a_29134_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.23864f
C3250 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C3251 a_3545_26914# a_3822_27060# 0.09983f
C3252 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[2\] 1.06971f
C3253 sar9b_0.net56 a_9450_17846# 0.26827f
C3254 tdc_0.RDY a_5331_16810# 0.26021f
C3255 sar9b_0.net2 sar9b_0.net5 0.0239f
C3256 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP a_62748_26999# 0.04592f
C3257 sar9b_0.net56 single_9b_cdac_1.SW[2] 0.31153f
C3258 a_8266_18445# sar9b_0.net5 0.04964f
C3259 sar9b_0.net10 sar9b_0.net36 0.03634f
C3260 a_10742_21091# a_11178_20806# 0.16939f
C3261 a_11658_22138# a_11842_22430# 0.44532f
C3262 a_2451_27234# a_2892_27039# 0.01819f
C3263 a_10932_25713# a_10937_25582# 0.44532f
C3264 a_7539_28566# uo_out[5] 0.40403f
C3265 a_11338_19178# sar9b_0.net61 0.24596f
C3266 sar9b_0.net32 a_12435_24802# 0.03774f
C3267 a_12618_23470# clk 0.0119f
C3268 a_7936_25137# sar9b_0.net54 0.03507f
C3269 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net62 0.03763f
C3270 uio_in[2] uio_in[1] 0.03102f
C3271 a_2931_28566# sar9b_0.net60 0.09891f
C3272 a_9258_21842# a_9782_21622# 0.04522f
C3273 a_8982_21902# a_9647_21523# 0.19065f
C3274 a_6534_17799# a_5322_17846# 0.07766f
C3275 a_11146_25483# a_10932_25713# 0.05022f
C3276 sar9b_0.net40 a_6562_25094# 0.02042f
C3277 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.02632f
C3278 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C3279 sar9b_0.net9 a_7188_22119# 0.22374f
C3280 a_8438_23755# sar9b_0.net54 0.02573f
C3281 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.02149f
C3282 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C3283 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.3196f
C3284 sar9b_0._07_ a_4072_19474# 0.1462f
C3285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.28523f
C3286 sar9b_0._07_ sar9b_0.net71 0.05408f
C3287 a_5460_28377# uo_out[6] 0.03666f
C3288 VDPWR a_4044_24776# 0.26952f
C3289 sar9b_0.net47 a_7193_22459# 0.10511f
C3290 a_10926_17021# sar9b_0.net48 0.19705f
C3291 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[0] 0.02165f
C3292 single_9b_cdac_0.SW[2] a_53154_26999# 0.28324f
C3293 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[5] 0.0313f
C3294 a_5633_20244# a_5481_20185# 0.22338f
C3295 sar9b_0.net31 sar9b_0.net12 0.61825f
C3296 sar9b_0.net48 a_6634_18206# 0.28205f
C3297 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.5604f
C3298 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.62443f
C3299 a_10607_25185# a_10218_24802# 0.06034f
C3300 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.84042f
C3301 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[3] 0.12359f
C3302 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.24223f
C3303 a_10644_16791# a_11436_17742# 0.01113f
C3304 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.02149f
C3305 sar9b_0._07_ a_4332_23043# 0.07997f
C3306 sar9b_0.net42 sar9b_0.net45 0.14568f
C3307 a_11338_19178# sar9b_0.net7 0.0556f
C3308 a_5441_22522# sar9b_0._12_ 0.04735f
C3309 single_9b_cdac_1.SW[3] th_dif_sw_0.VCN 0.09454f
C3310 sar9b_0.net38 a_8691_28566# 0.0583f
C3311 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.12358f
C3312 a_8031_26141# a_8340_26115# 0.07766f
C3313 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP a_38738_26999# 0.04592f
C3314 sar9b_0.net56 sar9b_0.net9 0.089f
C3315 VDPWR a_8691_28566# 0.50803f
C3316 a_11382_26138# a_11658_26134# 0.1263f
C3317 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.01198f
C3318 sar9b_0._10_ a_5196_19448# 0.10468f
C3319 single_9b_cdac_1.SW[4] sar9b_0.net2 0.03719f
C3320 a_8303_18859# sar9b_0.net61 0.03127f
C3321 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C3322 sar9b_0.net61 single_9b_cdac_1.SW[0] 0.03934f
C3323 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[0] 0.02149f
C3324 tdc_0.OUTP tdc_0.RDY 1.84081f
C3325 sar9b_0.net52 sar9b_0.net62 0.03789f
C3326 a_5322_27170# a_6282_27170# 0.03529f
C3327 sar9b_0.net56 sar9b_0.net61 0.16507f
C3328 sar9b_0.net59 uio_out[0] 0.11978f
C3329 a_10227_23490# sar9b_0.net54 0.18976f
C3330 sar9b_0.net13 sar9b_0.net35 0.02962f
C3331 a_16185_13034# tdc_0.phase_detector_0.pd_out_0.B 0.0174f
C3332 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.26707f
C3333 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C3334 sar9b_0.net58 a_6282_27170# 0.26031f
C3335 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.38397f
C3336 VDPWR a_11178_20806# 0.35985f
C3337 sar9b_0.net35 sar9b_0.cyclic_flag_0.FINAL 0.0808f
C3338 a_18214_3039# dw_17224_1400# 1.98311f
C3339 sar9b_0.net35 sar9b_0.net15 0.01154f
C3340 a_4922_20857# a_5083_21100# 0.19021f
C3341 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._12_ 0.12298f
C3342 a_6307_27584# sar9b_0.net60 0.03874f
C3343 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C3344 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C3345 sar9b_0.net58 sar9b_0.clknet_1_1__leaf_CLK 0.05967f
C3346 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.07517f
C3347 a_7338_24802# a_6378_24802# 0.03432f
C3348 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.12431f
C3349 a_11339_27039# sar9b_0.net52 0.07246f
C3350 a_12435_24802# sar9b_0.net12 0.22022f
C3351 sar9b_0.net8 a_10742_21091# 0.03386f
C3352 a_8512_27801# sar9b_0.cyclic_flag_0.FINAL 0.03823f
C3353 a_16331_9671# th_dif_sw_0.VCP 0.10881f
C3354 sar9b_0._03_ a_4698_25851# 0.11739f
C3355 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 3.27833f
C3356 a_10506_23174# sar9b_0.net38 0.02378f
C3357 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C3358 VDPWR a_10506_23174# 0.8367f
C3359 a_3206_22432# sar9b_0.net70 0.04299f
C3360 VDPWR sar9b_0.net33 0.38773f
C3361 th_dif_sw_0.VCN single_9b_cdac_0.cdac_sw_9b_0.S[3] 27.3302f
C3362 a_4210_22378# sar9b_0.clk_div_0.COUNT\[3\] 0.12081f
C3363 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[7] 0.24198f
C3364 a_8019_17910# sar9b_0.net35 0.16492f
C3365 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.clknet_0_CLK 0.08397f
C3366 sar9b_0.net26 sar9b_0.net73 0.02035f
C3367 sar9b_0.net7 sar9b_0.net56 0.25867f
C3368 single_9b_cdac_1.CF[2] th_dif_sw_0.VCN 0.09453f
C3369 a_8874_23470# sar9b_0.net37 0.02487f
C3370 sar9b_0.net38 a_9942_20810# 0.01655f
C3371 sar9b_0.net64 sar9b_0._07_ 0.04413f
C3372 VDPWR a_9942_20810# 0.29503f
C3373 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C3374 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.42509f
C3375 tdc_0.OUTP a_13011_16810# 0.01868f
C3376 a_8691_28566# a_8883_27466# 0.01221f
C3377 a_9939_28566# a_9323_28371# 0.03551f
C3378 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 2.81428f
C3379 sar9b_0.net36 a_10402_21098# 0.0105f
C3380 sar9b_0.net43 sar9b_0.net73 0.14358f
C3381 ua[0] single_9b_cdac_0.SW[0] 0.15351f
C3382 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.19266f
C3383 a_10402_25094# a_11178_24802# 0.3578f
C3384 sar9b_0.net21 a_7539_28566# 0.20381f
C3385 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.10499f
C3386 sar9b_0.net7 a_10803_18142# 0.01039f
C3387 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.42014f
C3388 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.01664f
C3389 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.10499f
C3390 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 a_54032_17740# 0.14695f
C3391 sar9b_0.net26 sar9b_0.net6 0.75213f
C3392 a_4467_24162# sar9b_0._15_ 0.11422f
C3393 sar9b_0.net41 a_11859_17910# 0.05709f
C3394 single_9b_cdac_0.cdac_sw_9b_0.S[5] a_39616_26990# 0.22512f
C3395 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[5] 17.8424f
C3396 a_2508_20780# a_2918_20140# 0.05315f
C3397 single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.10499f
C3398 sar9b_0.net43 a_10218_24802# 0.01463f
C3399 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36037f
C3400 sar9b_0.net68 a_5196_24776# 0.14653f
C3401 a_2931_28566# uio_out[1] 0.4065f
C3402 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.03488f
C3403 uo_out[0] ui_in[0] 0.0743f
C3404 a_6880_26815# a_6534_27123# 0.07649f
C3405 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.28523f
C3406 sar9b_0._11_ a_6636_20780# 0.02384f
C3407 sar9b_0.net8 a_8694_20570# 0.05489f
C3408 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.22879f
C3409 a_6346_23773# sar9b_0.net11 0.05901f
C3410 single_9b_cdac_0.SW[5] uo_out[0] 0.08425f
C3411 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] 1.15122f
C3412 a_10402_27758# a_10742_27751# 0.24088f
C3413 a_7914_27466# sar9b_0.net45 0.07701f
C3414 VDPWR a_11859_21906# 0.45768f
C3415 a_6307_27584# sar9b_0.net40 0.10226f
C3416 sar9b_0.net44 a_3156_26115# 0.23133f
C3417 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.SW[8] 0.17126f
C3418 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.03488f
C3419 sar9b_0.net8 sar9b_0.net38 0.02476f
C3420 a_21368_4076# th_dif_sw_0.VCP 0.18144f
C3421 sar9b_0.net43 a_9942_27470# 0.17078f
C3422 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_1.CF[3] 0.01346f
C3423 VDPWR sar9b_0.net8 1.26787f
C3424 sar9b_0.net49 sar9b_0.net39 0.01106f
C3425 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.10626f
C3426 single_9b_cdac_1.CF[1] clk 0.08196f
C3427 a_5628_19768# sar9b_0.net47 0.014f
C3428 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.30106f
C3429 a_5465_28246# sar9b_0.net45 0.02195f
C3430 a_5742_28392# a_5674_28147# 0.35559f
C3431 a_5628_19768# sar9b_0._07_ 0.03465f
C3432 sar9b_0.net10 a_7402_22441# 0.01467f
C3433 sar9b_0.net10 sar9b_0.net51 0.09304f
C3434 VDPWR a_7926_23234# 0.30357f
C3435 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.04988f
C3436 a_7289_21127# sar9b_0.net47 0.10682f
C3437 sar9b_0.net60 sar9b_0.net44 0.64939f
C3438 a_9730_24138# a_10070_24286# 0.24088f
C3439 sar9b_0.net73 a_11382_22142# 0.17249f
C3440 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 3.10626f
C3441 a_13011_19242# a_13216_18477# 0.01043f
C3442 th_dif_sw_0.CK sar9b_0.net73 0.16091f
C3443 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[4] 0.31534f
C3444 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.12431f
C3445 sar9b_0.net32 a_12182_26419# 0.01466f
C3446 sar9b_0.net42 sar9b_0.net31 0.08505f
C3447 a_8554_26437# sar9b_0.cyclic_flag_0.FINAL 0.06206f
C3448 sar9b_0.net3 sar9b_0.net17 0.49213f
C3449 sar9b_0.net8 sar9b_0.net1 0.02481f
C3450 sar9b_0.net13 a_13011_25902# 0.2478f
C3451 sar9b_0.net49 a_8982_21902# 0.22591f
C3452 single_9b_cdac_0.SW[6] single_9b_cdac_1.CF[7] 0.12064f
C3453 sar9b_0.net9 sar9b_0.net57 0.06836f
C3454 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[1] 1.55946f
C3455 sar9b_0._09_ sar9b_0.net16 0.56465f
C3456 sar9b_0.net4 sar9b_0.clk_div_0.COUNT\[1\] 0.02438f
C3457 sar9b_0.net33 sar9b_0.net29 0.01075f
C3458 sar9b_0.net26 sar9b_0.net50 0.09003f
C3459 single_9b_cdac_1.CF[7] clk 0.16146f
C3460 a_8303_18859# a_8438_18958# 0.35559f
C3461 a_2892_23070# sar9b_0.clk_div_0.COUNT\[1\] 0.01011f
C3462 sar9b_0._12_ a_5523_21528# 0.17627f
C3463 sar9b_0.net2 single_9b_cdac_1.SW[1] 0.77878f
C3464 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 2.82165f
C3465 a_9450_17846# a_9174_17906# 0.1263f
C3466 sar9b_0.net57 a_6922_23534# 0.06619f
C3467 sar9b_0.net57 sar9b_0.net61 0.18181f
C3468 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.02632f
C3469 single_9b_cdac_1.SW[2] a_9174_17906# 0.07801f
C3470 tdc_0.OUTP a_10644_16791# 0.07935f
C3471 a_10858_17113# a_10194_16784# 0.16939f
C3472 sar9b_0.net44 a_5506_26802# 0.08971f
C3473 a_7404_16784# sar9b_0.net6 0.01335f
C3474 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07579f
C3475 sar9b_0.net19 a_3540_27045# 0.04938f
C3476 a_7097_19795# a_7306_19777# 0.24088f
C3477 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C3478 a_7092_19455# a_6783_19481# 0.07766f
C3479 VDPWR a_14897_9355# 0.01057f
C3480 a_21684_3438# th_dif_sw_0.th_sw_1.CK 0.12114f
C3481 th_dif_sw_0.CK sar9b_0.net6 0.02947f
C3482 sar9b_0.net38 sar9b_0.net34 0.38358f
C3483 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.59531f
C3484 sar9b_0.net20 a_5151_28559# 0.06913f
C3485 a_5010_28495# a_5460_28377# 0.03432f
C3486 VDPWR sar9b_0.net34 0.38274f
C3487 a_13011_19242# sar9b_0.net42 0.22277f
C3488 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C3489 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.CF[3] 0.01346f
C3490 sar9b_0.net40 single_9b_cdac_1.SW[8] 0.02686f
C3491 a_4018_24235# a_3014_24136# 0.06302f
C3492 a_2931_28566# a_3156_27447# 0.01146f
C3493 a_10690_22806# a_11466_23174# 0.3578f
C3494 a_5711_17527# sar9b_0.net46 0.26531f
C3495 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS w_12795_1601# 0.38264f
C3496 sar9b_0.net53 clk 0.10487f
C3497 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.26942f
C3498 a_10895_22855# clk 0.0165f
C3499 sar9b_0.net63 sar9b_0.net35 0.03292f
C3500 a_10402_27758# a_10607_27849# 0.09983f
C3501 sar9b_0.net27 a_13216_19809# 0.01127f
C3502 sar9b_0.net41 sar9b_0.net74 0.02251f
C3503 VDPWR a_5322_27170# 0.86299f
C3504 sar9b_0.net51 a_7914_19178# 0.05227f
C3505 sar9b_0.net58 sar9b_0.net38 0.14084f
C3506 a_3206_22432# a_4011_22488# 0.29207f
C3507 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[6] 0.42014f
C3508 sar9b_0.net5 single_9b_cdac_1.SW[0] 0.03107f
C3509 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.6919f
C3510 a_8052_16791# sar9b_0.net27 0.01294f
C3511 VDPWR sar9b_0.net58 3.35769f
C3512 a_10378_27170# single_9b_cdac_0.SW[7] 0.01306f
C3513 single_9b_cdac_0.SW[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.24198f
C3514 sar9b_0.net55 a_6444_21738# 0.02142f
C3515 a_9138_27163# a_9593_26914# 0.3578f
C3516 a_9279_27227# a_9588_27045# 0.07766f
C3517 a_53154_26999# single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.59531f
C3518 a_9442_21474# sar9b_0.net57 0.0155f
C3519 sar9b_0.net58 a_4330_27170# 0.28291f
C3520 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26218f
C3521 sar9b_0.net56 sar9b_0.net5 1.07927f
C3522 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38715f
C3523 sar9b_0.net35 sar9b_0.net62 0.04291f
C3524 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.07579f
C3525 sar9b_0.net59 sar9b_0.net37 0.15299f
C3526 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.01751f
C3527 sar9b_0.net40 a_6922_23534# 0.01201f
C3528 sar9b_0.net40 sar9b_0.net61 0.03026f
C3529 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[6] 0.26427f
C3530 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.02149f
C3531 sar9b_0.net36 sar9b_0.net19 0.07564f
C3532 sar9b_0.net63 sar9b_0._14_ 0.30459f
C3533 sar9b_0.net40 sar9b_0.net44 0.06639f
C3534 a_12182_19759# sar9b_0.net6 0.02207f
C3535 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.6919f
C3536 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A 0.42784f
C3537 VDPWR a_6137_23791# 0.21454f
C3538 VDPWR a_6282_17846# 0.34765f
C3539 sar9b_0.net26 single_9b_cdac_1.CF[2] 0.03846f
C3540 sar9b_0.net58 a_3370_27769# 0.14413f
C3541 sar9b_0.net2 sar9b_0.net62 0.18559f
C3542 th_dif_sw_0.CK sar9b_0.net50 0.23424f
C3543 th_dif_sw_0.CK single_9b_cdac_1.SW[3] 0.69076f
C3544 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.17156f
C3545 VDPWR a_3370_26437# 0.20923f
C3546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3547 a_9730_24138# sar9b_0.net38 0.02314f
C3548 th_dif_sw_0.CK a_12618_18142# 0.06719f
C3549 a_9802_26815# sar9b_0.net59 0.17205f
C3550 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3551 VDPWR a_9730_24138# 0.22331f
C3552 sar9b_0.net23 a_8554_26437# 0.01362f
C3553 sar9b_0.net61 a_9174_17906# 0.04236f
C3554 sar9b_0.net46 sar9b_0.net4 0.06536f
C3555 sar9b_0.net45 a_7343_27849# 0.06174f
C3556 th_dif_sw_0.th_sw_1.CK a_10482_3438# 0.1221f
C3557 single_9b_cdac_1.CF[2] a_13011_20806# 0.01099f
C3558 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[3] 1.26495f
C3559 VDPWR a_7743_18149# 0.25964f
C3560 VDPWR single_9b_cdac_1.CF[0] 2.72978f
C3561 sar9b_0.net38 uo_out[3] 0.26142f
C3562 a_12684_20379# sar9b_0.net5 0.051f
C3563 VDPWR a_8057_17131# 0.24259f
C3564 VDPWR a_7138_27758# 0.2246f
C3565 a_11178_24802# a_10932_25713# 0.02278f
C3566 sar9b_0.net21 sar9b_0.net45 0.04091f
C3567 a_16222_11316# tdc_0.phase_detector_0.INP 0.02778f
C3568 VDPWR uo_out[3] 0.80535f
C3569 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[2] 0.01791f
C3570 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.1717f
C3571 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.02638f
C3572 sar9b_0.net27 single_9b_cdac_0.SW[0] 0.01491f
C3573 VDPWR a_12182_22423# 0.19338f
C3574 sar9b_0.net14 a_12531_28566# 0.05077f
C3575 a_12870_19603# sar9b_0.net27 0.0267f
C3576 sar9b_0.net13 a_10742_25087# 0.02523f
C3577 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.19266f
C3578 sar9b_0.net4 a_6378_24802# 0.2298f
C3579 a_11915_28371# sar9b_0.net14 0.20706f
C3580 clk th_dif_sw_0.VCP 1.62194f
C3581 sar9b_0.net31 sar9b_0.net74 0.23142f
C3582 sar9b_0.net24 sar9b_0.net34 0.14505f
C3583 a_5046_17906# sar9b_0.net46 0.41373f
C3584 single_9b_cdac_0.SW[2] clk 0.13337f
C3585 sar9b_0.net36 a_10607_21189# 0.02616f
C3586 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.CF[5] 0.12358f
C3587 a_24332_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.04592f
C3588 single_9b_cdac_0.cdac_sw_9b_0.S[0] ua[0] 1.19231f
C3589 VDPWR a_13011_20574# 0.42461f
C3590 a_12182_19759# sar9b_0.net50 0.14123f
C3591 sar9b_0.net7 sar9b_0.net40 0.02438f
C3592 sar9b_0.net47 sar9b_0._07_ 0.17483f
C3593 sar9b_0.net54 a_5753_24250# 0.09858f
C3594 a_2918_20140# a_3723_20140# 0.29221f
C3595 single_9b_cdac_1.SW[4] single_9b_cdac_1.SW[0] 0.02202f
C3596 a_8726_22954# clk 0.01799f
C3597 sar9b_0.net31 a_13216_22473# 0.28434f
C3598 sar9b_0.net36 a_10803_19474# 0.21894f
C3599 sar9b_0.clk_div_0.COUNT\[1\] sar9b_0.clknet_1_1__leaf_CLK 1.13184f
C3600 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] 1.15122f
C3601 VDPWR a_11842_23762# 0.2306f
C3602 single_9b_cdac_1.CF[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.26707f
C3603 VDPWR a_3425_20244# 0.10699f
C3604 a_10858_17113# sar9b_0.net27 0.025f
C3605 a_3994_19474# a_4072_19474# 0.01029f
C3606 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.SW[5] 0.02506f
C3607 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP ua[0] 1.15121f
C3608 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.02638f
C3609 VDPWR single_9b_cdac_0.SW[4] 2.61739f
C3610 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[1\] 0.02265f
C3611 a_3371_23106# sar9b_0.clknet_1_1__leaf_CLK 0.02302f
C3612 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.75853f
C3613 sar9b_0.net52 a_11842_26426# 0.09411f
C3614 sar9b_0._09_ sar9b_0._11_ 0.01658f
C3615 a_6880_26815# sar9b_0.net37 0.04911f
C3616 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.net65 0.16477f
C3617 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.95338f
C3618 sar9b_0.net46 a_3795_19512# 0.08659f
C3619 a_6678_27470# sar9b_0.net36 0.05745f
C3620 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.0303f
C3621 th_dif_sw_0.VCN single_9b_cdac_1.SW[7] 0.09453f
C3622 sar9b_0.net38 a_10528_20155# 0.31876f
C3623 a_4947_20140# a_5931_20140# 0.08669f
C3624 single_9b_cdac_1.cdac_sw_9b_0.S[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.3601f
C3625 VDPWR a_10528_20155# 0.20299f
C3626 sar9b_0.net63 sar9b_0._16_ 0.23068f
C3627 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.02149f
C3628 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net11 0.01289f
C3629 VDPWR a_11434_16874# 0.27783f
C3630 a_10553_18922# sar9b_0.net73 0.02068f
C3631 uio_out[0] ui_in[0] 0.06786f
C3632 a_10548_19053# a_10762_18823# 0.05022f
C3633 sar9b_0.net24 uo_out[3] 0.06521f
C3634 th_dif_sw_0.CK a_9132_7271# 0.69795f
C3635 a_7914_23470# sar9b_0.net62 0.02516f
C3636 sar9b_0.net29 single_9b_cdac_1.CF[0] 0.10817f
C3637 sar9b_0.net33 a_13216_26469# 0.30861f
C3638 a_7978_22202# sar9b_0.net62 0.01108f
C3639 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.45521f
C3640 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.3196f
C3641 sar9b_0.net27 a_12618_26134# 0.03607f
C3642 sar9b_0.net26 a_12618_22138# 0.02736f
C3643 a_8726_22954# a_9162_23174# 0.16939f
C3644 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.02149f
C3645 sar9b_0.net13 a_6902_25087# 0.05284f
C3646 a_5682_23444# a_6137_23791# 0.3578f
C3647 sar9b_0.net41 sar9b_0.net39 0.25189f
C3648 a_6132_23451# a_6346_23773# 0.04522f
C3649 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] 3.10215f
C3650 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.42015f
C3651 VDPWR a_5196_19448# 0.22579f
C3652 sar9b_0.net43 a_7347_24160# 0.03385f
C3653 VDPWR a_8031_26141# 0.26325f
C3654 VDPWR a_62748_26999# 1.81495f
C3655 a_8019_17910# sar9b_0.net56 0.06841f
C3656 single_9b_cdac_1.CF[3] th_dif_sw_0.VCN 0.09453f
C3657 a_7374_19685# sar9b_0.net35 0.01051f
C3658 a_16159_13315# tdc_0.RDY 0.14369f
C3659 a_7743_18149# sar9b_0.net48 0.03022f
C3660 VDPWR a_6444_21738# 0.29205f
C3661 a_4755_22138# a_5289_22527# 0.35097f
C3662 a_7638_19238# a_7914_19178# 0.1263f
C3663 a_5465_28246# uo_out[7] 0.0105f
C3664 sar9b_0.net29 a_13011_20574# 0.02075f
C3665 a_3161_26455# a_3370_26437# 0.24088f
C3666 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[4] 0.0313f
C3667 sar9b_0.net11 a_13011_24570# 0.22279f
C3668 a_6378_24802# a_5748_24381# 0.01007f
C3669 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 a_58824_17740# 0.14695f
C3670 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.62443f
C3671 single_9b_cdac_1.CF[4] single_9b_cdac_0.SW[0] 0.47599f
C3672 a_9546_24506# a_9935_24187# 0.05462f
C3673 a_9270_24566# a_9730_24138# 0.26257f
C3674 a_11718_23127# a_12064_22819# 0.07649f
C3675 sar9b_0.net42 sar9b_0.net10 0.04131f
C3676 sar9b_0.net56 a_8842_18206# 0.0572f
C3677 sar9b_0.net44 a_3156_27447# 0.236f
C3678 a_4125_25958# sar9b_0._03_ 0.1014f
C3679 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR 0.38716f
C3680 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.84426f
C3681 sar9b_0.net32 uo_out[0] 0.0917f
C3682 a_7404_17715# sar9b_0.net5 0.05199f
C3683 a_8052_18123# a_8266_18445# 0.04522f
C3684 single_9b_cdac_0.SW[4] sar9b_0.net29 0.07482f
C3685 a_3156_26115# a_2706_26108# 0.03471f
C3686 a_2508_26108# a_2847_26141# 0.07649f
C3687 sar9b_0.net52 sar9b_0.net11 0.15337f
C3688 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.28813f
C3689 a_5394_18116# a_5535_18149# 0.27388f
C3690 a_5844_18123# a_5849_18463# 0.44098f
C3691 a_7602_16784# a_8057_17131# 0.3578f
C3692 a_6346_23773# sar9b_0.net4 0.01825f
C3693 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[5] 1.95851f
C3694 a_2893_24992# sar9b_0.net68 0.07409f
C3695 a_6954_27466# a_7138_27758# 0.44532f
C3696 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP ua[0] 1.15121f
C3697 VDPWR a_4467_24162# 0.42883f
C3698 tdc_0.OUTN a_6867_16810# 0.28739f
C3699 a_10470_21795# sar9b_0.net38 0.02191f
C3700 VDPWR a_10470_21795# 0.2699f
C3701 a_3231_27227# a_3545_26914# 0.07826f
C3702 VDPWR a_10335_16817# 0.2584f
C3703 sar9b_0.clknet_1_0__leaf_CLK a_3425_20244# 0.0505f
C3704 a_11430_20935# a_11776_21141# 0.07649f
C3705 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.A 0.26382f
C3706 sar9b_0.net32 a_9939_28566# 0.04595f
C3707 a_11658_22138# a_12870_22267# 0.07766f
C3708 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.14972f
C3709 a_2892_27039# a_3090_27163# 0.06623f
C3710 a_10937_25582# a_11214_25728# 0.09983f
C3711 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.22879f
C3712 sar9b_0.net22 uo_out[5] 0.01216f
C3713 a_10690_22806# sar9b_0.net11 0.12946f
C3714 sar9b_0.net40 sar9b_0.net5 0.02461f
C3715 a_6767_25185# sar9b_0.net54 0.20328f
C3716 clk single_9b_cdac_1.SW[2] 0.17199f
C3717 a_10816_21487# a_10218_21842# 0.06623f
C3718 a_9442_21474# a_9647_21523# 0.09983f
C3719 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C3720 sar9b_0.net32 a_12491_27662# 0.02118f
C3721 sar9b_0.net13 a_10937_25582# 0.03829f
C3722 a_11146_25483# a_11214_25728# 0.35559f
C3723 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.84061f
C3724 a_6484_22845# clk 0.01293f
C3725 sar9b_0.net13 sar9b_0.net60 0.03465f
C3726 a_2835_24136# a_3262_24141# 0.04602f
C3727 a_8874_23470# sar9b_0.net54 0.09219f
C3728 a_5331_16810# sar9b_0.net4 0.1431f
C3729 a_7289_21127# a_6834_20780# 0.3578f
C3730 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C3731 VDPWR a_11382_26138# 0.29139f
C3732 single_9b_cdac_1.SW[1] single_9b_cdac_1.SW[0] 19.2136f
C3733 single_9b_cdac_1.CF[5] ua[0] 3.57763f
C3734 single_9b_cdac_1.cdac_sw_9b_0.S[5] th_dif_sw_0.VCP 6.58553f
C3735 sar9b_0.net57 a_5535_18149# 0.01663f
C3736 sar9b_0._17_ a_6444_21738# 0.02137f
C3737 a_11434_16874# sar9b_0.net48 0.19635f
C3738 a_54032_17740# single_9b_cdac_1.SW[2] 0.18991f
C3739 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.10499f
C3740 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.0303f
C3741 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[0] 0.0313f
C3742 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C3743 a_7188_22119# a_6879_22145# 0.07766f
C3744 VDPWR sar9b_0.clk_div_0.COUNT\[1\] 0.71891f
C3745 sar9b_0.net38 sar9b_0.net73 0.26685f
C3746 sar9b_0._08_ a_5196_19448# 0.06291f
C3747 VDPWR sar9b_0.net73 1.85779f
C3748 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN ua[0] 3.10215f
C3749 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.SW[5] 0.17355f
C3750 sar9b_0.net13 sar9b_0.net57 0.17396f
C3751 VDPWR sar9b_0.net17 0.77016f
C3752 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C3753 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.75815f
C3754 a_7890_26108# sar9b_0.net59 0.30461f
C3755 sar9b_0.net52 a_8098_23762# 0.0833f
C3756 clk a_14871_9671# 0.36908f
C3757 a_9760_22819# sar9b_0.net74 0.01641f
C3758 a_7188_22119# sar9b_0.net62 0.04051f
C3759 a_24332_26999# single_9b_cdac_0.SW[8] 0.28324f
C3760 single_9b_cdac_1.SW[8] clk 0.08196f
C3761 a_13011_24802# single_9b_cdac_1.CF[7] 0.05123f
C3762 th_dif_sw_0.CK a_11658_18142# 0.06562f
C3763 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C3764 sar9b_0.net1 sar9b_0.net73 0.94195f
C3765 a_10803_18142# single_9b_cdac_1.SW[1] 0.0113f
C3766 single_9b_cdac_0.cdac_sw_9b_0.S[7] a_29134_26999# 0.59531f
C3767 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.07517f
C3768 a_10218_24802# sar9b_0.net38 0.02016f
C3769 sar9b_0.net54 sar9b_0.net37 0.24974f
C3770 sar9b_0.net42 a_11382_19478# 0.02021f
C3771 a_10548_19053# sar9b_0.net42 0.05396f
C3772 a_10607_25185# sar9b_0.net52 0.19466f
C3773 VDPWR a_3371_23106# 0.3848f
C3774 a_6252_19074# a_5844_18123# 0.01266f
C3775 VDPWR a_10218_24802# 0.81345f
C3776 sar9b_0.net41 sar9b_0.net53 0.28496f
C3777 single_9b_cdac_0.SW[4] single_9b_cdac_0.SW[3] 12.7151f
C3778 single_9b_cdac_0.cdac_sw_9b_0.S[6] ua[0] 1.66285f
C3779 a_7602_18116# a_7404_18116# 0.06623f
C3780 a_5506_26802# a_5711_26851# 0.09983f
C3781 VDPWR a_6975_20813# 0.25935f
C3782 a_24332_26999# m2_23774_26966# 0.01541f
C3783 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 3.10626f
C3784 a_12064_22819# sar9b_0.net10 0.06469f
C3785 sar9b_0.net9 clk 0.02916f
C3786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C3787 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C3788 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.07579f
C3789 sar9b_0.net40 single_9b_cdac_1.SW[4] 0.1589f
C3790 tdc_0.OUTP th_dif_sw_0.CK 0.05462f
C3791 a_9942_27470# sar9b_0.net38 0.01957f
C3792 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.26427f
C3793 a_9942_27470# VDPWR 0.30254f
C3794 VDPWR sar9b_0.net6 2.96308f
C3795 sar9b_0._05_ sar9b_0.clknet_0_CLK 0.03678f
C3796 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[3] 0.12898f
C3797 a_8591_22855# sar9b_0.net11 0.05189f
C3798 a_8202_23174# sar9b_0.net54 0.18332f
C3799 a_5100_24375# sar9b_0.net39 0.0223f
C3800 a_5581_20992# sar9b_0._09_ 0.10212f
C3801 a_4136_25584# a_4365_25770# 0.18757f
C3802 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.69086f
C3803 sar9b_0.net56 sar9b_0.net62 0.01262f
C3804 a_11915_27039# single_9b_cdac_0.SW[4] 0.38596f
C3805 a_21684_3438# th_dif_sw_0.th_sw_1.CKB 0.03405f
C3806 a_5100_24375# a_5439_24563# 0.07649f
C3807 single_9b_cdac_1.SW[6] single_9b_cdac_1.SW[0] 0.02174f
C3808 sar9b_0.net1 sar9b_0.net6 0.06186f
C3809 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[0] 3.80682f
C3810 sar9b_0.net13 sar9b_0.net40 0.24488f
C3811 sar9b_0.net60 a_5674_28147# 0.02547f
C3812 a_7590_24931# a_6562_25094# 0.07826f
C3813 sar9b_0._16_ a_3747_25724# 0.02266f
C3814 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INP 0.06558f
C3815 a_10830_19068# sar9b_0.net36 0.02201f
C3816 single_9b_cdac_0.SW[5] a_38738_26999# 0.28324f
C3817 sar9b_0.net8 a_11178_20806# 0.05383f
C3818 sar9b_0.net14 uo_out[1] 0.127f
C3819 a_10335_16817# sar9b_0.net48 0.17419f
C3820 sar9b_0._03_ sar9b_0.clknet_1_1__leaf_CLK 0.23577f
C3821 VDPWR a_7498_21109# 0.19831f
C3822 a_11658_19474# single_9b_cdac_1.SW[8] 0.01298f
C3823 uio_in[7] uio_in[6] 0.03102f
C3824 a_7404_17715# a_8019_17910# 0.02256f
C3825 sar9b_0.net40 sar9b_0.net15 0.04777f
C3826 a_3561_22527# sar9b_0.clknet_1_1__leaf_CLK 0.04276f
C3827 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.84381f
C3828 sar9b_0._17_ sar9b_0.clk_div_0.COUNT\[1\] 0.15221f
C3829 a_2508_23444# sar9b_0.clknet_1_1__leaf_CLK 1.86751f
C3830 a_48343_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.23864f
C3831 single_9b_cdac_1.CF[3] a_13011_20806# 0.35649f
C3832 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.26942f
C3833 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07517f
C3834 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.0303f
C3835 sar9b_0.net68 sar9b_0.net39 0.01595f
C3836 single_9b_cdac_1.cdac_sw_9b_0.S[1] th_dif_sw_0.VCP 0.10984p
C3837 sar9b_0.net52 a_11658_26134# 0.18819f
C3838 VDPWR sar9b_0.net46 2.39016f
C3839 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C3840 th_dif_sw_0.CK sar9b_0.net28 0.15795f
C3841 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A 0.74663f
C3842 sar9b_0.net31 sar9b_0.net53 0.91386f
C3843 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C3844 VDPWR sar9b_0.net50 2.24819f
C3845 single_9b_cdac_0.SW[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.363f
C3846 a_9930_20510# a_10528_20155# 0.06623f
C3847 VDPWR single_9b_cdac_1.SW[3] 2.54341f
C3848 a_5126_20140# a_5374_20145# 0.05308f
C3849 a_4947_20140# a_5633_20244# 0.27693f
C3850 VDPWR a_12618_18142# 0.35481f
C3851 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.05472f
C3852 a_8694_20570# a_9154_20142# 0.26257f
C3853 a_8970_20510# a_9359_20191# 0.05462f
C3854 th_dif_sw_0.CKB tdc_0.RDY 0.6441f
C3855 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.11216f
C3856 a_9323_28371# a_9323_27662# 0.0246f
C3857 sar9b_0.net1 sar9b_0.net46 0.42025f
C3858 clk a_15151_10456# 0.19995f
C3859 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 2.71729f
C3860 a_10926_17021# a_11434_16874# 0.19065f
C3861 a_53154_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.23864f
C3862 a_5443_19074# a_5811_19178# 0.08134f
C3863 a_11430_24931# a_11178_24802# 0.27388f
C3864 a_5938_22378# a_5739_22488# 0.29821f
C3865 VDPWR a_6378_24802# 0.83745f
C3866 single_9b_cdac_1.CF[1] a_12435_20806# 0.35667f
C3867 sar9b_0.net48 sar9b_0.net73 0.46206f
C3868 VDPWR a_9154_20142# 0.24213f
C3869 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.05472f
C3870 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3871 a_3603_28156# sar9b_0.net60 0.28939f
C3872 sar9b_0.net49 sar9b_0.net61 0.13664f
C3873 a_9546_24506# sar9b_0.net12 0.21444f
C3874 a_6834_20780# sar9b_0.net47 0.26333f
C3875 sar9b_0.net8 a_9942_20810# 0.03985f
C3876 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDPWR 0.38716f
C3877 a_6252_20780# sar9b_0.net4 0.02886f
C3878 sar9b_0.net55 a_7347_24160# 0.19384f
C3879 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.71729f
C3880 a_12435_24802# single_9b_cdac_1.CF[7] 0.35432f
C3881 th_dif_sw_0.th_sw_1.CKB a_10482_3438# 0.0331f
C3882 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCN 1.01731f
C3883 a_9942_27470# sar9b_0.net24 0.01062f
C3884 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.22879f
C3885 sar9b_0.net1 a_9154_20142# 0.01157f
C3886 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.19266f
C3887 single_9b_cdac_1.SW[5] ua[0] 0.13353f
C3888 a_8595_17910# single_9b_cdac_1.SW[2] 0.09011f
C3889 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.12898f
C3890 sar9b_0.net40 a_12618_19474# 0.06297f
C3891 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.0303f
C3892 a_9996_16784# a_9450_17846# 0.0165f
C3893 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.84061f
C3894 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.38037f
C3895 a_6252_20780# sar9b_0._01_ 0.14179f
C3896 sar9b_0.net30 a_12047_26517# 0.02505f
C3897 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.10503f
C3898 a_10402_27758# a_11178_27466# 0.3578f
C3899 a_5823_23477# sar9b_0.net54 0.16953f
C3900 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.17533f
C3901 a_10378_27170# sar9b_0.net38 0.01469f
C3902 sar9b_0.net35 sar9b_0.net11 0.02957f
C3903 VDPWR a_10378_27170# 0.30084f
C3904 a_6307_27584# sar9b_0.net45 0.3888f
C3905 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C3906 sar9b_0.net43 sar9b_0.net52 0.08027f
C3907 sar9b_0.net48 sar9b_0.net6 1.12384f
C3908 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.45521f
C3909 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.38397f
C3910 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.42509f
C3911 single_9b_cdac_1.CF[5] sar9b_0.net27 0.03004f
C3912 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.36044f
C3913 sar9b_0.net2 sar9b_0.net11 0.02395f
C3914 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[3] 4.15101f
C3915 single_9b_cdac_0.SW[8] uo_out[1] 0.10947f
C3916 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[4] 0.06503f
C3917 a_3819_24136# a_4018_24235# 0.29821f
C3918 sar9b_0.net63 sar9b_0.net60 0.09293f
C3919 single_9b_cdac_1.CF[5] single_9b_cdac_0.SW[5] 1.8421f
C3920 a_7193_22459# a_7402_22441# 0.24088f
C3921 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.net4 0.02026f
C3922 sar9b_0.net32 a_12618_26134# 0.01453f
C3923 VDPWR single_9b_cdac_1.CF[2] 3.12459f
C3924 sar9b_0.net7 sar9b_0.net49 0.47708f
C3925 single_9b_cdac_0.SW[5] sar9b_0.net25 0.1111f
C3926 sar9b_0.net49 a_9442_21474# 0.10581f
C3927 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 3.04383f
C3928 single_9b_cdac_1.SW[4] a_13011_17910# 0.07172f
C3929 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.10626f
C3930 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.01751f
C3931 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[3] 1.55981f
C3932 sar9b_0.net40 sar9b_0._02_ 0.48012f
C3933 sar9b_0.net20 uo_out[5] 0.09694f
C3934 VDPWR a_11436_17742# 0.21601f
C3935 a_8098_18810# a_8874_19178# 0.3578f
C3936 sar9b_0.net13 a_6538_24506# 0.03555f
C3937 sar9b_0.net6 a_12047_19857# 0.01561f
C3938 sar9b_0.net38 a_10284_25707# 0.02385f
C3939 sar9b_0.net63 sar9b_0.net57 0.63977f
C3940 a_10858_17113# a_10649_17131# 0.24088f
C3941 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[8] 0.24288f
C3942 sar9b_0.net44 a_5846_26950# 0.05309f
C3943 sar9b_0.net10 sar9b_0.net39 0.16291f
C3944 a_7602_16784# sar9b_0.net6 0.04668f
C3945 sar9b_0.net36 sar9b_0.net37 0.0292f
C3946 VDPWR a_10284_25707# 0.20062f
C3947 sar9b_0._08_ sar9b_0.net46 0.2868f
C3948 sar9b_0._11_ sar9b_0.net10 0.01541f
C3949 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.07579f
C3950 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[6] 0.31534f
C3951 sar9b_0.net40 single_9b_cdac_1.SW[1] 0.10842f
C3952 sar9b_0.net59 single_9b_cdac_0.SW[5] 0.02001f
C3953 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.62443f
C3954 VDPWR a_9132_7271# 1.60705f
C3955 sar9b_0.net48 sar9b_0.net46 0.56511f
C3956 a_44418_17740# single_9b_cdac_1.SW[4] 0.18991f
C3957 sar9b_0.net20 a_5465_28246# 0.10985f
C3958 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.SW[2] 0.17157f
C3959 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C3960 sar9b_0.net48 sar9b_0.net50 0.03024f
C3961 sar9b_0.net57 sar9b_0.net62 0.5484f
C3962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 ua[0] 0.12344f
C3963 sar9b_0.net35 a_7338_24802# 0.03288f
C3964 a_8595_17910# sar9b_0.net61 0.0485f
C3965 a_9802_26815# sar9b_0.net36 0.06626f
C3966 a_11718_23127# sar9b_0.net53 0.17359f
C3967 sar9b_0._18_ a_3219_22860# 0.07732f
C3968 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS th_dif_sw_0.VCP 0.14643f
C3969 a_11030_22954# a_11466_23174# 0.16939f
C3970 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.CF[0] 0.10499f
C3971 sar9b_0.net56 a_8052_18123# 0.21417f
C3972 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.01003f
C3973 sar9b_0.net35 a_7443_21496# 0.01956f
C3974 sar9b_0.net55 a_6444_19448# 0.01836f
C3975 VDPWR a_5046_27230# 0.28883f
C3976 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C3977 a_5046_27230# a_4330_27170# 0.03811f
C3978 a_7743_16817# sar9b_0.net27 0.02921f
C3979 sar9b_0.net50 a_12047_19857# 0.22617f
C3980 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.47485f
C3981 a_9588_27045# a_9593_26914# 0.44532f
C3982 a_7602_16784# sar9b_0.net46 0.25599f
C3983 sar9b_0.net73 a_6634_18206# 0.17082f
C3984 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C3985 sar9b_0.net27 a_11842_22430# 0.01034f
C3986 VDPWR sar9b_0._03_ 0.5857f
C3987 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C3988 sar9b_0.net63 sar9b_0.net40 0.26974f
C3989 sar9b_0.net59 a_3540_27045# 0.0106f
C3990 VDPWR a_6346_23773# 0.20258f
C3991 VDPWR a_6880_17491# 0.19624f
C3992 a_3014_24136# sar9b_0.net68 0.11549f
C3993 sar9b_0.net40 a_6879_22145# 0.02015f
C3994 sar9b_0.net44 sar9b_0.net45 0.33602f
C3995 VDPWR a_3561_22527# 0.14464f
C3996 VDPWR a_2508_23444# 1.56828f
C3997 sar9b_0.clk_div_0.COUNT\[0\] a_4332_23043# 0.84737f
C3998 single_9b_cdac_1.CF[2] sar9b_0.net29 0.03358f
C3999 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.42784f
C4000 sar9b_0.net41 single_9b_cdac_1.SW[2] 0.0369f
C4001 th_dif_sw_0.CK a_12047_18525# 0.04966f
C4002 sar9b_0.net40 sar9b_0.net62 0.08027f
C4003 a_6880_17491# sar9b_0.net1 0.01138f
C4004 sar9b_0.net56 a_7284_20787# 0.21387f
C4005 single_9b_cdac_0.SW[7] uo_out[1] 0.04613f
C4006 VDPWR a_7347_24160# 0.44946f
C4007 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[7] 0.31534f
C4008 sar9b_0.net36 a_9323_27662# 0.03315f
C4009 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[4] 9.91576f
C4010 a_7914_23470# sar9b_0.net11 0.07548f
C4011 a_10926_17021# sar9b_0.net6 0.05497f
C4012 VDPWR a_8166_27595# 0.26961f
C4013 sar9b_0.net63 a_6861_22828# 0.16938f
C4014 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4015 a_3603_28156# uio_out[1] 0.013f
C4016 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.36044f
C4017 VDPWR a_5331_16810# 0.25165f
C4018 sar9b_0.net6 a_6634_18206# 0.09307f
C4019 VDPWR a_12618_22138# 0.32654f
C4020 a_6250_28502# a_5465_28246# 0.26257f
C4021 sar9b_0.net14 sar9b_0._06_ 0.04595f
C4022 sar9b_0.net13 a_11178_24802# 0.0805f
C4023 a_6102_24806# a_6562_25094# 0.26257f
C4024 VDPWR a_5460_28377# 0.81693f
C4025 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.0303f
C4026 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.clknet_1_1__leaf_CLK 0.19127f
C4027 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 2.82172f
C4028 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.28523f
C4029 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38397f
C4030 sar9b_0.net65 sar9b_0._05_ 0.31289f
C4031 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07579f
C4032 VDPWR a_38738_16877# 1.81495f
C4033 a_10548_19053# sar9b_0.net39 0.01144f
C4034 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.11907f
C4035 a_4755_22138# sar9b_0.net39 0.1069f
C4036 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.28575f
C4037 sar9b_0.net59 sar9b_0.net36 0.44441f
C4038 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.24207f
C4039 VDPWR a_12870_23599# 0.25929f
C4040 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.01402f
C4041 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C4042 a_10098_19171# sar9b_0.net36 0.0123f
C4043 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.A 0.10129f
C4044 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.CF[5] 0.01608f
C4045 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.71649f
C4046 a_5628_19768# a_5581_19664# 0.19021f
C4047 sar9b_0.net55 sar9b_0.clk_div_0.COUNT\[2\] 0.02107f
C4048 a_7097_19795# sar9b_0.net10 0.06701f
C4049 sar9b_0.net49 sar9b_0.net5 0.51189f
C4050 single_9b_cdac_1.SW[4] clk 0.09021f
C4051 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.07517f
C4052 VDPWR ua[4] 1.80222f
C4053 sar9b_0.net41 sar9b_0.net9 0.02887f
C4054 a_11658_23470# sar9b_0.net11 0.24021f
C4055 a_3027_22138# sar9b_0.clknet_1_1__leaf_CLK 0.03197f
C4056 sar9b_0.net60 a_4947_20140# 0.08548f
C4057 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.03484f
C4058 sar9b_0.net20 sar9b_0.net21 0.32153f
C4059 sar9b_0.net10 sar9b_0.net53 0.31214f
C4060 a_15400_11316# tdc_0.phase_detector_0.INN 0.02778f
C4061 a_7289_21127# sar9b_0.net51 0.06342f
C4062 a_3695_23038# sar9b_0.clknet_1_1__leaf_CLK 0.01667f
C4063 sar9b_0.net52 a_12870_26263# 0.17285f
C4064 VDPWR a_11658_18142# 0.82655f
C4065 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A 0.42509f
C4066 sar9b_0.net41 sar9b_0.net61 0.74807f
C4067 sar9b_0.net58 a_5322_27170# 0.17211f
C4068 a_5581_20992# a_5761_21100# 0.01239f
C4069 a_4044_24776# sar9b_0.clk_div_0.COUNT\[1\] 0.26612f
C4070 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.12431f
C4071 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4072 a_9930_20510# a_9154_20142# 0.3578f
C4073 a_7914_23470# a_8098_23762# 0.44532f
C4074 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.81434f
C4075 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.28523f
C4076 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C4077 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.22939f
C4078 a_5126_20140# a_6130_20239# 0.06302f
C4079 single_9b_cdac_0.SW[5] ua[0] 0.1911f
C4080 th_dif_sw_0.CKB th_dif_sw_0.VCN 0.12032f
C4081 sar9b_0.net7 a_10218_20806# 0.06569f
C4082 sar9b_0.net26 sar9b_0.net2 0.02343f
C4083 VDPWR tdc_0.OUTP 0.58425f
C4084 sar9b_0.net18 a_2508_27440# 0.28434f
C4085 a_3603_28156# a_3156_27447# 0.02744f
C4086 sar9b_0._09_ a_5481_20185# 0.02188f
C4087 a_10830_19068# a_10762_18823# 0.35559f
C4088 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 3.10626f
C4089 th_dif_sw_0.CK th_dif_sw_0.th_sw_1.CK 0.01565f
C4090 sar9b_0.net43 sar9b_0.net35 0.06071f
C4091 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.42784f
C4092 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.1588f
C4093 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_14871_9671# 0.18915f
C4094 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_0.SW[8] 0.15864f
C4095 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C4096 a_3438_26345# sar9b_0.net59 0.22622f
C4097 sar9b_0.net26 a_12047_22521# 0.01371f
C4098 a_5682_23444# a_6346_23773# 0.16939f
C4099 sar9b_0.net60 uo_out[6] 0.01362f
C4100 VDPWR a_6444_19448# 0.20267f
C4101 sar9b_0.net43 sar9b_0.net2 1.88515f
C4102 a_8345_26455# sar9b_0.net37 0.02763f
C4103 sar9b_0.net35 a_6132_23451# 0.01493f
C4104 tdc_0.phase_detector_0.pd_out_0.B tdc_0.RDY 0.0496f
C4105 VDPWR a_7470_22349# 0.26136f
C4106 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C4107 a_4934_22432# a_5938_22378# 0.06302f
C4108 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.10429f
C4109 a_8098_18810# a_7914_19178# 0.44098f
C4110 sar9b_0.net41 sar9b_0.net7 0.05595f
C4111 a_6538_24506# sar9b_0.net62 0.1665f
C4112 m2_23774_26966# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.26684f
C4113 VDPWR a_11722_25838# 0.30045f
C4114 a_10742_27751# sar9b_0.net45 0.02244f
C4115 sar9b_0.net41 a_9442_21474# 0.01846f
C4116 sar9b_0.net51 sar9b_0.net37 0.03332f
C4117 sar9b_0.net66 sar9b_0._04_ 0.02178f
C4118 a_5931_20140# sar9b_0.net4 0.01405f
C4119 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.SW[0] 0.22983f
C4120 single_9b_cdac_1.SW[3] a_48343_16877# 0.28324f
C4121 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP a_24332_16877# 0.04592f
C4122 a_3747_25724# a_4136_25584# 0.06302f
C4123 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02652f
C4124 a_10194_16784# sar9b_0.net27 0.05895f
C4125 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.0303f
C4126 a_8303_23853# a_8438_23755# 0.35559f
C4127 a_9472_23805# a_9126_23599# 0.07649f
C4128 a_11178_20806# sar9b_0.net73 0.01344f
C4129 VDPWR a_12531_28566# 0.45349f
C4130 a_10662_17799# a_9450_17846# 0.07766f
C4131 clk tdc_0.phase_detector_0.INP 0.18819f
C4132 a_3946_27530# a_3161_27787# 0.26257f
C4133 a_11915_28371# VDPWR 0.45787f
C4134 a_10662_17799# single_9b_cdac_1.SW[2] 0.03662f
C4135 VDPWR a_57946_16877# 1.81495f
C4136 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 3.10626f
C4137 sar9b_0.net35 a_7404_16784# 0.26643f
C4138 a_13011_17910# single_9b_cdac_1.SW[6] 0.35507f
C4139 a_7374_19685# sar9b_0.net40 0.01327f
C4140 a_2835_24136# sar9b_0.clknet_1_1__leaf_CLK 0.33556f
C4141 a_13011_19242# single_9b_cdac_1.SW[8] 0.01098f
C4142 VDPWR sar9b_0.net28 1.71321f
C4143 a_7092_19455# sar9b_0.net40 0.0376f
C4144 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[5] 0.01577f
C4145 sar9b_0.net33 a_11382_26138# 0.06166f
C4146 a_8595_17910# sar9b_0.net5 0.02485f
C4147 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.02638f
C4148 a_7602_18116# a_8057_18463# 0.3578f
C4149 a_2706_26108# a_2847_26141# 0.27388f
C4150 sar9b_0.net43 a_10758_24459# 0.03693f
C4151 a_12064_22819# a_11658_22138# 0.0165f
C4152 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[6] 0.02149f
C4153 a_5535_18149# a_5849_18463# 0.07826f
C4154 a_21368_4076# a_21684_3438# 0.62294f
C4155 a_5844_18123# a_6058_18445# 0.04522f
C4156 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96893f
C4157 VDPWR a_6252_20780# 0.26608f
C4158 VDPWR single_9b_cdac_1.SW[7] 2.36972f
C4159 a_6954_27466# a_8166_27595# 0.07766f
C4160 a_10707_23470# sar9b_0.net38 0.01005f
C4161 sar9b_0.net2 th_dif_sw_0.CK 0.02407f
C4162 a_10859_26330# sar9b_0.net36 0.01882f
C4163 sar9b_0.net67 a_3027_22138# 0.0723f
C4164 a_3822_27060# a_3754_26815# 0.35559f
C4165 VDPWR a_10707_23470# 0.26572f
C4166 sar9b_0.net56 a_9634_17478# 0.02665f
C4167 sar9b_0.net32 single_9b_cdac_1.CF[5] 0.011f
C4168 a_13011_23238# a_13216_23805# 0.01179f
C4169 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.18989f
C4170 sar9b_0.net43 a_9138_27163# 0.01333f
C4171 VDPWR a_9258_21842# 0.86858f
C4172 VDPWR a_9472_23805# 0.20106f
C4173 sar9b_0.net32 sar9b_0.net25 0.11681f
C4174 a_13011_20574# single_9b_cdac_1.CF[0] 0.36053f
C4175 sar9b_0._18_ sar9b_0.clknet_0_CLK 0.14719f
C4176 a_11842_22430# a_12870_22267# 0.07826f
C4177 a_11382_22142# a_12047_22521# 0.19065f
C4178 a_3090_27163# a_3231_27227# 0.27388f
C4179 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4180 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 1.50841f
C4181 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[2] 1.55949f
C4182 sar9b_0.net1 a_10707_23470# 0.25386f
C4183 a_11030_22954# sar9b_0.net11 0.0681f
C4184 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 a_58824_26990# 0.14695f
C4185 a_9546_24506# a_10506_24506# 0.03504f
C4186 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 a_25210_26990# 0.14695f
C4187 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.05279f
C4188 a_9647_21523# a_9782_21622# 0.35559f
C4189 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 3.27833f
C4190 a_13164_28398# uo_out[0] 0.0371f
C4191 a_9258_21842# sar9b_0.net1 0.01455f
C4192 a_8340_26115# a_9138_27163# 0.01342f
C4193 a_9472_23805# sar9b_0.net1 0.01959f
C4194 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.75853f
C4195 sar9b_0._02_ clk 0.01536f
C4196 a_3156_27447# a_2706_27440# 0.03471f
C4197 a_2508_27440# a_2847_27473# 0.07649f
C4198 sar9b_0.net70 a_3262_24141# 0.13578f
C4199 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.VCN 0.21849f
C4200 sar9b_0.net47 a_5581_19664# 0.07464f
C4201 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C4202 sar9b_0._14_ sar9b_0._15_ 0.01749f
C4203 VDPWR single_9b_cdac_1.CF[3] 2.76152f
C4204 single_9b_cdac_1.CF[4] ua[0] 3.57685f
C4205 sar9b_0._07_ a_5581_19664# 0.33323f
C4206 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38733f
C4207 single_9b_cdac_1.cdac_sw_9b_0.S[2] ua[0] 1.21558f
C4208 a_15151_10456# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.09051f
C4209 th_dif_sw_0.VCN single_9b_cdac_1.SW[0] 0.15316f
C4210 VDPWR sar9b_0.clk_div_0.COUNT\[2\] 1.36928f
C4211 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.28523f
C4212 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.62443f
C4213 sar9b_0.net47 a_7402_22441# 0.15391f
C4214 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.07517f
C4215 sar9b_0.net47 sar9b_0.net51 0.49323f
C4216 tdc_0.OUTP sar9b_0.net48 0.1166f
C4217 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.CF[3] 0.105f
C4218 sar9b_0.net45 a_10607_27849# 0.05607f
C4219 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.07852f
C4220 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[0] 18.6879f
C4221 a_11658_19474# a_12618_19474# 0.03432f
C4222 sar9b_0.net70 sar9b_0.net66 0.02815f
C4223 sar9b_0.net19 sar9b_0.net39 0.0141f
C4224 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.14695f
C4225 a_29134_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.23864f
C4226 sar9b_0.net52 a_9165_24988# 0.35265f
C4227 a_10662_17799# sar9b_0.net61 0.05961f
C4228 single_9b_cdac_1.SW[1] clk 0.99126f
C4229 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[0] 0.7639f
C4230 a_10607_25185# a_10742_25087# 0.35559f
C4231 a_8345_26455# sar9b_0.net59 0.08274f
C4232 sar9b_0.net52 a_9126_23599# 0.20232f
C4233 clk a_15265_9613# 0.01191f
C4234 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP a_43540_16877# 0.04592f
C4235 a_3166_20145# a_3273_20185# 0.14439f
C4236 th_dif_sw_0.CK a_11842_18434# 0.11252f
C4237 VDPWR a_3027_22138# 0.44684f
C4238 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.81428f
C4239 a_8554_26437# a_8340_26115# 0.04522f
C4240 a_7289_21127# a_7566_21017# 0.09983f
C4241 VDPWR a_13011_24570# 0.48259f
C4242 a_10194_16784# sar9b_0.net36 0.05607f
C4243 single_9b_cdac_1.cdac_sw_9b_0.S[4] ua[0] 1.94611f
C4244 a_8874_19178# sar9b_0.net61 0.01101f
C4245 sar9b_0.net29 sar9b_0.net28 1.82558f
C4246 single_9b_cdac_1.cdac_sw_9b_0.S[6] a_33936_16877# 0.59531f
C4247 sar9b_0.net8 sar9b_0.net73 0.02045f
C4248 VDPWR a_3695_23038# 0.22559f
C4249 a_6252_20780# sar9b_0._17_ 0.05545f
C4250 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN single_9b_cdac_1.SW[8] 0.1495f
C4251 a_13011_16810# sar9b_0.net40 0.21779f
C4252 VDPWR a_5938_22378# 0.38557f
C4253 sar9b_0.net16 a_4072_19474# 0.04195f
C4254 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_60565_29911# 0.01076f
C4255 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C4256 sar9b_0.net16 sar9b_0.net71 0.48375f
C4257 a_5711_26851# a_5846_26950# 0.35559f
C4258 sar9b_0.net30 a_12182_23755# 0.02293f
C4259 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[7] 0.02149f
C4260 a_24332_26999# VDPWR 1.81495f
C4261 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.10499f
C4262 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.11216f
C4263 single_9b_cdac_1.SW[5] a_39616_17740# 0.18991f
C4264 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.12358f
C4265 sar9b_0.net31 a_11430_24931# 0.0265f
C4266 sar9b_0.net52 sar9b_0.net38 0.0649f
C4267 a_16222_11316# tdc_0.phase_detector_0.pd_out_0.A 0.48692f
C4268 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[8] 0.363f
C4269 VDPWR sar9b_0.net52 3.91808f
C4270 sar9b_0.net63 clk 0.08413f
C4271 a_3561_22527# sar9b_0._12_ 0.03484f
C4272 a_4365_25770# a_4293_25852# 0.22517f
C4273 sar9b_0.clknet_0_CLK a_4332_23043# 1.32864f
C4274 a_4467_24162# sar9b_0.net58 0.09475f
C4275 a_11008_17491# a_10410_17846# 0.06623f
C4276 sar9b_0.net41 sar9b_0.net5 0.02649f
C4277 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.43767f
C4278 sar9b_0.net15 a_6252_19074# 0.25177f
C4279 a_7338_24802# a_6902_25087# 0.16939f
C4280 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 2.82222f
C4281 sar9b_0._07_ sar9b_0.clk_div_0.COUNT\[0\] 0.02059f
C4282 a_3372_25734# sar9b_0.net69 0.14523f
C4283 a_4136_25584# a_4698_25851# 0.05308f
C4284 sar9b_0.net42 a_11430_20935# 0.01027f
C4285 sar9b_0.net8 sar9b_0.net6 0.09366f
C4286 clk sar9b_0.net62 0.06683f
C4287 VDPWR a_6783_19481# 0.27053f
C4288 sar9b_0._17_ sar9b_0.clk_div_0.COUNT\[2\] 0.57711f
C4289 sar9b_0.net36 a_10410_17846# 0.02317f
C4290 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C4291 a_6678_27470# a_7343_27849# 0.19065f
C4292 single_9b_cdac_1.CF[3] sar9b_0.net29 0.47519f
C4293 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 3.10626f
C4294 a_11842_19766# single_9b_cdac_1.SW[8] 0.02175f
C4295 a_10166_3438# a_10482_3438# 0.62294f
C4296 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 2.82215f
C4297 VDPWR a_10690_22806# 0.22042f
C4298 single_9b_cdac_1.SW[6] clk 0.08446f
C4299 sar9b_0.net45 sar9b_0.cyclic_flag_0.FINAL 0.18011f
C4300 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[0] 0.27554f
C4301 a_6678_27470# sar9b_0.net21 0.01436f
C4302 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.01003f
C4303 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C4304 single_9b_cdac_1.SW[0] a_63626_17740# 0.18991f
C4305 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38702f
C4306 sar9b_0.net60 sar9b_0.net11 0.10348f
C4307 a_11338_19178# sar9b_0.net26 0.05306f
C4308 sar9b_0.net32 sar9b_0.net30 1.27934f
C4309 a_10227_23490# sar9b_0.net53 0.38452f
C4310 a_4749_27652# uo_out[7] 0.01802f
C4311 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[1] 17.5055f
C4312 a_5126_20140# a_5481_20185# 0.18752f
C4313 VDPWR a_12047_18525# 0.26725f
C4314 a_13011_21906# sar9b_0.net27 0.03613f
C4315 VDPWR a_2835_24136# 0.52652f
C4316 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0313f
C4317 sar9b_0._14_ sar9b_0.clknet_1_1__leaf_CLK 0.02074f
C4318 a_10926_17021# tdc_0.OUTP 0.06343f
C4319 sar9b_0.net35 sar9b_0.net55 0.02784f
C4320 th_dif_sw_0.CK th_dif_sw_0.CKB 0.08006f
C4321 sar9b_0.net58 sar9b_0.net17 0.01182f
C4322 a_5010_28495# sar9b_0.net60 0.06731f
C4323 a_11178_24802# a_11776_25137# 0.06623f
C4324 a_5811_19178# a_6252_19074# 0.0184f
C4325 a_3219_22860# sar9b_0._07_ 0.20806f
C4326 sar9b_0.net29 a_13011_24570# 0.02017f
C4327 sar9b_0.net28 single_9b_cdac_0.SW[3] 0.05131f
C4328 VDPWR a_9494_20290# 0.20426f
C4329 a_5289_22527# sar9b_0._07_ 0.01435f
C4330 sar9b_0.net57 sar9b_0.net11 0.86992f
C4331 single_9b_cdac_0.SW[8] uo_out[2] 0.10257f
C4332 sar9b_0.net3 a_2451_27234# 0.15641f
C4333 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.17533f
C4334 sar9b_0.net8 sar9b_0.net50 0.34359f
C4335 sar9b_0.clknet_0_CLK sar9b_0.net72 0.06286f
C4336 a_10762_18823# a_10098_19171# 0.16939f
C4337 single_9b_cdac_1.CF[8] ua[0] 5.00726f
C4338 a_9942_27470# sar9b_0.net34 0.03758f
C4339 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C4340 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.SW[7] 0.22983f
C4341 sar9b_0._18_ sar9b_0.net39 0.295f
C4342 a_10402_27758# single_9b_cdac_0.SW[7] 0.01715f
C4343 a_10182_20463# sar9b_0.net51 0.04388f
C4344 sar9b_0.net41 single_9b_cdac_1.SW[4] 0.24901f
C4345 sar9b_0.net1 a_9494_20290# 0.02028f
C4346 sar9b_0._11_ sar9b_0._18_ 0.03308f
C4347 sar9b_0.net64 sar9b_0.clknet_0_CLK 0.01151f
C4348 a_11008_17491# sar9b_0.net27 0.01194f
C4349 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.28523f
C4350 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.10429f
C4351 sar9b_0.net8 a_9154_20142# 0.01901f
C4352 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.02632f
C4353 a_10230_23234# sar9b_0.net36 0.01418f
C4354 a_11430_27595# a_11178_27466# 0.27388f
C4355 VDPWR a_4922_20857# 0.22486f
C4356 sar9b_0.net9 sar9b_0.net10 0.65359f
C4357 sar9b_0.net72 a_2893_24992# 0.03569f
C4358 a_7890_26108# a_8345_26455# 0.3578f
C4359 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y 0.07579f
C4360 sar9b_0.net36 sar9b_0.net27 0.4102f
C4361 a_7743_18149# sar9b_0.net73 0.09002f
C4362 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.28813f
C4363 sar9b_0.clknet_1_0__leaf_CLK a_3027_22138# 0.26938f
C4364 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.94957f
C4365 sar9b_0.net13 a_7590_24931# 0.04157f
C4366 a_6642_19448# sar9b_0.net47 0.33504f
C4367 sar9b_0.net41 sar9b_0.net13 0.0247f
C4368 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.05472f
C4369 a_10218_27466# sar9b_0.net59 0.16798f
C4370 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 1.56111f
C4371 a_6922_23534# sar9b_0.net10 0.17349f
C4372 sar9b_0.net10 sar9b_0.net61 0.02017f
C4373 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.11944f
C4374 VDPWR a_8591_22855# 0.29655f
C4375 single_9b_cdac_1.SW[1] a_58824_17740# 0.18991f
C4376 a_7566_21017# sar9b_0.net47 0.24689f
C4377 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C4378 a_13011_16810# a_13011_17910# 0.0246f
C4379 a_8386_22806# sar9b_0.net37 0.03128f
C4380 single_9b_cdac_1.CF[3] single_9b_cdac_0.SW[3] 1.96064f
C4381 sar9b_0._01_ a_5633_20244# 0.01113f
C4382 sar9b_0.net32 a_12047_26517# 0.01148f
C4383 sar9b_0.net2 a_10070_24286# 0.0649f
C4384 a_10482_3438# a_10254_2858# 0.11186f
C4385 sar9b_0.net49 a_9782_21622# 0.15031f
C4386 sar9b_0.net40 sar9b_0.net11 0.02451f
C4387 sar9b_0.net23 sar9b_0.net45 0.02681f
C4388 a_8438_18958# a_8874_19178# 0.16939f
C4389 sar9b_0.net57 a_8098_23762# 0.06831f
C4390 VDPWR a_5196_18116# 0.20215f
C4391 a_11859_21906# single_9b_cdac_1.CF[2] 0.35504f
C4392 VDPWR uo_out[1] 0.933f
C4393 ui_in[5] ui_in[4] 0.03102f
C4394 sar9b_0.net43 a_11030_22954# 0.01262f
C4395 sar9b_0.net52 a_9270_24566# 0.02178f
C4396 a_9174_17906# a_9634_17478# 0.26257f
C4397 a_9450_17846# a_9839_17527# 0.05462f
C4398 sar9b_0.net67 a_3454_22567# 0.1221f
C4399 sar9b_0.net2 a_10742_21091# 0.02055f
C4400 a_8202_23174# a_8386_22806# 0.43491f
C4401 single_9b_cdac_1.SW[2] a_9839_17527# 0.06063f
C4402 sar9b_0.net38 a_10623_25895# 0.02019f
C4403 sar9b_0.net30 sar9b_0.net12 0.09512f
C4404 sar9b_0.net56 a_9126_19131# 0.02432f
C4405 VDPWR a_10623_25895# 0.25685f
C4406 sar9b_0.net26 a_12684_20379# 0.01826f
C4407 a_7306_19777# a_7374_19685# 0.35559f
C4408 sar9b_0.net45 a_9593_26914# 0.02056f
C4409 a_5711_17527# sar9b_0.net56 0.06214f
C4410 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.19143f
C4411 a_7193_22459# sar9b_0.net39 0.17464f
C4412 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C4413 a_7092_19455# a_7306_19777# 0.04522f
C4414 VDPWR th_dif_sw_0.th_sw_1.CK 2.01535f
C4415 a_5753_24250# a_5962_24151# 0.24088f
C4416 single_9b_cdac_1.CF[1] single_9b_cdac_0.SW[0] 0.32684f
C4417 sar9b_0.net31 a_11214_25728# 0.01178f
C4418 a_9546_24506# sar9b_0.net53 0.19966f
C4419 sar9b_0._16_ sar9b_0.clknet_1_1__leaf_CLK 0.07072f
C4420 sar9b_0._18_ sar9b_0.net65 0.08636f
C4421 a_13011_21906# single_9b_cdac_1.CF[4] 0.35507f
C4422 a_6282_17846# sar9b_0.net46 0.32729f
C4423 sar9b_0.net12 a_9942_24806# 0.21789f
C4424 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 a_30012_26990# 0.14695f
C4425 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.19147f
C4426 th_dif_sw_0.CK th_dif_sw_0.th_sw_1.CKB 0.09539f
C4427 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C4428 sar9b_0.net13 sar9b_0.net31 0.02786f
C4429 VDPWR a_5931_20140# 0.09106f
C4430 sar9b_0.net23 a_9870_27060# 0.01769f
C4431 a_4332_23043# sar9b_0.net39 0.05206f
C4432 a_11466_23174# clk 0.02108f
C4433 single_9b_cdac_0.SW[7] uo_out[2] 0.69613f
C4434 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.12367f
C4435 th_dif_sw_0.CK single_9b_cdac_1.SW[0] 0.05143f
C4436 a_4922_20857# sar9b_0._17_ 0.32016f
C4437 a_5439_24563# a_5753_24250# 0.07826f
C4438 a_8874_19178# sar9b_0.net5 0.01167f
C4439 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.01608f
C4440 ua[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 3.10218f
C4441 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 1.71649f
C4442 a_10378_27170# sar9b_0.net34 0.01673f
C4443 VDPWR a_16159_13315# 0.22342f
C4444 a_12560_27128# sar9b_0.net27 0.02362f
C4445 sar9b_0.net53 a_11658_22138# 0.16567f
C4446 a_7743_18149# sar9b_0.net46 0.17277f
C4447 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[0] 1.12533f
C4448 a_9593_26914# a_9870_27060# 0.09983f
C4449 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[0] 0.06503f
C4450 a_8057_17131# sar9b_0.net46 0.08295f
C4451 single_9b_cdac_0.SW[2] a_12491_27662# 0.03543f
C4452 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[0] 0.37948f
C4453 sar9b_0.net27 a_12870_22267# 0.02852f
C4454 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0303f
C4455 single_9b_cdac_0.SW[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.15108f
C4456 a_4922_20857# sar9b_0._08_ 0.02439f
C4457 sar9b_0.net56 sar9b_0.net4 0.03241f
C4458 VDPWR a_3454_22567# 0.01572f
C4459 VDPWR a_8266_17113# 0.19893f
C4460 sar9b_0.net32 a_9323_28371# 0.22468f
C4461 VDPWR sar9b_0.net35 1.86196f
C4462 a_11915_27039# sar9b_0.net52 0.03127f
C4463 a_3603_28156# sar9b_0.net18 0.02874f
C4464 sar9b_0.net42 sar9b_0.net59 0.13366f
C4465 a_10548_19053# sar9b_0.net61 0.01669f
C4466 a_10803_18142# th_dif_sw_0.CK 0.095f
C4467 sar9b_0.net23 sar9b_0.net41 0.03354f
C4468 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[4] 0.06019f
C4469 sar9b_0.net61 a_9839_17527# 0.01999f
C4470 sar9b_0.net2 sar9b_0.net38 0.03026f
C4471 a_16331_9671# th_dif_sw_0.VCN 0.0647f
C4472 sar9b_0._12_ sar9b_0.clk_div_0.COUNT\[2\] 0.06165f
C4473 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C4474 VDPWR sar9b_0.net2 1.0982f
C4475 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[7] 0.19143f
C4476 a_10194_16784# a_10649_17131# 0.3578f
C4477 VDPWR a_8266_18445# 0.19813f
C4478 a_8940_24402# sar9b_0.net37 0.01757f
C4479 sar9b_0.net35 sar9b_0.net1 0.20023f
C4480 a_11434_16874# sar9b_0.net6 0.07229f
C4481 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.11216f
C4482 sar9b_0.net56 a_5046_17906# 0.13749f
C4483 sar9b_0.net34 a_10284_25707# 0.27185f
C4484 VDPWR a_8512_27801# 0.19986f
C4485 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.94202f
C4486 VDPWR a_13011_27234# 0.41846f
C4487 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.42784f
C4488 VDPWR sar9b_0._14_ 0.55641f
C4489 a_5739_22488# sar9b_0.net60 0.01946f
C4490 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22497f
C4491 VDPWR a_5235_27466# 0.38926f
C4492 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.7611f
C4493 sar9b_0.net65 a_4812_21738# 0.15545f
C4494 VDPWR a_12047_22521# 0.24932f
C4495 a_8266_18445# sar9b_0.net1 0.0136f
C4496 VDPWR a_5742_28392# 0.25649f
C4497 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.02666f
C4498 sar9b_0.net70 a_2892_23070# 0.01508f
C4499 sar9b_0.net41 single_9b_cdac_1.SW[1] 0.01957f
C4500 single_9b_cdac_1.CF[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.12898f
C4501 a_21684_3438# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.63339f
C4502 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[6] 14.2348f
C4503 a_3027_22138# sar9b_0._12_ 0.16198f
C4504 single_9b_cdac_1.CF[8] sar9b_0.net27 0.09104f
C4505 a_9414_23127# clk 0.01589f
C4506 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42509f
C4507 a_7539_28566# uo_out[6] 0.08058f
C4508 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[5] 0.01513f
C4509 sar9b_0.net43 sar9b_0.net60 0.02362f
C4510 VDPWR a_13216_23805# 0.20771f
C4511 a_11339_27039# sar9b_0.net45 0.10933f
C4512 a_5298_24499# sar9b_0.net60 0.011f
C4513 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.24199f
C4514 a_5938_22378# sar9b_0._12_ 0.07878f
C4515 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 2.81139f
C4516 single_9b_cdac_1.CF[2] single_9b_cdac_1.CF[0] 0.03575f
C4517 a_10548_19053# sar9b_0.net7 0.21355f
C4518 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A 2.29405f
C4519 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.26218f
C4520 VDPWR a_10758_24459# 0.26555f
C4521 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.28033f
C4522 sar9b_0.net32 sar9b_0.net27 0.2123f
C4523 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VDPWR 0.84061f
C4524 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.71649f
C4525 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 a_63626_17740# 0.14695f
C4526 sar9b_0.net32 single_9b_cdac_0.SW[5] 0.11624f
C4527 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.07579f
C4528 sar9b_0.net60 sar9b_0._10_ 0.38542f
C4529 a_9130_26198# sar9b_0.net41 0.17586f
C4530 a_4044_24776# sar9b_0.clk_div_0.COUNT\[2\] 0.01228f
C4531 a_43540_16877# single_9b_cdac_1.SW[4] 0.28324f
C4532 a_5322_27170# a_5046_27230# 0.1263f
C4533 sar9b_0.net43 sar9b_0.net57 0.05729f
C4534 VDPWR a_9138_27163# 0.37075f
C4535 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 0.24371f
C4536 VDPWR a_11842_18434# 0.23262f
C4537 a_8940_27039# sar9b_0.net37 0.05651f
C4538 sar9b_0.net58 a_5046_27230# 0.26485f
C4539 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0313f
C4540 a_11430_20935# sar9b_0.net39 0.02333f
C4541 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.31534f
C4542 a_9930_20510# a_9494_20290# 0.16939f
C4543 a_7914_23470# a_9126_23599# 0.07766f
C4544 a_7478_27751# sar9b_0.net36 0.06675f
C4545 sar9b_0.net35 sar9b_0._17_ 0.03063f
C4546 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 0.19266f
C4547 a_6738_22112# sar9b_0.net35 0.02157f
C4548 sar9b_0._07_ sar9b_0.clknet_0_CLK 0.16508f
C4549 sar9b_0.net57 a_6132_23451# 0.24363f
C4550 sar9b_0._07_ sar9b_0.net16 0.16722f
C4551 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[0] 0.01167f
C4552 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[5] 0.02021f
C4553 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.7611f
C4554 m2_23774_17236# single_9b_cdac_1.SW[8] 0.02037f
C4555 sar9b_0.net57 sar9b_0._10_ 0.02676f
C4556 sar9b_0.net7 a_10402_21098# 0.08721f
C4557 sar9b_0.net12 sar9b_0.net54 0.03647f
C4558 sar9b_0.net58 sar9b_0._03_ 0.03496f
C4559 a_10335_16817# sar9b_0.net6 0.04672f
C4560 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.84061f
C4561 VDPWR a_9363_20826# 0.44006f
C4562 sar9b_0.net18 a_2706_27440# 0.06755f
C4563 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[5] 7.94111f
C4564 sar9b_0.net4 a_5394_18116# 0.02958f
C4565 sar9b_0.net3 sar9b_0.net60 0.11243f
C4566 a_10553_18922# a_11338_19178# 0.26257f
C4567 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.26942f
C4568 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[6] 0.24288f
C4569 a_10995_28566# single_9b_cdac_0.SW[5] 0.01783f
C4570 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_15265_9613# 0.16728f
C4571 sar9b_0.net41 single_9b_cdac_1.SW[6] 0.01701f
C4572 sar9b_0.net40 sar9b_0.net26 0.02504f
C4573 single_9b_cdac_0.SW[6] uo_out[4] 0.02556f
C4574 a_3946_26198# sar9b_0.net59 0.24509f
C4575 sar9b_0.net35 sar9b_0.net48 0.03579f
C4576 a_13011_27234# sar9b_0.net29 0.01376f
C4577 a_9162_23174# a_9414_23127# 0.27388f
C4578 single_9b_cdac_1.CF[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.26707f
C4579 a_9363_20826# sar9b_0.net1 0.02566f
C4580 a_6137_23791# a_6346_23773# 0.24088f
C4581 a_6282_17846# a_6880_17491# 0.06623f
C4582 sar9b_0.net60 sar9b_0.net4 0.69419f
C4583 VDPWR a_8554_26437# 0.21407f
C4584 sar9b_0.net60 sar9b_0._15_ 0.04165f
C4585 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.CF[6] 0.03484f
C4586 a_3371_23106# sar9b_0.clk_div_0.COUNT\[1\] 0.10763f
C4587 sar9b_0.net13 a_6102_24806# 0.23362f
C4588 VDPWR a_7914_23470# 0.85718f
C4589 sar9b_0.net2 sar9b_0.net48 0.03105f
C4590 sar9b_0.net13 a_5580_24776# 0.01209f
C4591 VDPWR a_7978_22202# 0.29273f
C4592 a_8266_18445# sar9b_0.net48 0.02071f
C4593 VDPWR a_3946_27530# 0.29317f
C4594 a_4755_22138# a_5182_22567# 0.04602f
C4595 sar9b_0.net9 a_10218_21842# 0.02303f
C4596 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[3] 4.15032f
C4597 VDPWR sar9b_0._16_ 0.84748f
C4598 a_8438_18958# a_7914_19178# 0.04522f
C4599 VDPWR a_13011_25902# 0.47442f
C4600 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 2.824f
C4601 sar9b_0.net41 a_9782_21622# 0.02219f
C4602 sar9b_0.net43 sar9b_0.net40 0.02302f
C4603 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.22879f
C4604 a_10859_26330# sar9b_0.net42 0.04314f
C4605 sar9b_0._01_ sar9b_0.net60 0.26299f
C4606 single_9b_cdac_0.SW[2] a_54032_26990# 0.18991f
C4607 a_6484_22845# a_6744_23238# 0.17405f
C4608 sar9b_0.net40 a_10035_19474# 0.05886f
C4609 a_8595_17910# a_8052_18123# 0.0131f
C4610 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.S[0] 0.01492f
C4611 a_4125_25958# a_4136_25584# 0.54361f
C4612 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.28523f
C4613 sar9b_0.net29 a_13216_23805# 0.01558f
C4614 a_10649_17131# sar9b_0.net27 0.01161f
C4615 sar9b_0.net22 sar9b_0.cyclic_flag_0.FINAL 0.02996f
C4616 sar9b_0.net58 a_5460_28377# 0.15559f
C4617 sar9b_0.net6 sar9b_0.net73 0.44042f
C4618 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.22879f
C4619 VDPWR sar9b_0._06_ 0.47072f
C4620 sar9b_0.net57 sar9b_0.net4 0.32464f
C4621 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.02632f
C4622 a_2739_20140# a_2918_20140# 0.54426f
C4623 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C4624 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.12898f
C4625 a_8266_17113# a_7602_16784# 0.16939f
C4626 sar9b_0.net2 a_9270_24566# 0.03939f
C4627 a_8334_17021# a_8052_16791# 0.05462f
C4628 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[6] 0.17948f
C4629 sar9b_0.net40 a_6132_23451# 0.01344f
C4630 single_9b_cdac_0.SW[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.15242f
C4631 sar9b_0.net70 sar9b_0.clknet_1_1__leaf_CLK 0.27895f
C4632 a_7882_19538# sar9b_0.net40 0.04062f
C4633 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[4] 0.01525f
C4634 sar9b_0.net24 a_9138_27163# 0.03746f
C4635 single_9b_cdac_1.cdac_sw_9b_0.S[2] a_53154_16877# 0.59531f
C4636 sar9b_0.net21 sar9b_0.net37 0.06888f
C4637 single_9b_cdac_0.cdac_sw_9b_0.S[4] ua[0] 1.93763f
C4638 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[7] 0.0313f
C4639 sar9b_0._01_ sar9b_0.net57 0.02763f
C4640 a_21684_3438# a_18214_3039# 0.11186f
C4641 sar9b_0.net37 sar9b_0.net39 0.18921f
C4642 a_7138_27758# a_8166_27595# 0.07826f
C4643 single_9b_cdac_1.SW[0] a_9974_17626# 0.0138f
C4644 VDPWR a_3545_26914# 0.22169f
C4645 VDPWR th_dif_sw_0.CKB 1.43024f
C4646 tdc_0.OUTN a_7743_16817# 0.05748f
C4647 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.69086f
C4648 a_3545_26914# a_4330_27170# 0.26257f
C4649 VDPWR a_11658_23470# 0.84308f
C4650 a_6307_27584# a_6678_27470# 0.04761f
C4651 VDPWR a_2451_27234# 0.27934f
C4652 sar9b_0.net5 a_7914_19178# 0.20518f
C4653 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.3601f
C4654 sar9b_0.net23 a_7692_26108# 0.27877f
C4655 a_64331_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.01076f
C4656 single_9b_cdac_0.cdac_sw_9b_0.S[7] ua[0] 1.97045f
C4657 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.02149f
C4658 a_8982_21902# sar9b_0.net37 0.02238f
C4659 sar9b_0.net44 sar9b_0.net19 0.14271f
C4660 a_12182_22423# a_12618_22138# 0.16939f
C4661 sar9b_0.net40 th_dif_sw_0.CK 0.08068f
C4662 sar9b_0.net4 a_5443_19074# 0.31469f
C4663 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 1.71649f
C4664 VDPWR a_16222_11316# 0.52162f
C4665 sar9b_0.net46 sar9b_0.net73 0.14249f
C4666 sar9b_0.net36 sar9b_0.net51 0.02568f
C4667 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C4668 VDPWR a_5633_20244# 0.10568f
C4669 sar9b_0.net50 sar9b_0.net73 0.28503f
C4670 single_9b_cdac_1.SW[3] sar9b_0.net73 0.09966f
C4671 a_9442_21474# a_10218_21842# 0.3578f
C4672 single_9b_cdac_0.cdac_sw_9b_0.S[1] ua[0] 1.18579f
C4673 a_11339_27039# sar9b_0.net31 0.19953f
C4674 a_2706_27440# a_2847_27473# 0.27388f
C4675 a_3156_27447# a_3161_27787# 0.44098f
C4676 sar9b_0.net11 clk 0.17325f
C4677 sar9b_0.net40 sar9b_0.net4 0.05476f
C4678 a_13011_27234# single_9b_cdac_0.SW[3] 0.01848f
C4679 sar9b_0._09_ a_4947_20140# 0.01531f
C4680 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.03729f
C4681 sar9b_0.net45 uo_out[6] 0.06932f
C4682 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.12431f
C4683 sar9b_0.net30 a_12064_22819# 0.2744f
C4684 single_9b_cdac_0.SW[6] th_dif_sw_0.VCN 0.09468f
C4685 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.6919f
C4686 a_11842_19766# a_12618_19474# 0.3578f
C4687 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.02632f
C4688 a_13011_25902# sar9b_0.net29 0.01649f
C4689 sar9b_0.net60 a_6282_27170# 0.04032f
C4690 a_11842_23762# a_12870_23599# 0.07826f
C4691 VDPWR a_11338_19178# 0.29105f
C4692 sar9b_0.net19 a_3822_27060# 0.0307f
C4693 sar9b_0.net52 sar9b_0.net33 0.30065f
C4694 ua[3] th_dif_sw_0.VCN 3.30291f
C4695 sar9b_0.net30 sar9b_0.net74 0.03698f
C4696 sar9b_0.net8 single_9b_cdac_1.CF[3] 0.02324f
C4697 sar9b_0.net40 a_12182_19759# 0.06762f
C4698 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.04988f
C4699 clk th_dif_sw_0.VCN 2.08719f
C4700 sar9b_0.net46 sar9b_0.net6 0.09629f
C4701 a_2892_27039# sar9b_0.net19 0.29845f
C4702 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.93403f
C4703 sar9b_0.net50 sar9b_0.net6 0.16111f
C4704 sar9b_0._06_ sar9b_0.net29 0.03732f
C4705 single_9b_cdac_1.SW[8] a_13216_19809# 0.01788f
C4706 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.42784f
C4707 single_9b_cdac_1.SW[3] sar9b_0.net6 0.2526f
C4708 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.26427f
C4709 th_dif_sw_0.CK a_12870_18271# 0.06999f
C4710 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 ua[0] 0.12088f
C4711 a_12618_18142# sar9b_0.net6 0.01945f
C4712 sar9b_0.net63 a_5100_24375# 0.0166f
C4713 a_10816_21487# sar9b_0.net36 0.02497f
C4714 VDPWR sar9b_0._04_ 0.59309f
C4715 a_7289_21127# a_8074_20870# 0.26257f
C4716 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.CF[7] 0.12358f
C4717 a_3521_24240# a_3369_24181# 0.22338f
C4718 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.42784f
C4719 sar9b_0.net47 sar9b_0.net39 0.20215f
C4720 sar9b_0._07_ sar9b_0.net39 0.04027f
C4721 VDPWR a_10742_25087# 0.19934f
C4722 VDPWR a_7188_22119# 0.85695f
C4723 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[6] 0.01475f
C4724 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.10626f
C4725 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VDPWR 0.84061f
C4726 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C4727 sar9b_0.net32 a_12560_27128# 0.01666f
C4728 a_10506_23174# a_10690_22806# 0.44098f
C4729 sar9b_0._11_ sar9b_0._07_ 0.03254f
C4730 a_10239_19235# sar9b_0.net49 0.02293f
C4731 sar9b_0.net43 a_6538_24506# 0.03826f
C4732 sar9b_0.net63 a_5484_23444# 0.04251f
C4733 a_4211_19474# sar9b_0.net46 0.02075f
C4734 a_5506_26802# a_6282_27170# 0.3578f
C4735 a_10859_26330# sar9b_0.net74 0.1037f
C4736 sar9b_0.net67 sar9b_0.net70 0.05082f
C4737 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.03729f
C4738 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.03433f
C4739 a_10402_27758# sar9b_0.net38 0.02612f
C4740 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.363f
C4741 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C4742 a_10402_27758# VDPWR 0.22246f
C4743 single_9b_cdac_1.SW[5] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 0.36301f
C4744 sar9b_0.net36 sar9b_0.net12 0.02707f
C4745 a_8098_23762# clk 0.01832f
C4746 a_9162_23174# sar9b_0.net11 0.06676f
C4747 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.84423f
C4748 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.10499f
C4749 a_8386_22806# sar9b_0.net54 0.10034f
C4750 a_3454_22567# sar9b_0._12_ 0.02006f
C4751 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[8] 0.80778f
C4752 sar9b_0.net59 sar9b_0.net39 0.21806f
C4753 sar9b_0.net61 a_8052_16791# 0.07136f
C4754 sar9b_0.net63 sar9b_0.net68 0.09062f
C4755 a_6678_27470# sar9b_0.net44 0.04249f
C4756 VDPWR th_dif_sw_0.th_sw_1.CKB 3.04581f
C4757 single_9b_cdac_0.SW[1] ua[0] 0.14864f
C4758 sar9b_0.net32 a_12182_23755# 0.01954f
C4759 a_10858_17113# single_9b_cdac_1.SW[2] 0.02538f
C4760 sar9b_0.net7 a_10607_21189# 0.06928f
C4761 sar9b_0.net56 a_8694_20570# 0.01417f
C4762 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62538f
C4763 VDPWR a_8303_18859# 0.2747f
C4764 a_6767_25185# a_6562_25094# 0.09983f
C4765 a_4136_25584# sar9b_0.clknet_1_1__leaf_CLK 0.10289f
C4766 single_9b_cdac_0.SW[8] clk 0.42402f
C4767 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.05472f
C4768 VDPWR single_9b_cdac_1.SW[0] 3.84179f
C4769 a_10762_18823# sar9b_0.net36 0.01606f
C4770 single_9b_cdac_1.CF[6] ua[0] 3.57763f
C4771 a_8098_18810# sar9b_0.net37 0.01309f
C4772 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.95338f
C4773 a_12618_18142# sar9b_0.net50 0.26153f
C4774 VDPWR sar9b_0.net56 1.95434f
C4775 a_12870_19603# single_9b_cdac_1.SW[8] 0.01567f
C4776 a_3521_24240# a_3014_24136# 0.21226f
C4777 a_4934_22432# sar9b_0.net60 0.03501f
C4778 a_10482_3438# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.63339f
C4779 sar9b_0.net57 sar9b_0.net55 0.02755f
C4780 a_4011_22488# sar9b_0.clknet_1_1__leaf_CLK 0.06293f
C4781 VDPWR a_11030_22954# 0.20335f
C4782 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96907f
C4783 sar9b_0.net28 single_9b_cdac_1.CF[0] 0.0432f
C4784 single_9b_cdac_1.cdac_sw_9b_0.S[6] ua[0] 1.67132f
C4785 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C4786 a_13011_27234# a_13216_26469# 0.01043f
C4787 sar9b_0.net40 a_5748_24381# 0.02394f
C4788 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[5] 0.02038f
C4789 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 ua[0] 0.12076f
C4790 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[0] 0.03931f
C4791 sar9b_0.net40 a_6282_27170# 0.0332f
C4792 single_9b_cdac_1.cdac_sw_9b_0.S[3] single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.51772f
C4793 sar9b_0.net56 sar9b_0.net1 0.26215f
C4794 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[7] 1.10355f
C4795 a_11466_23174# sar9b_0.net31 0.017f
C4796 sar9b_0.net58 sar9b_0.clk_div_0.COUNT\[2\] 0.06301f
C4797 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.19266f
C4798 a_10803_18142# sar9b_0.net38 0.20613f
C4799 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C4800 sar9b_0._06_ single_9b_cdac_0.SW[3] 0.08528f
C4801 VDPWR a_10803_18142# 0.46102f
C4802 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.02618f
C4803 VDPWR sar9b_0.net70 0.75523f
C4804 sar9b_0.net16 a_4496_20468# 0.03603f
C4805 sar9b_0.net42 sar9b_0.net27 0.03289f
C4806 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.33229f
C4807 VDPWR a_12684_20379# 0.21989f
C4808 a_11434_16874# tdc_0.OUTP 0.04839f
C4809 sar9b_0.net42 single_9b_cdac_0.SW[5] 0.01977f
C4810 single_9b_cdac_1.CF[5] single_9b_cdac_1.CF[7] 0.02364f
C4811 a_6252_19074# a_6579_18832# 0.09203f
C4812 VDPWR a_6902_25087# 0.2038f
C4813 a_7188_22119# a_6738_22112# 0.03529f
C4814 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_0.SW[7] 0.17509f
C4815 a_11338_19178# sar9b_0.net48 0.20192f
C4816 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.22526f
C4817 a_9935_24187# sar9b_0.net12 0.01643f
C4818 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.31534f
C4819 sar9b_0.net55 a_5443_19074# 0.03144f
C4820 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 2.71729f
C4821 single_9b_cdac_1.CF[3] single_9b_cdac_1.CF[0] 0.04014f
C4822 a_2508_23444# sar9b_0.clk_div_0.COUNT\[1\] 0.06012f
C4823 a_11859_20574# sar9b_0.net51 0.08706f
C4824 sar9b_0.net52 sar9b_0.net34 0.06265f
C4825 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.01751f
C4826 a_11859_17910# sar9b_0.net27 0.05667f
C4827 sar9b_0.net40 sar9b_0.net55 1.09485f
C4828 sar9b_0.net21 a_6880_26815# 0.2711f
C4829 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.19266f
C4830 VDPWR uo_out[2] 0.90561f
C4831 sar9b_0._14_ a_4044_24776# 0.04883f
C4832 a_2893_24992# a_2940_25096# 0.19021f
C4833 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 3.10626f
C4834 sar9b_0.net27 a_4771_18260# 0.02095f
C4835 a_11178_27466# a_11776_27801# 0.06623f
C4836 a_6414_23681# sar9b_0.net54 0.20382f
C4837 tdc_0.phase_detector_0.INN tdc_0.phase_detector_0.INP 1.21226f
C4838 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._04_ 0.01564f
C4839 sar9b_0.net9 a_7193_22459# 0.01552f
C4840 sar9b_0.net13 a_7936_25137# 0.0469f
C4841 a_10227_18142# a_9634_17478# 0.01011f
C4842 a_7097_19795# sar9b_0.net47 0.13999f
C4843 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.28575f
C4844 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36044f
C4845 sar9b_0.net32 a_10995_28566# 0.04889f
C4846 a_8074_20870# sar9b_0.net47 0.22159f
C4847 a_54032_26990# single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22367f
C4848 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.0174f
C4849 sar9b_0.net63 sar9b_0.net10 0.04452f
C4850 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[7] 6.82494f
C4851 a_8726_22954# sar9b_0.net37 0.01269f
C4852 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.03729f
C4853 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.05472f
C4854 a_7936_25137# sar9b_0.cyclic_flag_0.FINAL 0.26867f
C4855 th_dif_sw_0.CK a_10166_3438# 0.0136f
C4856 w_17430_1606# dw_17224_1400# 9.71413f
C4857 sar9b_0.net26 clk 0.04511f
C4858 single_9b_cdac_0.SW[7] clk 1.04996f
C4859 sar9b_0.net57 a_9165_24988# 0.05719f
C4860 a_8303_18859# sar9b_0.net48 0.22623f
C4861 sar9b_0.net10 sar9b_0.net62 0.15663f
C4862 sar9b_0.net48 single_9b_cdac_1.SW[0] 0.1553f
C4863 VDPWR a_3156_26115# 0.78981f
C4864 VDPWR a_5394_18116# 0.35368f
C4865 sar9b_0.net56 sar9b_0.net48 0.26514f
C4866 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 ua[0] 0.1236f
C4867 a_8202_23174# a_8726_22954# 0.04522f
C4868 a_7926_23234# a_8591_22855# 0.19065f
C4869 sar9b_0.net43 clk 0.04165f
C4870 a_13011_25902# a_13216_26469# 0.01179f
C4871 VDPWR a_10937_25582# 0.2119f
C4872 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.12431f
C4873 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C4874 VDPWR sar9b_0.net60 2.99913f
C4875 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62573f
C4876 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.0303f
C4877 a_25210_26990# single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.22352f
C4878 a_4947_20140# a_5126_20140# 0.54426f
C4879 VDPWR a_11146_25483# 0.19884f
C4880 sar9b_0.net20 a_5674_28147# 0.06614f
C4881 a_5748_24381# a_6538_24506# 0.1263f
C4882 single_9b_cdac_1.cdac_sw_9b_0.S[3] a_48343_16877# 0.59531f
C4883 a_6132_23451# clk 0.01117f
C4884 sar9b_0.net42 sar9b_0.net36 0.59867f
C4885 a_11466_23174# a_11718_23127# 0.27388f
C4886 a_6880_17491# sar9b_0.net46 0.03742f
C4887 a_5182_22567# sar9b_0._18_ 0.01534f
C4888 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[1] 17.5055f
C4889 sar9b_0.net32 sar9b_0.net12 0.03166f
C4890 a_13011_23238# clk 0.0315f
C4891 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS th_dif_sw_0.VCN 0.14643f
C4892 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 3.26837f
C4893 uo_out[5] ui_in[0] 0.06786f
C4894 uo_out[6] uo_out[7] 2.95271f
C4895 single_9b_cdac_0.SW[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.36412f
C4896 sar9b_0.net24 uo_out[2] 0.09027f
C4897 sar9b_0.net16 sar9b_0.net27 0.02393f
C4898 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 ua[0] 0.12088f
C4899 VDPWR sar9b_0.net57 1.46403f
C4900 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[5] 0.02008f
C4901 a_10230_23234# sar9b_0.net74 0.2089f
C4902 VDPWR a_5506_26802# 0.2219f
C4903 a_9472_18823# sar9b_0.net5 0.02035f
C4904 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07517f
C4905 a_5581_20992# sar9b_0._07_ 0.02281f
C4906 VDPWR tdc_0.phase_detector_0.pd_out_0.B 1.26944f
C4907 sar9b_0.net70 sar9b_0.clknet_1_0__leaf_CLK 0.28843f
C4908 single_9b_cdac_0.SW[1] sar9b_0.net27 0.088f
C4909 sar9b_0.net53 a_11842_22430# 0.09838f
C4910 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[5] 0.01299f
C4911 sar9b_0.net49 sar9b_0.net26 0.02489f
C4912 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 0.69086f
C4913 VDPWR a_4136_25584# 0.84755f
C4914 tdc_0.OUTN sar9b_0.net27 0.2611f
C4915 single_9b_cdac_1.CF[6] sar9b_0.net27 0.05684f
C4916 sar9b_0.net27 a_13216_22473# 0.01241f
C4917 single_9b_cdac_1.CF[6] single_9b_cdac_0.SW[5] 0.09395f
C4918 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.28523f
C4919 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 2.71729f
C4920 sar9b_0.net52 single_9b_cdac_0.SW[4] 0.35739f
C4921 VDPWR a_7404_17715# 0.22602f
C4922 VDPWR a_48343_26999# 1.81495f
C4923 VDPWR a_4011_22488# 0.08627f
C4924 a_4812_28371# a_5010_28495# 0.06623f
C4925 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.26707f
C4926 sar9b_0.net41 a_9634_17478# 0.06387f
C4927 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 1.71649f
C4928 sar9b_0.net36 a_10482_25831# 0.02816f
C4929 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 0.42014f
C4930 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.75815f
C4931 a_3747_25724# a_3855_25792# 0.29821f
C4932 sar9b_0.net55 a_6538_24506# 0.0859f
C4933 a_8052_16791# sar9b_0.net5 0.21543f
C4934 sar9b_0.net43 sar9b_0.net49 0.0215f
C4935 a_10402_25094# a_9942_24806# 0.26257f
C4936 sar9b_0.net4 clk 0.04636f
C4937 single_9b_cdac_1.SW[5] single_9b_cdac_1.CF[7] 0.01475f
C4938 sar9b_0.net27 a_12618_23470# 0.02584f
C4939 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP a_48343_26999# 0.04592f
C4940 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C4941 a_16357_9613# th_dif_sw_0.VCN 0.10892f
C4942 sar9b_0.net41 sar9b_0.net11 0.07372f
C4943 a_7404_17715# sar9b_0.net1 0.27002f
C4944 sar9b_0._11_ a_4496_20468# 0.09559f
C4945 sar9b_0.net49 a_10035_19474# 0.26854f
C4946 VDPWR a_53154_26999# 1.81495f
C4947 a_10470_21795# a_9258_21842# 0.07766f
C4948 VDPWR a_5443_19074# 0.34039f
C4949 sar9b_0.net45 single_9b_cdac_0.SW[8] 0.08609f
C4950 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.05472f
C4951 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C4952 single_9b_cdac_1.CF[1] ua[0] 3.57763f
C4953 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.3196f
C4954 a_7638_23474# sar9b_0.net54 0.09716f
C4955 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C4956 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.03729f
C4957 tdc_0.OUTP sar9b_0.net6 0.49725f
C4958 sar9b_0.net60 sar9b_0._17_ 0.04099f
C4959 sar9b_0.net40 sar9b_0.net38 0.028f
C4960 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C4961 VDPWR sar9b_0.net40 1.99954f
C4962 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.0313f
C4963 sar9b_0.net30 sar9b_0.net53 0.04133f
C4964 a_5441_22522# sar9b_0.net60 0.01343f
C4965 a_4467_24162# sar9b_0.clk_div_0.COUNT\[2\] 0.16437f
C4966 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C4967 sar9b_0.net8 sar9b_0.net2 0.02074f
C4968 sar9b_0.net48 a_5394_18116# 0.26617f
C4969 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.42784f
C4970 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 ua[0] 0.13461f
C4971 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.06019f
C4972 sar9b_0._04_ sar9b_0._12_ 0.12021f
C4973 sar9b_0.net54 a_5962_24151# 0.14491f
C4974 a_24332_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.23864f
C4975 sar9b_0.net40 sar9b_0.net1 0.0276f
C4976 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.71729f
C4977 single_9b_cdac_1.CF[7] ua[0] 3.57763f
C4978 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.70254f
C4979 a_13011_21906# a_13216_22473# 0.01179f
C4980 sar9b_0._08_ sar9b_0.net60 0.18449f
C4981 a_11658_18142# sar9b_0.net50 0.17638f
C4982 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.42784f
C4983 VDPWR a_9174_17906# 0.28468f
C4984 single_9b_cdac_1.SW[3] a_11658_18142# 0.02689f
C4985 sar9b_0.net57 sar9b_0._17_ 0.02056f
C4986 a_11658_18142# a_12618_18142# 0.03432f
C4987 a_8115_28566# sar9b_0.net22 0.0346f
C4988 a_4083_28566# sar9b_0.net60 0.05402f
C4989 single_9b_cdac_1.SW[2] sar9b_0.net37 0.07696f
C4990 a_3161_26455# a_3156_26115# 0.44098f
C4991 VDPWR a_6861_22828# 0.14773f
C4992 a_10830_19068# sar9b_0.net7 0.01607f
C4993 sar9b_0.net49 th_dif_sw_0.CK 0.01033f
C4994 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 0.69086f
C4995 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.69086f
C4996 a_10218_27466# a_10995_28566# 0.01498f
C4997 a_7374_19685# sar9b_0.net10 0.04605f
C4998 sar9b_0.net60 a_5682_23444# 0.04812f
C4999 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A 0.11216f
C5000 a_7638_19238# sar9b_0.net51 0.03553f
C5001 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VDPWR 3.27795f
C5002 a_5439_24563# sar9b_0.net54 0.16847f
C5003 a_7590_24931# a_7338_24802# 0.27388f
C5004 a_7092_19455# sar9b_0.net10 0.25701f
C5005 sar9b_0.net38 a_9588_27045# 0.02021f
C5006 sar9b_0.net60 sar9b_0.clknet_1_0__leaf_CLK 0.04105f
C5007 tdc_0.OUTP single_9b_cdac_1.SW[3] 0.04678f
C5008 sar9b_0._08_ sar9b_0.net57 0.62749f
C5009 a_11466_23174# sar9b_0.net10 0.05039f
C5010 sar9b_0.net31 sar9b_0.net11 0.38707f
C5011 VDPWR a_9588_27045# 0.85382f
C5012 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 0.8438f
C5013 a_7566_21017# sar9b_0.net51 0.02936f
C5014 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02652f
C5015 a_8303_23853# sar9b_0.net54 0.0633f
C5016 a_9279_27227# sar9b_0.net37 0.07713f
C5017 VDPWR a_12870_18271# 0.27198f
C5018 sar9b_0.net36 sar9b_0.net74 0.21507f
C5019 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0.clk_div_0.COUNT\[1\] 0.12709f
C5020 a_11776_21141# sar9b_0.net39 0.01141f
C5021 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.06503f
C5022 a_7914_27466# sar9b_0.net36 0.06473f
C5023 VDPWR a_16331_9671# 0.67026f
C5024 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[4] 0.02005f
C5025 a_6954_27466# sar9b_0.net60 0.16181f
C5026 sar9b_0.net57 a_5682_23444# 0.06802f
C5027 a_11658_19474# a_12182_19759# 0.05022f
C5028 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C5029 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 0.3601f
C5030 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.38397f
C5031 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[4] 0.02215f
C5032 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.75853f
C5033 sar9b_0.net18 a_3161_27787# 0.01348f
C5034 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C5035 sar9b_0.net4 a_5849_18463# 0.01533f
C5036 dw_12589_1395# w_12795_1601# 9.86148f
C5037 single_9b_cdac_0.SW[5] a_13164_28398# 0.01688f
C5038 VDPWR uio_out[1] 1.23314f
C5039 a_40321_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.01076f
C5040 uio_in[6] uio_in[5] 0.03102f
C5041 sar9b_0.net35 sar9b_0.net58 0.03409f
C5042 sar9b_0.net40 sar9b_0._17_ 0.02904f
C5043 a_3371_23106# sar9b_0.clk_div_0.COUNT\[2\] 0.10533f
C5044 a_6738_22112# sar9b_0.net40 0.02168f
C5045 a_9414_23127# a_9760_22819# 0.07649f
C5046 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.24779f
C5047 a_9359_20191# sar9b_0.net51 0.07207f
C5048 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[4] 0.42014f
C5049 single_9b_cdac_0.SW[7] sar9b_0.net45 0.21976f
C5050 sar9b_0.net9 sar9b_0.net37 0.08996f
C5051 sar9b_0.net36 a_10506_24506# 0.0206f
C5052 a_3695_23038# sar9b_0.clk_div_0.COUNT\[1\] 0.07641f
C5053 a_8622_26345# sar9b_0.net37 0.01006f
C5054 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.26709f
C5055 a_9363_20826# sar9b_0.net8 0.03842f
C5056 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[2] 0.01297f
C5057 sar9b_0.net70 sar9b_0._12_ 0.02802f
C5058 sar9b_0.net52 a_11382_26138# 0.24197f
C5059 a_5235_27466# a_5322_27170# 0.01145f
C5060 sar9b_0.net64 a_5182_22567# 0.12016f
C5061 a_55773_29911# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C5062 sar9b_0.net58 sar9b_0._14_ 0.12417f
C5063 a_3438_26345# a_3946_26198# 0.19065f
C5064 sar9b_0.net61 sar9b_0.net37 0.52176f
C5065 sar9b_0.net44 sar9b_0.net37 0.76756f
C5066 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_1.CF[8] 0.01879f
C5067 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[7] 0.06912f
C5068 sar9b_0.net23 a_9939_28566# 0.20828f
C5069 a_6861_22828# sar9b_0._17_ 0.01915f
C5070 sar9b_0.net43 sar9b_0.net45 0.12328f
C5071 a_4125_25958# a_4293_25852# 0.27693f
C5072 sar9b_0.net40 sar9b_0.net48 0.10648f
C5073 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.19266f
C5074 sar9b_0.net58 a_5742_28392# 0.19468f
C5075 a_3922_20239# sar9b_0.net16 0.1201f
C5076 a_8019_17910# a_8052_16791# 0.03036f
C5077 a_10662_17799# a_9634_17478# 0.07826f
C5078 a_2918_20140# sar9b_0._00_ 0.27567f
C5079 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.84082f
C5080 sar9b_0.net2 a_9730_24138# 0.07985f
C5081 a_8842_16874# a_8052_16791# 0.1263f
C5082 a_8266_17113# a_8057_17131# 0.24088f
C5083 VDPWR a_6538_24506# 0.27686f
C5084 a_3371_23106# a_3695_23038# 0.15159f
C5085 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C5086 sar9b_0.net42 sar9b_0.net51 0.01622f
C5087 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[6] 1.94202f
C5088 th_dif_sw_0.VCP ua[0] 1.04697f
C5089 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[5] 0.19147f
C5090 single_9b_cdac_0.SW[2] ua[0] 0.15413f
C5091 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.07579f
C5092 a_8052_18123# a_7914_19178# 0.26288f
C5093 a_8202_23174# sar9b_0.net61 0.01019f
C5094 VDPWR a_13011_17910# 0.46728f
C5095 a_12618_19474# a_13216_19809# 0.06623f
C5096 sar9b_0.net48 a_9174_17906# 0.2009f
C5097 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[4] 0.28813f
C5098 sar9b_0.net55 clk 0.03649f
C5099 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C5100 sar9b_0.net22 uo_out[4] 0.11108f
C5101 a_5849_18463# a_6126_18353# 0.09983f
C5102 a_21368_4076# VDPWR 0.07949f
C5103 sar9b_0.net40 a_12047_19857# 0.04975f
C5104 a_7478_27751# a_7914_27466# 0.16939f
C5105 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C5106 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.07517f
C5107 single_9b_cdac_1.SW[3] single_9b_cdac_1.CF[3] 1.84733f
C5108 sar9b_0.net52 a_10218_24802# 0.16549f
C5109 a_10227_18142# th_dif_sw_0.CK 0.35616f
C5110 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.22875f
C5111 VDPWR a_3090_27163# 0.37894f
C5112 single_9b_cdac_0.SW[3] a_48343_26999# 0.28324f
C5113 a_5010_28495# uo_out[7] 0.02505f
C5114 sar9b_0.net43 a_9870_27060# 0.01268f
C5115 a_5484_23444# sar9b_0.net11 0.29424f
C5116 VDPWR a_9647_21523# 0.27298f
C5117 VDPWR a_3156_27447# 0.84513f
C5118 sar9b_0.net59 a_9279_27227# 0.1788f
C5119 a_9442_21474# sar9b_0.net37 0.01287f
C5120 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.28523f
C5121 a_12182_22423# a_12047_22521# 0.35559f
C5122 a_12870_22267# a_13216_22473# 0.07649f
C5123 sar9b_0.net4 a_6252_19074# 0.05708f
C5124 VDPWR a_16527_10454# 0.3789f
C5125 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C5126 a_3922_20239# a_3723_20140# 0.29821f
C5127 single_9b_cdac_1.CF[1] sar9b_0.net27 0.07881f
C5128 sar9b_0.net53 sar9b_0.net54 0.39148f
C5129 a_11718_23127# sar9b_0.net11 0.03005f
C5130 a_9730_24138# a_10758_24459# 0.07826f
C5131 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.42509f
C5132 a_10803_19474# single_9b_cdac_1.SW[1] 0.35106f
C5133 a_9782_21622# a_10218_21842# 0.16939f
C5134 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] 3.10218f
C5135 a_5151_28559# a_5465_28246# 0.07826f
C5136 single_9b_cdac_1.CF[2] sar9b_0.net28 0.04267f
C5137 a_9647_21523# sar9b_0.net1 0.02115f
C5138 a_2835_24136# sar9b_0.clk_div_0.COUNT\[1\] 0.02455f
C5139 sar9b_0.net60 a_5523_21528# 0.24769f
C5140 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 0.42015f
C5141 a_2847_27473# a_3161_27787# 0.07826f
C5142 a_3156_27447# a_3370_27769# 0.04522f
C5143 sar9b_0.net9 sar9b_0.net47 0.32405f
C5144 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[0] 0.26707f
C5145 sar9b_0.net41 sar9b_0.net26 0.02726f
C5146 sar9b_0._09_ sar9b_0._10_ 0.14294f
C5147 sar9b_0.net36 a_7343_27849# 0.04959f
C5148 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38317f
C5149 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02666f
C5150 sar9b_0.net47 sar9b_0.net61 0.15705f
C5151 sar9b_0.net63 a_6744_23238# 0.07362f
C5152 sar9b_0.net36 sar9b_0.net21 0.02863f
C5153 single_9b_cdac_1.CF[7] sar9b_0.net27 0.14896f
C5154 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C5155 sar9b_0.net60 a_6030_24396# 0.02375f
C5156 sar9b_0.net60 sar9b_0._12_ 0.23194f
C5157 a_12870_19603# a_12618_19474# 0.27388f
C5158 single_9b_cdac_0.SW[4] a_13011_27234# 0.05684f
C5159 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A 0.84042f
C5160 single_9b_cdac_1.CF[7] single_9b_cdac_0.SW[5] 0.02016f
C5161 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 2.7611f
C5162 sar9b_0.net31 a_11658_26134# 0.02303f
C5163 a_2828_22432# sar9b_0._05_ 0.01634f
C5164 sar9b_0.net43 sar9b_0.net41 0.34712f
C5165 sar9b_0.net13 a_5753_24250# 0.07055f
C5166 a_12182_23755# a_12618_23470# 0.16939f
C5167 sar9b_0.net36 sar9b_0.net39 0.02403f
C5168 sar9b_0.net42 sar9b_0.net12 0.02691f
C5169 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C5170 a_13011_24802# sar9b_0.net26 0.22283f
C5171 sar9b_0.net54 a_6562_25094# 0.07487f
C5172 a_8622_26345# sar9b_0.net59 0.24081f
C5173 sar9b_0.net41 a_10035_19474# 0.02751f
C5174 a_25210_26990# single_9b_cdac_0.SW[8] 0.18991f
C5175 VDPWR a_10166_3438# 0.07956f
C5176 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.22875f
C5177 a_3231_27227# sar9b_0.net19 0.04509f
C5178 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[8] 0.058f
C5179 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.17717f
C5180 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C5181 sar9b_0.net58 a_3946_27530# 0.24636f
C5182 a_12047_18525# sar9b_0.net6 0.01853f
C5183 sar9b_0.net59 sar9b_0.net44 0.32798f
C5184 single_9b_cdac_1.CF[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.26707f
C5185 sar9b_0.net63 sar9b_0._13_ 0.05991f
C5186 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[6] 0.02343f
C5187 single_9b_cdac_1.CF[3] single_9b_cdac_1.CF[2] 14.3503f
C5188 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.SW[3] 0.01382f
C5189 a_3521_24240# a_3819_24136# 0.02614f
C5190 sar9b_0.net57 sar9b_0._12_ 0.01983f
C5191 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C5192 single_9b_cdac_1.CF[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.0313f
C5193 sar9b_0.net18 sar9b_0.net3 0.04914f
C5194 VDPWR a_11178_24802# 0.33967f
C5195 a_10230_23234# sar9b_0.net53 0.22171f
C5196 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.01751f
C5197 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VDPWR 3.27795f
C5198 sar9b_0.net16 a_5581_19664# 0.01792f
C5199 a_10506_23174# a_11030_22954# 0.04522f
C5200 a_10230_23234# a_10895_22855# 0.19065f
C5201 sar9b_0.clk_div_0.COUNT\[3\] a_4236_21738# 0.02104f
C5202 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95338f
C5203 a_11842_26426# a_12182_26419# 0.24088f
C5204 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A 0.0303f
C5205 a_5846_26950# a_6282_27170# 0.16939f
C5206 sar9b_0.net30 a_12047_23853# 0.03166f
C5207 sar9b_0.net53 sar9b_0.net27 0.03024f
C5208 sar9b_0.net20 uo_out[6] 0.34847f
C5209 single_9b_cdac_0.cdac_sw_9b_0.S[6] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24779f
C5210 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.26625f
C5211 sar9b_0.net32 single_9b_cdac_1.CF[6] 0.03698f
C5212 a_5083_21100# sar9b_0._18_ 0.10881f
C5213 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN 2.82223f
C5214 sar9b_0.net20 a_8115_28566# 0.21703f
C5215 sar9b_0.net56 a_9942_20810# 0.04264f
C5216 a_11430_27595# VDPWR 0.26904f
C5217 single_9b_cdac_0.SW[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.36512f
C5218 sar9b_0.net31 sar9b_0.net26 0.03062f
C5219 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.42784f
C5220 single_9b_cdac_0.cdac_sw_9b_0.S[4] a_43540_26999# 0.59531f
C5221 sar9b_0._09_ sar9b_0._01_ 0.03554f
C5222 a_9760_22819# sar9b_0.net11 0.04919f
C5223 a_8726_22954# sar9b_0.net54 0.14f
C5224 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[2] 0.22004f
C5225 a_4011_22488# sar9b_0._12_ 0.04991f
C5226 VDPWR a_4018_24235# 0.3802f
C5227 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.38397f
C5228 single_9b_cdac_0.SW[6] a_34814_26990# 0.18991f
C5229 sar9b_0._07_ a_5481_20185# 0.02028f
C5230 sar9b_0.net58 a_3545_26914# 0.10032f
C5231 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.17533f
C5232 sar9b_0.net32 a_12618_23470# 0.0684f
C5233 a_4293_25852# sar9b_0.clknet_1_1__leaf_CLK 0.04421f
C5234 sar9b_0.net63 sar9b_0.net69 0.04307f
C5235 a_12047_18525# sar9b_0.net50 0.22675f
C5236 VDPWR a_7306_19777# 0.20423f
C5237 single_9b_cdac_0.SW[6] sar9b_0.net38 0.16268f
C5238 single_9b_cdac_1.SW[3] a_12047_18525# 0.01367f
C5239 sar9b_0.net49 a_10742_21091# 0.13511f
C5240 a_7478_27751# a_7343_27849# 0.35559f
C5241 a_2547_28132# a_2931_28566# 0.09678f
C5242 single_9b_cdac_0.SW[6] VDPWR 2.34024f
C5243 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0.clknet_1_1__leaf_CLK 0.04637f
C5244 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN 2.82223f
C5245 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[4] 0.02164f
C5246 sar9b_0.net38 clk 0.04449f
C5247 VDPWR ua[3] 1.80857f
C5248 sar9b_0.net10 sar9b_0.net11 0.2401f
C5249 VDPWR clk 4.0924f
C5250 a_10858_17113# single_9b_cdac_1.SW[1] 0.01467f
C5251 single_9b_cdac_1.SW[2] ua[0] 0.14772f
C5252 a_10402_25094# sar9b_0.net36 0.0133f
C5253 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[8] 0.04036f
C5254 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.84427f
C5255 sar9b_0.net56 sar9b_0.net8 0.13034f
C5256 sar9b_0._09_ a_3795_19512# 0.09292f
C5257 a_9154_20142# a_9494_20290# 0.24088f
C5258 sar9b_0.net1 clk 0.04871f
C5259 a_4467_24162# sar9b_0._14_ 0.11012f
C5260 VDPWR a_10254_2858# 0.51112f
C5261 sar9b_0.net22 single_9b_cdac_0.SW[8] 0.02541f
C5262 sar9b_0._09_ a_3180_19448# 0.26014f
C5263 sar9b_0.net66 sar9b_0._05_ 0.18138f
C5264 sar9b_0.clk_div_0.COUNT\[2\] sar9b_0._03_ 0.03884f
C5265 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C5266 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62538f
C5267 sar9b_0.clknet_0_CLK sar9b_0.clk_div_0.COUNT\[0\] 0.86907f
C5268 single_9b_cdac_0.SW[2] sar9b_0.net27 0.06976f
C5269 single_9b_cdac_1.CF[4] single_9b_cdac_1.CF[7] 0.02091f
C5270 sar9b_0.net59 a_4749_27652# 0.27144f
C5271 single_9b_cdac_0.SW[2] single_9b_cdac_0.SW[5] 0.02056f
C5272 a_12435_24802# sar9b_0.net26 0.09225f
C5273 sar9b_0.net5 sar9b_0.net37 0.14722f
C5274 a_6250_28502# uo_out[6] 0.02897f
C5275 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.04988f
C5276 a_2508_23444# sar9b_0.clk_div_0.COUNT\[2\] 0.03301f
C5277 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.12367f
C5278 sar9b_0.net52 a_10284_25707# 0.02758f
C5279 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C5280 sar9b_0.net31 a_11382_22142# 0.03867f
C5281 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP ua[0] 1.1512f
C5282 single_9b_cdac_0.SW[4] sar9b_0._06_ 0.22289f
C5283 single_9b_cdac_1.CF[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.06503f
C5284 sar9b_0.net55 a_6252_19074# 0.17527f
C5285 m2_23774_17236# a_24332_16877# 0.01541f
C5286 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP a_33936_16877# 0.04592f
C5287 sar9b_0.net38 a_7539_28566# 0.05709f
C5288 a_10402_27758# sar9b_0.net34 0.01319f
C5289 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C5290 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C5291 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.03488f
C5292 VDPWR a_7539_28566# 0.41703f
C5293 sar9b_0.net35 sar9b_0.clk_div_0.COUNT\[1\] 0.03758f
C5294 sar9b_0.net74 sar9b_0.net12 0.05557f
C5295 a_11658_23470# a_11842_23762# 0.44532f
C5296 sar9b_0.net26 a_12435_20806# 0.0353f
C5297 sar9b_0.net35 sar9b_0.net73 0.26229f
C5298 single_9b_cdac_1.SW[8] ua[0] 0.13942f
C5299 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 0.6919f
C5300 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.28523f
C5301 a_10194_16784# a_9450_17846# 0.01861f
C5302 VDPWR a_6636_20780# 0.20851f
C5303 sar9b_0.net36 sar9b_0.net53 0.06691f
C5304 a_10895_22855# sar9b_0.net36 0.01323f
C5305 sar9b_0.net49 a_8694_20570# 0.22589f
C5306 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.SW[5] 0.244f
C5307 sar9b_0.net2 sar9b_0.net73 0.03106f
C5308 a_33936_16877# single_9b_cdac_1.SW[6] 0.28324f
C5309 a_3561_22527# a_3027_22138# 0.35097f
C5310 VDPWR a_11658_19474# 0.84186f
C5311 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 ua[0] 0.13178f
C5312 a_8266_18445# sar9b_0.net73 0.05509f
C5313 sar9b_0.net46 a_5196_18116# 0.01474f
C5314 a_11382_18146# sar9b_0.net39 0.01041f
C5315 sar9b_0.net49 sar9b_0.net38 0.54905f
C5316 sar9b_0._14_ sar9b_0.clk_div_0.COUNT\[1\] 0.03517f
C5317 sar9b_0.net13 a_6767_25185# 0.07236f
C5318 a_3713_22522# sar9b_0.net65 0.02109f
C5319 VDPWR tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.45583f
C5320 a_10742_27751# sar9b_0.net59 0.14619f
C5321 VDPWR sar9b_0.net49 2.96485f
C5322 VDPWR a_9162_23174# 0.37599f
C5323 sar9b_0.net43 a_5100_24375# 0.27992f
C5324 sar9b_0.net10 a_7443_21496# 0.02366f
C5325 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07517f
C5326 a_5100_24375# a_5298_24499# 0.06623f
C5327 a_6879_22145# a_7193_22459# 0.07826f
C5328 sar9b_0._17_ clk 0.03014f
C5329 sar9b_0.net49 sar9b_0.net1 0.10608f
C5330 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A 0.28523f
C5331 a_8266_17113# sar9b_0.net6 0.01365f
C5332 sar9b_0.net1 a_9162_23174# 0.01832f
C5333 m2_23774_17236# single_9b_cdac_1.cdac_sw_9b_0.S[8] 0.58106f
C5334 sar9b_0.net35 sar9b_0.net6 0.53411f
C5335 sar9b_0._13_ a_4811_23656# 0.11957f
C5336 single_9b_cdac_0.cdac_sw_9b_0.S[2] ua[0] 1.2071f
C5337 a_10239_19235# a_10548_19053# 0.07766f
C5338 sar9b_0.net29 clk 0.03602f
C5339 uio_in[1] uio_in[0] 0.03102f
C5340 a_8874_19178# a_9126_19131# 0.27388f
C5341 VDPWR a_2847_26141# 0.31739f
C5342 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5343 VDPWR a_5849_18463# 0.21922f
C5344 a_7193_22459# sar9b_0.net62 0.02169f
C5345 a_9634_17478# a_9839_17527# 0.09983f
C5346 a_9450_17846# a_10410_17846# 0.03493f
C5347 sar9b_0.net2 sar9b_0.net6 0.19883f
C5348 single_9b_cdac_1.SW[2] a_10410_17846# 0.06269f
C5349 a_4811_23656# a_5002_23764# 0.01358f
C5350 a_5506_17478# a_5711_17527# 0.09983f
C5351 a_11915_28371# a_12531_28566# 0.03551f
C5352 a_6282_17846# sar9b_0.net56 0.06691f
C5353 a_7402_22441# sar9b_0.net39 0.03886f
C5354 sar9b_0.net51 sar9b_0.net39 0.01895f
C5355 a_5126_20140# sar9b_0._10_ 0.06232f
C5356 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[4] 1.64863f
C5357 a_6030_24396# a_6538_24506# 0.19065f
C5358 sar9b_0.net13 sar9b_0.net37 0.03945f
C5359 a_5682_23444# clk 0.01117f
C5360 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.03488f
C5361 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 2.81428f
C5362 single_9b_cdac_1.CF[0] single_9b_cdac_1.SW[0] 1.83507f
C5363 a_9935_24187# sar9b_0.net53 0.2035f
C5364 a_8334_17021# sar9b_0.net27 0.06035f
C5365 a_10830_19068# single_9b_cdac_1.SW[1] 0.01619f
C5366 sar9b_0.net42 a_10482_25831# 0.02488f
C5367 sar9b_0.cyclic_flag_0.FINAL sar9b_0.net37 0.17246f
C5368 a_8266_17113# sar9b_0.net46 0.13705f
C5369 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.3186f
C5370 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[4] 0.01997f
C5371 sar9b_0.net35 sar9b_0.net46 0.32715f
C5372 single_9b_cdac_1.cdac_sw_9b_0.S[2] th_dif_sw_0.VCP 54.8348f
C5373 a_17125_9355# th_dif_sw_0.VCP 0.05474f
C5374 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VDPWR 0.38397f
C5375 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[1] 0.0147f
C5376 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.7611f
C5377 VDPWR a_5846_26950# 0.20642f
C5378 sar9b_0.net26 a_11842_19766# 0.02027f
C5379 clk rst_n 0.03102f
C5380 sar9b_0.net28 single_9b_cdac_1.SW[7] 0.0883f
C5381 a_5100_24375# sar9b_0._15_ 0.06016f
C5382 a_5711_26851# sar9b_0.net37 0.0259f
C5383 a_2835_24136# a_2508_23444# 0.01422f
C5384 sar9b_0.net53 a_12870_22267# 0.17311f
C5385 a_8266_18445# sar9b_0.net46 0.14299f
C5386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 a_34814_26990# 0.14695f
C5387 a_11466_23174# a_11658_22138# 0.01821f
C5388 sar9b_0.net59 a_10607_27849# 0.21965f
C5389 VDPWR a_4293_25852# 0.10504f
C5390 sar9b_0.net2 single_9b_cdac_1.SW[3] 0.19941f
C5391 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C5392 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.25152f
C5393 a_5812_21028# sar9b_0._11_ 0.06033f
C5394 a_6867_16810# a_7404_16784# 0.01177f
C5395 a_5506_17478# sar9b_0.net4 0.03413f
C5396 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.19266f
C5397 a_43540_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.23864f
C5398 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 a_25210_17740# 0.14695f
C5399 sar9b_0.net8 sar9b_0.net57 0.16844f
C5400 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_1.CF[8] 0.26707f
C5401 VDPWR a_8595_17910# 0.49252f
C5402 a_11842_18434# sar9b_0.net6 0.02355f
C5403 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[5] 0.01482f
C5404 sar9b_0.net63 sar9b_0.net72 0.26712f
C5405 single_9b_cdac_1.CF[8] single_9b_cdac_1.CF[7] 3.85504f
C5406 VDPWR sar9b_0.clk_div_0.COUNT\[3\] 0.34467f
C5407 a_5010_28495# sar9b_0.net20 0.08006f
C5408 a_8019_17910# sar9b_0.net37 0.20475f
C5409 sar9b_0.net57 a_7926_23234# 0.01631f
C5410 sar9b_0.net53 a_12182_23755# 0.14448f
C5411 a_7602_18116# sar9b_0.net5 0.04179f
C5412 sar9b_0.net41 a_9974_17626# 0.06988f
C5413 VDPWR a_9996_16784# 0.1892f
C5414 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[3] 0.026f
C5415 a_10218_20806# a_10742_21091# 0.05022f
C5416 a_3855_25792# a_4125_25958# 0.08669f
C5417 sar9b_0._16_ sar9b_0.clk_div_0.COUNT\[1\] 0.1686f
C5418 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.71729f
C5419 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[5] 4.15352f
C5420 single_9b_cdac_1.cdac_sw_9b_0.S[4] th_dif_sw_0.VCP 13.5521f
C5421 a_10284_25707# a_10623_25895# 0.07649f
C5422 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.71729f
C5423 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.69086f
C5424 sar9b_0.net61 a_10410_17846# 0.05361f
C5425 single_9b_cdac_1.CF[3] sar9b_0.net28 0.03461f
C5426 sar9b_0.net27 single_9b_cdac_1.SW[2] 0.12181f
C5427 sar9b_0._01_ a_5126_20140# 0.2535f
C5428 sar9b_0.net49 sar9b_0.net48 0.59286f
C5429 VDPWR a_6252_19074# 0.21971f
C5430 single_9b_cdac_0.SW[3] clk 0.13418f
C5431 a_10227_18142# sar9b_0.net38 0.06078f
C5432 a_5506_17478# a_5046_17906# 0.26257f
C5433 a_5711_17527# a_5322_17846# 0.05462f
C5434 a_11658_26134# a_12182_26419# 0.05022f
C5435 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.SW[7] 0.17154f
C5436 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0.net39 0.07149f
C5437 sar9b_0.net32 single_9b_cdac_1.CF[7] 0.01485f
C5438 VDPWR a_10227_18142# 0.43915f
C5439 a_2508_20780# sar9b_0.clknet_0_CLK 0.47881f
C5440 sar9b_0.net49 a_9900_19047# 0.01024f
C5441 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.05472f
C5442 a_6954_27466# a_7539_28566# 0.03399f
C5443 a_8842_18206# sar9b_0.net37 0.01698f
C5444 a_6922_23534# sar9b_0.net54 0.26015f
C5445 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.07579f
C5446 a_12684_20379# a_13011_20574# 0.08132f
C5447 a_9132_7271# th_dif_sw_0.th_sw_1.CK 2.28032f
C5448 sar9b_0.net26 sar9b_0.net10 0.0815f
C5449 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.S[5] 0.27713f
C5450 a_5196_24776# sar9b_0.net39 0.03191f
C5451 sar9b_0.net38 sar9b_0.net45 0.14791f
C5452 a_11658_19474# a_12047_19857# 0.06034f
C5453 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.95338f
C5454 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5455 VDPWR sar9b_0.net45 1.95717f
C5456 sar9b_0.net58 a_3156_26115# 0.01128f
C5457 uo_out[3] uo_out[2] 3.18986f
C5458 sar9b_0.net59 a_2706_26108# 0.26567f
C5459 sar9b_0.net48 a_5849_18463# 0.10592f
C5460 VDPWR th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.17946f
C5461 a_6102_24806# sar9b_0.net4 0.02847f
C5462 sar9b_0.net42 sar9b_0.net74 0.61827f
C5463 sar9b_0.net43 sar9b_0.net10 0.02603f
C5464 a_5580_24776# sar9b_0._15_ 0.26726f
C5465 a_11842_18434# sar9b_0.net50 0.09528f
C5466 sar9b_0.net47 sar9b_0.net15 0.02183f
C5467 single_9b_cdac_1.SW[3] a_11842_18434# 0.10099f
C5468 sar9b_0.net58 sar9b_0.net60 0.88421f
C5469 sar9b_0.net8 sar9b_0.net40 0.02953f
C5470 a_11658_18142# a_12047_18525# 0.06034f
C5471 a_11842_18434# a_12618_18142# 0.3578f
C5472 sar9b_0.net27 single_9b_cdac_1.SW[8] 0.0444f
C5473 sar9b_0.net32 sar9b_0.net53 0.15479f
C5474 sar9b_0.net17 a_2451_27234# 0.0211f
C5475 a_11722_25838# sar9b_0.net52 0.22698f
C5476 a_3161_26455# a_2847_26141# 0.07826f
C5477 a_3370_26437# a_3156_26115# 0.04522f
C5478 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[5] 0.31534f
C5479 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.6919f
C5480 a_6783_19481# a_6444_19448# 0.07649f
C5481 sar9b_0.net23 sar9b_0.net37 0.02446f
C5482 a_7882_19538# sar9b_0.net10 0.05509f
C5483 a_11436_17742# sar9b_0.net2 0.28173f
C5484 sar9b_0.net60 a_6137_23791# 0.02305f
C5485 a_8098_18810# sar9b_0.net51 0.0158f
C5486 a_5322_17846# sar9b_0.net4 0.02133f
C5487 a_5289_22527# sar9b_0.net39 0.0302f
C5488 a_7338_24802# a_7936_25137# 0.06623f
C5489 sar9b_0.net9 a_10230_23234# 0.03894f
C5490 a_13011_23238# sar9b_0.net10 0.22279f
C5491 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.02666f
C5492 sar9b_0.net59 sar9b_0.cyclic_flag_0.FINAL 0.74539f
C5493 a_7097_19795# sar9b_0.net51 0.02536f
C5494 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[6] 0.0313f
C5495 sar9b_0.net9 sar9b_0.net27 0.03863f
C5496 a_5322_27170# a_5506_26802# 0.43491f
C5497 VDPWR a_9870_27060# 0.26408f
C5498 a_8074_20870# sar9b_0.net51 0.06285f
C5499 a_10182_20463# sar9b_0.net5 0.04725f
C5500 VDPWR sar9b_0._09_ 0.86773f
C5501 sar9b_0.net38 a_10218_20806# 0.01292f
C5502 sar9b_0.net42 a_10506_24506# 0.01765f
C5503 sar9b_0.net58 a_5506_26802# 0.08623f
C5504 VDPWR a_4812_28371# 0.19653f
C5505 a_8098_23762# a_8438_23755# 0.24088f
C5506 VDPWR a_10218_20806# 0.83839f
C5507 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.22497f
C5508 VDPWR sar9b_0.net18 1.35357f
C5509 sar9b_0.net61 sar9b_0.net27 0.12915f
C5510 VDPWR a_16357_9613# 0.18873f
C5511 a_6307_27584# sar9b_0.net36 0.04789f
C5512 a_5322_17846# a_5046_17906# 0.1263f
C5513 a_7138_27758# sar9b_0.net60 0.0875f
C5514 sar9b_0.net58 a_4136_25584# 0.04102f
C5515 sar9b_0.net57 a_6137_23791# 0.07535f
C5516 a_11842_19766# a_12182_19759# 0.24088f
C5517 a_7289_21127# sar9b_0.net62 0.02399f
C5518 sar9b_0.net10 a_11382_22142# 0.06561f
C5519 sar9b_0.net47 a_5811_19178# 0.01123f
C5520 a_9802_26815# a_9593_26914# 0.24088f
C5521 single_9b_cdac_0.SW[7] a_29134_26999# 0.28324f
C5522 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.0303f
C5523 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.S[3] 0.22939f
C5524 sar9b_0.net65 sar9b_0.clk_div_0.COUNT\[0\] 0.08053f
C5525 sar9b_0.net18 a_3370_27769# 0.02082f
C5526 a_11338_19178# sar9b_0.net73 0.01335f
C5527 a_10402_25094# sar9b_0.net12 0.10692f
C5528 sar9b_0.net14 uo_out[0] 0.26202f
C5529 single_9b_cdac_1.CF[8] single_9b_cdac_0.SW[2] 0.01637f
C5530 sar9b_0._12_ clk 0.1358f
C5531 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 a_30012_17740# 0.14695f
C5532 VDPWR single_9b_cdac_1.cdac_sw_9b_0.S[1] 4.14969f
C5533 a_3695_23038# sar9b_0.clk_div_0.COUNT\[2\] 0.21948f
C5534 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45521f
C5535 sar9b_0.net36 single_9b_cdac_1.SW[2] 0.1913f
C5536 sar9b_0.net45 a_8883_27466# 0.30828f
C5537 sar9b_0.net41 sar9b_0.net38 0.17261f
C5538 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 2.71729f
C5539 sar9b_0.net24 sar9b_0.net45 0.03105f
C5540 VDPWR a_7590_24931# 0.27042f
C5541 VDPWR sar9b_0.net41 1.4128f
C5542 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.0303f
C5543 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[2] 0.01297f
C5544 single_9b_cdac_1.SW[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.17209f
C5545 sar9b_0.net49 a_9930_20510# 0.25469f
C5546 a_3561_22527# a_3454_22567# 0.14439f
C5547 a_9130_26198# sar9b_0.net37 0.01529f
C5548 a_4210_22378# sar9b_0.clknet_0_CLK 0.03169f
C5549 single_9b_cdac_1.cdac_sw_9b_0.S[2] single_9b_cdac_1.SW[2] 0.22543f
C5550 a_10227_18142# sar9b_0.net48 0.02398f
C5551 a_10548_19053# sar9b_0.net26 0.06094f
C5552 a_4755_22138# a_5739_22488# 0.08669f
C5553 a_9126_19131# a_7914_19178# 0.07766f
C5554 a_13011_21906# sar9b_0.net9 0.22439f
C5555 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y 0.07517f
C5556 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A a_40321_15495# 0.01076f
C5557 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.28523f
C5558 sar9b_0.net41 sar9b_0.net1 0.90489f
C5559 sar9b_0.net40 sar9b_0.net58 0.01707f
C5560 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INN 0.06563f
C5561 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.02632f
C5562 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36044f
C5563 sar9b_0.net7 sar9b_0.net27 0.06127f
C5564 sar9b_0.net68 sar9b_0.clknet_1_1__leaf_CLK 0.02176f
C5565 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.12359f
C5566 sar9b_0.net44 a_3540_27045# 0.27099f
C5567 uo_out[0] th_dif_sw_0.VCN 0.08774f
C5568 th_dif_sw_0.th_sw_1.CK ua[4] 0.42268f
C5569 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN ua[0] 3.10217f
C5570 sar9b_0.net35 a_7347_24160# 0.03326f
C5571 VDPWR a_13011_24802# 0.4961f
C5572 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[4] 10.6485f
C5573 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.27803f
C5574 a_3855_25792# sar9b_0.clknet_1_1__leaf_CLK 0.07223f
C5575 sar9b_0.net40 a_6137_23791# 0.01879f
C5576 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_1.CF[4] 0.10499f
C5577 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.04988f
C5578 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.03729f
C5579 a_10218_24802# a_10742_25087# 0.05022f
C5580 a_4811_23656# sar9b_0.net72 0.2012f
C5581 sar9b_0.net62 sar9b_0.net37 0.04598f
C5582 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.03436f
C5583 sar9b_0.net13 sar9b_0.net30 0.0911f
C5584 sar9b_0.net12 sar9b_0.net53 0.44449f
C5585 single_9b_cdac_1.CF[5] single_9b_cdac_1.SW[1] 0.22097f
C5586 VDPWR a_2918_20140# 0.90101f
C5587 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VDPWR 0.38397f
C5588 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5589 sar9b_0._09_ sar9b_0._17_ 0.04079f
C5590 a_8057_18463# a_8334_18353# 0.09983f
C5591 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.02632f
C5592 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01003f
C5593 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[3] 0.01887f
C5594 a_6058_18445# a_6126_18353# 0.35559f
C5595 a_5849_18463# a_6634_18206# 0.26257f
C5596 a_18214_3039# VDPWR 0.51112f
C5597 sar9b_0.net23 sar9b_0.net59 1.32079f
C5598 a_8166_27595# a_8512_27801# 0.07649f
C5599 VDPWR a_3754_26815# 0.20695f
C5600 sar9b_0.net56 sar9b_0.net73 0.05473f
C5601 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.62443f
C5602 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38317f
C5603 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[6] 0.02056f
C5604 sar9b_0.net9 sar9b_0.net36 0.33969f
C5605 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 0.0115f
C5606 sar9b_0.net13 a_9942_24806# 0.08367f
C5607 a_11008_17491# sar9b_0.net61 0.03855f
C5608 single_9b_cdac_0.SW[2] a_13067_27662# 0.3597f
C5609 a_8202_23174# sar9b_0.net62 0.02827f
C5610 sar9b_0._09_ sar9b_0._08_ 0.0865f
C5611 a_3540_27045# a_3822_27060# 0.06034f
C5612 a_9942_27470# a_10402_27758# 0.26257f
C5613 VDPWR sar9b_0.net31 1.59832f
C5614 a_6954_27466# sar9b_0.net45 0.02051f
C5615 VDPWR a_2847_27473# 0.29759f
C5616 single_9b_cdac_1.SW[4] ua[0] 0.13619f
C5617 single_9b_cdac_1.cdac_sw_9b_0.S[5] single_9b_cdac_1.cdac_sw_9b_0.S[7] 1.06635f
C5618 a_5581_20992# a_5812_21028# 0.10754f
C5619 sar9b_0.net51 a_5844_18123# 0.01122f
C5620 sar9b_0.net59 a_9593_26914# 0.11113f
C5621 sar9b_0.net9 single_9b_cdac_1.CF[4] 0.01701f
C5622 sar9b_0.net42 sar9b_0.net39 1.25124f
C5623 VDPWR tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.45581f
C5624 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.42014f
C5625 a_5235_27466# a_5460_28377# 0.01146f
C5626 sar9b_0.net36 sar9b_0.net61 0.03284f
C5627 sar9b_0.net44 sar9b_0.net36 0.21739f
C5628 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 1.55982f
C5629 a_4083_28566# a_4812_28371# 0.01209f
C5630 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.05472f
C5631 a_11338_19178# sar9b_0.net50 0.01132f
C5632 a_5460_28377# a_5742_28392# 0.06034f
C5633 sar9b_0.net18 a_4083_28566# 0.2051f
C5634 a_3603_28156# sar9b_0.net59 0.32304f
C5635 sar9b_0.net70 sar9b_0.clk_div_0.COUNT\[1\] 0.23038f
C5636 single_9b_cdac_0.SW[8] uo_out[0] 0.10191f
C5637 sar9b_0.net42 a_11382_23474# 0.02429f
C5638 a_12531_28566# uo_out[1] 0.38317f
C5639 a_10803_18142# sar9b_0.net73 0.13298f
C5640 a_11915_28371# uo_out[1] 0.04028f
C5641 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.02545f
C5642 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5643 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.3196f
C5644 tdc_0.OUTP a_16159_13315# 0.05276f
C5645 sar9b_0.net6 single_9b_cdac_1.SW[0] 0.10368f
C5646 a_7890_26108# sar9b_0.cyclic_flag_0.FINAL 0.083f
C5647 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.01751f
C5648 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 a_34814_17740# 0.14695f
C5649 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A 0.42784f
C5650 sar9b_0.net56 sar9b_0.net6 0.14505f
C5651 sar9b_0._05_ a_4236_21738# 0.27985f
C5652 a_11859_17910# sar9b_0.net39 0.20696f
C5653 sar9b_0.net57 a_5196_19448# 0.01615f
C5654 ui_in[4] ui_in[3] 0.03102f
C5655 sar9b_0.net66 sar9b_0.net69 0.14538f
C5656 sar9b_0.net47 a_6879_22145# 0.17478f
C5657 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP 3.27788f
C5658 a_7638_19238# a_8098_18810# 0.26257f
C5659 a_12182_23755# a_12047_23853# 0.35559f
C5660 a_12870_23599# a_13216_23805# 0.07649f
C5661 sar9b_0.net70 a_3371_23106# 0.01159f
C5662 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 3.27832f
C5663 VDPWR a_13011_19242# 0.48316f
C5664 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[6] 0.06019f
C5665 a_9130_26198# sar9b_0.net59 0.27842f
C5666 sar9b_0.net41 sar9b_0.net48 0.33991f
C5667 sar9b_0.net7 a_11008_17491# 0.27173f
C5668 a_10858_17113# a_10644_16791# 0.04522f
C5669 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.02545f
C5670 VDPWR th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.17946f
C5671 sar9b_0.net47 sar9b_0.net62 0.38866f
C5672 a_6642_19448# a_7097_19795# 0.3578f
C5673 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[4] 0.17948f
C5674 a_13011_24802# sar9b_0.net29 0.01443f
C5675 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN 0.02519f
C5676 sar9b_0.net41 a_9900_19047# 0.01957f
C5677 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.01175f
C5678 a_11915_27039# sar9b_0.net45 0.10003f
C5679 sar9b_0.net7 sar9b_0.net36 0.02886f
C5680 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[8] 0.23119f
C5681 a_7566_21017# a_8074_20870# 0.19065f
C5682 tdc_0.OUTP sar9b_0.net2 0.24126f
C5683 single_9b_cdac_1.CF[6] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.06503f
C5684 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C5685 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.17533f
C5686 sar9b_0._18_ sar9b_0.net66 0.0125f
C5687 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.6919f
C5688 VDPWR a_12435_24802# 0.45648f
C5689 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A 0.12431f
C5690 sar9b_0.net41 a_9270_24566# 0.01466f
C5691 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02778f
C5692 sar9b_0.net63 a_5823_23477# 0.05368f
C5693 a_11842_26426# a_12618_26134# 0.3578f
C5694 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.28523f
C5695 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 ua[0] 0.12344f
C5696 single_9b_cdac_1.SW[3] single_9b_cdac_1.SW[0] 0.0223f
C5697 sar9b_0.net56 sar9b_0.net46 2.24988f
C5698 a_10506_23174# clk 0.01873f
C5699 VDPWR a_10662_17799# 0.26449f
C5700 sar9b_0.net60 a_4583_20468# 0.01054f
C5701 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.SW[4] 0.17303f
C5702 a_53154_16877# single_9b_cdac_1.SW[2] 0.28324f
C5703 VDPWR uo_out[7] 1.05965f
C5704 a_11776_27801# VDPWR 0.20399f
C5705 VDPWR a_12435_20806# 0.43957f
C5706 a_3206_22432# a_3713_22522# 0.21226f
C5707 sar9b_0.net12 a_10932_25713# 0.01703f
C5708 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 ua[0] 0.12378f
C5709 a_8057_18463# sar9b_0.net61 0.01568f
C5710 sar9b_0.net42 a_10402_25094# 0.01861f
C5711 sar9b_0.net31 sar9b_0.net29 0.0246f
C5712 sar9b_0.clk_div_0.COUNT\[3\] sar9b_0._12_ 0.05952f
C5713 VDPWR a_5100_24375# 0.1934f
C5714 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.42509f
C5715 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.69086f
C5716 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.95338f
C5717 sar9b_0.net56 a_9154_20142# 0.01042f
C5718 sar9b_0.net36 a_4749_27652# 0.07973f
C5719 sar9b_0.net58 a_3090_27163# 0.26444f
C5720 VDPWR a_8874_19178# 0.41712f
C5721 a_11658_18142# a_11842_18434# 0.44532f
C5722 sar9b_0.clknet_1_0__leaf_CLK a_2918_20140# 0.12018f
C5723 th_dif_sw_0.VCN single_9b_cdac_0.SW[0] 0.09453f
C5724 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.45521f
C5725 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.17533f
C5726 VDPWR a_5484_23444# 0.19999f
C5727 VDPWR a_5506_17478# 0.21624f
C5728 sar9b_0.net27 sar9b_0.net5 0.07039f
C5729 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[1\] 0.02478f
C5730 single_9b_cdac_1.cdac_sw_9b_0.S[7] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.25152f
C5731 sar9b_0.net21 uo_out[5] 0.07619f
C5732 VDPWR a_7692_26108# 0.20712f
C5733 sar9b_0.net58 a_3156_27447# 0.17605f
C5734 sar9b_0.clknet_0_CLK sar9b_0.net39 0.08885f
C5735 sar9b_0.net49 a_11178_20806# 0.26056f
C5736 VDPWR a_5126_20140# 0.84448f
C5737 a_10803_18142# single_9b_cdac_1.SW[3] 0.3509f
C5738 sar9b_0.net17 sar9b_0.net60 0.14205f
C5739 sar9b_0.net50 a_12684_20379# 0.11466f
C5740 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.31534f
C5741 VDPWR a_11718_23127# 0.26767f
C5742 sar9b_0.net23 a_7890_26108# 0.05346f
C5743 single_9b_cdac_0.SW[7] uo_out[0] 0.04546f
C5744 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.28523f
C5745 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[1] 0.2176f
C5746 a_7289_21127# a_7284_20787# 0.44098f
C5747 a_10218_20806# a_9930_20510# 0.01059f
C5748 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[8] 2.12011f
C5749 sar9b_0.net16 a_2603_17006# 0.22549f
C5750 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.69086f
C5751 VDPWR sar9b_0.net68 0.48583f
C5752 VDPWR a_6867_16810# 0.26271f
C5753 a_8052_18123# sar9b_0.net37 0.01856f
C5754 VDPWR a_43540_16877# 1.81495f
C5755 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[1\] 0.01596f
C5756 sar9b_0.net13 sar9b_0.net54 1.09911f
C5757 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C5758 a_11859_20574# single_9b_cdac_1.SW[8] 0.35377f
C5759 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[5] 0.01887f
C5760 a_6378_24802# a_6902_25087# 0.05022f
C5761 sar9b_0.net42 sar9b_0.net53 0.62196f
C5762 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 0.42014f
C5763 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 2.7611f
C5764 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN 2.81718f
C5765 VDPWR a_3855_25792# 0.09015f
C5766 a_11382_23474# sar9b_0.net74 0.18434f
C5767 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_41357_15501# 0.01076f
C5768 sar9b_0._09_ a_3991_19768# 0.01296f
C5769 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN ua[0] 3.10218f
C5770 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.0303f
C5771 single_9b_cdac_1.CF[2] single_9b_cdac_1.SW[0] 0.22502f
C5772 sar9b_0.cyclic_flag_0.FINAL sar9b_0.net54 0.09984f
C5773 sar9b_0.net1 a_6867_16810# 0.1431f
C5774 a_11382_18146# sar9b_0.net61 0.02131f
C5775 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.6919f
C5776 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C5777 a_2739_20140# a_3166_20145# 0.04602f
C5778 sar9b_0.net52 a_10623_25895# 0.21039f
C5779 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.45521f
C5780 a_7926_23234# clk 0.01904f
C5781 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.3196f
C5782 sar9b_0.net35 sar9b_0.clk_div_0.COUNT\[2\] 0.02371f
C5783 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y single_9b_cdac_1.CF[6] 0.12898f
C5784 VDPWR a_6102_24806# 0.29526f
C5785 sar9b_0.net41 a_9930_20510# 0.02662f
C5786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.42509f
C5787 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 2.81428f
C5788 single_9b_cdac_1.SW[1] ua[0] 0.15672f
C5789 sar9b_0.net38 sar9b_0.net22 0.04437f
C5790 VDPWR a_5580_24776# 0.24626f
C5791 sar9b_0.net49 a_9942_20810# 0.28171f
C5792 a_7404_17715# sar9b_0.net73 0.12657f
C5793 sar9b_0.net57 a_10218_24802# 0.2148f
C5794 VDPWR sar9b_0.net22 0.53629f
C5795 a_4755_22138# sar9b_0.clknet_1_1__leaf_CLK 0.22079f
C5796 single_9b_cdac_1.SW[8] sar9b_0.net51 0.0423f
C5797 a_11658_23470# a_12870_23599# 0.07766f
C5798 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[0] 0.01887f
C5799 a_9132_7271# th_dif_sw_0.th_sw_1.CKB 0.01594f
C5800 single_9b_cdac_1.SW[4] sar9b_0.net27 0.46877f
C5801 VDPWR a_5761_21100# 0.01372f
C5802 a_10649_17131# single_9b_cdac_1.SW[2] 0.0163f
C5803 sar9b_0._14_ sar9b_0.clk_div_0.COUNT\[2\] 0.02642f
C5804 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5805 a_8345_26455# a_8622_26345# 0.09983f
C5806 VDPWR a_5322_17846# 0.85398f
C5807 a_3454_22567# a_3027_22138# 0.04602f
C5808 sar9b_0.net67 sar9b_0._05_ 0.21501f
C5809 VDPWR a_11842_19766# 0.23652f
C5810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.10626f
C5811 a_9472_18823# sar9b_0.net26 0.27337f
C5812 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C5813 sar9b_0.net9 sar9b_0.net51 0.02854f
C5814 a_10662_17799# sar9b_0.net48 0.1748f
C5815 a_7374_19685# sar9b_0.net47 0.29639f
C5816 sar9b_0.net40 sar9b_0.clk_div_0.COUNT\[1\] 0.0227f
C5817 a_11178_27466# sar9b_0.net59 0.26568f
C5818 sar9b_0.net65 sar9b_0.clknet_0_CLK 0.2446f
C5819 VDPWR a_9760_22819# 0.20965f
C5820 sar9b_0.net40 sar9b_0.net73 0.05965f
C5821 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[1] 2.07974f
C5822 sar9b_0._07_ a_4947_20140# 0.02502f
C5823 sar9b_0.net13 sar9b_0.net27 0.04207f
C5824 a_7092_19455# sar9b_0.net47 0.18759f
C5825 single_9b_cdac_1.SW[5] single_9b_cdac_1.SW[6] 8.40786f
C5826 a_4018_24235# sar9b_0.net58 0.01775f
C5827 a_14897_9355# clk 0.02917f
C5828 a_7470_22349# a_7978_22202# 0.19065f
C5829 sar9b_0.net61 sar9b_0.net51 0.06277f
C5830 sar9b_0.net3 sar9b_0.net19 0.0315f
C5831 sar9b_0.clk_div_0.COUNT\[0\] a_6484_22845# 0.24895f
C5832 sar9b_0.net7 a_11382_18146# 0.05241f
C5833 a_7404_17715# sar9b_0.net6 0.01668f
C5834 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[6] 0.02011f
C5835 a_57946_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.04592f
C5836 sar9b_0.net31 a_11915_27039# 0.03331f
C5837 sar9b_0.net8 a_11658_19474# 0.2065f
C5838 sar9b_0.net36 sar9b_0.net5 0.02542f
C5839 sar9b_0.net1 a_9760_22819# 0.0139f
C5840 a_8874_19178# sar9b_0.net48 0.29136f
C5841 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 0.17533f
C5842 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31753_29911# 0.01076f
C5843 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A 0.84061f
C5844 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP ua[0] 1.15121f
C5845 a_10402_25094# sar9b_0.net74 0.02019f
C5846 a_10548_19053# a_10553_18922# 0.44532f
C5847 sar9b_0.net8 sar9b_0.net49 0.4261f
C5848 a_4755_22138# a_4934_22432# 0.54361f
C5849 a_9126_19131# a_9472_18823# 0.07649f
C5850 tdc_0.OUTP th_dif_sw_0.CKB 0.30524f
C5851 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C5852 sar9b_0.net60 a_6378_24802# 0.01004f
C5853 a_6861_22828# sar9b_0.clk_div_0.COUNT\[1\] 0.05496f
C5854 VDPWR a_6058_18445# 0.20217f
C5855 sar9b_0.net43 a_9546_24506# 0.06524f
C5856 a_9839_17527# a_9974_17626# 0.35559f
C5857 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A a_49926_15495# 0.01076f
C5858 single_9b_cdac_0.SW[1] single_9b_cdac_1.CF[7] 0.02109f
C5859 a_9363_20826# a_9258_21842# 0.02481f
C5860 a_8386_22806# a_8726_22954# 0.24088f
C5861 a_8202_23174# a_9414_23127# 0.07766f
C5862 sar9b_0.net57 sar9b_0.net46 0.19212f
C5863 a_5484_23444# a_5682_23444# 0.06623f
C5864 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.26942f
C5865 a_5711_17527# a_5846_17626# 0.35559f
C5866 sar9b_0.net10 sar9b_0.net38 0.02721f
C5867 a_6975_20813# sar9b_0.net40 0.01008f
C5868 sar9b_0.net52 sar9b_0.net2 0.02335f
C5869 a_12531_28566# sar9b_0._06_ 0.02926f
C5870 VDPWR sar9b_0.net10 3.17323f
C5871 single_9b_cdac_1.CF[6] single_9b_cdac_1.CF[7] 5.94919f
C5872 a_6880_17491# sar9b_0.net56 0.0197f
C5873 single_9b_cdac_1.SW[6] ua[0] 0.13161f
C5874 a_13216_23805# a_13011_24570# 0.01043f
C5875 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.03729f
C5876 sar9b_0.net40 sar9b_0.net6 0.05038f
C5877 a_10816_21487# sar9b_0.net9 0.31769f
C5878 VDPWR a_3027_21906# 0.29917f
C5879 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.SW[0] 0.17156f
C5880 sar9b_0.net22 a_8883_27466# 0.02815f
C5881 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.CF[7] 0.0174f
C5882 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN 0.12358f
C5883 a_6137_23791# clk 0.01311f
C5884 sar9b_0.net1 sar9b_0.net10 0.02729f
C5885 VDPWR sar9b_0._05_ 0.50167f
C5886 a_8842_16874# sar9b_0.net27 0.08083f
C5887 a_8303_23853# a_7638_23474# 0.19065f
C5888 a_7404_17715# sar9b_0.net46 0.03295f
C5889 sar9b_0.net7 sar9b_0.net51 0.02342f
C5890 a_10649_17131# sar9b_0.net61 0.01074f
C5891 sar9b_0.net6 a_9174_17906# 0.18423f
C5892 a_7284_20787# sar9b_0.net47 0.17237f
C5893 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04988f
C5894 a_21177_7457# th_dif_sw_0.VCP 0.0867f
C5895 sar9b_0.net74 sar9b_0.net53 0.63719f
C5896 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN single_9b_cdac_1.CF[0] 0.12358f
C5897 a_10895_22855# sar9b_0.net74 0.02448f
C5898 single_9b_cdac_0.SW[6] uo_out[3] 0.30173f
C5899 VDPWR a_12182_26419# 0.20236f
C5900 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN ua[0] 3.10207f
C5901 single_9b_cdac_1.CF[0] clk 0.08196f
C5902 sar9b_0.net27 a_12618_19474# 0.02681f
C5903 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_1.SW[0] 0.12586f
C5904 sar9b_0.net70 a_2508_23444# 0.08416f
C5905 single_9b_cdac_0.cdac_sw_9b_0.S[8] single_9b_cdac_0.cdac_sw_9b_0.S[6] 1.08672f
C5906 a_8052_18123# a_7602_18116# 0.03471f
C5907 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C5908 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A 0.95338f
C5909 sar9b_0.net17 uio_out[1] 0.1629f
C5910 a_5439_24563# sar9b_0.net39 0.01949f
C5911 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A a_64331_15495# 0.01076f
C5912 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[4] 1.90184f
C5913 sar9b_0.net63 a_2940_25096# 0.02555f
C5914 single_9b_cdac_0.cdac_sw_9b_0.S[0] th_dif_sw_0.VCN 0.21769p
C5915 sar9b_0.net40 sar9b_0.net50 0.30217f
C5916 th_dif_sw_0.th_sw_1.CKB ua[4] 0.08416f
C5917 sar9b_0.net40 single_9b_cdac_1.SW[3] 0.03187f
C5918 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[1] 0.84424f
C5919 sar9b_0.net53 a_12618_23470# 0.26167f
C5920 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y 0.3196f
C5921 a_8057_18463# sar9b_0.net5 0.10125f
C5922 sar9b_0.net40 a_12618_18142# 0.01397f
C5923 a_10402_21098# a_10742_21091# 0.24088f
C5924 a_10218_20806# a_11178_20806# 0.03432f
C5925 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.2428f
C5926 a_11382_22142# a_11658_22138# 0.1263f
C5927 a_10482_25831# a_10932_25713# 0.03432f
C5928 sar9b_0.net53 a_10506_24506# 0.24393f
C5929 a_11842_23762# clk 0.01052f
C5930 sar9b_0.net13 sar9b_0.net36 0.024f
C5931 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.22879f
C5932 VDPWR a_7914_19178# 0.75628f
C5933 VDPWR a_29134_26999# 1.81495f
C5934 a_11658_26134# a_12618_26134# 0.03432f
C5935 sar9b_0.net40 a_6378_24802# 0.0119f
C5936 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.3196f
C5937 single_9b_cdac_0.SW[6] single_9b_cdac_0.SW[4] 0.03895f
C5938 sar9b_0.net10 sar9b_0._17_ 0.01904f
C5939 sar9b_0.net36 sar9b_0.cyclic_flag_0.FINAL 0.23039f
C5940 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.05632f
C5941 single_9b_cdac_0.cdac_sw_9b_0.S[4] a_44418_26990# 0.22513f
C5942 single_9b_cdac_0.SW[4] clk 0.1627f
C5943 a_7188_22119# a_7470_22349# 0.05462f
C5944 a_11842_19766# a_12047_19857# 0.09983f
C5945 a_2892_23070# sar9b_0.net69 0.01085f
C5946 a_48343_26999# single_9b_cdac_0.cdac_sw_9b_0.S[3] 0.59531f
C5947 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 0.26707f
C5948 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.SW[4] 0.22983f
C5949 sar9b_0.net48 a_6058_18445# 0.14602f
C5950 a_10548_19053# sar9b_0.net38 0.01246f
C5951 single_9b_cdac_1.SW[1] sar9b_0.net27 0.17807f
C5952 tdc_0.OUTP single_9b_cdac_1.SW[0] 0.86423f
C5953 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A 0.01751f
C5954 sar9b_0.net54 sar9b_0.net62 0.89973f
C5955 single_9b_cdac_0.SW[1] single_9b_cdac_0.SW[2] 16.8504f
C5956 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.22875f
C5957 VDPWR a_11382_19478# 0.30104f
C5958 VDPWR a_10548_19053# 0.83308f
C5959 VDPWR a_4755_22138# 0.4525f
C5960 a_12870_18271# sar9b_0.net50 0.17284f
C5961 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 0.19266f
C5962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP a_48343_16877# 0.04592f
C5963 sar9b_0.net52 a_7914_23470# 0.15191f
C5964 VDPWR a_9839_17527# 0.25186f
C5965 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38397f
C5966 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[6] 0.02024f
C5967 a_12870_18271# a_12618_18142# 0.27388f
C5968 a_11842_18434# a_12047_18525# 0.09983f
C5969 a_9942_20810# a_10218_20806# 0.1263f
C5970 VDPWR tdc_0.phase_detector_0.INN 0.51155f
C5971 single_9b_cdac_1.CF[2] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.12898f
C5972 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_1.CF[5] 0.06503f
C5973 sar9b_0.net60 sar9b_0._03_ 0.02848f
C5974 a_2892_23070# sar9b_0._18_ 0.28345f
C5975 single_9b_cdac_1.cdac_sw_9b_0.S[6] th_dif_sw_0.VCP 3.33405f
C5976 sar9b_0.net11 sar9b_0.net37 0.02799f
C5977 a_6540_22112# sar9b_0.net39 0.30426f
C5978 single_9b_cdac_1.CF[4] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.06503f
C5979 sar9b_0._10_ sar9b_0.net71 0.01246f
C5980 sar9b_0._11_ sar9b_0.net65 0.09114f
C5981 a_45123_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A 0.01076f
C5982 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.05472f
C5983 sar9b_0.net43 a_5753_24250# 0.01111f
C5984 a_5046_27230# a_5506_26802# 0.26257f
C5985 a_5322_27170# a_5846_26950# 0.04522f
C5986 a_5298_24499# a_5753_24250# 0.3578f
C5987 sar9b_0.clknet_1_0__leaf_CLK a_3027_21906# 0.01945f
C5988 a_11859_20574# sar9b_0.net5 0.03891f
C5989 sar9b_0.net20 sar9b_0.net38 0.02978f
C5990 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C5991 sar9b_0.net38 a_10402_21098# 0.0282f
C5992 sar9b_0.net42 a_11104_24151# 0.30428f
C5993 sar9b_0.net58 a_5846_26950# 0.13488f
C5994 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A 0.84061f
C5995 single_9b_cdac_0.SW[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.14962f
C5996 VDPWR sar9b_0.net20 0.27201f
C5997 a_8098_23762# a_8874_23470# 0.3578f
C5998 VDPWR a_10402_21098# 0.21902f
C5999 sar9b_0.net74 a_10932_25713# 0.06691f
C6000 sar9b_0.clknet_1_0__leaf_CLK sar9b_0._05_ 0.03201f
C6001 sar9b_0.net41 a_9942_20810# 0.01321f
C6002 a_8202_23174# sar9b_0.net11 0.26859f
C6003 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 ua[0] 0.12077f
C6004 a_8166_27595# sar9b_0.net60 0.17093f
C6005 sar9b_0.net57 a_6346_23773# 0.03377f
C6006 a_10378_27170# a_9588_27045# 0.1263f
C6007 a_4136_25584# sar9b_0._03_ 0.29527f
C6008 sar9b_0.net60 a_5460_28377# 0.02635f
C6009 a_33936_26999# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.23864f
C6010 a_11430_24931# sar9b_0.net12 0.07831f
C6011 single_9b_cdac_1.SW[0] single_9b_cdac_1.SW[7] 0.02168f
C6012 sar9b_0.net8 a_10218_20806# 0.04227f
C6013 sar9b_0.net5 sar9b_0.net51 1.21471f
C6014 a_7188_22119# sar9b_0.clk_div_0.COUNT\[2\] 0.01175f
C6015 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN ua[0] 3.10215f
C6016 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[7] 0.06019f
C6017 sar9b_0.net45 sar9b_0.net34 0.19873f
C6018 sar9b_0.net53 sar9b_0.net39 0.01835f
C6019 VDPWR a_7936_25137# 0.20887f
C6020 a_6880_17491# a_7404_17715# 0.01194f
C6021 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A 0.12431f
C6022 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 2.7611f
C6023 sar9b_0.net23 sar9b_0.net36 0.02152f
C6024 clk ena 0.03102f
C6025 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_50962_15501# 0.01076f
C6026 single_9b_cdac_0.cdac_sw_9b_0.S[8] ua[0] 16.2797f
C6027 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A 0.28523f
C6028 sar9b_0.net48 a_7914_19178# 0.17382f
C6029 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A 0.38397f
C6030 VDPWR a_8438_23755# 0.20949f
C6031 a_11382_23474# sar9b_0.net53 0.25588f
C6032 a_10830_19068# sar9b_0.net26 0.04966f
C6033 a_8098_23762# sar9b_0.net37 0.01305f
C6034 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A 0.84059f
C6035 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A 0.04988f
C6036 sar9b_0.net14 sar9b_0.net25 0.2521f
C6037 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.3196f
C6038 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[7] 0.01887f
C6039 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP 1.55985f
C6040 VDPWR a_33936_26999# 1.81495f
C6041 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.SW[0] 0.08409f
C6042 a_13011_16810# single_9b_cdac_1.SW[5] 0.35162f
C6043 a_4755_22138# a_5441_22522# 0.27693f
C6044 sar9b_0.net36 a_9593_26914# 0.11605f
C6045 sar9b_0.net31 sar9b_0.net33 0.02107f
C6046 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26942f
C6047 sar9b_0.net9 sar9b_0.net42 0.01827f
C6048 single_9b_cdac_1.CF[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C6049 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 a_49221_17740# 0.14695f
C6050 sar9b_0.net58 sar9b_0.net45 0.10292f
C6051 sar9b_0.net4 a_5753_24250# 0.02172f
C6052 sar9b_0.net41 sar9b_0.net8 0.02515f
C6053 a_8970_20510# a_8694_20570# 0.1263f
C6054 single_9b_cdac_1.CF[3] single_9b_cdac_1.SW[0] 0.2246f
C6055 a_11339_27039# single_9b_cdac_0.SW[5] 0.36476f
C6056 single_9b_cdac_1.CF[1] single_9b_cdac_1.CF[7] 0.01994f
C6057 sar9b_0.net36 single_9b_cdac_1.SW[1] 0.03305f
C6058 sar9b_0._15_ a_5753_24250# 0.05531f
C6059 sar9b_0.net69 sar9b_0.clknet_1_1__leaf_CLK 0.08399f
C6060 sar9b_0.net42 sar9b_0.net61 0.08366f
C6061 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A 0.45521f
C6062 a_10218_24802# a_11178_24802# 0.03432f
C6063 single_9b_cdac_1.CF[4] single_9b_cdac_1.SW[1] 0.22097f
C6064 a_5289_22527# a_5182_22567# 0.14439f
C6065 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.75899f
C6066 VDPWR a_8970_20510# 0.9047f
C6067 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.02778f
C6068 sar9b_0.net34 a_9870_27060# 0.01531f
C6069 a_10548_19053# sar9b_0.net48 0.16225f
C6070 a_6250_28502# sar9b_0.net38 0.16677f
C6071 sar9b_0.net48 a_9839_17527# 0.2029f
C6072 single_9b_cdac_1.CF[8] sar9b_0.net13 0.01097f
C6073 a_8057_18463# a_8842_18206# 0.26257f
C6074 single_9b_cdac_1.CF[5] th_dif_sw_0.VCN 0.09453f
C6075 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A 0.95338f
C6076 VDPWR a_6250_28502# 0.29018f
C6077 a_10239_19235# a_10098_19171# 0.27388f
C6078 single_9b_cdac_0.cdac_sw_9b_0.S[4] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.28033f
C6079 m2_23774_17236# VDPWR 0.19016f
C6080 sar9b_0.net68 a_4044_24776# 0.041f
C6081 sar9b_0.net52 a_10742_25087# 0.12673f
C6082 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A 0.03729f
C6083 a_10218_21842# sar9b_0.net38 0.02659f
C6084 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_65367_15501# 0.01076f
C6085 a_10227_23490# sar9b_0.net38 0.02331f
C6086 sar9b_0._18_ sar9b_0.clknet_1_1__leaf_CLK 0.02875f
C6087 sar9b_0.net32 sar9b_0.net13 0.02694f
C6088 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62553f
C6089 clk sar9b_0.clk_div_0.COUNT\[1\] 0.08722f
C6090 single_9b_cdac_1.cdac_sw_9b_0.S[8] ua[0] 16.2977f
C6091 sar9b_0.net30 a_11842_26426# 0.01579f
C6092 a_5823_23477# sar9b_0.net11 0.05916f
C6093 VDPWR a_10218_21842# 0.36269f
C6094 a_3795_19512# a_4072_19474# 0.26693f
C6095 a_10218_27466# a_10742_27751# 0.05022f
C6096 VDPWR a_10227_23490# 0.4365f
C6097 a_7138_27758# sar9b_0.net45 0.01918f
C6098 single_9b_cdac_0.cdac_sw_9b_0.S[0] single_9b_cdac_0.cdac_sw_9b_0.S[5] 0.33229f
C6099 a_5581_20992# sar9b_0._11_ 0.06877f
C6100 a_11382_19478# a_12047_19857# 0.19065f
C6101 sar9b_0.net71 a_3795_19512# 0.03166f
C6102 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.24399f
C6103 a_10742_21091# a_10607_21189# 0.35559f
C6104 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[2] 0.31534f
C6105 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.95338f
C6106 a_3231_27227# a_3540_27045# 0.07766f
C6107 a_4812_28371# sar9b_0.net58 0.02979f
C6108 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.S[5] 1.56015f
C6109 sar9b_0.net18 sar9b_0.net58 0.33351f
C6110 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A 0.95338f
C6111 a_10227_23490# sar9b_0.net1 0.13989f
C6112 a_11722_25838# a_10937_25582# 0.26257f
C6113 a_3161_27787# a_3438_27677# 0.09983f
C6114 sar9b_0._06_ uo_out[1] 0.0432f
C6115 a_9546_24506# a_10070_24286# 0.04522f
C6116 sar9b_0.net2 a_10758_24459# 0.07084f
C6117 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A a_54737_15495# 0.01076f
C6118 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.02638f
C6119 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C6120 sar9b_0.net7 sar9b_0.net42 0.12319f
C6121 single_9b_cdac_0.cdac_sw_9b_0.S[2] single_9b_cdac_0.cdac_sw_9b_0.S[1] 16.8012f
C6122 single_9b_cdac_1.CF[1] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 0.42014f
C6123 sar9b_0.net74 a_11104_24151# 0.01447f
C6124 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B 0.36961f
C6125 a_8345_26455# sar9b_0.cyclic_flag_0.FINAL 0.12177f
C6126 a_10470_21795# sar9b_0.net49 0.17598f
C6127 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[2] 0.01297f
C6128 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y 0.07579f
C6129 single_9b_cdac_0.cdac_sw_9b_0.S[6] th_dif_sw_0.VCN 3.33405f
C6130 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP ua[0] 1.17995f
C6131 single_9b_cdac_1.CF[5] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.0313f
C6132 sar9b_0.net47 a_7443_21496# 0.31185f
C6133 sar9b_0.net70 a_3027_22138# 0.03062f
C6134 sar9b_0.net15 sar9b_0.net51 0.14145f
C6135 VDPWR uo_out[0] 0.86559f
C6136 sar9b_0.net64 sar9b_0.net4 0.04411f
C6137 VDPWR sar9b_0.net19 0.3982f
C6138 a_9323_27662# single_9b_cdac_0.SW[8] 0.35813f
C6139 sar9b_0.net19 a_4330_27170# 0.04522f
C6140 a_11178_27466# single_9b_cdac_0.SW[5] 0.03553f
C6141 a_4934_22432# sar9b_0._18_ 0.02193f
C6142 sar9b_0.net45 single_9b_cdac_0.SW[4] 0.24467f
C6143 sar9b_0._05_ sar9b_0._12_ 0.12977f
C6144 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y 0.07517f
C6145 a_6252_20780# sar9b_0.net60 0.02523f
C6146 a_5628_19768# sar9b_0._10_ 0.06416f
C6147 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C6148 a_9939_28566# sar9b_0.net38 0.04052f
C6149 a_5748_24381# a_5753_24250# 0.44532f
C6150 a_10506_24506# a_11104_24151# 0.06623f
C6151 sar9b_0.net22 a_8691_28566# 0.2096f
C6152 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.26625f
C6153 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN ua[0] 3.10045f
C6154 a_9939_28566# VDPWR 0.44769f
C6155 VDPWR a_6744_23238# 0.16029f
C6156 a_6922_23534# a_6414_23681# 0.19065f
C6157 a_10895_22855# sar9b_0.net53 0.2218f
C6158 a_3369_24181# a_3014_24136# 0.18752f
C6159 sar9b_0.net49 sar9b_0.net73 0.10388f
C6160 a_10690_22806# a_11030_22954# 0.24088f
C6161 a_10506_23174# a_11718_23127# 0.07766f
C6162 sar9b_0.net41 a_9730_24138# 0.02215f
C6163 sar9b_0.net26 sar9b_0.net37 0.22151f
C6164 a_11842_26426# a_12047_26517# 0.09983f
C6165 a_12870_26263# a_12618_26134# 0.27388f
C6166 single_9b_cdac_0.cdac_sw_9b_0.S[5] a_38738_26999# 0.59531f
C6167 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP 0.19266f
C6168 a_6282_27170# a_6534_27123# 0.27388f
C6169 tdc_0.OUTP sar9b_0.net40 0.02274f
C6170 VDPWR a_12491_27662# 0.49074f
C6171 a_3946_26198# sar9b_0.net44 0.05662f
C6172 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN single_9b_cdac_1.CF[4] 0.03478f
C6173 sar9b_0.net9 sar9b_0.net74 0.10219f
C6174 a_10218_27466# a_10607_27849# 0.06034f
C6175 sar9b_0.net38 a_10607_21189# 0.01344f
C6176 sar9b_0.net30 sar9b_0.net11 0.14416f
C6177 a_6636_20780# a_6975_20813# 0.07649f
C6178 a_7284_20787# a_6834_20780# 0.03471f
C6179 a_7638_19238# sar9b_0.net5 0.03793f
C6180 sar9b_0.net51 a_5811_19178# 0.11557f
C6181 VDPWR a_10607_21189# 0.26776f
C6182 a_3206_22432# a_4210_22378# 0.06302f
C6183 a_9414_23127# sar9b_0.net54 0.18588f
C6184 sar9b_0.net40 a_6444_19448# 0.30912f
C6185 a_3206_22432# sar9b_0.clknet_0_CLK 0.01173f
C6186 VDPWR sar9b_0._13_ 0.47588f
C6187 tdc_0.RDY sar9b_0.net27 0.05081f
C6188 sar9b_0.net43 sar9b_0.net37 0.04982f
C6189 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.03488f
C6190 a_8940_27039# a_9279_27227# 0.07649f
C6191 single_9b_cdac_1.cdac_sw_9b_0.S[0] ua[0] 1.20078f
C6192 VDPWR a_10803_19474# 0.44387f
C6193 a_9258_21842# sar9b_0.net57 0.22486f
C6194 single_9b_cdac_1.SW[3] clk 0.10355f
C6195 sar9b_0.net58 a_3754_26815# 0.14463f
C6196 sar9b_0.net13 sar9b_0.net12 0.39165f
C6197 sar9b_0.net60 sar9b_0.clk_div_0.COUNT\[2\] 0.03174f
C6198 sar9b_0.net61 tdc_0.OUTN 0.01037f
C6199 a_5633_20244# a_5931_20140# 0.02614f
C6200 sar9b_0._14_ sar9b_0._16_ 0.12248f
C6201 single_9b_cdac_0.SW[2] single_9b_cdac_1.CF[7] 0.02052f
C6202 VDPWR a_9472_18823# 0.21089f
C6203 a_11658_18142# a_12870_18271# 0.07766f
C6204 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP 0.02666f
C6205 VDPWR a_5846_17626# 0.19864f
C6206 sar9b_0.net32 sar9b_0.net23 0.04971f
C6207 a_9126_19131# sar9b_0.net37 0.058f
C6208 sar9b_0.net58 a_2847_27473# 0.17334f
C6209 a_3922_20239# a_2739_20140# 0.0649f
C6210 a_13011_27234# sar9b_0._06_ 0.21168f
C6211 sar9b_0.net8 a_12435_20806# 0.08962f
C6212 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.02149f
C6213 a_8340_26115# sar9b_0.net37 0.02741f
C6214 sar9b_0.net43 a_9802_26815# 0.01853f
C6215 single_9b_cdac_1.CF[1] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN 0.12358f
C6216 single_9b_cdac_1.CF[8] single_9b_cdac_1.SW[1] 0.2162f
C6217 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6218 uo_out[6] ui_in[0] 0.06786f
C6219 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A single_9b_cdac_1.CF[4] 0.02149f
C6220 a_9472_18823# sar9b_0.net1 0.01552f
C6221 VDPWR a_9546_24506# 0.86145f
C6222 a_2835_24136# sar9b_0.net70 0.06896f
C6223 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.95338f
C6224 sar9b_0.net57 sar9b_0.clk_div_0.COUNT\[2\] 0.01818f
C6225 VDPWR a_13216_19809# 0.21451f
C6226 a_10644_16791# a_10194_16784# 0.03493f
C6227 a_9996_16784# a_10335_16817# 0.07649f
C6228 sar9b_0.net40 sar9b_0.net28 0.10374f
C6229 single_9b_cdac_1.SW[5] th_dif_sw_0.VCN 0.09453f
C6230 VDPWR a_8052_16791# 0.86212f
C6231 VDPWR a_6678_27470# 0.2784f
C6232 single_9b_cdac_1.CF[0] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A 0.0313f
C6233 sar9b_0.net5 a_9359_20191# 0.0567f
C6234 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.CF[0] 0.01887f
C6235 a_5938_22378# sar9b_0.net60 0.01049f
C6236 sar9b_0.net6 a_5849_18463# 0.01813f
C6237 a_4934_22432# a_4332_23043# 0.01428f
C6238 a_4755_22138# sar9b_0._12_ 0.15278f
C6239 VDPWR sar9b_0.net69 1.21061f
C6240 sar9b_0.net40 single_9b_cdac_1.SW[7] 0.05122f
C6241 sar9b_0._09_ a_5196_19448# 0.04256f
C6242 VDPWR a_11658_22138# 0.83163f
C6243 a_9939_28566# sar9b_0.net24 0.05176f
C6244 a_6744_23238# sar9b_0._17_ 0.03116f
C6245 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.06503f
C6246 sar9b_0.net72 sar9b_0.clknet_1_1__leaf_CLK 0.02825f
C6247 a_11658_19474# sar9b_0.net50 0.19816f
C6248 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.12223f
C6249 sar9b_0._00_ a_3166_20145# 0.13532f
C6250 a_2739_20140# a_3273_20185# 0.35097f
C6251 a_2918_20140# a_3425_20244# 0.21226f
C6252 sar9b_0.net52 a_10937_25582# 0.11747f
C6253 sar9b_0.net31 a_12182_22423# 0.02073f
C6254 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 ua[0] 0.12069f
C6255 a_11146_25483# sar9b_0.net52 0.17111f
C6256 single_9b_cdac_1.CF[2] clk 0.09194f
C6257 th_dif_sw_0.VCN ua[0] 0.86465f
C6258 a_12491_27662# sar9b_0.net29 0.22249f
C6259 VDPWR sar9b_0._18_ 1.75124f
C6260 a_11382_23474# a_12047_23853# 0.19065f
C6261 sar9b_0.net43 a_9323_27662# 0.04771f
C6262 sar9b_0.net42 sar9b_0.net5 0.01903f
C6263 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.CKB 4.72443f
C6264 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VDPWR 0.62443f
C6265 a_10644_16791# a_10410_17846# 0.01861f
C6266 sar9b_0.net59 single_9b_cdac_0.SW[7] 0.07361f
C6267 sar9b_0.net49 a_9154_20142# 0.09704f
C6268 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[2] 0.24301f
C6269 VDPWR single_9b_cdac_0.SW[0] 3.07511f
C6270 a_8345_26455# a_9130_26198# 0.26257f
C6271 sar9b_0.net40 sar9b_0.clk_div_0.COUNT\[2\] 0.02492f
C6272 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 1.71649f
C6273 a_4011_22488# a_3027_22138# 0.08669f
C6274 VDPWR a_12870_19603# 0.27172f
C6275 a_10098_19171# sar9b_0.net26 0.06434f
C6276 sar9b_0.net52 sar9b_0.net57 0.87251f
C6277 a_10227_18142# sar9b_0.net73 0.11717f
C6278 a_13011_23238# single_9b_cdac_1.CF[5] 0.35518f
C6279 sar9b_0.net58 uo_out[7] 0.13384f
C6280 VDPWR a_33936_16877# 1.81495f
C6281 a_10607_25185# a_9942_24806# 0.19065f
C6282 a_7882_19538# sar9b_0.net47 0.23112f
C6283 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 2.7611f
C6284 a_9930_20510# a_8970_20510# 0.03529f
C6285 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6286 sar9b_0._07_ sar9b_0._10_ 0.0757f
C6287 a_6922_23534# a_7638_23474# 0.03811f
C6288 a_4922_20857# a_4886_21124# 0.01114f
C6289 sar9b_0.net43 sar9b_0.net59 0.30303f
C6290 sar9b_0.clk_div_0.COUNT\[0\] sar9b_0._02_ 0.06001f
C6291 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN single_9b_cdac_0.cdac_sw_9b_0.S[4] 0.84427f
C6292 a_8595_17910# sar9b_0.net6 0.03608f
C6293 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_55773_15501# 0.01076f
C6294 a_10803_19474# sar9b_0.net48 0.02063f
C6295 sar9b_0.net8 a_11842_19766# 0.02187f
C6296 a_10649_17131# single_9b_cdac_1.SW[1] 0.0197f
C6297 a_6861_22828# sar9b_0.clk_div_0.COUNT\[2\] 0.04796f
C6298 a_9996_16784# sar9b_0.net6 0.05001f
C6299 uio_in[5] uio_in[4] 0.03102f
C6300 a_9472_18823# sar9b_0.net48 0.04471f
C6301 VDPWR a_10858_17113# 0.19951f
C6302 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.cdac_sw_9b_0.S[6] 17.8424f
C6303 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 3.27795f
C6304 a_11430_24931# sar9b_0.net74 0.01382f
C6305 sar9b_0.net29 a_13216_19809# 0.27892f
C6306 a_10553_18922# a_10830_19068# 0.09983f
C6307 a_8340_26115# sar9b_0.net59 0.17782f
C6308 a_4934_22432# sar9b_0.net64 0.25605f
C6309 a_9472_18823# a_9900_19047# 0.01872f
C6310 sar9b_0.net33 a_12182_26419# 0.06698f
C6311 sar9b_0.net51 sar9b_0.net62 0.49495f
C6312 single_9b_cdac_0.SW[8] ua[0] 0.20384f
C6313 sar9b_0.net63 a_7483_23174# 0.01409f
C6314 a_9634_17478# a_10410_17846# 0.3578f
C6315 sar9b_0.net27 a_11842_26426# 0.01173f
C6316 sar9b_0.net9 sar9b_0.net39 0.52789f
C6317 sar9b_0.net26 a_11842_22430# 0.02923f
C6318 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y 0.07579f
C6319 a_6132_23451# a_5823_23477# 0.07766f
C6320 a_5506_17478# a_6282_17846# 0.3578f
C6321 VDPWR a_4072_19474# 0.11411f
C6322 sar9b_0.net44 sar9b_0.net21 0.03003f
C6323 uo_out[2] uo_out[1] 3.05143f
C6324 uo_out[4] ui_in[0] 0.06786f
C6325 VDPWR sar9b_0.net71 0.30617f
C6326 sar9b_0.net30 a_11658_26134# 0.01536f
C6327 sar9b_0.net58 sar9b_0.net68 0.02945f
C6328 sar9b_0.net61 sar9b_0.net39 0.42188f
C6329 sar9b_0.net44 sar9b_0.net39 0.24822f
C6330 VDPWR a_7193_22459# 0.22562f
C6331 VDPWR a_4812_21738# 0.27108f
C6332 a_10166_3438# ua[4] 0.65763f
C6333 sar9b_0.net56 sar9b_0.net35 0.5676f
C6334 sar9b_0.net47 sar9b_0.net4 0.03459f
C6335 a_9942_27470# sar9b_0.net45 0.08179f
C6336 sar9b_0._07_ sar9b_0.net4 0.13017f
C6337 sar9b_0.net11 sar9b_0.net54 0.36694f
C6338 sar9b_0._18_ sar9b_0._17_ 0.19231f
C6339 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 1.71649f
C6340 a_9546_24506# a_9270_24566# 0.1263f
C6341 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A 0.62443f
C6342 a_12491_27662# single_9b_cdac_0.SW[3] 0.38351f
C6343 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A 0.10429f
C6344 single_9b_cdac_1.CF[7] single_9b_cdac_1.SW[2] 0.01297f
C6345 sar9b_0.net18 sar9b_0.net17 0.03659f
C6346 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.CF[6] 0.0313f
C6347 a_3521_24240# sar9b_0.clknet_1_1__leaf_CLK 0.04554f
C6348 VDPWR uio_out[0] 0.76516f
C6349 a_11030_22954# sar9b_0.net2 0.01198f
C6350 dw_12589_1395# a_10482_3438# 0.05479f
C6351 VDPWR a_5753_24250# 0.21444f
C6352 a_30717_29917# single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A 0.01076f
C6353 VDPWR a_4332_23043# 1.38139f
C6354 sar9b_0._01_ sar9b_0._07_ 0.14158f
C6355 sar9b_0.net13 sar9b_0.net42 0.02401f
C6356 a_6783_19481# sar9b_0.net40 0.05886f
C6357 VDPWR a_12618_26134# 0.35483f
C6358 a_11859_17910# single_9b_cdac_1.SW[4] 0.35232f
C6359 VDPWR a_6534_27123# 0.27103f
C6360 a_6282_27170# sar9b_0.net37 0.06133f
C6361 sar9b_0._08_ sar9b_0._18_ 0.02837f
C6362 single_9b_cdac_1.CF[1] single_9b_cdac_1.SW[8] 0.03927f
C6363 a_8052_18123# a_8057_18463# 0.44098f
C6364 sar9b_0.net29 single_9b_cdac_0.SW[0] 0.03951f
C6365 sar9b_0.net30 sar9b_0.net26 0.11005f
C6366 a_5196_18116# a_5394_18116# 0.06623f
C6367 sar9b_0.net63 sar9b_0.clk_div_0.COUNT\[0\] 0.2165f
C6368 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.08121f
C6369 a_7404_16784# a_7743_16817# 0.07649f
C6370 a_8052_16791# a_7602_16784# 0.03471f
C6371 a_6678_27470# a_6954_27466# 0.1263f
C6372 sar9b_0.net35 a_6902_25087# 0.0142f
C6373 sar9b_0.net2 a_10803_18142# 0.0218f
C6374 single_9b_cdac_1.cdac_sw_9b_0.S[8] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.22655f
C6375 sar9b_0.net41 sar9b_0.net73 0.0295f
C6376 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[0] 0.36674f
C6377 sar9b_0.net7 sar9b_0.net39 0.0839f
C6378 sar9b_0.net53 a_12047_23853# 0.22582f
C6379 sar9b_0.net57 a_8591_22855# 0.01229f
C6380 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.69086f
C6381 a_10402_21098# a_11178_20806# 0.3578f
C6382 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.12431f
C6383 a_11382_22142# a_11842_22430# 0.26257f
C6384 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C6385 a_10623_25895# a_10937_25582# 0.07826f
C6386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A 0.42509f
C6387 a_7338_24802# sar9b_0.net54 0.26564f
C6388 a_10230_23234# sar9b_0.net11 0.04733f
C6389 a_6282_17846# a_5322_17846# 0.03529f
C6390 a_9258_21842# a_9647_21523# 0.05462f
C6391 a_8982_21902# a_9442_21474# 0.26257f
C6392 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP ua[0] 1.14952f
C6393 a_11658_26134# a_12047_26517# 0.06034f
C6394 a_10859_26330# single_9b_cdac_0.SW[7] 0.37246f
C6395 single_9b_cdac_0.SW[5] sar9b_0.net14 0.06325f
C6396 sar9b_0.net27 sar9b_0.net11 0.03459f
C6397 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 2.7611f
C6398 a_8098_23762# sar9b_0.net54 0.02919f
C6399 sar9b_0._07_ a_3795_19512# 0.11659f
C6400 sar9b_0.net57 a_5196_18116# 0.09147f
C6401 sar9b_0.net43 a_9942_24806# 0.01787f
C6402 a_6738_22112# a_7193_22459# 0.3578f
C6403 a_7188_22119# a_7978_22202# 0.1263f
C6404 VDPWR sar9b_0.net72 0.65198f
C6405 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[8] 1.41793f
C6406 a_10858_17113# sar9b_0.net48 0.12168f
C6407 single_9b_cdac_0.SW[7] ua[0] 0.25507f
C6408 a_5374_20145# a_5481_20185# 0.14439f
C6409 sar9b_0.net41 sar9b_0.net6 0.02799f
C6410 sar9b_0.net31 a_11382_26138# 0.01042f
C6411 sar9b_0._08_ a_4072_19474# 0.09389f
C6412 a_10254_2858# ua[4] 0.12559f
C6413 a_9323_28371# single_9b_cdac_0.SW[8] 0.0233f
C6414 sar9b_0._09_ sar9b_0.net46 0.01177f
C6415 sar9b_0._08_ sar9b_0.net71 0.35019f
C6416 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A 0.42509f
C6417 ui_in[0] th_dif_sw_0.VCN 0.22659f
C6418 VDPWR a_10830_19068# 0.26619f
C6419 a_3206_22432# sar9b_0.net65 0.02448f
C6420 VDPWR sar9b_0.net64 0.46487f
C6421 sar9b_0.net56 a_9363_20826# 0.12663f
C6422 single_9b_cdac_0.SW[5] th_dif_sw_0.VCN 0.09454f
C6423 a_10644_16791# a_11008_17491# 0.0165f
C6424 a_9942_20810# a_10402_21098# 0.26257f
C6425 a_10378_27170# sar9b_0.net45 0.05318f
C6426 a_7890_26108# a_8340_26115# 0.03529f
C6427 a_8031_26141# a_7692_26108# 0.07649f
C6428 single_9b_cdac_0.cdac_sw_9b_0.S[5] ua[0] 1.56372f
C6429 sar9b_0.net17 a_2847_27473# 0.02024f
C6430 a_8074_20870# sar9b_0.net9 0.16977f
C6431 a_8098_18810# sar9b_0.net61 0.02618f
C6432 sar9b_0.net9 sar9b_0.net53 0.14548f
C6433 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VDPWR 0.62443f
C6434 sar9b_0.net8 a_11382_19478# 0.03762f
C6435 single_9b_cdac_0.SW[3] single_9b_cdac_0.SW[0] 0.01042f
C6436 single_9b_cdac_1.SW[5] th_dif_sw_0.CK 0.23096f
C6437 sar9b_0.net35 sar9b_0.net60 0.02971f
C6438 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[0] 4.151f
C6439 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_1.CF[3] 0.31534f
C6440 a_8074_20870# sar9b_0.net61 0.0249f
C6441 a_4083_28566# uio_out[0] 0.37232f
C6442 a_7092_19455# sar9b_0.net51 0.02272f
C6443 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[6] 0.01482f
C6444 a_16159_13315# tdc_0.phase_detector_0.pd_out_0.B 0.38171f
C6445 sar9b_0._07_ sar9b_0.clknet_1_1__leaf_CLK 0.02605f
C6446 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.27795f
C6447 a_9126_23599# a_8874_23470# 0.27388f
C6448 VDPWR a_11430_20935# 0.27331f
C6449 sar9b_0.net74 a_11214_25728# 0.06877f
C6450 sar9b_0.net41 single_9b_cdac_1.SW[3] 0.03054f
C6451 single_9b_cdac_1.cdac_sw_9b_0.S[0] single_9b_cdac_1.cdac_sw_9b_0.S[2] 0.70254f
C6452 a_21684_3438# dw_17224_1400# 0.05479f
C6453 sar9b_0.net13 sar9b_0.net74 0.34392f
C6454 a_10378_27170# a_9870_27060# 0.19065f
C6455 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A 0.62443f
C6456 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 single_9b_cdac_1.SW[4] 0.24199f
C6457 a_5100_24375# a_4467_24162# 0.01351f
C6458 sar9b_0.net35 sar9b_0.net57 0.03434f
C6459 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 3.27833f
C6460 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 ua[0] 0.12358f
C6461 a_7590_24931# a_6378_24802# 0.07766f
C6462 sar9b_0.net60 a_5742_28392# 0.06229f
C6463 a_33936_16877# single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 0.23864f
C6464 sar9b_0.net47 sar9b_0.net55 0.03364f
C6465 a_11776_25137# sar9b_0.net12 0.07772f
C6466 sar9b_0._07_ sar9b_0.net55 0.01037f
C6467 single_9b_cdac_0.SW[5] single_9b_cdac_0.SW[8] 0.05858f
C6468 sar9b_0.net41 a_9154_20142# 0.02308f
C6469 sar9b_0.net8 a_10402_21098# 0.16495f
C6470 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A 0.69086f
C6471 VDPWR a_5628_19768# 0.19326f
C6472 a_14871_9671# th_dif_sw_0.VCP 0.07081f
C6473 single_9b_cdac_0.cdac_sw_9b_0.S[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 0.84427f
C6474 VDPWR a_7289_21127# 0.22771f
C6475 th_dif_sw_0.CKB single_9b_cdac_1.SW[0] 0.0171f
C6476 sar9b_0.net28 clk 0.52609f
C6477 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A 0.95338f
C6478 VDPWR a_6767_25185# 0.26598f
C6479 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.7611f
C6480 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y 0.07517f
C6481 sar9b_0.net36 sar9b_0.net11 0.02201f
C6482 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP 0.19266f
C6483 a_9165_24988# sar9b_0.net37 0.01216f
C6484 ui_in[0] ui_in[1] 0.03102f
C6485 sar9b_0._12_ sar9b_0.net69 0.23206f
C6486 a_7404_17715# sar9b_0.net35 0.03641f
C6487 VDPWR a_8874_23470# 0.39649f
C6488 sar9b_0.net64 sar9b_0._17_ 0.0131f
C6489 clk single_9b_cdac_1.SW[7] 0.08277f
C6490 single_9b_cdac_1.cdac_sw_9b_0.S[4] single_9b_cdac_1.cdac_sw_9b_0.S[0] 0.43767f
C6491 a_9126_23599# sar9b_0.net37 0.02665f
C6492 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A 0.75849f
C6493 a_4934_22432# sar9b_0._07_ 0.01085f
C6494 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.45521f
C6495 a_4018_24235# sar9b_0.clk_div_0.COUNT\[2\] 0.15815f
C6496 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 0.02618f
C6497 VDPWR a_3521_24240# 0.10938f
C6498 sar9b_0._10_ a_4496_20468# 0.16691f
C6499 a_7284_20787# sar9b_0.net51 0.07994f
C6500 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 0.19266f
C6501 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C6502 a_12588_16784# a_13011_16810# 0.05125f
C6503 VDPWR a_38738_26999# 1.81495f
C6504 sar9b_0.net5 sar9b_0.net39 0.02145f
C6505 a_10858_17113# a_10926_17021# 0.35559f
C6506 single_9b_cdac_1.CF[2] single_9b_cdac_1.cdac_sw_9b_0.S[1] 0.01515f
C6507 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN 2.82172f
C6508 a_30012_17740# single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.22513f
C6509 a_10402_25094# a_11430_24931# 0.07826f
C6510 sar9b_0._18_ sar9b_0._12_ 0.02191f
C6511 a_10830_19068# sar9b_0.net48 0.22344f
C6512 sar9b_0.net40 sar9b_0.net35 0.52689f
C6513 a_8694_20570# sar9b_0.net37 0.01919f
C6514 single_9b_cdac_1.CF[4] th_dif_sw_0.VCN 0.09453f
C6515 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A single_9b_cdac_1.CF[5] 0.06019f
C6516 single_9b_cdac_0.SW[2] single_9b_cdac_0.cdac_sw_9b_0.S[2] 0.22543f
C6517 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP 0.10499f
C6518 sar9b_0.cyclic_flag_0.FINAL a_8940_27039# 0.01546f
C6519 a_10553_18922# a_10098_19171# 0.3578f
C6520 single_9b_cdac_1.CF[3] clk 0.109f
C6521 sar9b_0.net43 sar9b_0.net54 0.53075f
C6522 a_5298_24499# sar9b_0.net54 0.25564f
C6523 sar9b_0.net41 a_11436_17742# 0.07436f
C6524 sar9b_0.net40 sar9b_0.net2 0.02933f
C6525 sar9b_0.clk_div_0.COUNT\[2\] clk 0.11336f
C6526 VDPWR sar9b_0.net37 2.42386f
C6527 a_2508_20780# a_2739_20140# 0.01678f
C6528 single_9b_cdac_1.cdac_sw_9b_0.S[5] a_38738_16877# 0.59531f
C6529 sar9b_0.net52 a_11178_24802# 0.24274f
C6530 a_6880_26815# a_6282_27170# 0.06623f
C6531 a_4330_27170# sar9b_0.net37 0.17592f
C6532 sar9b_0.net8 a_8970_20510# 0.23591f
C6533 a_4072_19474# a_3991_19768# 0.03072f
C6534 a_3795_19512# a_4292_19768# 0.02251f
C6535 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 0.02813f
C6536 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C6537 a_10218_27466# a_11178_27466# 0.03432f
C6538 a_6132_23451# sar9b_0.net54 0.17758f
C6539 a_8166_27595# sar9b_0.net45 0.03834f
C6540 VDPWR a_3438_27677# 0.25451f
C6541 single_9b_cdac_1.CF[3] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17948f
C6542 sar9b_0.net68 sar9b_0.clk_div_0.COUNT\[1\] 0.35672f
C6543 sar9b_0.net1 sar9b_0.net37 0.27714f
C6544 sar9b_0.net6 a_12435_20806# 0.19538f
C6545 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP single_9b_cdac_1.CF[2] 0.19321f
C6546 VDPWR a_9802_26815# 0.20303f
C6547 sar9b_0.net20 sar9b_0.net58 0.46059f
C6548 a_5465_28246# a_5674_28147# 0.24088f
C6549 a_5460_28377# sar9b_0.net45 0.20577f
C6550 single_9b_cdac_1.SW[3] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP 0.17185f
C6551 VDPWR a_8202_23174# 0.87317f
C6552 a_3370_27769# a_3438_27677# 0.35559f
C6553 sar9b_0.net32 a_11842_26426# 0.01684f
C6554 sar9b_0.net42 a_11339_27039# 0.01795f
C6555 a_10607_25185# sar9b_0.net36 0.02216f
C6556 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP 3.27843f
C6557 sar9b_0.net3 a_2547_28132# 0.27678f
C6558 sar9b_0.net36 single_9b_cdac_0.SW[8] 0.07497f
C6559 sar9b_0.net49 a_9258_21842# 0.19249f
C6560 sar9b_0.net26 sar9b_0.net27 0.67638f
C6561 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C6562 single_9b_cdac_0.SW[7] single_9b_cdac_0.SW[5] 0.11961f
C6563 single_9b_cdac_1.SW[4] sar9b_0.net39 0.01225f
C6564 a_8098_18810# a_8438_18958# 0.24088f
C6565 sar9b_0.net57 a_7914_23470# 0.22944f
C6566 sar9b_0.net57 a_7978_22202# 0.01265f
C6567 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 2.7611f
C6568 single_9b_cdac_1.SW[2] a_9450_17846# 0.01334f
C6569 sar9b_0.net27 a_13011_20806# 0.04065f
C6570 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A 0.12431f
C6571 sar9b_0.net52 clk 0.01379f
C6572 single_9b_cdac_0.SW[7] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 0.36542f
C6573 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.62443f
C6574 sar9b_0.net54 sar9b_0.net4 0.17203f
C6575 sar9b_0.net56 single_9b_cdac_1.SW[0] 0.04752f
C6576 single_9b_cdac_0.cdac_sw_9b_0.S[5] single_9b_cdac_0.SW[5] 0.22549f
C6577 a_9942_20810# a_10607_21189# 0.19065f
C6578 sar9b_0._15_ sar9b_0.net54 0.08938f
C6579 single_9b_cdac_1.CF[6] single_9b_cdac_1.SW[1] 0.22097f
C6580 VDPWR single_9b_cdac_1.CF[5] 2.58659f
C6581 a_7092_19455# a_6642_19448# 0.03471f
C6582 single_9b_cdac_1.CF[8] single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y 0.12898f
C6583 a_21368_4076# th_dif_sw_0.th_sw_1.CK 0.0478f
C6584 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08121f
C6585 a_5010_28495# a_5151_28559# 0.27388f
C6586 a_5753_24250# a_6030_24396# 0.09983f
C6587 VDPWR sar9b_0.net25 0.46378f
C6588 VDPWR a_9323_27662# 0.45921f
C6589 VDPWR sar9b_0.net47 2.56257f
C6590 a_4018_24235# a_2835_24136# 0.0649f
C6591 a_3819_24136# a_3014_24136# 0.29221f
C6592 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 single_9b_cdac_1.SW[7] 0.363f
C6593 VDPWR sar9b_0._07_ 0.94013f
C6594 sar9b_0.net24 sar9b_0.net37 0.25988f
C6595 a_5506_17478# sar9b_0.net46 0.1904f
C6596 a_13011_23238# sar9b_0.net27 0.04162f
C6597 sar9b_0.net63 a_6414_23681# 0.04702f
C6598 a_12618_26134# a_13216_26469# 0.06623f
C6599 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 single_9b_cdac_0.cdac_sw_9b_0.S[6] 0.36006f
C6600 a_8334_17021# sar9b_0.net61 0.06633f
C6601 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 2.82172f
C6602 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP single_9b_cdac_1.CF[2] 0.10503f
C6603 a_10690_22806# clk 0.02916f
C6604 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.CF[5] 0.42014f
C6605 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y single_9b_cdac_1.CF[7] 0.17948f
C6606 single_9b_cdac_0.cdac_sw_9b_0.S[6] a_34814_26990# 0.22352f
C6607 a_8098_18810# sar9b_0.net5 0.01301f
C6608 sar9b_0.net51 a_6579_18832# 0.26023f
C6609 sar9b_0.net58 a_6250_28502# 0.20323f
C6610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A 0.12431f
C6611 sar9b_0.net24 a_9802_26815# 0.01411f
C6612 a_7404_16784# sar9b_0.net27 0.02142f
C6613 a_8334_18353# sar9b_0.net61 0.02726f
C6614 sar9b_0.net59 sar9b_0.net38 0.05434f
C6615 single_9b_cdac_1.SW[8] single_9b_cdac_1.SW[2] 0.21903f
C6616 a_9138_27163# a_9588_27045# 0.03432f
C6617 VDPWR sar9b_0.net59 4.515f
C6618 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 1.71649f
C6619 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN 0.17533f
C6620 a_10098_19171# sar9b_0.net38 0.02641f
C6621 sar9b_0.net48 sar9b_0.net37 0.18456f
C6622 th_dif_sw_0.CK sar9b_0.net27 0.02592f
C6623 sar9b_0.net63 a_2893_24992# 0.0883f
C6624 VDPWR a_10098_19171# 0.35321f
C6625 a_6307_27584# sar9b_0.net44 0.23235f
C6626 a_11842_19766# sar9b_0.net6 0.01376f
C6627 a_11842_18434# a_12870_18271# 0.07826f
C6628 sar9b_0.net3 ui_in[0] 0.05952f
C6629 a_13011_21906# a_13011_20806# 0.0246f
C6630 sar9b_0.net32 sar9b_0.net14 0.14467f
C6631 VDPWR single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.62555f
C6632 VDPWR single_9b_cdac_0.cdac_sw_9b_0.S[6] 4.16175f
C6633 VDPWR a_5823_23477# 0.26508f
C6634 a_9900_19047# sar9b_0.net37 0.27085f
C6635 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C6636 sar9b_0.net32 sar9b_0.net11 0.02514f
C6637 a_8940_24402# sar9b_0.net62 0.23108f
C6638 sar9b_0.net10 sar9b_0.net73 0.07697f
C6639 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.12223f
C6640 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP single_9b_cdac_1.CF[6] 0.10499f
C6641 sar9b_0.net8 a_10607_21189# 0.01911f
C6642 sar9b_0.net27 sar9b_0.net4 0.23295f
C6643 VDPWR single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A 0.38397f
C6644 single_9b_cdac_1.CF[8] th_dif_sw_0.VCN 0.09453f
C6645 sar9b_0.net64 a_5523_21528# 0.03232f
C6646 sar9b_0.net61 a_9450_17846# 0.04773f
C6647 sar9b_0.net12 a_11842_26426# 0.02738f
C6648 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP 1.56037f
C6649 a_7566_21017# a_7284_20787# 0.05462f
C6650 th_dif_sw_0.th_sw_1.CK a_10166_3438# 0.04891f
C6651 sar9b_0.net61 single_9b_cdac_1.SW[2] 0.04325f
C6652 a_10644_16791# a_10649_17131# 0.43869f
C6653 single_9b_cdac_1.SW[4] single_9b_cdac_1.CF[7] 0.01482f
C6654 VDPWR a_7602_18116# 0.3287f
C6655 sar9b_0.net26 sar9b_0.net36 0.0273f
C6656 single_9b_cdac_0.SW[7] sar9b_0.net36 0.33484f
C6657 VDPWR a_7743_16817# 0.26065f
C6658 single_9b_cdac_1.SW[6] single_9b_cdac_1.CF[6] 2.01497f
C6659 a_15400_11316# tdc_0.phase_detector_0.INP 0.02415f
C6660 sar9b_0.net64 sar9b_0._12_ 0.3293f
C6661 a_11466_23174# sar9b_0.net42 0.01972f
C6662 sar9b_0.net19 a_5322_27170# 0.02142f
C6663 VDPWR a_11842_22430# 0.22622f
C6664 a_6975_20813# sar9b_0.net10 0.03184f
C6665 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A 0.11216f
C6666 sar9b_0.net13 a_10402_25094# 0.01895f
C6667 a_7602_18116# sar9b_0.net1 0.03058f
C6668 single_9b_cdac_1.cdac_sw_9b_0.S[6] single_9b_cdac_1.SW[6] 0.22497f
C6669 a_6102_24806# a_6378_24802# 0.1263f
C6670 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A 0.42784f
C6671 a_8883_27466# a_9323_27662# 0.03138f
C6672 sar9b_0.net58 sar9b_0.net19 0.19557f
C6673 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN single_9b_cdac_1.cdac_sw_9b_0.S[7] 0.84426f
C6674 a_5322_17846# sar9b_0.net46 0.23175f
C6675 single_9b_cdac_1.CF[5] sar9b_0.net29 0.09978f
C6676 single_9b_cdac_1.CF[0] single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A 0.02149f
C6677 sar9b_0.net43 sar9b_0.net36 0.11895f
C6678 sar9b_0._07_ sar9b_0._17_ 0.02418f
C6679 a_11842_19766# sar9b_0.net50 0.10082f
C6680 a_6738_22112# sar9b_0.net47 0.26419f
C6681 sar9b_0.net54 a_5748_24381# 0.18387f
C6682 a_2739_20140# a_3723_20140# 0.08669f
C6683 sar9b_0._00_ a_3273_20185# 0.04988f
C6684 a_8591_22855# clk 0.02075f
C6685 sar9b_0.net31 a_12618_22138# 0.06744f
C6686 sar9b_0.net36 a_10035_19474# 0.01195f
C6687 a_5441_22522# sar9b_0._07_ 0.02011f
C6688 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.6919f
C6689 VDPWR a_3166_20145# 0.02403f
C6690 a_7188_22119# sar9b_0.net57 0.01211f
C6691 sar9b_0._02_ sar9b_0.net39 0.04135f
C6692 ua[1] VGND 0.14595f
C6693 ua[2] VGND 0.14595f
C6694 ua[5] VGND 0.14595f
C6695 ua[6] VGND 0.14595f
C6696 ua[7] VGND 0.14595f
C6697 ena VGND 0.06982f
C6698 rst_n VGND 0.04231f
C6699 ui_in[1] VGND 0.04231f
C6700 ui_in[2] VGND 0.04231f
C6701 ui_in[3] VGND 0.04231f
C6702 ui_in[4] VGND 0.04231f
C6703 ui_in[5] VGND 0.04231f
C6704 ui_in[6] VGND 0.04231f
C6705 ui_in[7] VGND 0.04231f
C6706 uio_in[0] VGND 0.04231f
C6707 uio_in[1] VGND 0.04231f
C6708 uio_in[2] VGND 0.04231f
C6709 uio_in[3] VGND 0.04231f
C6710 uio_in[4] VGND 0.04231f
C6711 uio_in[5] VGND 0.04231f
C6712 uio_in[6] VGND 0.04231f
C6713 uio_in[7] VGND 0.04264f
C6714 ua[3] VGND 13.5574f
C6715 ua[4] VGND 13.4686f
C6716 clk VGND 28.193f
C6717 ui_in[0] VGND 17.1737f
C6718 uo_out[7] VGND 5.41879f
C6719 uo_out[1] VGND 4.49964f
C6720 uo_out[0] VGND 6.32256f
C6721 uo_out[2] VGND 4.375f
C6722 uo_out[3] VGND 4.4898f
C6723 uo_out[4] VGND 4.97269f
C6724 uo_out[6] VGND 5.39467f
C6725 uo_out[5] VGND 5.08381f
C6726 uio_out[0] VGND 5.71643f
C6727 uio_out[1] VGND 7.50245f
C6728 ua[0] VGND 0.11733p
C6729 VDPWR VGND 0.97985p
C6730 m2_23774_17236# VGND 0.24462f
C6731 m2_23774_26966# VGND 0.24462f
C6732 a_18214_3039# VGND 1.49705f $ **FLOATING
C6733 a_21684_3438# VGND 4.00493f $ **FLOATING
C6734 a_21368_4076# VGND 15.5335f $ **FLOATING
C6735 a_10254_2858# VGND 1.4958f $ **FLOATING
C6736 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VGND 3.32878f $ **FLOATING
C6737 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VGND 3.32496f $ **FLOATING
C6738 a_10482_3438# VGND 4.00493f $ **FLOATING
C6739 a_10166_3438# VGND 16.0184f $ **FLOATING
C6740 th_dif_sw_0.th_sw_1.CKB VGND 8.08199f $ **FLOATING
C6741 th_dif_sw_0.th_sw_1.CK VGND 9.07818f $ **FLOATING
C6742 a_21177_7457# VGND 2.80515f $ **FLOATING
C6743 a_9132_7271# VGND 2.80492f $ **FLOATING
C6744 a_17125_9355# VGND 0.09476f $ **FLOATING
C6745 a_14897_9355# VGND 0.09476f $ **FLOATING
C6746 th_dif_sw_0.VCP VGND 55.6678f $ **FLOATING
C6747 th_dif_sw_0.VCN VGND 67.3957f $ **FLOATING
C6748 a_16357_9613# VGND 0.05938f $ **FLOATING
C6749 a_15265_9613# VGND 0.05938f $ **FLOATING
C6750 a_16331_9671# VGND 0.82151f $ **FLOATING
C6751 a_14871_9671# VGND 0.82187f $ **FLOATING
C6752 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VGND 0.66688f $ **FLOATING
C6753 a_16881_10256# VGND 0.01123f $ **FLOATING
C6754 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VGND 0.66603f $ **FLOATING
C6755 a_15197_10290# VGND 0.01123f $ **FLOATING
C6756 a_16527_10454# VGND 0.18095f $ **FLOATING
C6757 a_15151_10456# VGND 0.18103f $ **FLOATING
C6758 a_16222_11316# VGND 0.04271f $ **FLOATING
C6759 a_15400_11316# VGND 0.04271f $ **FLOATING
C6760 tdc_0.phase_detector_0.INP VGND 1.24598f $ **FLOATING
C6761 tdc_0.phase_detector_0.INN VGND 1.87249f $ **FLOATING
C6762 a_16970_11404# VGND 0.20846f $ **FLOATING
C6763 a_15052_11404# VGND 0.20846f $ **FLOATING
C6764 tdc_0.phase_detector_0.pd_out_0.A VGND 2.40659f $ **FLOATING
C6765 tdc_0.phase_detector_0.pd_out_0.B VGND 1.65957f $ **FLOATING
C6766 a_16159_13315# VGND 0.26136f $ **FLOATING
C6767 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6768 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.41378f $ **FLOATING
C6769 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6770 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.45426f $ **FLOATING
C6771 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6772 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND 1.60512f $ **FLOATING
C6773 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND 1.57322f $ **FLOATING
C6774 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.39423f $ **FLOATING
C6775 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6776 a_63626_17740# VGND 0.89497f $ **FLOATING
C6777 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND 2.68117f $ **FLOATING
C6778 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6779 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6780 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6781 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6782 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6783 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND 3.19276f $ **FLOATING
C6784 a_62748_16877# VGND 0.16243f $ **FLOATING
C6785 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6786 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6787 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND 4.52812f $ **FLOATING
C6788 single_9b_cdac_1.cdac_sw_9b_0.S[0] VGND 94.0914f $ **FLOATING
C6789 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6790 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6791 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND 6.36367f $ **FLOATING
C6792 a_58824_17740# VGND 0.89548f $ **FLOATING
C6793 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND 2.66663f $ **FLOATING
C6794 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6795 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.405f $ **FLOATING
C6796 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6797 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44881f $ **FLOATING
C6798 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6799 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND 3.16257f $ **FLOATING
C6800 a_57946_16877# VGND 0.16243f $ **FLOATING
C6801 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND 1.58431f $ **FLOATING
C6802 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND 1.56057f $ **FLOATING
C6803 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND 4.51086f $ **FLOATING
C6804 single_9b_cdac_1.cdac_sw_9b_0.S[1] VGND 47.9165f $ **FLOATING
C6805 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37225f $ **FLOATING
C6806 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6807 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND 6.34714f $ **FLOATING
C6808 a_54032_17740# VGND 0.89543f $ **FLOATING
C6809 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND 2.66664f $ **FLOATING
C6810 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6811 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40542f $ **FLOATING
C6812 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6813 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44912f $ **FLOATING
C6814 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6815 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND 3.16256f $ **FLOATING
C6816 a_53154_16877# VGND 0.16243f $ **FLOATING
C6817 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND 1.58193f $ **FLOATING
C6818 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND 1.56099f $ **FLOATING
C6819 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND 4.51373f $ **FLOATING
C6820 single_9b_cdac_1.cdac_sw_9b_0.S[2] VGND 30.3253f $ **FLOATING
C6821 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37352f $ **FLOATING
C6822 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6823 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND 6.34762f $ **FLOATING
C6824 a_49221_17740# VGND 0.89502f $ **FLOATING
C6825 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND 2.66535f $ **FLOATING
C6826 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6827 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40525f $ **FLOATING
C6828 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6829 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44899f $ **FLOATING
C6830 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6831 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND 3.16312f $ **FLOATING
C6832 a_48343_16877# VGND 0.16243f $ **FLOATING
C6833 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND 1.58513f $ **FLOATING
C6834 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND 1.56081f $ **FLOATING
C6835 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND 4.51233f $ **FLOATING
C6836 single_9b_cdac_1.cdac_sw_9b_0.S[3] VGND 21.4947f $ **FLOATING
C6837 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37301f $ **FLOATING
C6838 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6839 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND 6.3477f $ **FLOATING
C6840 a_44418_17740# VGND 0.89497f $ **FLOATING
C6841 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND 2.665f $ **FLOATING
C6842 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6843 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6844 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6845 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6846 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6847 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND 3.16281f $ **FLOATING
C6848 a_43540_16877# VGND 0.16243f $ **FLOATING
C6849 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6850 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6851 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND 4.51195f $ **FLOATING
C6852 single_9b_cdac_1.cdac_sw_9b_0.S[4] VGND 20.61f $ **FLOATING
C6853 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6854 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6855 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6856 a_39616_17740# VGND 0.89497f $ **FLOATING
C6857 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND 2.66616f $ **FLOATING
C6858 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6859 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6860 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6861 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6862 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6863 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6864 a_38738_16877# VGND 0.16243f $ **FLOATING
C6865 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6866 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6867 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND 4.51201f $ **FLOATING
C6868 single_9b_cdac_1.cdac_sw_9b_0.S[5] VGND 16.1449f $ **FLOATING
C6869 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6870 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6871 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6872 a_34814_17740# VGND 0.89548f $ **FLOATING
C6873 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND 2.66683f $ **FLOATING
C6874 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6875 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6876 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6877 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6878 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6879 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6880 a_33936_16877# VGND 0.16243f $ **FLOATING
C6881 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6882 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6883 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND 4.51252f $ **FLOATING
C6884 single_9b_cdac_1.cdac_sw_9b_0.S[6] VGND 15.6371f $ **FLOATING
C6885 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6886 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6887 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND 6.3475f $ **FLOATING
C6888 a_30012_17740# VGND 0.89497f $ **FLOATING
C6889 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND 2.66498f $ **FLOATING
C6890 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C6891 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C6892 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C6893 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C6894 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C6895 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND 3.16277f $ **FLOATING
C6896 a_29134_16877# VGND 0.16243f $ **FLOATING
C6897 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C6898 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C6899 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND 4.51193f $ **FLOATING
C6900 single_9b_cdac_1.cdac_sw_9b_0.S[7] VGND 14.5496f $ **FLOATING
C6901 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37294f $ **FLOATING
C6902 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C6903 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND 6.34748f $ **FLOATING
C6904 a_25210_17740# VGND 0.89548f $ **FLOATING
C6905 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND 2.68106f $ **FLOATING
C6906 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND 3.16216f $ **FLOATING
C6907 a_24332_16877# VGND 0.16243f $ **FLOATING
C6908 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND 4.71828f $ **FLOATING
C6909 single_9b_cdac_1.SW[5] VGND 6.60196f $ **FLOATING
C6910 a_13011_16810# VGND 0.63654f $ **FLOATING
C6911 tdc_0.OUTP VGND 3.42864f $ **FLOATING
C6912 a_12588_16784# VGND 0.3641f $ **FLOATING
C6913 a_11434_16874# VGND 0.16615f $ **FLOATING
C6914 a_10926_17021# VGND 0.17322f $ **FLOATING
C6915 a_10858_17113# VGND 0.13557f $ **FLOATING
C6916 a_10649_17131# VGND 0.93597f $ **FLOATING
C6917 a_10335_16817# VGND 0.30597f $ **FLOATING
C6918 a_10194_16784# VGND 0.35867f $ **FLOATING
C6919 a_10644_16791# VGND 0.61756f $ **FLOATING
C6920 a_9996_16784# VGND 0.3018f $ **FLOATING
C6921 a_8842_16874# VGND 0.13599f $ **FLOATING
C6922 a_8334_17021# VGND 0.17338f $ **FLOATING
C6923 a_8266_17113# VGND 0.13376f $ **FLOATING
C6924 a_8057_17131# VGND 0.92848f $ **FLOATING
C6925 a_7743_16817# VGND 0.30616f $ **FLOATING
C6926 a_7602_16784# VGND 0.36252f $ **FLOATING
C6927 a_8052_16791# VGND 0.6075f $ **FLOATING
C6928 a_7404_16784# VGND 0.30035f $ **FLOATING
C6929 a_6867_16810# VGND 0.38007f $ **FLOATING
C6930 tdc_0.OUTN VGND 5.01507f $ **FLOATING
C6931 a_5331_16810# VGND 0.38321f $ **FLOATING
C6932 tdc_0.RDY VGND 6.15869f $ **FLOATING
C6933 th_dif_sw_0.CKB VGND 16.3637f $ **FLOATING
C6934 a_2603_17006# VGND 0.67873f $ **FLOATING
C6935 single_9b_cdac_1.cdac_sw_9b_0.S[8] VGND 13.6188f $ **FLOATING
C6936 single_9b_cdac_1.SW[6] VGND 6.72589f $ **FLOATING
C6937 a_13011_17910# VGND 0.63061f $ **FLOATING
C6938 single_9b_cdac_1.SW[4] VGND 6.88153f $ **FLOATING
C6939 a_11859_17910# VGND 0.6882f $ **FLOATING
C6940 a_11436_17742# VGND 0.33062f $ **FLOATING
C6941 a_11008_17491# VGND 0.27893f $ **FLOATING
C6942 a_10662_17799# VGND 0.29366f $ **FLOATING
C6943 a_10410_17846# VGND 0.34331f $ **FLOATING
C6944 a_9974_17626# VGND 0.1176f $ **FLOATING
C6945 a_9839_17527# VGND 0.15642f $ **FLOATING
C6946 a_9634_17478# VGND 0.88707f $ **FLOATING
C6947 a_9174_17906# VGND 0.1327f $ **FLOATING
C6948 a_9450_17846# VGND 0.59308f $ **FLOATING
C6949 single_9b_cdac_1.SW[0] VGND 15.1733f $ **FLOATING
C6950 single_9b_cdac_1.SW[2] VGND 7.72854f $ **FLOATING
C6951 a_8595_17910# VGND 0.5964f $ **FLOATING
C6952 a_8019_17910# VGND 0.60315f $ **FLOATING
C6953 a_7404_17715# VGND 0.24299f $ **FLOATING
C6954 a_6880_17491# VGND 0.29519f $ **FLOATING
C6955 a_6534_17799# VGND 0.31348f $ **FLOATING
C6956 a_6282_17846# VGND 0.36418f $ **FLOATING
C6957 a_5846_17626# VGND 0.1724f $ **FLOATING
C6958 a_5711_17527# VGND 0.19862f $ **FLOATING
C6959 a_5506_17478# VGND 0.95291f $ **FLOATING
C6960 a_5046_17906# VGND 0.14415f $ **FLOATING
C6961 a_5322_17846# VGND 0.6425f $ **FLOATING
C6962 single_9b_cdac_1.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND 6.37641f $ **FLOATING
C6963 a_12047_18525# VGND 0.1897f $ **FLOATING
C6964 a_13216_18477# VGND 0.28599f $ **FLOATING
C6965 a_12618_18142# VGND 0.35255f $ **FLOATING
C6966 a_12870_18271# VGND 0.29854f $ **FLOATING
C6967 a_12182_18427# VGND 0.1325f $ **FLOATING
C6968 a_11842_18434# VGND 0.9417f $ **FLOATING
C6969 a_11658_18142# VGND 0.67802f $ **FLOATING
C6970 a_11382_18146# VGND 0.1608f $ **FLOATING
C6971 single_9b_cdac_1.SW[3] VGND 8.35662f $ **FLOATING
C6972 th_dif_sw_0.CK VGND 10.2695f $ **FLOATING
C6973 a_10803_18142# VGND 0.61263f $ **FLOATING
C6974 a_10227_18142# VGND 0.62055f $ **FLOATING
C6975 a_8842_18206# VGND 0.12267f $ **FLOATING
C6976 a_8334_18353# VGND 0.15504f $ **FLOATING
C6977 a_8266_18445# VGND 0.11469f $ **FLOATING
C6978 a_8057_18463# VGND 0.88109f $ **FLOATING
C6979 a_7743_18149# VGND 0.29328f $ **FLOATING
C6980 a_7602_18116# VGND 0.33292f $ **FLOATING
C6981 a_8052_18123# VGND 0.56532f $ **FLOATING
C6982 a_7404_18116# VGND 0.27413f $ **FLOATING
C6983 a_6634_18206# VGND 0.15117f $ **FLOATING
C6984 a_6126_18353# VGND 0.19104f $ **FLOATING
C6985 a_6058_18445# VGND 0.16799f $ **FLOATING
C6986 a_5849_18463# VGND 0.98369f $ **FLOATING
C6987 a_5535_18149# VGND 0.31139f $ **FLOATING
C6988 a_5394_18116# VGND 0.39633f $ **FLOATING
C6989 a_5844_18123# VGND 0.62179f $ **FLOATING
C6990 a_5196_18116# VGND 0.28271f $ **FLOATING
C6991 a_4771_18260# VGND 0.50939f $ **FLOATING
C6992 single_9b_cdac_1.SW[7] VGND 6.05886f $ **FLOATING
C6993 a_13011_19242# VGND 0.63648f $ **FLOATING
C6994 a_11338_19178# VGND 0.17146f $ **FLOATING
C6995 a_10762_18823# VGND 0.12318f $ **FLOATING
C6996 a_10830_19068# VGND 0.1661f $ **FLOATING
C6997 a_10553_18922# VGND 0.91659f $ **FLOATING
C6998 a_10548_19053# VGND 0.59692f $ **FLOATING
C6999 a_10239_19235# VGND 0.2919f $ **FLOATING
C7000 a_10098_19171# VGND 0.34247f $ **FLOATING
C7001 a_9900_19047# VGND 0.28365f $ **FLOATING
C7002 a_9472_18823# VGND 0.27623f $ **FLOATING
C7003 a_9126_19131# VGND 0.29177f $ **FLOATING
C7004 a_8874_19178# VGND 0.34094f $ **FLOATING
C7005 a_8438_18958# VGND 0.13218f $ **FLOATING
C7006 a_8303_18859# VGND 0.17139f $ **FLOATING
C7007 a_8098_18810# VGND 0.9231f $ **FLOATING
C7008 a_7638_19238# VGND 0.13759f $ **FLOATING
C7009 a_7914_19178# VGND 0.58482f $ **FLOATING
C7010 a_6579_18832# VGND 0.45588f $ **FLOATING
C7011 a_6252_19074# VGND 0.32141f $ **FLOATING
C7012 a_5811_19178# VGND 0.27961f $ **FLOATING
C7013 a_5443_19074# VGND 0.44526f $ **FLOATING
C7014 a_12047_19857# VGND 0.19066f $ **FLOATING
C7015 a_13216_19809# VGND 0.29524f $ **FLOATING
C7016 a_12618_19474# VGND 0.35239f $ **FLOATING
C7017 a_12870_19603# VGND 0.29287f $ **FLOATING
C7018 a_12182_19759# VGND 0.13111f $ **FLOATING
C7019 a_11842_19766# VGND 0.96526f $ **FLOATING
C7020 a_11658_19474# VGND 0.62067f $ **FLOATING
C7021 a_11382_19478# VGND 0.17055f $ **FLOATING
C7022 single_9b_cdac_1.SW[1] VGND 7.77706f $ **FLOATING
C7023 sar9b_0.net48 VGND 3.00596f $ **FLOATING
C7024 a_10803_19474# VGND 0.61976f $ **FLOATING
C7025 a_10035_19474# VGND 0.62781f $ **FLOATING
C7026 a_7882_19538# VGND 0.1244f $ **FLOATING
C7027 a_7374_19685# VGND 0.15921f $ **FLOATING
C7028 a_7306_19777# VGND 0.1167f $ **FLOATING
C7029 a_5761_19487# VGND 0.01222f $ **FLOATING
C7030 a_7097_19795# VGND 0.88857f $ **FLOATING
C7031 a_6783_19481# VGND 0.29276f $ **FLOATING
C7032 a_6642_19448# VGND 0.34651f $ **FLOATING
C7033 a_5628_19768# VGND 0.01308f $ **FLOATING
C7034 a_7092_19455# VGND 0.59664f $ **FLOATING
C7035 a_6444_19448# VGND 0.28777f $ **FLOATING
C7036 a_5581_19664# VGND 0.29099f $ **FLOATING
C7037 a_5196_19448# VGND 0.34938f $ **FLOATING
C7038 a_4072_19474# VGND 0.47181f $ **FLOATING
C7039 a_3795_19512# VGND 0.2312f $ **FLOATING
C7040 sar9b_0.net46 VGND 3.29711f $ **FLOATING
C7041 sar9b_0.net71 VGND 0.32339f $ **FLOATING
C7042 a_3180_19448# VGND 0.35853f $ **FLOATING
C7043 sar9b_0.net50 VGND 1.2487f $ **FLOATING
C7044 a_13011_20574# VGND 0.61397f $ **FLOATING
C7045 sar9b_0.net5 VGND 1.48438f $ **FLOATING
C7046 a_12684_20379# VGND 0.25006f $ **FLOATING
C7047 single_9b_cdac_1.SW[8] VGND 6.02413f $ **FLOATING
C7048 a_11859_20574# VGND 0.71415f $ **FLOATING
C7049 a_10528_20155# VGND 0.29045f $ **FLOATING
C7050 a_10182_20463# VGND 0.30322f $ **FLOATING
C7051 a_9930_20510# VGND 0.34846f $ **FLOATING
C7052 a_9494_20290# VGND 0.13056f $ **FLOATING
C7053 a_9359_20191# VGND 0.16916f $ **FLOATING
C7054 a_9154_20142# VGND 0.92156f $ **FLOATING
C7055 a_8694_20570# VGND 0.13812f $ **FLOATING
C7056 a_8970_20510# VGND 0.66102f $ **FLOATING
C7057 sar9b_0.net15 VGND 0.46616f $ **FLOATING
C7058 a_6130_20239# VGND 0.46131f $ **FLOATING
C7059 a_5931_20140# VGND 0.28737f $ **FLOATING
C7060 a_5481_20185# VGND 0.15828f $ **FLOATING
C7061 a_5633_20244# VGND 0.20547f $ **FLOATING
C7062 a_5374_20145# VGND 0.01758f $ **FLOATING
C7063 a_4496_20468# VGND 0.17016f $ **FLOATING
C7064 sar9b_0._10_ VGND 0.37869f $ **FLOATING
C7065 a_5126_20140# VGND 0.71166f $ **FLOATING
C7066 a_4947_20140# VGND 1.23378f $ **FLOATING
C7067 sar9b_0.net16 VGND 1.53593f $ **FLOATING
C7068 a_3922_20239# VGND 0.41543f $ **FLOATING
C7069 a_3723_20140# VGND 0.24243f $ **FLOATING
C7070 a_3273_20185# VGND 0.15798f $ **FLOATING
C7071 a_3425_20244# VGND 0.18716f $ **FLOATING
C7072 a_3166_20145# VGND 0.02072f $ **FLOATING
C7073 sar9b_0._00_ VGND 0.34642f $ **FLOATING
C7074 a_2918_20140# VGND 0.66229f $ **FLOATING
C7075 a_2739_20140# VGND 1.25389f $ **FLOATING
C7076 a_10607_21189# VGND 0.16031f $ **FLOATING
C7077 a_13011_20806# VGND 0.62155f $ **FLOATING
C7078 a_12435_20806# VGND 0.63677f $ **FLOATING
C7079 sar9b_0.net6 VGND 1.99773f $ **FLOATING
C7080 a_11776_21141# VGND 0.31771f $ **FLOATING
C7081 a_11178_20806# VGND 0.34832f $ **FLOATING
C7082 a_11430_20935# VGND 0.29503f $ **FLOATING
C7083 a_10742_21091# VGND 0.11828f $ **FLOATING
C7084 a_10402_21098# VGND 0.89532f $ **FLOATING
C7085 a_10218_20806# VGND 0.58532f $ **FLOATING
C7086 a_9942_20810# VGND 0.14176f $ **FLOATING
C7087 a_9363_20826# VGND 0.45753f $ **FLOATING
C7088 sar9b_0.net56 VGND 1.44734f $ **FLOATING
C7089 a_8074_20870# VGND 0.14861f $ **FLOATING
C7090 a_7566_21017# VGND 0.17208f $ **FLOATING
C7091 a_7498_21109# VGND 0.13435f $ **FLOATING
C7092 a_5183_20819# VGND 0.01178f $ **FLOATING
C7093 a_7289_21127# VGND 0.92471f $ **FLOATING
C7094 a_6975_20813# VGND 0.30878f $ **FLOATING
C7095 a_6834_20780# VGND 0.37224f $ **FLOATING
C7096 sar9b_0._01_ VGND 0.97665f $ **FLOATING
C7097 a_7284_20787# VGND 0.60133f $ **FLOATING
C7098 a_6636_20780# VGND 0.29286f $ **FLOATING
C7099 sar9b_0._11_ VGND 0.67367f $ **FLOATING
C7100 a_6252_20780# VGND 0.39203f $ **FLOATING
C7101 a_5812_21028# VGND 0.3166f $ **FLOATING
C7102 sar9b_0._08_ VGND 0.57215f $ **FLOATING
C7103 sar9b_0._09_ VGND 0.59924f $ **FLOATING
C7104 a_5581_20992# VGND 0.30562f $ **FLOATING
C7105 a_4922_20857# VGND 0.24594f $ **FLOATING
C7106 a_2508_20780# VGND 2.7729f $ **FLOATING
C7107 a_13011_21906# VGND 0.63044f $ **FLOATING
C7108 a_11859_21906# VGND 0.72107f $ **FLOATING
C7109 sar9b_0.net7 VGND 1.24263f $ **FLOATING
C7110 a_10816_21487# VGND 0.30071f $ **FLOATING
C7111 a_10470_21795# VGND 0.3024f $ **FLOATING
C7112 a_10218_21842# VGND 0.34969f $ **FLOATING
C7113 a_9782_21622# VGND 0.13363f $ **FLOATING
C7114 a_9647_21523# VGND 0.17263f $ **FLOATING
C7115 a_9442_21474# VGND 0.92619f $ **FLOATING
C7116 a_8982_21902# VGND 0.13981f $ **FLOATING
C7117 a_9258_21842# VGND 0.60132f $ **FLOATING
C7118 sar9b_0.net49 VGND 2.18775f $ **FLOATING
C7119 sar9b_0.net8 VGND 3.73402f $ **FLOATING
C7120 a_7443_21496# VGND 0.49853f $ **FLOATING
C7121 sar9b_0.net51 VGND 2.5769f $ **FLOATING
C7122 a_6444_21738# VGND 0.39129f $ **FLOATING
C7123 a_5523_21528# VGND 0.30787f $ **FLOATING
C7124 a_4812_21738# VGND 0.38426f $ **FLOATING
C7125 a_4236_21738# VGND 0.35329f $ **FLOATING
C7126 a_3027_21906# VGND 0.35644f $ **FLOATING
C7127 a_12047_22521# VGND 0.20349f $ **FLOATING
C7128 a_13216_22473# VGND 0.29599f $ **FLOATING
C7129 a_12618_22138# VGND 0.36248f $ **FLOATING
C7130 a_12870_22267# VGND 0.30878f $ **FLOATING
C7131 a_12182_22423# VGND 0.1466f $ **FLOATING
C7132 a_11842_22430# VGND 0.97398f $ **FLOATING
C7133 a_11658_22138# VGND 0.64577f $ **FLOATING
C7134 a_11382_22142# VGND 0.15492f $ **FLOATING
C7135 sar9b_0.net73 VGND 2.09299f $ **FLOATING
C7136 sar9b_0.net61 VGND 3.33314f $ **FLOATING
C7137 a_7978_22202# VGND 0.12351f $ **FLOATING
C7138 a_7470_22349# VGND 0.15862f $ **FLOATING
C7139 a_7402_22441# VGND 0.11773f $ **FLOATING
C7140 a_7193_22459# VGND 0.888f $ **FLOATING
C7141 a_6879_22145# VGND 0.29152f $ **FLOATING
C7142 sar9b_0.net47 VGND 2.48893f $ **FLOATING
C7143 a_6738_22112# VGND 0.33464f $ **FLOATING
C7144 a_5739_22488# VGND 0.25938f $ **FLOATING
C7145 a_5182_22567# VGND 0.01826f $ **FLOATING
C7146 a_7188_22119# VGND 0.58869f $ **FLOATING
C7147 a_6540_22112# VGND 0.2837f $ **FLOATING
C7148 a_5938_22378# VGND 0.43981f $ **FLOATING
C7149 a_5289_22527# VGND 0.1531f $ **FLOATING
C7150 a_5441_22522# VGND 0.18149f $ **FLOATING
C7151 sar9b_0.net64 VGND 1.22538f $ **FLOATING
C7152 a_4934_22432# VGND 0.65617f $ **FLOATING
C7153 a_4755_22138# VGND 1.27206f $ **FLOATING
C7154 sar9b_0.clk_div_0.COUNT\[3\] VGND 0.68828f $ **FLOATING
C7155 a_4011_22488# VGND 0.2324f $ **FLOATING
C7156 a_3454_22567# VGND 0.01679f $ **FLOATING
C7157 a_4210_22378# VGND 0.40953f $ **FLOATING
C7158 a_3561_22527# VGND 0.15284f $ **FLOATING
C7159 a_3713_22522# VGND 0.18104f $ **FLOATING
C7160 sar9b_0.net67 VGND 0.81321f $ **FLOATING
C7161 a_3206_22432# VGND 0.66139f $ **FLOATING
C7162 sar9b_0._05_ VGND 0.79927f $ **FLOATING
C7163 sar9b_0._04_ VGND 0.78117f $ **FLOATING
C7164 a_3027_22138# VGND 1.2701f $ **FLOATING
C7165 sar9b_0.clknet_1_0__leaf_CLK VGND 1.92116f $ **FLOATING
C7166 a_13011_23238# VGND 0.6362f $ **FLOATING
C7167 a_12064_22819# VGND 0.32582f $ **FLOATING
C7168 a_11718_23127# VGND 0.32104f $ **FLOATING
C7169 a_11466_23174# VGND 0.37219f $ **FLOATING
C7170 a_11030_22954# VGND 0.1247f $ **FLOATING
C7171 a_10895_22855# VGND 0.16542f $ **FLOATING
C7172 a_10690_22806# VGND 0.91522f $ **FLOATING
C7173 a_10230_23234# VGND 0.13716f $ **FLOATING
C7174 a_10506_23174# VGND 0.64615f $ **FLOATING
C7175 sar9b_0.net9 VGND 2.28378f $ **FLOATING
C7176 a_9760_22819# VGND 0.28806f $ **FLOATING
C7177 a_9414_23127# VGND 0.2958f $ **FLOATING
C7178 a_9162_23174# VGND 0.35069f $ **FLOATING
C7179 a_8726_22954# VGND 0.12072f $ **FLOATING
C7180 a_8591_22855# VGND 0.15931f $ **FLOATING
C7181 a_8386_22806# VGND 0.90687f $ **FLOATING
C7182 a_7926_23234# VGND 0.13601f $ **FLOATING
C7183 a_8202_23174# VGND 0.60825f $ **FLOATING
C7184 a_7597_23174# VGND 0.01081f $ **FLOATING
C7185 sar9b_0._17_ VGND 0.54536f $ **FLOATING
C7186 a_6744_23238# VGND 0.27119f $ **FLOATING
C7187 sar9b_0._02_ VGND 0.50023f $ **FLOATING
C7188 a_6861_22828# VGND 0.22749f $ **FLOATING
C7189 a_6484_22845# VGND 0.38938f $ **FLOATING
C7190 sar9b_0._12_ VGND 2.03947f $ **FLOATING
C7191 a_4332_23043# VGND 2.49415f $ **FLOATING
C7192 sar9b_0.clk_div_0.COUNT\[0\] VGND 0.5303f $ **FLOATING
C7193 sar9b_0._07_ VGND 3.63856f $ **FLOATING
C7194 sar9b_0.net66 VGND 0.36733f $ **FLOATING
C7195 sar9b_0.net65 VGND 1.04893f $ **FLOATING
C7196 a_3695_23038# VGND 0.27588f $ **FLOATING
C7197 a_3219_22860# VGND 0.23516f $ **FLOATING
C7198 a_3371_23106# VGND 0.25044f $ **FLOATING
C7199 sar9b_0._18_ VGND 0.52436f $ **FLOATING
C7200 a_2892_23070# VGND 0.3304f $ **FLOATING
C7201 a_12047_23853# VGND 0.20399f $ **FLOATING
C7202 a_13216_23805# VGND 0.29598f $ **FLOATING
C7203 a_12618_23470# VGND 0.36236f $ **FLOATING
C7204 a_12870_23599# VGND 0.3087f $ **FLOATING
C7205 a_12182_23755# VGND 0.14911f $ **FLOATING
C7206 a_11842_23762# VGND 0.97787f $ **FLOATING
C7207 a_11658_23470# VGND 0.66469f $ **FLOATING
C7208 a_11382_23474# VGND 0.15995f $ **FLOATING
C7209 a_10707_23470# VGND 0.36843f $ **FLOATING
C7210 sar9b_0.net1 VGND 2.40289f $ **FLOATING
C7211 a_10227_23490# VGND 0.467f $ **FLOATING
C7212 a_8303_23853# VGND 0.16637f $ **FLOATING
C7213 a_9472_23805# VGND 0.29613f $ **FLOATING
C7214 a_8874_23470# VGND 0.35331f $ **FLOATING
C7215 a_9126_23599# VGND 0.29994f $ **FLOATING
C7216 a_8438_23755# VGND 0.13265f $ **FLOATING
C7217 a_8098_23762# VGND 0.9183f $ **FLOATING
C7218 a_7914_23470# VGND 0.6159f $ **FLOATING
C7219 a_7638_23474# VGND 0.11866f $ **FLOATING
C7220 sar9b_0.net10 VGND 1.74489f $ **FLOATING
C7221 a_6922_23534# VGND 0.11783f $ **FLOATING
C7222 a_6414_23681# VGND 0.16683f $ **FLOATING
C7223 a_6346_23773# VGND 0.12324f $ **FLOATING
C7224 a_6137_23791# VGND 0.93229f $ **FLOATING
C7225 a_5823_23477# VGND 0.31555f $ **FLOATING
C7226 a_5682_23444# VGND 0.37293f $ **FLOATING
C7227 a_6132_23451# VGND 0.58878f $ **FLOATING
C7228 a_5484_23444# VGND 0.29255f $ **FLOATING
C7229 a_4811_23656# VGND 0.28975f $ **FLOATING
C7230 sar9b_0.clknet_0_CLK VGND 2.22837f $ **FLOATING
C7231 a_2508_23444# VGND 2.77512f $ **FLOATING
C7232 a_13011_24570# VGND 0.62981f $ **FLOATING
C7233 sar9b_0.net11 VGND 3.57213f $ **FLOATING
C7234 a_11104_24151# VGND 0.30915f $ **FLOATING
C7235 a_10758_24459# VGND 0.303f $ **FLOATING
C7236 a_10506_24506# VGND 0.35537f $ **FLOATING
C7237 a_10070_24286# VGND 0.13107f $ **FLOATING
C7238 a_9935_24187# VGND 0.16193f $ **FLOATING
C7239 a_9730_24138# VGND 0.91556f $ **FLOATING
C7240 a_9270_24566# VGND 0.1136f $ **FLOATING
C7241 a_9546_24506# VGND 0.60387f $ **FLOATING
C7242 sar9b_0.net2 VGND 1.31622f $ **FLOATING
C7243 a_8940_24402# VGND 0.33197f $ **FLOATING
C7244 a_7347_24160# VGND 0.51748f $ **FLOATING
C7245 sar9b_0.net55 VGND 1.13897f $ **FLOATING
C7246 sar9b_0.net62 VGND 1.27467f $ **FLOATING
C7247 a_6538_24506# VGND 0.1602f $ **FLOATING
C7248 a_5962_24151# VGND 0.17011f $ **FLOATING
C7249 a_6030_24396# VGND 0.20052f $ **FLOATING
C7250 a_5753_24250# VGND 0.95497f $ **FLOATING
C7251 a_5748_24381# VGND 0.60642f $ **FLOATING
C7252 a_5439_24563# VGND 0.30942f $ **FLOATING
C7253 a_4467_24162# VGND 0.1655f $ **FLOATING
C7254 sar9b_0._13_ VGND 0.30005f $ **FLOATING
C7255 a_5298_24499# VGND 0.38655f $ **FLOATING
C7256 a_5100_24375# VGND 0.29673f $ **FLOATING
C7257 a_4018_24235# VGND 0.41892f $ **FLOATING
C7258 a_3819_24136# VGND 0.2435f $ **FLOATING
C7259 a_3369_24181# VGND 0.15303f $ **FLOATING
C7260 a_3521_24240# VGND 0.18898f $ **FLOATING
C7261 a_3262_24141# VGND 0.02073f $ **FLOATING
C7262 sar9b_0.net70 VGND 0.58889f $ **FLOATING
C7263 a_3014_24136# VGND 0.63058f $ **FLOATING
C7264 a_2835_24136# VGND 1.26692f $ **FLOATING
C7265 a_10607_25185# VGND 0.16691f $ **FLOATING
C7266 a_13011_24802# VGND 0.62905f $ **FLOATING
C7267 sar9b_0.net26 VGND 2.14803f $ **FLOATING
C7268 a_12435_24802# VGND 0.64526f $ **FLOATING
C7269 a_11776_25137# VGND 0.32738f $ **FLOATING
C7270 a_11178_24802# VGND 0.35816f $ **FLOATING
C7271 a_11430_24931# VGND 0.30602f $ **FLOATING
C7272 a_10742_25087# VGND 0.13219f $ **FLOATING
C7273 a_10402_25094# VGND 0.91973f $ **FLOATING
C7274 a_10218_24802# VGND 0.5916f $ **FLOATING
C7275 sar9b_0.net57 VGND 2.74111f $ **FLOATING
C7276 a_9942_24806# VGND 0.1549f $ **FLOATING
C7277 sar9b_0.net53 VGND 2.57915f $ **FLOATING
C7278 a_6767_25185# VGND 0.17399f $ **FLOATING
C7279 a_9165_24988# VGND 0.47483f $ **FLOATING
C7280 a_7936_25137# VGND 0.3013f $ **FLOATING
C7281 a_7338_24802# VGND 0.35928f $ **FLOATING
C7282 a_7590_24931# VGND 0.30299f $ **FLOATING
C7283 a_6902_25087# VGND 0.1354f $ **FLOATING
C7284 a_6562_25094# VGND 0.92936f $ **FLOATING
C7285 a_6378_24802# VGND 0.661f $ **FLOATING
C7286 sar9b_0.net4 VGND 1.56917f $ **FLOATING
C7287 a_6102_24806# VGND 0.15486f $ **FLOATING
C7288 sar9b_0.net54 VGND 2.72635f $ **FLOATING
C7289 sar9b_0._15_ VGND 0.7538f $ **FLOATING
C7290 a_5580_24776# VGND 0.35113f $ **FLOATING
C7291 sar9b_0.clk_div_0.COUNT\[2\] VGND 0.9962f $ **FLOATING
C7292 a_5196_24776# VGND 0.33541f $ **FLOATING
C7293 a_4044_24776# VGND 0.344f $ **FLOATING
C7294 sar9b_0.net68 VGND 0.89917f $ **FLOATING
C7295 sar9b_0._14_ VGND 0.97587f $ **FLOATING
C7296 a_2893_24992# VGND 0.22912f $ **FLOATING
C7297 sar9b_0.net72 VGND 1.71102f $ **FLOATING
C7298 sar9b_0.net63 VGND 1.46347f $ **FLOATING
C7299 a_13011_25902# VGND 0.63761f $ **FLOATING
C7300 a_11722_25838# VGND 0.17423f $ **FLOATING
C7301 sar9b_0.net13 VGND 1.83091f $ **FLOATING
C7302 a_11146_25483# VGND 0.13526f $ **FLOATING
C7303 a_11214_25728# VGND 0.17226f $ **FLOATING
C7304 a_10937_25582# VGND 0.93944f $ **FLOATING
C7305 a_10932_25713# VGND 0.63975f $ **FLOATING
C7306 a_10623_25895# VGND 0.30445f $ **FLOATING
C7307 a_10482_25831# VGND 0.35993f $ **FLOATING
C7308 a_10284_25707# VGND 0.30192f $ **FLOATING
C7309 sar9b_0.clknet_1_1__leaf_CLK VGND 1.99526f $ **FLOATING
C7310 a_4698_25851# VGND 0.02231f $ **FLOATING
C7311 sar9b_0._03_ VGND 0.34487f $ **FLOATING
C7312 a_4293_25852# VGND 0.18854f $ **FLOATING
C7313 a_4365_25770# VGND 0.16167f $ **FLOATING
C7314 a_4136_25584# VGND 0.6886f $ **FLOATING
C7315 sar9b_0.clk_div_0.COUNT\[1\] VGND 1.70819f $ **FLOATING
C7316 sar9b_0.net69 VGND 1.15997f $ **FLOATING
C7317 a_4125_25958# VGND 1.27131f $ **FLOATING
C7318 a_3855_25792# VGND 0.24272f $ **FLOATING
C7319 a_3747_25724# VGND 0.41638f $ **FLOATING
C7320 sar9b_0._16_ VGND 0.40855f $ **FLOATING
C7321 a_3372_25734# VGND 0.33769f $ **FLOATING
C7322 a_12047_26517# VGND 0.19151f $ **FLOATING
C7323 a_13216_26469# VGND 0.28884f $ **FLOATING
C7324 a_12618_26134# VGND 0.35065f $ **FLOATING
C7325 a_12870_26263# VGND 0.29813f $ **FLOATING
C7326 a_12182_26419# VGND 0.13385f $ **FLOATING
C7327 a_11842_26426# VGND 0.96869f $ **FLOATING
C7328 a_11658_26134# VGND 0.62093f $ **FLOATING
C7329 sar9b_0.net12 VGND 1.66742f $ **FLOATING
C7330 a_11382_26138# VGND 0.14597f $ **FLOATING
C7331 sar9b_0.net74 VGND 1.58493f $ **FLOATING
C7332 sar9b_0.net33 VGND 1.05333f $ **FLOATING
C7333 a_10859_26330# VGND 0.61787f $ **FLOATING
C7334 sar9b_0.net41 VGND 2.17416f $ **FLOATING
C7335 a_9130_26198# VGND 0.15692f $ **FLOATING
C7336 a_8622_26345# VGND 0.17118f $ **FLOATING
C7337 a_8554_26437# VGND 0.13269f $ **FLOATING
C7338 a_8345_26455# VGND 0.92555f $ **FLOATING
C7339 a_8031_26141# VGND 0.30485f $ **FLOATING
C7340 a_7890_26108# VGND 0.35529f $ **FLOATING
C7341 a_8340_26115# VGND 0.61091f $ **FLOATING
C7342 a_7692_26108# VGND 0.30296f $ **FLOATING
C7343 sar9b_0.net35 VGND 2.44446f $ **FLOATING
C7344 a_3946_26198# VGND 0.15782f $ **FLOATING
C7345 a_3438_26345# VGND 0.17121f $ **FLOATING
C7346 a_3370_26437# VGND 0.13251f $ **FLOATING
C7347 a_3161_26455# VGND 0.9217f $ **FLOATING
C7348 a_2847_26141# VGND 0.3046f $ **FLOATING
C7349 a_2706_26108# VGND 0.36022f $ **FLOATING
C7350 a_3156_26115# VGND 0.59376f $ **FLOATING
C7351 a_2508_26108# VGND 0.30075f $ **FLOATING
C7352 a_63626_26990# VGND 0.89497f $ **FLOATING
C7353 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLK0 VGND 2.68117f $ **FLOATING
C7354 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.CLKB0 VGND 3.19275f $ **FLOATING
C7355 a_62748_26999# VGND 0.16243f $ **FLOATING
C7356 single_9b_cdac_0.SW[0] VGND 11.0253f $ **FLOATING
C7357 a_58824_26990# VGND 0.89548f $ **FLOATING
C7358 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLK0 VGND 2.66663f $ **FLOATING
C7359 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWN VGND 6.36459f $ **FLOATING
C7360 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.39423f $ **FLOATING
C7361 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7362 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.45426f $ **FLOATING
C7363 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7364 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x8.A VGND 1.57322f $ **FLOATING
C7365 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x1.A VGND 1.60512f $ **FLOATING
C7366 single_9b_cdac_0.cdac_sw_9b_0.S[0] VGND 94.5927f $ **FLOATING
C7367 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.CLKB0 VGND 3.16256f $ **FLOATING
C7368 a_57946_26999# VGND 0.16243f $ **FLOATING
C7369 a_54032_26990# VGND 0.89543f $ **FLOATING
C7370 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VGND 2.66664f $ **FLOATING
C7371 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWN VGND 6.34807f $ **FLOATING
C7372 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7373 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7374 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7375 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7376 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.tg_sw_3_3.SWP VGND 4.52773f $ **FLOATING
C7377 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7378 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7379 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.41378f $ **FLOATING
C7380 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7381 single_9b_cdac_0.cdac_sw_9b_0.S[1] VGND 47.9165f $ **FLOATING
C7382 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VGND 3.16255f $ **FLOATING
C7383 a_53154_26999# VGND 0.16243f $ **FLOATING
C7384 a_49221_26990# VGND 0.89502f $ **FLOATING
C7385 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLK0 VGND 2.66535f $ **FLOATING
C7386 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWN VGND 6.34853f $ **FLOATING
C7387 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37221f $ **FLOATING
C7388 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7389 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44881f $ **FLOATING
C7390 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7391 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.tg_sw_3_3.SWP VGND 4.51045f $ **FLOATING
C7392 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VGND 1.56057f $ **FLOATING
C7393 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7394 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7395 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VGND 1.58431f $ **FLOATING
C7396 single_9b_cdac_0.cdac_sw_9b_0.S[2] VGND 30.3253f $ **FLOATING
C7397 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.CLKB0 VGND 3.16311f $ **FLOATING
C7398 a_48343_26999# VGND 0.16243f $ **FLOATING
C7399 a_44418_26990# VGND 0.89497f $ **FLOATING
C7400 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLK0 VGND 2.665f $ **FLOATING
C7401 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWN VGND 6.34862f $ **FLOATING
C7402 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37348f $ **FLOATING
C7403 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7404 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44912f $ **FLOATING
C7405 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7406 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.tg_sw_3_3.SWP VGND 4.51335f $ **FLOATING
C7407 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x8.A VGND 1.56099f $ **FLOATING
C7408 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7409 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.405f $ **FLOATING
C7410 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x1.A VGND 1.58193f $ **FLOATING
C7411 single_9b_cdac_0.cdac_sw_9b_0.S[3] VGND 21.4947f $ **FLOATING
C7412 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.CLKB0 VGND 3.16279f $ **FLOATING
C7413 a_43540_26999# VGND 0.16243f $ **FLOATING
C7414 a_39616_26990# VGND 0.89497f $ **FLOATING
C7415 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLK0 VGND 2.66616f $ **FLOATING
C7416 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWN VGND 6.34842f $ **FLOATING
C7417 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.37296f $ **FLOATING
C7418 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7419 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44899f $ **FLOATING
C7420 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7421 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.tg_sw_3_3.SWP VGND 4.51193f $ **FLOATING
C7422 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x8.A VGND 1.56081f $ **FLOATING
C7423 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7424 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40542f $ **FLOATING
C7425 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x1.A VGND 1.58513f $ **FLOATING
C7426 single_9b_cdac_0.cdac_sw_9b_0.S[4] VGND 20.61f $ **FLOATING
C7427 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7428 a_38738_26999# VGND 0.16243f $ **FLOATING
C7429 a_34814_26990# VGND 0.89548f $ **FLOATING
C7430 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLK0 VGND 2.66683f $ **FLOATING
C7431 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWN VGND 6.34843f $ **FLOATING
C7432 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7433 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7434 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7435 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7436 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.tg_sw_3_3.SWP VGND 4.51156f $ **FLOATING
C7437 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7438 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7439 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40525f $ **FLOATING
C7440 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7441 single_9b_cdac_0.cdac_sw_9b_0.S[5] VGND 16.1449f $ **FLOATING
C7442 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7443 a_33936_26999# VGND 0.16243f $ **FLOATING
C7444 a_30012_26990# VGND 0.89497f $ **FLOATING
C7445 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLK0 VGND 2.66498f $ **FLOATING
C7446 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWN VGND 6.34843f $ **FLOATING
C7447 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7448 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7449 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7450 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7451 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.tg_sw_3_3.SWP VGND 4.51162f $ **FLOATING
C7452 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7453 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7454 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7455 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7456 single_9b_cdac_0.cdac_sw_9b_0.S[6] VGND 15.6371f $ **FLOATING
C7457 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.CLKB0 VGND 3.16276f $ **FLOATING
C7458 a_29134_26999# VGND 0.16243f $ **FLOATING
C7459 single_9b_cdac_0.SW[7] VGND 7.22415f $ **FLOATING
C7460 a_25210_26990# VGND 0.89548f $ **FLOATING
C7461 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLK0 VGND 2.68106f $ **FLOATING
C7462 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWN VGND 6.3484f $ **FLOATING
C7463 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7464 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7465 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7466 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7467 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.tg_sw_3_3.SWP VGND 4.51212f $ **FLOATING
C7468 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7469 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7470 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7471 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7472 single_9b_cdac_0.cdac_sw_9b_0.S[7] VGND 14.5496f $ **FLOATING
C7473 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.CLKB0 VGND 3.17698f $ **FLOATING
C7474 a_24332_26999# VGND 0.16243f $ **FLOATING
C7475 single_9b_cdac_0.SW[1] VGND 7.88723f $ **FLOATING
C7476 a_12647_27128# VGND 0.01049f $ **FLOATING
C7477 a_12560_27128# VGND 0.18115f $ **FLOATING
C7478 a_13011_27234# VGND 0.59986f $ **FLOATING
C7479 sar9b_0.net27 VGND 1.75655f $ **FLOATING
C7480 single_9b_cdac_0.SW[4] VGND 7.53235f $ **FLOATING
C7481 single_9b_cdac_0.SW[5] VGND 7.99262f $ **FLOATING
C7482 sar9b_0.net52 VGND 3.396f $ **FLOATING
C7483 sar9b_0.net30 VGND 0.98276f $ **FLOATING
C7484 a_11915_27039# VGND 0.68615f $ **FLOATING
C7485 sar9b_0.net31 VGND 0.75736f $ **FLOATING
C7486 a_11339_27039# VGND 0.62214f $ **FLOATING
C7487 sar9b_0.net42 VGND 1.35212f $ **FLOATING
C7488 a_10378_27170# VGND 0.13252f $ **FLOATING
C7489 a_9802_26815# VGND 0.11561f $ **FLOATING
C7490 a_9870_27060# VGND 0.16016f $ **FLOATING
C7491 a_9593_26914# VGND 0.89305f $ **FLOATING
C7492 a_9588_27045# VGND 0.60592f $ **FLOATING
C7493 a_9279_27227# VGND 0.28615f $ **FLOATING
C7494 a_9138_27163# VGND 0.33078f $ **FLOATING
C7495 a_8940_27039# VGND 0.28409f $ **FLOATING
C7496 a_6880_26815# VGND 0.30246f $ **FLOATING
C7497 a_6534_27123# VGND 0.29776f $ **FLOATING
C7498 a_6282_27170# VGND 0.35829f $ **FLOATING
C7499 a_5846_26950# VGND 0.15475f $ **FLOATING
C7500 a_5711_26851# VGND 0.20102f $ **FLOATING
C7501 a_5506_26802# VGND 0.94424f $ **FLOATING
C7502 a_5046_27230# VGND 0.11169f $ **FLOATING
C7503 a_5322_27170# VGND 0.61739f $ **FLOATING
C7504 sar9b_0.net39 VGND 5.04702f $ **FLOATING
C7505 sar9b_0.net37 VGND 3.30771f $ **FLOATING
C7506 a_4330_27170# VGND 0.1075f $ **FLOATING
C7507 a_3754_26815# VGND 0.11452f $ **FLOATING
C7508 a_3822_27060# VGND 0.15534f $ **FLOATING
C7509 a_3545_26914# VGND 0.88258f $ **FLOATING
C7510 a_3540_27045# VGND 0.57229f $ **FLOATING
C7511 a_3231_27227# VGND 0.28633f $ **FLOATING
C7512 a_3090_27163# VGND 0.3281f $ **FLOATING
C7513 a_2892_27039# VGND 0.27715f $ **FLOATING
C7514 a_2451_27234# VGND 0.36326f $ **FLOATING
C7515 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWN VGND 6.37207f $ **FLOATING
C7516 single_9b_cdac_0.SW[2] VGND 7.79108f $ **FLOATING
C7517 single_9b_cdac_0.SW[3] VGND 7.69147f $ **FLOATING
C7518 a_10607_27849# VGND 0.17037f $ **FLOATING
C7519 sar9b_0.net28 VGND 2.13028f $ **FLOATING
C7520 a_13067_27662# VGND 0.62659f $ **FLOATING
C7521 sar9b_0.net29 VGND 1.17448f $ **FLOATING
C7522 a_12491_27662# VGND 0.63745f $ **FLOATING
C7523 a_11776_27801# VGND 0.33209f $ **FLOATING
C7524 a_11178_27466# VGND 0.37061f $ **FLOATING
C7525 a_11430_27595# VGND 0.30882f $ **FLOATING
C7526 a_10742_27751# VGND 0.13782f $ **FLOATING
C7527 a_10402_27758# VGND 0.92755f $ **FLOATING
C7528 a_10218_27466# VGND 0.65521f $ **FLOATING
C7529 a_9942_27470# VGND 0.15547f $ **FLOATING
C7530 sar9b_0.net43 VGND 2.18762f $ **FLOATING
C7531 single_9b_cdac_0.SW[8] VGND 9.42114f $ **FLOATING
C7532 a_7343_27849# VGND 0.16308f $ **FLOATING
C7533 sar9b_0.net34 VGND 0.84365f $ **FLOATING
C7534 a_9323_27662# VGND 0.63074f $ **FLOATING
C7535 a_8883_27466# VGND 0.45025f $ **FLOATING
C7536 sar9b_0.cyclic_flag_0.FINAL VGND 1.13968f $ **FLOATING
C7537 a_8512_27801# VGND 0.28448f $ **FLOATING
C7538 a_7914_27466# VGND 0.34106f $ **FLOATING
C7539 a_8166_27595# VGND 0.29361f $ **FLOATING
C7540 a_7478_27751# VGND 0.12296f $ **FLOATING
C7541 a_7138_27758# VGND 0.91809f $ **FLOATING
C7542 a_6954_27466# VGND 0.61234f $ **FLOATING
C7543 a_6678_27470# VGND 0.11676f $ **FLOATING
C7544 sar9b_0.net40 VGND 4.42282f $ **FLOATING
C7545 a_6307_27584# VGND 0.41924f $ **FLOATING
C7546 a_5235_27466# VGND 0.61697f $ **FLOATING
C7547 sar9b_0.net19 VGND 1.72645f $ **FLOATING
C7548 a_4749_27652# VGND 0.44592f $ **FLOATING
C7549 sar9b_0.net36 VGND 3.44267f $ **FLOATING
C7550 sar9b_0.net44 VGND 1.32306f $ **FLOATING
C7551 a_3946_27530# VGND 0.1577f $ **FLOATING
C7552 a_3438_27677# VGND 0.1683f $ **FLOATING
C7553 a_3370_27769# VGND 0.13183f $ **FLOATING
C7554 a_3161_27787# VGND 0.91973f $ **FLOATING
C7555 a_2847_27473# VGND 0.30295f $ **FLOATING
C7556 a_2706_27440# VGND 0.35511f $ **FLOATING
C7557 a_3156_27447# VGND 0.60874f $ **FLOATING
C7558 a_2508_27440# VGND 0.29951f $ **FLOATING
C7559 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VGND 1.3729f $ **FLOATING
C7560 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x10.A VGND 1.39185f $ **FLOATING
C7561 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VGND 0.44898f $ **FLOATING
C7562 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x6.A VGND 0.47224f $ **FLOATING
C7563 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.tg_sw_3_3.SWP VGND 4.51154f $ **FLOATING
C7564 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x8.A VGND 1.56079f $ **FLOATING
C7565 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7566 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7567 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x1.A VGND 1.58505f $ **FLOATING
C7568 single_9b_cdac_0.cdac_sw_9b_0.S[8] VGND 13.6188f $ **FLOATING
C7569 sar9b_0._06_ VGND 0.51759f $ **FLOATING
C7570 a_13164_28398# VGND 0.35538f $ **FLOATING
C7571 a_12531_28566# VGND 0.66182f $ **FLOATING
C7572 sar9b_0.net25 VGND 0.48263f $ **FLOATING
C7573 sar9b_0.net14 VGND 0.57635f $ **FLOATING
C7574 a_11915_28371# VGND 0.69798f $ **FLOATING
C7575 a_10995_28566# VGND 0.63419f $ **FLOATING
C7576 sar9b_0.net24 VGND 1.19162f $ **FLOATING
C7577 a_9939_28566# VGND 0.66415f $ **FLOATING
C7578 sar9b_0.net23 VGND 0.45975f $ **FLOATING
C7579 single_9b_cdac_0.SW[6] VGND 7.61708f $ **FLOATING
C7580 sar9b_0.net32 VGND 2.57466f $ **FLOATING
C7581 a_9323_28371# VGND 0.65565f $ **FLOATING
C7582 a_8691_28566# VGND 0.6426f $ **FLOATING
C7583 sar9b_0.net22 VGND 0.37611f $ **FLOATING
C7584 a_8115_28566# VGND 0.63526f $ **FLOATING
C7585 a_7539_28566# VGND 0.63297f $ **FLOATING
C7586 sar9b_0.net21 VGND 0.59997f $ **FLOATING
C7587 sar9b_0.net38 VGND 1.58614f $ **FLOATING
C7588 a_6250_28502# VGND 0.14552f $ **FLOATING
C7589 sar9b_0.net45 VGND 1.28036f $ **FLOATING
C7590 a_5674_28147# VGND 0.15778f $ **FLOATING
C7591 a_5742_28392# VGND 0.21088f $ **FLOATING
C7592 a_5465_28246# VGND 0.95941f $ **FLOATING
C7593 a_5460_28377# VGND 0.66988f $ **FLOATING
C7594 a_5151_28559# VGND 0.30729f $ **FLOATING
C7595 sar9b_0.net58 VGND 3.01825f $ **FLOATING
C7596 sar9b_0.net20 VGND 1.32881f $ **FLOATING
C7597 a_5010_28495# VGND 0.36594f $ **FLOATING
C7598 a_4812_28371# VGND 0.29879f $ **FLOATING
C7599 sar9b_0.net59 VGND 2.86651f $ **FLOATING
C7600 a_4083_28566# VGND 0.64865f $ **FLOATING
C7601 sar9b_0.net18 VGND 0.41648f $ **FLOATING
C7602 a_3603_28156# VGND 0.47335f $ **FLOATING
C7603 sar9b_0.net60 VGND 3.34485f $ **FLOATING
C7604 a_2931_28566# VGND 0.64119f $ **FLOATING
C7605 sar9b_0.net17 VGND 0.6804f $ **FLOATING
C7606 a_2547_28132# VGND 0.43769f $ **FLOATING
C7607 sar9b_0.net3 VGND 0.60828f $ **FLOATING
C7608 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.tg_sw_3_3.SWP VGND 4.71478f $ **FLOATING
C7609 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x4.A VGND 0.42464f $ **FLOATING
C7610 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VGND 0.40523f $ **FLOATING
C7611 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_2.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7612 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_1.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7613 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7614 single_9b_cdac_1.CF[0] VGND 15.8339f $ **FLOATING
C7615 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_4.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7616 single_9b_cdac_1.CF[1] VGND 11.5306f $ **FLOATING
C7617 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_3.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7618 single_9b_cdac_1.CF[2] VGND 11.2901f $ **FLOATING
C7619 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_5.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7620 single_9b_cdac_1.CF[3] VGND 10.9802f $ **FLOATING
C7621 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_6.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7622 single_9b_cdac_1.CF[4] VGND 10.9973f $ **FLOATING
C7623 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_7.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7624 single_9b_cdac_1.CF[5] VGND 10.4191f $ **FLOATING
C7625 single_9b_cdac_0.cdac_sw_9b_0.cdac_sw_3_8.nooverlap_clk_0.x3.Y VGND 0.35827f $ **FLOATING
C7626 single_9b_cdac_1.CF[6] VGND 10.1217f $ **FLOATING
C7627 single_9b_cdac_1.CF[7] VGND 10.1149f $ **FLOATING
C7628 single_9b_cdac_1.CF[8] VGND 8.83586f $ **FLOATING
C7629 dw_17224_1400# VGND 27.9938f $ **FLOATING
C7630 dw_12589_1395# VGND 28.2006f $ **FLOATING
.ends
