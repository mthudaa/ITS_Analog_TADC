magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< pwell >>
rect -184 -95 184 157
<< nmos >>
rect -100 -69 100 131
<< ndiff >>
rect -158 116 -100 131
rect -158 82 -146 116
rect -112 82 -100 116
rect -158 48 -100 82
rect -158 14 -146 48
rect -112 14 -100 48
rect -158 -20 -100 14
rect -158 -54 -146 -20
rect -112 -54 -100 -20
rect -158 -69 -100 -54
rect 100 116 158 131
rect 100 82 112 116
rect 146 82 158 116
rect 100 48 158 82
rect 100 14 112 48
rect 146 14 158 48
rect 100 -20 158 14
rect 100 -54 112 -20
rect 146 -54 158 -20
rect 100 -69 158 -54
<< ndiffc >>
rect -146 82 -112 116
rect -146 14 -112 48
rect -146 -54 -112 -20
rect 112 82 146 116
rect 112 14 146 48
rect 112 -54 146 -20
<< poly >>
rect -100 131 100 157
rect -100 -107 100 -69
rect -100 -124 -17 -107
rect -58 -141 -17 -124
rect 17 -124 100 -107
rect 17 -141 58 -124
rect -58 -157 58 -141
<< polycont >>
rect -17 -141 17 -107
<< locali >>
rect -146 116 -112 135
rect -146 48 -112 50
rect -146 12 -112 14
rect -146 -73 -112 -54
rect 112 116 146 135
rect 112 48 146 50
rect 112 12 146 14
rect 112 -73 146 -54
rect -58 -141 -17 -107
rect 17 -141 58 -107
<< viali >>
rect -146 82 -112 84
rect -146 50 -112 82
rect -146 -20 -112 12
rect -146 -22 -112 -20
rect 112 82 146 84
rect 112 50 146 82
rect 112 -20 146 12
rect 112 -22 146 -20
rect -17 -141 17 -107
<< metal1 >>
rect -152 84 -106 131
rect -152 50 -146 84
rect -112 50 -106 84
rect -152 12 -106 50
rect -152 -22 -146 12
rect -112 -22 -106 12
rect -152 -69 -106 -22
rect 106 84 152 131
rect 106 50 112 84
rect 146 50 152 84
rect 106 12 152 50
rect 106 -22 112 12
rect 146 -22 152 12
rect 106 -69 152 -22
rect -54 -107 54 -101
rect -54 -141 -17 -107
rect 17 -141 54 -107
rect -54 -147 54 -141
<< end >>
