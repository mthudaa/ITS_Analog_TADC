magic
tech sky130A
magscale 1 2
timestamp 1757911661
<< viali >>
rect 12223 14450 12257 14484
rect 2143 14376 2177 14410
rect 3295 14376 3329 14410
rect 3967 14376 4001 14410
rect 6751 14376 6785 14410
rect 7327 14376 7361 14410
rect 7903 14376 7937 14410
rect 8767 14376 8801 14410
rect 9151 14376 9185 14410
rect 10207 14376 10241 14410
rect 11359 14376 11393 14410
rect 11743 14376 11777 14410
rect 2719 14302 2753 14336
rect 2911 14302 2945 14336
rect 5599 14302 5633 14336
rect 12415 14302 12449 14336
rect 1759 14228 1793 14262
rect 1855 14228 1889 14262
rect 3391 14228 3425 14262
rect 5983 14228 6017 14262
rect 7423 14228 7457 14262
rect 7999 14228 8033 14262
rect 11263 14228 11297 14262
rect 2239 14154 2273 14188
rect 6847 14154 6881 14188
rect 8479 14154 8513 14188
rect 9247 14154 9281 14188
rect 10303 14154 10337 14188
rect 11839 14154 11873 14188
rect 1759 13858 1793 13892
rect 4543 13858 4577 13892
rect 7807 13858 7841 13892
rect 8479 13858 8513 13892
rect 11071 13858 11105 13892
rect 4063 13710 4097 13744
rect 8191 13710 8225 13744
rect 3295 13636 3329 13670
rect 4255 13636 4289 13670
rect 5519 13636 5553 13670
rect 6175 13636 6209 13670
rect 9439 13636 9473 13670
rect 3679 13562 3713 13596
rect 4447 13562 4481 13596
rect 5599 13562 5633 13596
rect 5791 13562 5825 13596
rect 8095 13562 8129 13596
rect 8767 13562 8801 13596
rect 9055 13562 9089 13596
rect 11935 13562 11969 13596
rect 12511 13562 12545 13596
rect 11647 13414 11681 13448
rect 12223 13414 12257 13448
rect 1855 13192 1889 13226
rect 2047 13192 2081 13226
rect 6175 13192 6209 13226
rect 8095 13192 8129 13226
rect 10495 13192 10529 13226
rect 11647 13192 11681 13226
rect 12031 13192 12065 13226
rect 11071 13118 11105 13152
rect 4063 13044 4097 13078
rect 10783 13044 10817 13078
rect 11359 13044 11393 13078
rect 11839 13044 11873 13078
rect 12223 13044 12257 13078
rect 1567 12970 1601 13004
rect 3679 12970 3713 13004
rect 4543 12970 4577 13004
rect 9727 12970 9761 13004
rect 10111 12970 10145 13004
rect 4159 12896 4193 12930
rect 12511 12748 12545 12782
rect 1759 12526 1793 12560
rect 6943 12526 6977 12560
rect 10207 12526 10241 12560
rect 3295 12304 3329 12338
rect 8479 12304 8513 12338
rect 10879 12304 10913 12338
rect 3679 12230 3713 12264
rect 8863 12230 8897 12264
rect 10303 12230 10337 12264
rect 10495 12230 10529 12264
rect 12511 12156 12545 12190
rect 9439 11860 9473 11894
rect 11455 11712 11489 11746
rect 12223 11712 12257 11746
rect 2623 11638 2657 11672
rect 4351 11638 4385 11672
rect 11071 11638 11105 11672
rect 2431 11564 2465 11598
rect 3967 11564 4001 11598
rect 12511 11564 12545 11598
rect 2815 11416 2849 11450
rect 1951 11194 1985 11228
rect 4639 11194 4673 11228
rect 7231 11194 7265 11228
rect 12511 11194 12545 11228
rect 10975 11120 11009 11154
rect 2335 10972 2369 11006
rect 3295 10972 3329 11006
rect 4447 10972 4481 11006
rect 4831 10972 4865 11006
rect 5599 10972 5633 11006
rect 8671 10972 8705 11006
rect 9439 10972 9473 11006
rect 1663 10898 1697 10932
rect 1855 10898 1889 10932
rect 2623 10898 2657 10932
rect 4255 10898 4289 10932
rect 5215 10898 5249 10932
rect 8479 10898 8513 10932
rect 9055 10898 9089 10932
rect 11647 10898 11681 10932
rect 12223 10898 12257 10932
rect 1855 10824 1889 10858
rect 3103 10750 3137 10784
rect 11935 10750 11969 10784
rect 3775 10528 3809 10562
rect 12223 10380 12257 10414
rect 1951 10306 1985 10340
rect 3775 10306 3809 10340
rect 3871 10306 3905 10340
rect 5887 10306 5921 10340
rect 6463 10306 6497 10340
rect 8287 10306 8321 10340
rect 8767 10306 8801 10340
rect 2335 10232 2369 10266
rect 4063 10232 4097 10266
rect 6271 10232 6305 10266
rect 6655 10232 6689 10266
rect 8383 10232 8417 10266
rect 3487 10084 3521 10118
rect 4255 10084 4289 10118
rect 7999 10084 8033 10118
rect 10399 10084 10433 10118
rect 12511 10084 12545 10118
rect 3871 9862 3905 9896
rect 8767 9862 8801 9896
rect 12415 9862 12449 9896
rect 9535 9714 9569 9748
rect 3391 9640 3425 9674
rect 4063 9640 4097 9674
rect 6271 9640 6305 9674
rect 7135 9640 7169 9674
rect 9343 9640 9377 9674
rect 9823 9640 9857 9674
rect 10879 9640 10913 9674
rect 4255 9566 4289 9600
rect 6655 9566 6689 9600
rect 6751 9566 6785 9600
rect 10495 9566 10529 9600
rect 4639 9492 4673 9526
rect 10111 9418 10145 9452
rect 2527 9196 2561 9230
rect 11359 9196 11393 9230
rect 12511 9196 12545 9230
rect 5599 9048 5633 9082
rect 6271 9048 6305 9082
rect 6559 9048 6593 9082
rect 6655 9048 6689 9082
rect 6751 9048 6785 9082
rect 9343 9048 9377 9082
rect 12223 9048 12257 9082
rect 2239 8974 2273 9008
rect 2335 8974 2369 9008
rect 2911 8974 2945 9008
rect 3007 8974 3041 9008
rect 3199 8974 3233 9008
rect 5215 8974 5249 9008
rect 5311 8974 5345 9008
rect 5503 8974 5537 9008
rect 7423 8974 7457 9008
rect 9727 8974 9761 9008
rect 7039 8900 7073 8934
rect 6463 8826 6497 8860
rect 1951 8752 1985 8786
rect 5407 8752 5441 8786
rect 9055 8752 9089 8786
rect 5407 8530 5441 8564
rect 12415 8530 12449 8564
rect 1567 8308 1601 8342
rect 1759 8308 1793 8342
rect 1855 8308 1889 8342
rect 2047 8308 2081 8342
rect 2143 8308 2177 8342
rect 3871 8308 3905 8342
rect 7327 8308 7361 8342
rect 10879 8308 10913 8342
rect 2527 8234 2561 8268
rect 4255 8234 4289 8268
rect 7711 8234 7745 8268
rect 10495 8234 10529 8268
rect 1663 8086 1697 8120
rect 1951 8086 1985 8120
rect 3679 8086 3713 8120
rect 5695 8086 5729 8120
rect 2431 7864 2465 7898
rect 3295 7864 3329 7898
rect 5503 7864 5537 7898
rect 12511 7864 12545 7898
rect 5023 7790 5057 7824
rect 10111 7790 10145 7824
rect 6751 7716 6785 7750
rect 11071 7716 11105 7750
rect 12223 7716 12257 7750
rect 2143 7642 2177 7676
rect 3487 7642 3521 7676
rect 4063 7642 4097 7676
rect 4639 7642 4673 7676
rect 4831 7642 4865 7676
rect 5791 7642 5825 7676
rect 6559 7642 6593 7676
rect 8479 7642 8513 7676
rect 3871 7568 3905 7602
rect 8095 7568 8129 7602
rect 11359 7568 11393 7602
rect 4543 7124 4577 7158
rect 5887 7124 5921 7158
rect 7807 7050 7841 7084
rect 8671 7050 8705 7084
rect 12511 7050 12545 7084
rect 3391 6976 3425 7010
rect 4351 6976 4385 7010
rect 4831 6976 4865 7010
rect 5503 6976 5537 7010
rect 7423 6976 7457 7010
rect 8479 6976 8513 7010
rect 9439 6976 9473 7010
rect 3871 6902 3905 6936
rect 5215 6902 5249 6936
rect 9055 6902 9089 6936
rect 11647 6902 11681 6936
rect 12223 6902 12257 6936
rect 11935 6828 11969 6862
rect 4639 6754 4673 6788
rect 5311 6754 5345 6788
rect 11071 6754 11105 6788
rect 3679 6532 3713 6566
rect 3967 6532 4001 6566
rect 9823 6532 9857 6566
rect 3775 6384 3809 6418
rect 4447 6384 4481 6418
rect 7807 6384 7841 6418
rect 11071 6384 11105 6418
rect 12223 6384 12257 6418
rect 1855 6310 1889 6344
rect 4063 6310 4097 6344
rect 8191 6310 8225 6344
rect 11935 6310 11969 6344
rect 2239 6236 2273 6270
rect 12511 6236 12545 6270
rect 11743 6162 11777 6196
rect 3391 6088 3425 6122
rect 5599 6088 5633 6122
rect 11359 6088 11393 6122
rect 2239 5866 2273 5900
rect 4639 5866 4673 5900
rect 10495 5718 10529 5752
rect 12511 5718 12545 5752
rect 2527 5644 2561 5678
rect 3007 5644 3041 5678
rect 4447 5644 4481 5678
rect 4831 5644 4865 5678
rect 7231 5644 7265 5678
rect 7615 5644 7649 5678
rect 10879 5644 10913 5678
rect 3295 5570 3329 5604
rect 4255 5570 4289 5604
rect 5311 5570 5345 5604
rect 9247 5570 9281 5604
rect 10015 5570 10049 5604
rect 3391 5496 3425 5530
rect 3679 5496 3713 5530
rect 5599 5422 5633 5456
rect 9535 5422 9569 5456
rect 10303 5422 10337 5456
rect 5311 5200 5345 5234
rect 9055 5200 9089 5234
rect 12511 5200 12545 5234
rect 5215 5126 5249 5160
rect 8767 5126 8801 5160
rect 4735 5052 4769 5086
rect 5887 5052 5921 5086
rect 12223 5052 12257 5086
rect 5023 4978 5057 5012
rect 5599 4978 5633 5012
rect 5695 4978 5729 5012
rect 7135 4978 7169 5012
rect 10687 4978 10721 5012
rect 4639 4904 4673 4938
rect 6751 4904 6785 4938
rect 11071 4904 11105 4938
rect 10495 4386 10529 4420
rect 5983 4312 6017 4346
rect 8191 4312 8225 4346
rect 10879 4312 10913 4346
rect 4063 4238 4097 4272
rect 6367 4238 6401 4272
rect 8575 4238 8609 4272
rect 9439 4238 9473 4272
rect 10015 4238 10049 4272
rect 12511 4238 12545 4272
rect 3967 4090 4001 4124
rect 4351 4090 4385 4124
rect 6559 4090 6593 4124
rect 9727 4090 9761 4124
rect 10303 4090 10337 4124
rect 6463 3868 6497 3902
rect 10303 3868 10337 3902
rect 12511 3868 12545 3902
rect 6175 3794 6209 3828
rect 10495 3794 10529 3828
rect 4159 3720 4193 3754
rect 7231 3720 7265 3754
rect 7807 3720 7841 3754
rect 11071 3720 11105 3754
rect 12223 3720 12257 3754
rect 4543 3646 4577 3680
rect 6751 3646 6785 3680
rect 8671 3646 8705 3680
rect 10687 3646 10721 3680
rect 8287 3572 8321 3606
rect 11359 3572 11393 3606
rect 7519 3424 7553 3458
rect 8095 3424 8129 3458
rect 4735 3202 4769 3236
rect 6271 3202 6305 3236
rect 6559 3202 6593 3236
rect 9247 3202 9281 3236
rect 12511 3202 12545 3236
rect 11167 3054 11201 3088
rect 11647 3054 11681 3088
rect 4447 2980 4481 3014
rect 6079 2980 6113 3014
rect 8191 2980 8225 3014
rect 10783 2980 10817 3014
rect 11839 2980 11873 3014
rect 2047 2906 2081 2940
rect 8575 2906 8609 2940
rect 12223 2906 12257 2940
rect 1759 2758 1793 2792
<< metal1 >>
rect 1152 14678 13056 14700
rect 1152 14626 4966 14678
rect 5018 14626 5030 14678
rect 5082 14626 5094 14678
rect 5146 14626 5158 14678
rect 5210 14626 5222 14678
rect 5274 14626 5286 14678
rect 5338 14626 10966 14678
rect 11018 14626 11030 14678
rect 11082 14626 11094 14678
rect 11146 14626 11158 14678
rect 11210 14626 11222 14678
rect 11274 14626 11286 14678
rect 11338 14626 13056 14678
rect 1152 14604 13056 14626
rect 11536 14555 11542 14567
rect 8770 14527 11542 14555
rect 5602 14453 7358 14481
rect 1840 14367 1846 14419
rect 1898 14407 1904 14419
rect 2131 14410 2189 14416
rect 2131 14407 2143 14410
rect 1898 14379 2143 14407
rect 1898 14367 1904 14379
rect 2131 14376 2143 14379
rect 2177 14376 2189 14410
rect 2131 14370 2189 14376
rect 3280 14367 3286 14419
rect 3338 14367 3344 14419
rect 3955 14410 4013 14416
rect 3955 14376 3967 14410
rect 4001 14407 4013 14410
rect 5602 14407 5630 14453
rect 4001 14379 5630 14407
rect 4001 14376 4013 14379
rect 3955 14370 4013 14376
rect 6160 14367 6166 14419
rect 6218 14407 6224 14419
rect 7330 14416 7358 14453
rect 6739 14410 6797 14416
rect 6739 14407 6751 14410
rect 6218 14379 6751 14407
rect 6218 14367 6224 14379
rect 6739 14376 6751 14379
rect 6785 14376 6797 14410
rect 6739 14370 6797 14376
rect 7315 14410 7373 14416
rect 7315 14376 7327 14410
rect 7361 14376 7373 14410
rect 7315 14370 7373 14376
rect 7888 14367 7894 14419
rect 7946 14367 7952 14419
rect 8770 14416 8798 14527
rect 11536 14515 11542 14527
rect 11594 14515 11600 14567
rect 12211 14484 12269 14490
rect 12211 14481 12223 14484
rect 11362 14453 12223 14481
rect 8755 14410 8813 14416
rect 8755 14376 8767 14410
rect 8801 14376 8813 14410
rect 8755 14370 8813 14376
rect 9136 14367 9142 14419
rect 9194 14367 9200 14419
rect 9328 14367 9334 14419
rect 9386 14407 9392 14419
rect 11362 14416 11390 14453
rect 12211 14450 12223 14453
rect 12257 14450 12269 14484
rect 12211 14444 12269 14450
rect 10195 14410 10253 14416
rect 10195 14407 10207 14410
rect 9386 14379 10207 14407
rect 9386 14367 9392 14379
rect 10195 14376 10207 14379
rect 10241 14376 10253 14410
rect 10195 14370 10253 14376
rect 11347 14410 11405 14416
rect 11347 14376 11359 14410
rect 11393 14376 11405 14410
rect 11731 14410 11789 14416
rect 11731 14407 11743 14410
rect 11347 14370 11405 14376
rect 11458 14379 11743 14407
rect 2707 14336 2765 14342
rect 2707 14302 2719 14336
rect 2753 14302 2765 14336
rect 2707 14296 2765 14302
rect 2899 14336 2957 14342
rect 2899 14302 2911 14336
rect 2945 14333 2957 14336
rect 2945 14305 3998 14333
rect 2945 14302 2957 14305
rect 2899 14296 2957 14302
rect 1744 14219 1750 14271
rect 1802 14219 1808 14271
rect 1843 14262 1901 14268
rect 1843 14228 1855 14262
rect 1889 14259 1901 14262
rect 2722 14259 2750 14296
rect 3970 14271 3998 14305
rect 5584 14293 5590 14345
rect 5642 14293 5648 14345
rect 5680 14293 5686 14345
rect 5738 14333 5744 14345
rect 5738 14305 7454 14333
rect 5738 14293 5744 14305
rect 1889 14231 2750 14259
rect 1889 14228 1901 14231
rect 1843 14222 1901 14228
rect 1936 14145 1942 14197
rect 1994 14185 2000 14197
rect 2227 14188 2285 14194
rect 2227 14185 2239 14188
rect 1994 14157 2239 14185
rect 1994 14145 2000 14157
rect 2227 14154 2239 14157
rect 2273 14154 2285 14188
rect 2722 14185 2750 14231
rect 3376 14219 3382 14271
rect 3434 14219 3440 14271
rect 3952 14219 3958 14271
rect 4010 14219 4016 14271
rect 4048 14219 4054 14271
rect 4106 14259 4112 14271
rect 7426 14268 7454 14305
rect 11056 14293 11062 14345
rect 11114 14333 11120 14345
rect 11458 14333 11486 14379
rect 11731 14376 11743 14379
rect 11777 14376 11789 14410
rect 12304 14407 12310 14419
rect 11731 14370 11789 14376
rect 11842 14379 12310 14407
rect 11114 14305 11486 14333
rect 11114 14293 11120 14305
rect 5971 14262 6029 14268
rect 4106 14231 4464 14259
rect 4106 14219 4112 14231
rect 5971 14228 5983 14262
rect 6017 14259 6029 14262
rect 7411 14262 7469 14268
rect 6017 14231 7214 14259
rect 6017 14228 6029 14231
rect 5971 14222 6029 14228
rect 2722 14157 5726 14185
rect 2227 14148 2285 14154
rect 5698 14123 5726 14157
rect 6544 14145 6550 14197
rect 6602 14185 6608 14197
rect 6835 14188 6893 14194
rect 6835 14185 6847 14188
rect 6602 14157 6847 14185
rect 6602 14145 6608 14157
rect 6835 14154 6847 14157
rect 6881 14154 6893 14188
rect 6835 14148 6893 14154
rect 5680 14071 5686 14123
rect 5738 14071 5744 14123
rect 7186 14111 7214 14231
rect 7411 14228 7423 14262
rect 7457 14228 7469 14262
rect 7411 14222 7469 14228
rect 7984 14219 7990 14271
rect 8042 14219 8048 14271
rect 11251 14262 11309 14268
rect 11251 14228 11263 14262
rect 11297 14259 11309 14262
rect 11842 14259 11870 14379
rect 12304 14367 12310 14379
rect 12362 14367 12368 14419
rect 12016 14293 12022 14345
rect 12074 14333 12080 14345
rect 12403 14336 12461 14342
rect 12403 14333 12415 14336
rect 12074 14305 12415 14333
rect 12074 14293 12080 14305
rect 12403 14302 12415 14305
rect 12449 14302 12461 14336
rect 12403 14296 12461 14302
rect 11297 14231 11870 14259
rect 11297 14228 11309 14231
rect 11251 14222 11309 14228
rect 8467 14188 8525 14194
rect 8467 14154 8479 14188
rect 8513 14185 8525 14188
rect 8656 14185 8662 14197
rect 8513 14157 8662 14185
rect 8513 14154 8525 14157
rect 8467 14148 8525 14154
rect 8656 14145 8662 14157
rect 8714 14145 8720 14197
rect 8848 14145 8854 14197
rect 8906 14185 8912 14197
rect 9235 14188 9293 14194
rect 9235 14185 9247 14188
rect 8906 14157 9247 14185
rect 8906 14145 8912 14157
rect 9235 14154 9247 14157
rect 9281 14154 9293 14188
rect 9235 14148 9293 14154
rect 10000 14145 10006 14197
rect 10058 14185 10064 14197
rect 10291 14188 10349 14194
rect 10291 14185 10303 14188
rect 10058 14157 10303 14185
rect 10058 14145 10064 14157
rect 10291 14154 10303 14157
rect 10337 14154 10349 14188
rect 10291 14148 10349 14154
rect 11440 14145 11446 14197
rect 11498 14185 11504 14197
rect 11827 14188 11885 14194
rect 11827 14185 11839 14188
rect 11498 14157 11839 14185
rect 11498 14145 11504 14157
rect 11827 14154 11839 14157
rect 11873 14154 11885 14188
rect 11827 14148 11885 14154
rect 9616 14111 9622 14123
rect 7186 14083 9622 14111
rect 9616 14071 9622 14083
rect 9674 14071 9680 14123
rect 1152 14012 13056 14034
rect 1152 13960 1966 14012
rect 2018 13960 2030 14012
rect 2082 13960 2094 14012
rect 2146 13960 2158 14012
rect 2210 13960 2222 14012
rect 2274 13960 2286 14012
rect 2338 13960 7966 14012
rect 8018 13960 8030 14012
rect 8082 13960 8094 14012
rect 8146 13960 8158 14012
rect 8210 13960 8222 14012
rect 8274 13960 8286 14012
rect 8338 13960 13056 14012
rect 1152 13938 13056 13960
rect 1747 13892 1805 13898
rect 1747 13858 1759 13892
rect 1793 13889 1805 13892
rect 3280 13889 3286 13901
rect 1793 13861 3286 13889
rect 1793 13858 1805 13861
rect 1747 13852 1805 13858
rect 3280 13849 3286 13861
rect 3338 13849 3344 13901
rect 4240 13849 4246 13901
rect 4298 13889 4304 13901
rect 4531 13892 4589 13898
rect 4531 13889 4543 13892
rect 4298 13861 4543 13889
rect 4298 13849 4304 13861
rect 4531 13858 4543 13861
rect 4577 13858 4589 13892
rect 4531 13852 4589 13858
rect 7795 13892 7853 13898
rect 7795 13858 7807 13892
rect 7841 13889 7853 13892
rect 7888 13889 7894 13901
rect 7841 13861 7894 13889
rect 7841 13858 7853 13861
rect 7795 13852 7853 13858
rect 7888 13849 7894 13861
rect 7946 13849 7952 13901
rect 8467 13892 8525 13898
rect 8467 13858 8479 13892
rect 8513 13889 8525 13892
rect 8560 13889 8566 13901
rect 8513 13861 8566 13889
rect 8513 13858 8525 13861
rect 8467 13852 8525 13858
rect 8560 13849 8566 13861
rect 8618 13849 8624 13901
rect 11056 13849 11062 13901
rect 11114 13849 11120 13901
rect 5584 13815 5590 13827
rect 5410 13787 5590 13815
rect 4048 13741 4054 13753
rect 3504 13713 4054 13741
rect 4048 13701 4054 13713
rect 4106 13701 4112 13753
rect 3283 13670 3341 13676
rect 3283 13636 3295 13670
rect 3329 13667 3341 13670
rect 3568 13667 3574 13679
rect 3329 13639 3574 13667
rect 3329 13636 3341 13639
rect 3283 13630 3341 13636
rect 3568 13627 3574 13639
rect 3626 13627 3632 13679
rect 4240 13627 4246 13679
rect 4298 13627 4304 13679
rect 3667 13596 3725 13602
rect 3667 13562 3679 13596
rect 3713 13562 3725 13596
rect 3667 13556 3725 13562
rect 3682 13519 3710 13556
rect 3952 13553 3958 13605
rect 4010 13593 4016 13605
rect 4258 13593 4286 13627
rect 4010 13565 4286 13593
rect 4010 13553 4016 13565
rect 4432 13553 4438 13605
rect 4490 13553 4496 13605
rect 5410 13593 5438 13787
rect 5584 13775 5590 13787
rect 5642 13815 5648 13827
rect 5642 13787 8222 13815
rect 5642 13775 5648 13787
rect 5680 13701 5686 13753
rect 5738 13741 5744 13753
rect 8194 13750 8222 13787
rect 9238 13753 9290 13759
rect 8179 13744 8237 13750
rect 5738 13713 6000 13741
rect 5738 13701 5744 13713
rect 8179 13710 8191 13744
rect 8225 13710 8237 13744
rect 8179 13704 8237 13710
rect 5488 13627 5494 13679
rect 5546 13676 5552 13679
rect 5546 13670 5565 13676
rect 5553 13667 5565 13670
rect 6163 13670 6221 13676
rect 6163 13667 6175 13670
rect 5553 13639 6175 13667
rect 5553 13636 5565 13639
rect 5546 13630 5565 13636
rect 6163 13636 6175 13639
rect 6209 13636 6221 13670
rect 8194 13667 8222 13704
rect 9238 13695 9290 13701
rect 9427 13670 9485 13676
rect 9427 13667 9439 13670
rect 8194 13639 9439 13667
rect 6163 13630 6221 13636
rect 9427 13636 9439 13639
rect 9473 13667 9485 13670
rect 9473 13639 9854 13667
rect 9473 13636 9485 13639
rect 9427 13630 9485 13636
rect 5546 13627 5552 13630
rect 5587 13596 5645 13602
rect 5587 13593 5599 13596
rect 5410 13565 5599 13593
rect 5587 13562 5599 13565
rect 5633 13562 5645 13596
rect 5587 13556 5645 13562
rect 5776 13553 5782 13605
rect 5834 13553 5840 13605
rect 7792 13553 7798 13605
rect 7850 13593 7856 13605
rect 8083 13596 8141 13602
rect 8083 13593 8095 13596
rect 7850 13565 8095 13593
rect 7850 13553 7856 13565
rect 8083 13562 8095 13565
rect 8129 13562 8141 13596
rect 8083 13556 8141 13562
rect 8755 13596 8813 13602
rect 8755 13562 8767 13596
rect 8801 13562 8813 13596
rect 8755 13556 8813 13562
rect 8656 13519 8662 13531
rect 3682 13491 8662 13519
rect 8656 13479 8662 13491
rect 8714 13479 8720 13531
rect 8770 13519 8798 13556
rect 8944 13553 8950 13605
rect 9002 13593 9008 13605
rect 9043 13596 9101 13602
rect 9043 13593 9055 13596
rect 9002 13565 9055 13593
rect 9002 13553 9008 13565
rect 9043 13562 9055 13565
rect 9089 13562 9101 13596
rect 9043 13556 9101 13562
rect 8770 13491 9470 13519
rect 9442 13457 9470 13491
rect 9826 13457 9854 13639
rect 11923 13596 11981 13602
rect 11923 13562 11935 13596
rect 11969 13593 11981 13596
rect 12400 13593 12406 13605
rect 11969 13565 12406 13593
rect 11969 13562 11981 13565
rect 11923 13556 11981 13562
rect 12400 13553 12406 13565
rect 12458 13553 12464 13605
rect 12499 13596 12557 13602
rect 12499 13562 12511 13596
rect 12545 13593 12557 13596
rect 12784 13593 12790 13605
rect 12545 13565 12790 13593
rect 12545 13562 12557 13565
rect 12499 13556 12557 13562
rect 12784 13553 12790 13565
rect 12842 13553 12848 13605
rect 9424 13405 9430 13457
rect 9482 13405 9488 13457
rect 9808 13405 9814 13457
rect 9866 13405 9872 13457
rect 11635 13448 11693 13454
rect 11635 13414 11647 13448
rect 11681 13445 11693 13448
rect 11824 13445 11830 13457
rect 11681 13417 11830 13445
rect 11681 13414 11693 13417
rect 11635 13408 11693 13414
rect 11824 13405 11830 13417
rect 11882 13405 11888 13457
rect 12211 13448 12269 13454
rect 12211 13414 12223 13448
rect 12257 13445 12269 13448
rect 12400 13445 12406 13457
rect 12257 13417 12406 13445
rect 12257 13414 12269 13417
rect 12211 13408 12269 13414
rect 12400 13405 12406 13417
rect 12458 13405 12464 13457
rect 1152 13346 13056 13368
rect 1152 13294 4966 13346
rect 5018 13294 5030 13346
rect 5082 13294 5094 13346
rect 5146 13294 5158 13346
rect 5210 13294 5222 13346
rect 5274 13294 5286 13346
rect 5338 13294 10966 13346
rect 11018 13294 11030 13346
rect 11082 13294 11094 13346
rect 11146 13294 11158 13346
rect 11210 13294 11222 13346
rect 11274 13294 11286 13346
rect 11338 13294 13056 13346
rect 1152 13272 13056 13294
rect 1744 13183 1750 13235
rect 1802 13223 1808 13235
rect 1843 13226 1901 13232
rect 1843 13223 1855 13226
rect 1802 13195 1855 13223
rect 1802 13183 1808 13195
rect 1843 13192 1855 13195
rect 1889 13192 1901 13226
rect 1843 13186 1901 13192
rect 2035 13226 2093 13232
rect 2035 13192 2047 13226
rect 2081 13223 2093 13226
rect 4432 13223 4438 13235
rect 2081 13195 4438 13223
rect 2081 13192 2093 13195
rect 2035 13186 2093 13192
rect 4432 13183 4438 13195
rect 4490 13183 4496 13235
rect 6160 13183 6166 13235
rect 6218 13183 6224 13235
rect 8083 13226 8141 13232
rect 8083 13192 8095 13226
rect 8129 13223 8141 13226
rect 9328 13223 9334 13235
rect 8129 13195 9334 13223
rect 8129 13192 8141 13195
rect 8083 13186 8141 13192
rect 9328 13183 9334 13195
rect 9386 13183 9392 13235
rect 10483 13226 10541 13232
rect 10483 13192 10495 13226
rect 10529 13223 10541 13226
rect 10672 13223 10678 13235
rect 10529 13195 10678 13223
rect 10529 13192 10541 13195
rect 10483 13186 10541 13192
rect 10672 13183 10678 13195
rect 10730 13183 10736 13235
rect 11635 13226 11693 13232
rect 11635 13223 11647 13226
rect 10786 13195 11647 13223
rect 8464 13149 8470 13161
rect 4066 13121 8470 13149
rect 4066 13084 4094 13121
rect 8464 13109 8470 13121
rect 8522 13109 8528 13161
rect 8656 13109 8662 13161
rect 8714 13149 8720 13161
rect 10000 13149 10006 13161
rect 8714 13121 10006 13149
rect 8714 13109 8720 13121
rect 10000 13109 10006 13121
rect 10058 13109 10064 13161
rect 10786 13149 10814 13195
rect 11635 13192 11647 13195
rect 11681 13192 11693 13226
rect 11635 13186 11693 13192
rect 12016 13183 12022 13235
rect 12074 13183 12080 13235
rect 12304 13183 12310 13235
rect 12362 13183 12368 13235
rect 10690 13121 10814 13149
rect 11059 13152 11117 13158
rect 10690 13087 10718 13121
rect 11059 13118 11071 13152
rect 11105 13149 11117 13152
rect 12322 13149 12350 13183
rect 11105 13121 12350 13149
rect 11105 13118 11117 13121
rect 11059 13112 11117 13118
rect 4051 13078 4109 13084
rect 4051 13044 4063 13078
rect 4097 13044 4109 13078
rect 5488 13075 5494 13087
rect 4051 13038 4109 13044
rect 4162 13047 5494 13075
rect 784 12961 790 13013
rect 842 13001 848 13013
rect 1555 13004 1613 13010
rect 1555 13001 1567 13004
rect 842 12973 1567 13001
rect 842 12961 848 12973
rect 1555 12970 1567 12973
rect 1601 12970 1613 13004
rect 1555 12964 1613 12970
rect 3568 12961 3574 13013
rect 3626 13001 3632 13013
rect 3667 13004 3725 13010
rect 3667 13001 3679 13004
rect 3626 12973 3679 13001
rect 3626 12961 3632 12973
rect 3667 12970 3679 12973
rect 3713 13001 3725 13004
rect 4162 13001 4190 13047
rect 4432 13001 4438 13013
rect 3713 12973 4190 13001
rect 4258 12973 4438 13001
rect 3713 12970 3725 12973
rect 3667 12964 3725 12970
rect 4147 12930 4205 12936
rect 3874 12853 3902 12913
rect 4147 12896 4159 12930
rect 4193 12927 4205 12930
rect 4258 12927 4286 12973
rect 4432 12961 4438 12973
rect 4490 12961 4496 13013
rect 4546 13010 4574 13047
rect 5488 13035 5494 13047
rect 5546 13035 5552 13087
rect 9808 13035 9814 13087
rect 9866 13075 9872 13087
rect 9866 13047 10334 13075
rect 9866 13035 9872 13047
rect 4531 13004 4589 13010
rect 4531 12970 4543 13004
rect 4577 12970 4589 13004
rect 4531 12964 4589 12970
rect 9715 13004 9773 13010
rect 9715 12970 9727 13004
rect 9761 13001 9773 13004
rect 9826 13001 9854 13035
rect 9761 12973 9854 13001
rect 10099 13004 10157 13010
rect 9761 12970 9773 12973
rect 9715 12964 9773 12970
rect 10099 12970 10111 13004
rect 10145 13001 10157 13004
rect 10192 13001 10198 13013
rect 10145 12973 10198 13001
rect 10145 12970 10157 12973
rect 10099 12964 10157 12970
rect 10192 12961 10198 12973
rect 10250 12961 10256 13013
rect 10306 13001 10334 13047
rect 10672 13035 10678 13087
rect 10730 13035 10736 13087
rect 10768 13035 10774 13087
rect 10826 13035 10832 13087
rect 11347 13078 11405 13084
rect 11347 13044 11359 13078
rect 11393 13075 11405 13078
rect 11440 13075 11446 13087
rect 11393 13047 11446 13075
rect 11393 13044 11405 13047
rect 11347 13038 11405 13044
rect 11440 13035 11446 13047
rect 11498 13035 11504 13087
rect 11827 13078 11885 13084
rect 11827 13044 11839 13078
rect 11873 13044 11885 13078
rect 11827 13038 11885 13044
rect 11842 13001 11870 13038
rect 12208 13035 12214 13087
rect 12266 13035 12272 13087
rect 10306 12973 11870 13001
rect 4193 12899 4286 12927
rect 4193 12896 4205 12899
rect 4147 12890 4205 12896
rect 4048 12853 4054 12865
rect 3874 12825 4054 12853
rect 4048 12813 4054 12825
rect 4106 12853 4112 12865
rect 4354 12853 4382 12913
rect 8752 12887 8758 12939
rect 8810 12887 8816 12939
rect 4106 12825 4382 12853
rect 8770 12853 8798 12887
rect 9232 12853 9238 12865
rect 8770 12825 9238 12853
rect 4106 12813 4112 12825
rect 9232 12813 9238 12825
rect 9290 12813 9296 12865
rect 12496 12739 12502 12791
rect 12554 12739 12560 12791
rect 1152 12680 13056 12702
rect 1152 12628 1966 12680
rect 2018 12628 2030 12680
rect 2082 12628 2094 12680
rect 2146 12628 2158 12680
rect 2210 12628 2222 12680
rect 2274 12628 2286 12680
rect 2338 12628 7966 12680
rect 8018 12628 8030 12680
rect 8082 12628 8094 12680
rect 8146 12628 8158 12680
rect 8210 12628 8222 12680
rect 8274 12628 8286 12680
rect 8338 12628 13056 12680
rect 1152 12606 13056 12628
rect 1747 12560 1805 12566
rect 1747 12526 1759 12560
rect 1793 12557 1805 12560
rect 1840 12557 1846 12569
rect 1793 12529 1846 12557
rect 1793 12526 1805 12529
rect 1747 12520 1805 12526
rect 1840 12517 1846 12529
rect 1898 12517 1904 12569
rect 6931 12560 6989 12566
rect 6931 12526 6943 12560
rect 6977 12557 6989 12560
rect 9136 12557 9142 12569
rect 6977 12529 9142 12557
rect 6977 12526 6989 12529
rect 6931 12520 6989 12526
rect 9136 12517 9142 12529
rect 9194 12517 9200 12569
rect 9904 12517 9910 12569
rect 9962 12557 9968 12569
rect 10195 12560 10253 12566
rect 10195 12557 10207 12560
rect 9962 12529 10207 12557
rect 9962 12517 9968 12529
rect 10195 12526 10207 12529
rect 10241 12526 10253 12560
rect 10195 12520 10253 12526
rect 8752 12483 8758 12495
rect 7330 12455 8758 12483
rect 4240 12409 4246 12421
rect 3504 12381 4246 12409
rect 4240 12369 4246 12381
rect 4298 12409 4304 12421
rect 7330 12409 7358 12455
rect 8752 12443 8758 12455
rect 8810 12443 8816 12495
rect 4298 12395 7358 12409
rect 10678 12421 10730 12427
rect 4298 12381 7344 12395
rect 4298 12369 4304 12381
rect 10678 12363 10730 12369
rect 3283 12338 3341 12344
rect 3283 12304 3295 12338
rect 3329 12335 3341 12338
rect 3568 12335 3574 12347
rect 3329 12307 3574 12335
rect 3329 12304 3341 12307
rect 3283 12298 3341 12304
rect 3568 12295 3574 12307
rect 3626 12295 3632 12347
rect 7216 12295 7222 12347
rect 7274 12335 7280 12347
rect 7792 12335 7798 12347
rect 7274 12307 7798 12335
rect 7274 12295 7280 12307
rect 7792 12295 7798 12307
rect 7850 12335 7856 12347
rect 8467 12338 8525 12344
rect 8467 12335 8479 12338
rect 7850 12307 8479 12335
rect 7850 12295 7856 12307
rect 8467 12304 8479 12307
rect 8513 12304 8525 12338
rect 8467 12298 8525 12304
rect 10864 12295 10870 12347
rect 10922 12295 10928 12347
rect 3667 12264 3725 12270
rect 3667 12230 3679 12264
rect 3713 12261 3725 12264
rect 6544 12261 6550 12273
rect 3713 12233 6550 12261
rect 3713 12230 3725 12233
rect 3667 12224 3725 12230
rect 6544 12221 6550 12233
rect 6602 12221 6608 12273
rect 8851 12264 8909 12270
rect 8851 12230 8863 12264
rect 8897 12261 8909 12264
rect 8944 12261 8950 12273
rect 8897 12233 8950 12261
rect 8897 12230 8909 12233
rect 8851 12224 8909 12230
rect 8944 12221 8950 12233
rect 9002 12221 9008 12273
rect 10291 12264 10349 12270
rect 10291 12230 10303 12264
rect 10337 12230 10349 12264
rect 10291 12224 10349 12230
rect 10306 12187 10334 12224
rect 10480 12221 10486 12273
rect 10538 12221 10544 12273
rect 12499 12190 12557 12196
rect 12499 12187 12511 12190
rect 10306 12159 12511 12187
rect 12499 12156 12511 12159
rect 12545 12156 12557 12190
rect 12499 12150 12557 12156
rect 1152 12014 13056 12036
rect 1152 11962 4966 12014
rect 5018 11962 5030 12014
rect 5082 11962 5094 12014
rect 5146 11962 5158 12014
rect 5210 11962 5222 12014
rect 5274 11962 5286 12014
rect 5338 11962 10966 12014
rect 11018 11962 11030 12014
rect 11082 11962 11094 12014
rect 11146 11962 11158 12014
rect 11210 11962 11222 12014
rect 11274 11962 11286 12014
rect 11338 11962 13056 12014
rect 1152 11940 13056 11962
rect 9424 11851 9430 11903
rect 9482 11851 9488 11903
rect 10480 11703 10486 11755
rect 10538 11743 10544 11755
rect 11443 11746 11501 11752
rect 11443 11743 11455 11746
rect 10538 11715 11455 11743
rect 10538 11703 10544 11715
rect 11443 11712 11455 11715
rect 11489 11712 11501 11746
rect 11443 11706 11501 11712
rect 12211 11746 12269 11752
rect 12211 11712 12223 11746
rect 12257 11712 12269 11746
rect 12211 11706 12269 11712
rect 2608 11629 2614 11681
rect 2666 11629 2672 11681
rect 2800 11629 2806 11681
rect 2858 11669 2864 11681
rect 4339 11672 4397 11678
rect 4339 11669 4351 11672
rect 2858 11641 4351 11669
rect 2858 11629 2864 11641
rect 4339 11638 4351 11641
rect 4385 11638 4397 11672
rect 4339 11632 4397 11638
rect 10960 11629 10966 11681
rect 11018 11669 11024 11681
rect 11059 11672 11117 11678
rect 11059 11669 11071 11672
rect 11018 11641 11071 11669
rect 11018 11629 11024 11641
rect 11059 11638 11071 11641
rect 11105 11669 11117 11672
rect 12226 11669 12254 11706
rect 11105 11641 12254 11669
rect 11105 11638 11117 11641
rect 11059 11632 11117 11638
rect 1744 11555 1750 11607
rect 1802 11595 1808 11607
rect 2419 11598 2477 11604
rect 2419 11595 2431 11598
rect 1802 11567 2431 11595
rect 1802 11555 1808 11567
rect 2419 11564 2431 11567
rect 2465 11564 2477 11598
rect 2419 11558 2477 11564
rect 3955 11598 4013 11604
rect 3955 11564 3967 11598
rect 4001 11595 4013 11598
rect 4624 11595 4630 11607
rect 4001 11567 4630 11595
rect 4001 11564 4013 11567
rect 3955 11558 4013 11564
rect 4624 11555 4630 11567
rect 4682 11555 4688 11607
rect 9922 11521 9950 11581
rect 12496 11555 12502 11607
rect 12554 11555 12560 11607
rect 10672 11521 10678 11533
rect 9922 11493 10678 11521
rect 2704 11407 2710 11459
rect 2762 11447 2768 11459
rect 2803 11450 2861 11456
rect 2803 11447 2815 11450
rect 2762 11419 2815 11447
rect 2762 11407 2768 11419
rect 2803 11416 2815 11419
rect 2849 11416 2861 11450
rect 2803 11410 2861 11416
rect 8464 11407 8470 11459
rect 8522 11447 8528 11459
rect 9922 11447 9950 11493
rect 10672 11481 10678 11493
rect 10730 11481 10736 11533
rect 8522 11419 9950 11447
rect 8522 11407 8528 11419
rect 1152 11348 13056 11370
rect 1152 11296 1966 11348
rect 2018 11296 2030 11348
rect 2082 11296 2094 11348
rect 2146 11296 2158 11348
rect 2210 11296 2222 11348
rect 2274 11296 2286 11348
rect 2338 11296 7966 11348
rect 8018 11296 8030 11348
rect 8082 11296 8094 11348
rect 8146 11296 8158 11348
rect 8210 11296 8222 11348
rect 8274 11296 8286 11348
rect 8338 11296 13056 11348
rect 1152 11274 13056 11296
rect 1939 11228 1997 11234
rect 1939 11194 1951 11228
rect 1985 11225 1997 11228
rect 2608 11225 2614 11237
rect 1985 11197 2614 11225
rect 1985 11194 1997 11197
rect 1939 11188 1997 11194
rect 2608 11185 2614 11197
rect 2666 11185 2672 11237
rect 4624 11185 4630 11237
rect 4682 11185 4688 11237
rect 7216 11185 7222 11237
rect 7274 11185 7280 11237
rect 12499 11228 12557 11234
rect 12499 11194 12511 11228
rect 12545 11225 12557 11228
rect 12976 11225 12982 11237
rect 12545 11197 12982 11225
rect 12545 11194 12557 11197
rect 12499 11188 12557 11194
rect 12976 11185 12982 11197
rect 13034 11185 13040 11237
rect 10960 11151 10966 11163
rect 8386 11123 10966 11151
rect 4144 11077 4150 11089
rect 1666 11049 4150 11077
rect 1666 10938 1694 11049
rect 4144 11037 4150 11049
rect 4202 11037 4208 11089
rect 7216 11077 7222 11089
rect 6768 11049 7222 11077
rect 7216 11037 7222 11049
rect 7274 11037 7280 11089
rect 2323 11006 2381 11012
rect 2323 10972 2335 11006
rect 2369 10972 2381 11006
rect 2323 10966 2381 10972
rect 1651 10932 1709 10938
rect 1651 10898 1663 10932
rect 1697 10898 1709 10932
rect 1843 10932 1901 10938
rect 1843 10929 1855 10932
rect 1651 10892 1709 10898
rect 1762 10901 1855 10929
rect 1762 10781 1790 10901
rect 1843 10898 1855 10901
rect 1889 10898 1901 10932
rect 1843 10892 1901 10898
rect 1843 10858 1901 10864
rect 1843 10824 1855 10858
rect 1889 10855 1901 10858
rect 2338 10855 2366 10966
rect 2704 10963 2710 11015
rect 2762 11003 2768 11015
rect 3283 11006 3341 11012
rect 3283 11003 3295 11006
rect 2762 10975 3295 11003
rect 2762 10963 2768 10975
rect 3283 10972 3295 10975
rect 3329 10972 3341 11006
rect 3283 10966 3341 10972
rect 3376 10963 3382 11015
rect 3434 11003 3440 11015
rect 4435 11006 4493 11012
rect 4435 11003 4447 11006
rect 3434 10975 4447 11003
rect 3434 10963 3440 10975
rect 4435 10972 4447 10975
rect 4481 10972 4493 11006
rect 4435 10966 4493 10972
rect 4816 10963 4822 11015
rect 4874 10963 4880 11015
rect 5488 10963 5494 11015
rect 5546 11003 5552 11015
rect 5587 11006 5645 11012
rect 5587 11003 5599 11006
rect 5546 10975 5599 11003
rect 5546 10963 5552 10975
rect 5587 10972 5599 10975
rect 5633 10972 5645 11006
rect 8386 11003 8414 11123
rect 10960 11111 10966 11123
rect 11018 11111 11024 11163
rect 8464 11037 8470 11089
rect 8522 11077 8528 11089
rect 8522 11049 9264 11077
rect 8522 11037 8528 11049
rect 5587 10966 5645 10972
rect 5794 10975 8414 11003
rect 5794 10941 5822 10975
rect 8656 10963 8662 11015
rect 8714 10963 8720 11015
rect 9427 11006 9485 11012
rect 9427 11003 9439 11006
rect 8770 10975 9439 11003
rect 2611 10932 2669 10938
rect 2611 10898 2623 10932
rect 2657 10929 2669 10932
rect 4243 10932 4301 10938
rect 4243 10929 4255 10932
rect 2657 10901 4255 10929
rect 2657 10898 2669 10901
rect 2611 10892 2669 10898
rect 4243 10898 4255 10901
rect 4289 10898 4301 10932
rect 4243 10892 4301 10898
rect 5203 10932 5261 10938
rect 5203 10898 5215 10932
rect 5249 10929 5261 10932
rect 5776 10929 5782 10941
rect 5249 10901 5782 10929
rect 5249 10898 5261 10901
rect 5203 10892 5261 10898
rect 5776 10889 5782 10901
rect 5834 10889 5840 10941
rect 8464 10889 8470 10941
rect 8522 10889 8528 10941
rect 1889 10827 3902 10855
rect 1889 10824 1901 10827
rect 1843 10818 1901 10824
rect 3874 10793 3902 10827
rect 3091 10784 3149 10790
rect 3091 10781 3103 10784
rect 1762 10753 3103 10781
rect 3091 10750 3103 10753
rect 3137 10781 3149 10784
rect 3568 10781 3574 10793
rect 3137 10753 3574 10781
rect 3137 10750 3149 10753
rect 3091 10744 3149 10750
rect 3568 10741 3574 10753
rect 3626 10741 3632 10793
rect 3856 10741 3862 10793
rect 3914 10741 3920 10793
rect 7504 10741 7510 10793
rect 7562 10781 7568 10793
rect 8770 10781 8798 10975
rect 9427 10972 9439 10975
rect 9473 10972 9485 11006
rect 9427 10966 9485 10972
rect 9040 10889 9046 10941
rect 9098 10929 9104 10941
rect 10864 10929 10870 10941
rect 9098 10901 10870 10929
rect 9098 10889 9104 10901
rect 10864 10889 10870 10901
rect 10922 10929 10928 10941
rect 11635 10932 11693 10938
rect 11635 10929 11647 10932
rect 10922 10901 11647 10929
rect 10922 10889 10928 10901
rect 11635 10898 11647 10901
rect 11681 10898 11693 10932
rect 11635 10892 11693 10898
rect 11728 10889 11734 10941
rect 11786 10929 11792 10941
rect 12211 10932 12269 10938
rect 12211 10929 12223 10932
rect 11786 10901 12223 10929
rect 11786 10889 11792 10901
rect 12211 10898 12223 10901
rect 12257 10898 12269 10932
rect 12211 10892 12269 10898
rect 7562 10753 8798 10781
rect 7562 10741 7568 10753
rect 11920 10741 11926 10793
rect 11978 10741 11984 10793
rect 1152 10682 13056 10704
rect 1152 10630 4966 10682
rect 5018 10630 5030 10682
rect 5082 10630 5094 10682
rect 5146 10630 5158 10682
rect 5210 10630 5222 10682
rect 5274 10630 5286 10682
rect 5338 10630 10966 10682
rect 11018 10630 11030 10682
rect 11082 10630 11094 10682
rect 11146 10630 11158 10682
rect 11210 10630 11222 10682
rect 11274 10630 11286 10682
rect 11338 10630 13056 10682
rect 1152 10608 13056 10630
rect 3763 10562 3821 10568
rect 3763 10528 3775 10562
rect 3809 10559 3821 10562
rect 4048 10559 4054 10571
rect 3809 10531 4054 10559
rect 3809 10528 3821 10531
rect 3763 10522 3821 10528
rect 4048 10519 4054 10531
rect 4106 10519 4112 10571
rect 4816 10519 4822 10571
rect 4874 10519 4880 10571
rect 5776 10519 5782 10571
rect 5834 10519 5840 10571
rect 1939 10340 1997 10346
rect 1939 10306 1951 10340
rect 1985 10337 1997 10340
rect 2800 10337 2806 10349
rect 1985 10309 2806 10337
rect 1985 10306 1997 10309
rect 1939 10300 1997 10306
rect 2800 10297 2806 10309
rect 2858 10297 2864 10349
rect 3760 10297 3766 10349
rect 3818 10297 3824 10349
rect 3856 10297 3862 10349
rect 3914 10297 3920 10349
rect 4834 10337 4862 10519
rect 4066 10309 4862 10337
rect 5794 10337 5822 10519
rect 7120 10445 7126 10497
rect 7178 10485 7184 10497
rect 9136 10485 9142 10497
rect 7178 10457 9142 10485
rect 7178 10445 7184 10457
rect 9136 10445 9142 10457
rect 9194 10445 9200 10497
rect 10096 10411 10102 10423
rect 6082 10383 6686 10411
rect 5875 10340 5933 10346
rect 5875 10337 5887 10340
rect 5794 10309 5887 10337
rect 2323 10266 2381 10272
rect 2323 10232 2335 10266
rect 2369 10263 2381 10266
rect 2416 10263 2422 10275
rect 2369 10235 2422 10263
rect 2369 10232 2381 10235
rect 2323 10226 2381 10232
rect 2416 10223 2422 10235
rect 2474 10223 2480 10275
rect 4066 10272 4094 10309
rect 5875 10306 5887 10309
rect 5921 10306 5933 10340
rect 5875 10300 5933 10306
rect 4051 10266 4109 10272
rect 4051 10232 4063 10266
rect 4097 10232 4109 10266
rect 6082 10249 6110 10383
rect 6451 10340 6509 10346
rect 6451 10337 6463 10340
rect 6178 10309 6463 10337
rect 4051 10226 4109 10232
rect 5680 10149 5686 10201
rect 5738 10189 5744 10201
rect 6178 10189 6206 10309
rect 6451 10306 6463 10309
rect 6497 10306 6509 10340
rect 6451 10300 6509 10306
rect 6658 10272 6686 10383
rect 8290 10383 10102 10411
rect 8290 10346 8318 10383
rect 10096 10371 10102 10383
rect 10154 10371 10160 10423
rect 10960 10371 10966 10423
rect 11018 10411 11024 10423
rect 12211 10414 12269 10420
rect 12211 10411 12223 10414
rect 11018 10383 12223 10411
rect 11018 10371 11024 10383
rect 12211 10380 12223 10383
rect 12257 10380 12269 10414
rect 12211 10374 12269 10380
rect 8275 10340 8333 10346
rect 8275 10306 8287 10340
rect 8321 10306 8333 10340
rect 8275 10300 8333 10306
rect 8755 10340 8813 10346
rect 8755 10306 8767 10340
rect 8801 10337 8813 10340
rect 9040 10337 9046 10349
rect 8801 10309 9046 10337
rect 8801 10306 8813 10309
rect 8755 10300 8813 10306
rect 9040 10297 9046 10309
rect 9098 10297 9104 10349
rect 6259 10266 6317 10272
rect 6259 10232 6271 10266
rect 6305 10232 6317 10266
rect 6259 10226 6317 10232
rect 6643 10266 6701 10272
rect 6643 10232 6655 10266
rect 6689 10263 6701 10266
rect 7216 10263 7222 10275
rect 6689 10235 7222 10263
rect 6689 10232 6701 10235
rect 6643 10226 6701 10232
rect 5738 10161 6206 10189
rect 6274 10189 6302 10226
rect 7216 10223 7222 10235
rect 7274 10223 7280 10275
rect 8371 10266 8429 10272
rect 8371 10263 8383 10266
rect 8002 10235 8383 10263
rect 6274 10161 7358 10189
rect 5738 10149 5744 10161
rect 7330 10127 7358 10161
rect 3376 10075 3382 10127
rect 3434 10115 3440 10127
rect 3475 10118 3533 10124
rect 3475 10115 3487 10118
rect 3434 10087 3487 10115
rect 3434 10075 3440 10087
rect 3475 10084 3487 10087
rect 3521 10084 3533 10118
rect 3475 10078 3533 10084
rect 4243 10118 4301 10124
rect 4243 10084 4255 10118
rect 4289 10115 4301 10118
rect 7120 10115 7126 10127
rect 4289 10087 7126 10115
rect 4289 10084 4301 10087
rect 4243 10078 4301 10084
rect 7120 10075 7126 10087
rect 7178 10075 7184 10127
rect 7312 10075 7318 10127
rect 7370 10115 7376 10127
rect 8002 10124 8030 10235
rect 8371 10232 8383 10235
rect 8417 10232 8429 10266
rect 8371 10226 8429 10232
rect 9520 10223 9526 10275
rect 9578 10223 9584 10275
rect 9136 10149 9142 10201
rect 9194 10189 9200 10201
rect 10288 10189 10294 10201
rect 9194 10161 10294 10189
rect 9194 10149 9200 10161
rect 10288 10149 10294 10161
rect 10346 10149 10352 10201
rect 7987 10118 8045 10124
rect 7987 10115 7999 10118
rect 7370 10087 7999 10115
rect 7370 10075 7376 10087
rect 7987 10084 7999 10087
rect 8033 10084 8045 10118
rect 7987 10078 8045 10084
rect 10192 10075 10198 10127
rect 10250 10115 10256 10127
rect 10387 10118 10445 10124
rect 10387 10115 10399 10118
rect 10250 10087 10399 10115
rect 10250 10075 10256 10087
rect 10387 10084 10399 10087
rect 10433 10115 10445 10118
rect 10576 10115 10582 10127
rect 10433 10087 10582 10115
rect 10433 10084 10445 10087
rect 10387 10078 10445 10084
rect 10576 10075 10582 10087
rect 10634 10075 10640 10127
rect 12496 10075 12502 10127
rect 12554 10075 12560 10127
rect 1152 10016 13056 10038
rect 1152 9964 1966 10016
rect 2018 9964 2030 10016
rect 2082 9964 2094 10016
rect 2146 9964 2158 10016
rect 2210 9964 2222 10016
rect 2274 9964 2286 10016
rect 2338 9964 7966 10016
rect 8018 9964 8030 10016
rect 8082 9964 8094 10016
rect 8146 9964 8158 10016
rect 8210 9964 8222 10016
rect 8274 9964 8286 10016
rect 8338 9964 13056 10016
rect 1152 9942 13056 9964
rect 3760 9853 3766 9905
rect 3818 9893 3824 9905
rect 3859 9896 3917 9902
rect 3859 9893 3871 9896
rect 3818 9865 3871 9893
rect 3818 9853 3824 9865
rect 3859 9862 3871 9865
rect 3905 9862 3917 9896
rect 3859 9856 3917 9862
rect 8755 9896 8813 9902
rect 8755 9862 8767 9896
rect 8801 9893 8813 9896
rect 9040 9893 9046 9905
rect 8801 9865 9046 9893
rect 8801 9862 8813 9865
rect 8755 9856 8813 9862
rect 9040 9853 9046 9865
rect 9098 9853 9104 9905
rect 11536 9853 11542 9905
rect 11594 9893 11600 9905
rect 12403 9896 12461 9902
rect 12403 9893 12415 9896
rect 11594 9865 12415 9893
rect 11594 9853 11600 9865
rect 12403 9862 12415 9865
rect 12449 9862 12461 9896
rect 12403 9856 12461 9862
rect 7216 9819 7222 9831
rect 6466 9791 7222 9819
rect 2800 9705 2806 9757
rect 2858 9705 2864 9757
rect 6466 9731 6494 9791
rect 7216 9779 7222 9791
rect 7274 9819 7280 9831
rect 7274 9791 8606 9819
rect 7274 9779 7280 9791
rect 8464 9745 8470 9757
rect 8304 9717 8470 9745
rect 8464 9705 8470 9717
rect 8522 9705 8528 9757
rect 8578 9683 8606 9791
rect 10678 9757 10730 9763
rect 8656 9705 8662 9757
rect 8714 9745 8720 9757
rect 9520 9745 9526 9757
rect 8714 9717 9526 9745
rect 8714 9705 8720 9717
rect 9520 9705 9526 9717
rect 9578 9745 9584 9757
rect 9578 9717 10678 9745
rect 9578 9705 9584 9717
rect 10678 9699 10730 9705
rect 3379 9674 3437 9680
rect 3379 9640 3391 9674
rect 3425 9671 3437 9674
rect 3472 9671 3478 9683
rect 3425 9643 3478 9671
rect 3425 9640 3437 9643
rect 3379 9634 3437 9640
rect 3472 9631 3478 9643
rect 3530 9631 3536 9683
rect 3568 9631 3574 9683
rect 3626 9671 3632 9683
rect 4051 9674 4109 9680
rect 4051 9671 4063 9674
rect 3626 9643 4063 9671
rect 3626 9631 3632 9643
rect 4051 9640 4063 9643
rect 4097 9640 4109 9674
rect 4051 9634 4109 9640
rect 4528 9631 4534 9683
rect 4586 9671 4592 9683
rect 6259 9674 6317 9680
rect 6259 9671 6271 9674
rect 4586 9643 6271 9671
rect 4586 9631 4592 9643
rect 6259 9640 6271 9643
rect 6305 9671 6317 9674
rect 7123 9674 7181 9680
rect 7123 9671 7135 9674
rect 6305 9643 7135 9671
rect 6305 9640 6317 9643
rect 6259 9634 6317 9640
rect 7123 9640 7135 9643
rect 7169 9671 7181 9674
rect 7504 9671 7510 9683
rect 7169 9643 7510 9671
rect 7169 9640 7181 9643
rect 7123 9634 7181 9640
rect 7504 9631 7510 9643
rect 7562 9631 7568 9683
rect 8560 9631 8566 9683
rect 8618 9671 8624 9683
rect 9331 9674 9389 9680
rect 9331 9671 9343 9674
rect 8618 9643 9343 9671
rect 8618 9631 8624 9643
rect 9331 9640 9343 9643
rect 9377 9640 9389 9674
rect 9331 9634 9389 9640
rect 9811 9674 9869 9680
rect 9811 9640 9823 9674
rect 9857 9640 9869 9674
rect 9811 9634 9869 9640
rect 10867 9674 10925 9680
rect 10867 9640 10879 9674
rect 10913 9671 10925 9674
rect 10960 9671 10966 9683
rect 10913 9643 10966 9671
rect 10913 9640 10925 9643
rect 10867 9634 10925 9640
rect 4144 9557 4150 9609
rect 4202 9597 4208 9609
rect 4243 9600 4301 9606
rect 4243 9597 4255 9600
rect 4202 9569 4255 9597
rect 4202 9557 4208 9569
rect 4243 9566 4255 9569
rect 4289 9597 4301 9600
rect 5776 9597 5782 9609
rect 4289 9569 5782 9597
rect 4289 9566 4301 9569
rect 4243 9560 4301 9566
rect 5776 9557 5782 9569
rect 5834 9557 5840 9609
rect 6640 9557 6646 9609
rect 6698 9557 6704 9609
rect 6739 9600 6797 9606
rect 6739 9566 6751 9600
rect 6785 9597 6797 9600
rect 6785 9569 7454 9597
rect 6785 9566 6797 9569
rect 6739 9560 6797 9566
rect 4627 9526 4685 9532
rect 4627 9492 4639 9526
rect 4673 9523 4685 9526
rect 6754 9523 6782 9560
rect 4673 9495 6782 9523
rect 4673 9492 4685 9495
rect 4627 9486 4685 9492
rect 7426 9461 7454 9569
rect 8752 9557 8758 9609
rect 8810 9597 8816 9609
rect 9826 9597 9854 9634
rect 10960 9631 10966 9643
rect 11018 9631 11024 9683
rect 10480 9597 10486 9609
rect 8810 9569 9854 9597
rect 10114 9569 10486 9597
rect 8810 9557 8816 9569
rect 10114 9461 10142 9569
rect 10480 9557 10486 9569
rect 10538 9557 10544 9609
rect 7408 9409 7414 9461
rect 7466 9409 7472 9461
rect 10096 9409 10102 9461
rect 10154 9409 10160 9461
rect 1152 9350 13056 9372
rect 1152 9298 4966 9350
rect 5018 9298 5030 9350
rect 5082 9298 5094 9350
rect 5146 9298 5158 9350
rect 5210 9298 5222 9350
rect 5274 9298 5286 9350
rect 5338 9298 10966 9350
rect 11018 9298 11030 9350
rect 11082 9298 11094 9350
rect 11146 9298 11158 9350
rect 11210 9298 11222 9350
rect 11274 9298 11286 9350
rect 11338 9298 13056 9350
rect 1152 9276 13056 9298
rect 2515 9230 2573 9236
rect 2515 9196 2527 9230
rect 2561 9227 2573 9230
rect 4624 9227 4630 9239
rect 2561 9199 4630 9227
rect 2561 9196 2573 9199
rect 2515 9190 2573 9196
rect 4624 9187 4630 9199
rect 4682 9187 4688 9239
rect 10864 9187 10870 9239
rect 10922 9187 10928 9239
rect 11344 9187 11350 9239
rect 11402 9187 11408 9239
rect 12496 9187 12502 9239
rect 12554 9187 12560 9239
rect 2704 9153 2710 9165
rect 2338 9125 2710 9153
rect 2338 9014 2366 9125
rect 2704 9113 2710 9125
rect 2762 9153 2768 9165
rect 2762 9125 6590 9153
rect 2762 9113 2768 9125
rect 5392 9079 5398 9091
rect 4930 9051 5398 9079
rect 2227 9008 2285 9014
rect 2227 8974 2239 9008
rect 2273 8974 2285 9008
rect 2227 8968 2285 8974
rect 2323 9008 2381 9014
rect 2323 8974 2335 9008
rect 2369 8974 2381 9008
rect 2323 8968 2381 8974
rect 2899 9008 2957 9014
rect 2899 8974 2911 9008
rect 2945 8974 2957 9008
rect 2899 8968 2957 8974
rect 1840 8743 1846 8795
rect 1898 8783 1904 8795
rect 1939 8786 1997 8792
rect 1939 8783 1951 8786
rect 1898 8755 1951 8783
rect 1898 8743 1904 8755
rect 1939 8752 1951 8755
rect 1985 8752 1997 8786
rect 2242 8783 2270 8968
rect 2914 8857 2942 8968
rect 2992 8965 2998 9017
rect 3050 8965 3056 9017
rect 3187 9008 3245 9014
rect 3187 8974 3199 9008
rect 3233 9005 3245 9008
rect 4930 9005 4958 9051
rect 5392 9039 5398 9051
rect 5450 9079 5456 9091
rect 5587 9082 5645 9088
rect 5587 9079 5599 9082
rect 5450 9051 5599 9079
rect 5450 9039 5456 9051
rect 5587 9048 5599 9051
rect 5633 9048 5645 9082
rect 5587 9042 5645 9048
rect 5776 9039 5782 9091
rect 5834 9079 5840 9091
rect 6562 9088 6590 9125
rect 7408 9113 7414 9165
rect 7466 9153 7472 9165
rect 10882 9153 10910 9187
rect 7466 9125 10910 9153
rect 7466 9113 7472 9125
rect 6259 9082 6317 9088
rect 6259 9079 6271 9082
rect 5834 9051 6271 9079
rect 5834 9039 5840 9051
rect 6259 9048 6271 9051
rect 6305 9048 6317 9082
rect 6259 9042 6317 9048
rect 6547 9082 6605 9088
rect 6547 9048 6559 9082
rect 6593 9048 6605 9082
rect 6547 9042 6605 9048
rect 6643 9082 6701 9088
rect 6643 9048 6655 9082
rect 6689 9048 6701 9082
rect 6643 9042 6701 9048
rect 6739 9082 6797 9088
rect 6739 9048 6751 9082
rect 6785 9048 6797 9082
rect 6739 9042 6797 9048
rect 3233 8977 4958 9005
rect 3233 8974 3245 8977
rect 3187 8968 3245 8974
rect 5200 8965 5206 9017
rect 5258 8965 5264 9017
rect 5296 8965 5302 9017
rect 5354 8965 5360 9017
rect 5491 9008 5549 9014
rect 5491 8974 5503 9008
rect 5537 9005 5549 9008
rect 5794 9005 5822 9039
rect 5537 8977 5822 9005
rect 6274 9005 6302 9042
rect 6658 9005 6686 9042
rect 6274 8977 6686 9005
rect 5537 8974 5549 8977
rect 5491 8968 5549 8974
rect 3472 8891 3478 8943
rect 3530 8891 3536 8943
rect 6754 8931 6782 9042
rect 7426 9014 7454 9113
rect 9331 9082 9389 9088
rect 9331 9048 9343 9082
rect 9377 9079 9389 9082
rect 10096 9079 10102 9091
rect 9377 9051 10102 9079
rect 9377 9048 9389 9051
rect 9331 9042 9389 9048
rect 10096 9039 10102 9051
rect 10154 9039 10160 9091
rect 10960 9039 10966 9091
rect 11018 9079 11024 9091
rect 12211 9082 12269 9088
rect 12211 9079 12223 9082
rect 11018 9051 12223 9079
rect 11018 9039 11024 9051
rect 12211 9048 12223 9051
rect 12257 9048 12269 9082
rect 12211 9042 12269 9048
rect 7411 9008 7469 9014
rect 7411 8974 7423 9008
rect 7457 8974 7469 9008
rect 7411 8968 7469 8974
rect 9715 9008 9773 9014
rect 9715 8974 9727 9008
rect 9761 9005 9773 9008
rect 9808 9005 9814 9017
rect 9761 8977 9814 9005
rect 9761 8974 9773 8977
rect 9715 8968 9773 8974
rect 9808 8965 9814 8977
rect 9866 8965 9872 9017
rect 8566 8943 8618 8949
rect 4834 8903 6782 8931
rect 7027 8934 7085 8940
rect 3376 8857 3382 8869
rect 2914 8829 3382 8857
rect 3376 8817 3382 8829
rect 3434 8857 3440 8869
rect 4834 8857 4862 8903
rect 7027 8900 7039 8934
rect 7073 8931 7085 8934
rect 7120 8931 7126 8943
rect 7073 8903 7126 8931
rect 7073 8900 7085 8903
rect 7027 8894 7085 8900
rect 7120 8891 7126 8903
rect 7178 8891 7184 8943
rect 10672 8891 10678 8943
rect 10730 8891 10736 8943
rect 8566 8885 8618 8891
rect 3434 8829 4862 8857
rect 3434 8817 3440 8829
rect 5584 8817 5590 8869
rect 5642 8857 5648 8869
rect 6451 8860 6509 8866
rect 6451 8857 6463 8860
rect 5642 8829 6463 8857
rect 5642 8817 5648 8829
rect 6451 8826 6463 8829
rect 6497 8826 6509 8860
rect 6451 8820 6509 8826
rect 4336 8783 4342 8795
rect 2242 8755 4342 8783
rect 1939 8746 1997 8752
rect 4336 8743 4342 8755
rect 4394 8743 4400 8795
rect 5395 8786 5453 8792
rect 5395 8752 5407 8786
rect 5441 8783 5453 8786
rect 5776 8783 5782 8795
rect 5441 8755 5782 8783
rect 5441 8752 5453 8755
rect 5395 8746 5453 8752
rect 5776 8743 5782 8755
rect 5834 8743 5840 8795
rect 9040 8743 9046 8795
rect 9098 8743 9104 8795
rect 1152 8684 13056 8706
rect 1152 8632 1966 8684
rect 2018 8632 2030 8684
rect 2082 8632 2094 8684
rect 2146 8632 2158 8684
rect 2210 8632 2222 8684
rect 2274 8632 2286 8684
rect 2338 8632 7966 8684
rect 8018 8632 8030 8684
rect 8082 8632 8094 8684
rect 8146 8632 8158 8684
rect 8210 8632 8222 8684
rect 8274 8632 8286 8684
rect 8338 8632 13056 8684
rect 1152 8610 13056 8632
rect 1840 8521 1846 8573
rect 1898 8521 1904 8573
rect 5392 8521 5398 8573
rect 5450 8521 5456 8573
rect 10768 8521 10774 8573
rect 10826 8561 10832 8573
rect 12403 8564 12461 8570
rect 12403 8561 12415 8564
rect 10826 8533 12415 8561
rect 10826 8521 10832 8533
rect 12403 8530 12415 8533
rect 12449 8530 12461 8564
rect 12403 8524 12461 8530
rect 1858 8413 1886 8521
rect 6640 8447 6646 8499
rect 6698 8487 6704 8499
rect 6698 8459 9950 8487
rect 6698 8447 6704 8459
rect 6742 8425 6794 8431
rect 1858 8385 2078 8413
rect 1555 8342 1613 8348
rect 1555 8308 1567 8342
rect 1601 8308 1613 8342
rect 1555 8302 1613 8308
rect 1570 8265 1598 8302
rect 1744 8299 1750 8351
rect 1802 8299 1808 8351
rect 2050 8348 2078 8385
rect 6742 8367 6794 8373
rect 1843 8342 1901 8348
rect 1843 8308 1855 8342
rect 1889 8308 1901 8342
rect 1843 8302 1901 8308
rect 2035 8342 2093 8348
rect 2035 8308 2047 8342
rect 2081 8308 2093 8342
rect 2035 8302 2093 8308
rect 2131 8342 2189 8348
rect 2131 8308 2143 8342
rect 2177 8339 2189 8342
rect 2416 8339 2422 8351
rect 2177 8311 2422 8339
rect 2177 8308 2189 8311
rect 2131 8302 2189 8308
rect 1858 8265 1886 8302
rect 2416 8299 2422 8311
rect 2474 8299 2480 8351
rect 2800 8299 2806 8351
rect 2858 8339 2864 8351
rect 3859 8342 3917 8348
rect 3859 8339 3871 8342
rect 2858 8311 3871 8339
rect 2858 8299 2864 8311
rect 3859 8308 3871 8311
rect 3905 8308 3917 8342
rect 3859 8302 3917 8308
rect 7315 8342 7373 8348
rect 7315 8308 7327 8342
rect 7361 8339 7373 8342
rect 7792 8339 7798 8351
rect 7361 8311 7798 8339
rect 7361 8308 7373 8311
rect 7315 8302 7373 8308
rect 7792 8299 7798 8311
rect 7850 8339 7856 8351
rect 9808 8339 9814 8351
rect 7850 8311 9814 8339
rect 7850 8299 7856 8311
rect 9808 8299 9814 8311
rect 9866 8299 9872 8351
rect 9922 8339 9950 8459
rect 10678 8425 10730 8431
rect 10678 8367 10730 8373
rect 10867 8342 10925 8348
rect 10867 8339 10879 8342
rect 9922 8311 10879 8339
rect 10867 8308 10879 8311
rect 10913 8339 10925 8342
rect 10960 8339 10966 8351
rect 10913 8311 10966 8339
rect 10913 8308 10925 8311
rect 10867 8302 10925 8308
rect 10960 8299 10966 8311
rect 11018 8299 11024 8351
rect 1570 8237 1886 8265
rect 1858 8191 1886 8237
rect 2512 8225 2518 8277
rect 2570 8225 2576 8277
rect 4240 8225 4246 8277
rect 4298 8225 4304 8277
rect 7696 8225 7702 8277
rect 7754 8225 7760 8277
rect 10480 8225 10486 8277
rect 10538 8225 10544 8277
rect 5296 8191 5302 8203
rect 1858 8163 5302 8191
rect 5296 8151 5302 8163
rect 5354 8151 5360 8203
rect 1648 8077 1654 8129
rect 1706 8077 1712 8129
rect 1936 8077 1942 8129
rect 1994 8077 2000 8129
rect 3664 8077 3670 8129
rect 3722 8077 3728 8129
rect 4432 8077 4438 8129
rect 4490 8117 4496 8129
rect 5683 8120 5741 8126
rect 5683 8117 5695 8120
rect 4490 8089 5695 8117
rect 4490 8077 4496 8089
rect 5683 8086 5695 8089
rect 5729 8117 5741 8120
rect 10672 8117 10678 8129
rect 5729 8089 10678 8117
rect 5729 8086 5741 8089
rect 5683 8080 5741 8086
rect 10672 8077 10678 8089
rect 10730 8077 10736 8129
rect 1152 8018 13056 8040
rect 1152 7966 4966 8018
rect 5018 7966 5030 8018
rect 5082 7966 5094 8018
rect 5146 7966 5158 8018
rect 5210 7966 5222 8018
rect 5274 7966 5286 8018
rect 5338 7966 10966 8018
rect 11018 7966 11030 8018
rect 11082 7966 11094 8018
rect 11146 7966 11158 8018
rect 11210 7966 11222 8018
rect 11274 7966 11286 8018
rect 11338 7966 13056 8018
rect 1152 7944 13056 7966
rect 1648 7855 1654 7907
rect 1706 7855 1712 7907
rect 1936 7855 1942 7907
rect 1994 7855 2000 7907
rect 2320 7855 2326 7907
rect 2378 7895 2384 7907
rect 2419 7898 2477 7904
rect 2419 7895 2431 7898
rect 2378 7867 2431 7895
rect 2378 7855 2384 7867
rect 2419 7864 2431 7867
rect 2465 7864 2477 7898
rect 2419 7858 2477 7864
rect 2512 7855 2518 7907
rect 2570 7895 2576 7907
rect 3283 7898 3341 7904
rect 3283 7895 3295 7898
rect 2570 7867 3295 7895
rect 2570 7855 2576 7867
rect 3283 7864 3295 7867
rect 3329 7864 3341 7898
rect 3283 7858 3341 7864
rect 3664 7855 3670 7907
rect 3722 7855 3728 7907
rect 4240 7855 4246 7907
rect 4298 7895 4304 7907
rect 5491 7898 5549 7904
rect 5491 7895 5503 7898
rect 4298 7867 5503 7895
rect 4298 7855 4304 7867
rect 5491 7864 5503 7867
rect 5537 7864 5549 7898
rect 5491 7858 5549 7864
rect 12499 7898 12557 7904
rect 12499 7864 12511 7898
rect 12545 7895 12557 7898
rect 12880 7895 12886 7907
rect 12545 7867 12886 7895
rect 12545 7864 12557 7867
rect 12499 7858 12557 7864
rect 12880 7855 12886 7867
rect 12938 7855 12944 7907
rect 1666 7673 1694 7855
rect 1954 7747 1982 7855
rect 1954 7719 2894 7747
rect 2131 7676 2189 7682
rect 2131 7673 2143 7676
rect 1666 7645 2143 7673
rect 2131 7642 2143 7645
rect 2177 7642 2189 7676
rect 2866 7673 2894 7719
rect 3475 7676 3533 7682
rect 3475 7673 3487 7676
rect 2866 7645 3487 7673
rect 2131 7636 2189 7642
rect 3475 7642 3487 7645
rect 3521 7642 3533 7676
rect 3682 7673 3710 7855
rect 4816 7781 4822 7833
rect 4874 7781 4880 7833
rect 5011 7824 5069 7830
rect 5011 7790 5023 7824
rect 5057 7821 5069 7824
rect 5392 7821 5398 7833
rect 5057 7793 5398 7821
rect 5057 7790 5069 7793
rect 5011 7784 5069 7790
rect 5392 7781 5398 7793
rect 5450 7781 5456 7833
rect 9808 7781 9814 7833
rect 9866 7821 9872 7833
rect 10099 7824 10157 7830
rect 10099 7821 10111 7824
rect 9866 7793 10111 7821
rect 9866 7781 9872 7793
rect 10099 7790 10111 7793
rect 10145 7821 10157 7824
rect 10145 7793 12254 7821
rect 10145 7790 10157 7793
rect 10099 7784 10157 7790
rect 4051 7676 4109 7682
rect 4051 7673 4063 7676
rect 3682 7645 4063 7673
rect 3475 7636 3533 7642
rect 4051 7642 4063 7645
rect 4097 7642 4109 7676
rect 4051 7636 4109 7642
rect 4624 7633 4630 7685
rect 4682 7633 4688 7685
rect 4834 7682 4862 7781
rect 6736 7707 6742 7759
rect 6794 7707 6800 7759
rect 10384 7707 10390 7759
rect 10442 7747 10448 7759
rect 12226 7756 12254 7793
rect 11059 7750 11117 7756
rect 11059 7747 11071 7750
rect 10442 7719 11071 7747
rect 10442 7707 10448 7719
rect 11059 7716 11071 7719
rect 11105 7716 11117 7750
rect 11059 7710 11117 7716
rect 12211 7750 12269 7756
rect 12211 7716 12223 7750
rect 12257 7716 12269 7750
rect 12211 7710 12269 7716
rect 4819 7676 4877 7682
rect 4819 7642 4831 7676
rect 4865 7673 4877 7676
rect 5008 7673 5014 7685
rect 4865 7645 5014 7673
rect 4865 7642 4877 7645
rect 4819 7636 4877 7642
rect 5008 7633 5014 7645
rect 5066 7633 5072 7685
rect 5776 7633 5782 7685
rect 5834 7633 5840 7685
rect 6547 7676 6605 7682
rect 6547 7642 6559 7676
rect 6593 7673 6605 7676
rect 7120 7673 7126 7685
rect 6593 7645 7126 7673
rect 6593 7642 6605 7645
rect 6547 7636 6605 7642
rect 7120 7633 7126 7645
rect 7178 7633 7184 7685
rect 7504 7633 7510 7685
rect 7562 7673 7568 7685
rect 8467 7676 8525 7682
rect 8467 7673 8479 7676
rect 7562 7645 8479 7673
rect 7562 7633 7568 7645
rect 8467 7642 8479 7645
rect 8513 7642 8525 7676
rect 8467 7636 8525 7642
rect 2992 7559 2998 7611
rect 3050 7599 3056 7611
rect 3856 7599 3862 7611
rect 3050 7571 3862 7599
rect 3050 7559 3056 7571
rect 3856 7559 3862 7571
rect 3914 7559 3920 7611
rect 7888 7559 7894 7611
rect 7946 7599 7952 7611
rect 8083 7602 8141 7608
rect 8083 7599 8095 7602
rect 7946 7571 8095 7599
rect 7946 7559 7952 7571
rect 8083 7568 8095 7571
rect 8129 7568 8141 7602
rect 8083 7562 8141 7568
rect 9424 7559 9430 7611
rect 9482 7559 9488 7611
rect 11347 7602 11405 7608
rect 11347 7568 11359 7602
rect 11393 7599 11405 7602
rect 12304 7599 12310 7611
rect 11393 7571 12310 7599
rect 11393 7568 11405 7571
rect 11347 7562 11405 7568
rect 12304 7559 12310 7571
rect 12362 7559 12368 7611
rect 1152 7352 13056 7374
rect 1152 7300 1966 7352
rect 2018 7300 2030 7352
rect 2082 7300 2094 7352
rect 2146 7300 2158 7352
rect 2210 7300 2222 7352
rect 2274 7300 2286 7352
rect 2338 7300 7966 7352
rect 8018 7300 8030 7352
rect 8082 7300 8094 7352
rect 8146 7300 8158 7352
rect 8210 7300 8222 7352
rect 8274 7300 8286 7352
rect 8338 7300 13056 7352
rect 1152 7278 13056 7300
rect 6640 7229 6646 7241
rect 5890 7201 6646 7229
rect 4336 7115 4342 7167
rect 4394 7155 4400 7167
rect 5890 7164 5918 7201
rect 6640 7189 6646 7201
rect 6698 7189 6704 7241
rect 4531 7158 4589 7164
rect 4531 7155 4543 7158
rect 4394 7127 4543 7155
rect 4394 7115 4400 7127
rect 4531 7124 4543 7127
rect 4577 7124 4589 7158
rect 4531 7118 4589 7124
rect 5875 7158 5933 7164
rect 5875 7124 5887 7158
rect 5921 7124 5933 7158
rect 9424 7155 9430 7167
rect 5875 7118 5933 7124
rect 8674 7127 9430 7155
rect 2416 7041 2422 7093
rect 2474 7041 2480 7093
rect 4354 7053 5630 7081
rect 3379 7010 3437 7016
rect 3379 6976 3391 7010
rect 3425 7007 3437 7010
rect 3472 7007 3478 7019
rect 3425 6979 3478 7007
rect 3425 6976 3437 6979
rect 3379 6970 3437 6976
rect 3472 6967 3478 6979
rect 3530 6967 3536 7019
rect 4354 7016 4382 7053
rect 5602 7019 5630 7053
rect 6736 7041 6742 7093
rect 6794 7041 6800 7093
rect 7792 7041 7798 7093
rect 7850 7041 7856 7093
rect 8674 7090 8702 7127
rect 9424 7115 9430 7127
rect 9482 7115 9488 7167
rect 8659 7084 8717 7090
rect 7906 7053 8606 7081
rect 4339 7010 4397 7016
rect 4339 6976 4351 7010
rect 4385 6976 4397 7010
rect 4339 6970 4397 6976
rect 4432 6967 4438 7019
rect 4490 7007 4496 7019
rect 4819 7010 4877 7016
rect 4819 7007 4831 7010
rect 4490 6979 4831 7007
rect 4490 6967 4496 6979
rect 4819 6976 4831 6979
rect 4865 6976 4877 7010
rect 5491 7010 5549 7016
rect 5491 7007 5503 7010
rect 4819 6970 4877 6976
rect 4930 6979 5503 7007
rect 3856 6893 3862 6945
rect 3914 6893 3920 6945
rect 3952 6893 3958 6945
rect 4010 6933 4016 6945
rect 4930 6933 4958 6979
rect 5491 6976 5503 6979
rect 5537 6976 5549 7010
rect 5491 6970 5549 6976
rect 5584 6967 5590 7019
rect 5642 6967 5648 7019
rect 7411 7010 7469 7016
rect 7411 6976 7423 7010
rect 7457 7007 7469 7010
rect 7906 7007 7934 7053
rect 8578 7019 8606 7053
rect 8659 7050 8671 7084
rect 8705 7050 8717 7084
rect 9442 7067 9470 7115
rect 8659 7044 8717 7050
rect 12496 7041 12502 7093
rect 12554 7041 12560 7093
rect 7457 6979 7934 7007
rect 8467 7010 8525 7016
rect 7457 6976 7469 6979
rect 7411 6970 7469 6976
rect 8467 6976 8479 7010
rect 8513 6976 8525 7010
rect 8467 6970 8525 6976
rect 4010 6905 4958 6933
rect 4010 6893 4016 6905
rect 5008 6893 5014 6945
rect 5066 6933 5072 6945
rect 5203 6936 5261 6942
rect 5203 6933 5215 6936
rect 5066 6905 5215 6933
rect 5066 6893 5072 6905
rect 5203 6902 5215 6905
rect 5249 6902 5261 6936
rect 5203 6896 5261 6902
rect 7120 6893 7126 6945
rect 7178 6933 7184 6945
rect 8482 6933 8510 6970
rect 8560 6967 8566 7019
rect 8618 7007 8624 7019
rect 9427 7010 9485 7016
rect 9427 7007 9439 7010
rect 8618 6979 9439 7007
rect 8618 6967 8624 6979
rect 9427 6976 9439 6979
rect 9473 6976 9485 7010
rect 9427 6970 9485 6976
rect 9043 6936 9101 6942
rect 7178 6905 8606 6933
rect 7178 6893 7184 6905
rect 4336 6819 4342 6871
rect 4394 6859 4400 6871
rect 5026 6859 5054 6893
rect 8578 6871 8606 6905
rect 9043 6902 9055 6936
rect 9089 6933 9101 6936
rect 10384 6933 10390 6945
rect 9089 6905 10390 6933
rect 9089 6902 9101 6905
rect 9043 6896 9101 6902
rect 10384 6893 10390 6905
rect 10442 6893 10448 6945
rect 11632 6893 11638 6945
rect 11690 6893 11696 6945
rect 12211 6936 12269 6942
rect 12211 6902 12223 6936
rect 12257 6902 12269 6936
rect 12211 6896 12269 6902
rect 4394 6831 5054 6859
rect 4394 6819 4400 6831
rect 8560 6819 8566 6871
rect 8618 6819 8624 6871
rect 11920 6819 11926 6871
rect 11978 6819 11984 6871
rect 4624 6745 4630 6797
rect 4682 6745 4688 6797
rect 4816 6745 4822 6797
rect 4874 6785 4880 6797
rect 5299 6788 5357 6794
rect 5299 6785 5311 6788
rect 4874 6757 5311 6785
rect 4874 6745 4880 6757
rect 5299 6754 5311 6757
rect 5345 6754 5357 6788
rect 5299 6748 5357 6754
rect 7888 6745 7894 6797
rect 7946 6785 7952 6797
rect 10864 6785 10870 6797
rect 7946 6757 10870 6785
rect 7946 6745 7952 6757
rect 10864 6745 10870 6757
rect 10922 6785 10928 6797
rect 11059 6788 11117 6794
rect 11059 6785 11071 6788
rect 10922 6757 11071 6785
rect 10922 6745 10928 6757
rect 11059 6754 11071 6757
rect 11105 6785 11117 6788
rect 12226 6785 12254 6896
rect 11105 6757 12254 6785
rect 11105 6754 11117 6757
rect 11059 6748 11117 6754
rect 1152 6686 13056 6708
rect 1152 6634 4966 6686
rect 5018 6634 5030 6686
rect 5082 6634 5094 6686
rect 5146 6634 5158 6686
rect 5210 6634 5222 6686
rect 5274 6634 5286 6686
rect 5338 6634 10966 6686
rect 11018 6634 11030 6686
rect 11082 6634 11094 6686
rect 11146 6634 11158 6686
rect 11210 6634 11222 6686
rect 11274 6634 11286 6686
rect 11338 6634 13056 6686
rect 1152 6612 13056 6634
rect 3667 6566 3725 6572
rect 3667 6532 3679 6566
rect 3713 6532 3725 6566
rect 3667 6526 3725 6532
rect 3682 6489 3710 6526
rect 3952 6523 3958 6575
rect 4010 6523 4016 6575
rect 4336 6523 4342 6575
rect 4394 6523 4400 6575
rect 4816 6563 4822 6575
rect 4450 6535 4822 6563
rect 4354 6489 4382 6523
rect 3682 6461 4382 6489
rect 3763 6418 3821 6424
rect 3763 6384 3775 6418
rect 3809 6415 3821 6418
rect 4336 6415 4342 6427
rect 3809 6387 4342 6415
rect 3809 6384 3821 6387
rect 3763 6378 3821 6384
rect 4336 6375 4342 6387
rect 4394 6375 4400 6427
rect 4450 6424 4478 6535
rect 4816 6523 4822 6535
rect 4874 6523 4880 6575
rect 9616 6523 9622 6575
rect 9674 6563 9680 6575
rect 9811 6566 9869 6572
rect 9811 6563 9823 6566
rect 9674 6535 9823 6563
rect 9674 6523 9680 6535
rect 9811 6532 9823 6535
rect 9857 6532 9869 6566
rect 9811 6526 9869 6532
rect 4435 6418 4493 6424
rect 4435 6384 4447 6418
rect 4481 6384 4493 6418
rect 4435 6378 4493 6384
rect 7696 6375 7702 6427
rect 7754 6415 7760 6427
rect 7795 6418 7853 6424
rect 7795 6415 7807 6418
rect 7754 6387 7807 6415
rect 7754 6375 7760 6387
rect 7795 6384 7807 6387
rect 7841 6384 7853 6418
rect 7795 6378 7853 6384
rect 10288 6375 10294 6427
rect 10346 6415 10352 6427
rect 11059 6418 11117 6424
rect 11059 6415 11071 6418
rect 10346 6387 11071 6415
rect 10346 6375 10352 6387
rect 11059 6384 11071 6387
rect 11105 6384 11117 6418
rect 11059 6378 11117 6384
rect 12211 6418 12269 6424
rect 12211 6384 12223 6418
rect 12257 6384 12269 6418
rect 12211 6378 12269 6384
rect 1843 6344 1901 6350
rect 1843 6310 1855 6344
rect 1889 6341 1901 6344
rect 2416 6341 2422 6353
rect 1889 6313 2422 6341
rect 1889 6310 1901 6313
rect 1843 6304 1901 6310
rect 2416 6301 2422 6313
rect 2474 6341 2480 6353
rect 4051 6344 4109 6350
rect 4051 6341 4063 6344
rect 2474 6313 4063 6341
rect 2474 6301 2480 6313
rect 4051 6310 4063 6313
rect 4097 6310 4109 6344
rect 4051 6304 4109 6310
rect 7888 6301 7894 6353
rect 7946 6341 7952 6353
rect 8179 6344 8237 6350
rect 8179 6341 8191 6344
rect 7946 6313 8191 6341
rect 7946 6301 7952 6313
rect 8179 6310 8191 6313
rect 8225 6310 8237 6344
rect 8179 6304 8237 6310
rect 8560 6301 8566 6353
rect 8618 6341 8624 6353
rect 11923 6344 11981 6350
rect 11923 6341 11935 6344
rect 8618 6313 11935 6341
rect 8618 6301 8624 6313
rect 11923 6310 11935 6313
rect 11969 6310 11981 6344
rect 11923 6304 11981 6310
rect 2227 6270 2285 6276
rect 2227 6236 2239 6270
rect 2273 6267 2285 6270
rect 9424 6267 9430 6279
rect 2273 6239 2462 6267
rect 9360 6239 9430 6267
rect 2273 6236 2285 6239
rect 2227 6230 2285 6236
rect 2434 6205 2462 6239
rect 9424 6227 9430 6239
rect 9482 6227 9488 6279
rect 12226 6267 12254 6378
rect 9538 6239 12254 6267
rect 2416 6153 2422 6205
rect 2474 6153 2480 6205
rect 8560 6153 8566 6205
rect 8618 6193 8624 6205
rect 9538 6193 9566 6239
rect 12496 6227 12502 6279
rect 12554 6227 12560 6279
rect 11731 6196 11789 6202
rect 11731 6193 11743 6196
rect 8618 6165 9566 6193
rect 10786 6165 11743 6193
rect 8618 6153 8624 6165
rect 10786 6131 10814 6165
rect 11731 6162 11743 6165
rect 11777 6162 11789 6196
rect 11731 6156 11789 6162
rect 3376 6079 3382 6131
rect 3434 6079 3440 6131
rect 5584 6079 5590 6131
rect 5642 6079 5648 6131
rect 10768 6079 10774 6131
rect 10826 6079 10832 6131
rect 11344 6079 11350 6131
rect 11402 6079 11408 6131
rect 1152 6020 13056 6042
rect 1152 5968 1966 6020
rect 2018 5968 2030 6020
rect 2082 5968 2094 6020
rect 2146 5968 2158 6020
rect 2210 5968 2222 6020
rect 2274 5968 2286 6020
rect 2338 5968 7966 6020
rect 8018 5968 8030 6020
rect 8082 5968 8094 6020
rect 8146 5968 8158 6020
rect 8210 5968 8222 6020
rect 8274 5968 8286 6020
rect 8338 5968 13056 6020
rect 1152 5946 13056 5968
rect 2227 5900 2285 5906
rect 2227 5866 2239 5900
rect 2273 5897 2285 5900
rect 2416 5897 2422 5909
rect 2273 5869 2422 5897
rect 2273 5866 2285 5869
rect 2227 5860 2285 5866
rect 2416 5857 2422 5869
rect 2474 5857 2480 5909
rect 4336 5857 4342 5909
rect 4394 5897 4400 5909
rect 4627 5900 4685 5906
rect 4627 5897 4639 5900
rect 4394 5869 4639 5897
rect 4394 5857 4400 5869
rect 4627 5866 4639 5869
rect 4673 5866 4685 5900
rect 4627 5860 4685 5866
rect 4624 5749 4630 5761
rect 2530 5721 4630 5749
rect 2530 5684 2558 5721
rect 4624 5709 4630 5721
rect 4682 5709 4688 5761
rect 6736 5709 6742 5761
rect 6794 5709 6800 5761
rect 10480 5709 10486 5761
rect 10538 5709 10544 5761
rect 10768 5709 10774 5761
rect 10826 5709 10832 5761
rect 12499 5752 12557 5758
rect 12499 5718 12511 5752
rect 12545 5749 12557 5752
rect 12592 5749 12598 5761
rect 12545 5721 12598 5749
rect 12545 5718 12557 5721
rect 12499 5712 12557 5718
rect 12592 5709 12598 5721
rect 12650 5709 12656 5761
rect 2515 5678 2573 5684
rect 2515 5644 2527 5678
rect 2561 5644 2573 5678
rect 2515 5638 2573 5644
rect 2995 5678 3053 5684
rect 2995 5644 3007 5678
rect 3041 5644 3053 5678
rect 2995 5638 3053 5644
rect 3010 5527 3038 5638
rect 3376 5635 3382 5687
rect 3434 5675 3440 5687
rect 4435 5678 4493 5684
rect 4435 5675 4447 5678
rect 3434 5647 4447 5675
rect 3434 5635 3440 5647
rect 4435 5644 4447 5647
rect 4481 5644 4493 5678
rect 4435 5638 4493 5644
rect 4720 5635 4726 5687
rect 4778 5675 4784 5687
rect 4819 5678 4877 5684
rect 4819 5675 4831 5678
rect 4778 5647 4831 5675
rect 4778 5635 4784 5647
rect 4819 5644 4831 5647
rect 4865 5644 4877 5678
rect 4819 5638 4877 5644
rect 3283 5604 3341 5610
rect 3283 5570 3295 5604
rect 3329 5601 3341 5604
rect 4243 5604 4301 5610
rect 4243 5601 4255 5604
rect 3329 5573 4255 5601
rect 3329 5570 3341 5573
rect 3283 5564 3341 5570
rect 4243 5570 4255 5573
rect 4289 5570 4301 5604
rect 4243 5564 4301 5570
rect 5299 5604 5357 5610
rect 5299 5570 5311 5604
rect 5345 5601 5357 5604
rect 6754 5601 6782 5709
rect 7219 5678 7277 5684
rect 7219 5644 7231 5678
rect 7265 5644 7277 5678
rect 7219 5638 7277 5644
rect 5345 5573 6782 5601
rect 5345 5570 5357 5573
rect 5299 5564 5357 5570
rect 3379 5530 3437 5536
rect 3010 5499 3326 5527
rect 3298 5465 3326 5499
rect 3379 5496 3391 5530
rect 3425 5496 3437 5530
rect 3379 5490 3437 5496
rect 3667 5530 3725 5536
rect 3667 5496 3679 5530
rect 3713 5527 3725 5530
rect 4432 5527 4438 5539
rect 3713 5499 4438 5527
rect 3713 5496 3725 5499
rect 3667 5490 3725 5496
rect 3280 5413 3286 5465
rect 3338 5413 3344 5465
rect 3394 5453 3422 5490
rect 4432 5487 4438 5499
rect 4490 5487 4496 5539
rect 6640 5487 6646 5539
rect 6698 5527 6704 5539
rect 7234 5527 7262 5638
rect 7312 5635 7318 5687
rect 7370 5675 7376 5687
rect 7603 5678 7661 5684
rect 7603 5675 7615 5678
rect 7370 5647 7615 5675
rect 7370 5635 7376 5647
rect 7603 5644 7615 5647
rect 7649 5644 7661 5678
rect 7603 5638 7661 5644
rect 10864 5635 10870 5687
rect 10922 5635 10928 5687
rect 9235 5604 9293 5610
rect 9235 5570 9247 5604
rect 9281 5601 9293 5604
rect 9424 5601 9430 5613
rect 9281 5573 9430 5601
rect 9281 5570 9293 5573
rect 9235 5564 9293 5570
rect 9424 5561 9430 5573
rect 9482 5561 9488 5613
rect 10000 5561 10006 5613
rect 10058 5561 10064 5613
rect 6698 5499 7262 5527
rect 7906 5499 12254 5527
rect 6698 5487 6704 5499
rect 4144 5453 4150 5465
rect 3394 5425 4150 5453
rect 4144 5413 4150 5425
rect 4202 5413 4208 5465
rect 5587 5456 5645 5462
rect 5587 5422 5599 5456
rect 5633 5453 5645 5456
rect 5776 5453 5782 5465
rect 5633 5425 5782 5453
rect 5633 5422 5645 5425
rect 5587 5416 5645 5422
rect 5776 5413 5782 5425
rect 5834 5453 5840 5465
rect 7906 5453 7934 5499
rect 12226 5465 12254 5499
rect 5834 5425 7934 5453
rect 5834 5413 5840 5425
rect 9520 5413 9526 5465
rect 9578 5413 9584 5465
rect 10288 5413 10294 5465
rect 10346 5413 10352 5465
rect 12208 5413 12214 5465
rect 12266 5413 12272 5465
rect 1152 5354 13056 5376
rect 1152 5302 4966 5354
rect 5018 5302 5030 5354
rect 5082 5302 5094 5354
rect 5146 5302 5158 5354
rect 5210 5302 5222 5354
rect 5274 5302 5286 5354
rect 5338 5302 10966 5354
rect 11018 5302 11030 5354
rect 11082 5302 11094 5354
rect 11146 5302 11158 5354
rect 11210 5302 11222 5354
rect 11274 5302 11286 5354
rect 11338 5302 13056 5354
rect 1152 5280 13056 5302
rect 3280 5191 3286 5243
rect 3338 5231 3344 5243
rect 4720 5231 4726 5243
rect 3338 5203 4726 5231
rect 3338 5191 3344 5203
rect 4720 5191 4726 5203
rect 4778 5191 4784 5243
rect 5296 5191 5302 5243
rect 5354 5231 5360 5243
rect 5680 5231 5686 5243
rect 5354 5203 5686 5231
rect 5354 5191 5360 5203
rect 5680 5191 5686 5203
rect 5738 5191 5744 5243
rect 7120 5191 7126 5243
rect 7178 5191 7184 5243
rect 8368 5191 8374 5243
rect 8426 5231 8432 5243
rect 9043 5234 9101 5240
rect 9043 5231 9055 5234
rect 8426 5203 9055 5231
rect 8426 5191 8432 5203
rect 9043 5200 9055 5203
rect 9089 5200 9101 5234
rect 9043 5194 9101 5200
rect 12496 5191 12502 5243
rect 12554 5191 12560 5243
rect 5203 5160 5261 5166
rect 5203 5126 5215 5160
rect 5249 5157 5261 5160
rect 7138 5157 7166 5191
rect 5249 5129 7166 5157
rect 8755 5160 8813 5166
rect 5249 5126 5261 5129
rect 5203 5120 5261 5126
rect 4720 5043 4726 5095
rect 4778 5083 4784 5095
rect 5488 5083 5494 5095
rect 4778 5055 5494 5083
rect 4778 5043 4784 5055
rect 5488 5043 5494 5055
rect 5546 5043 5552 5095
rect 5011 5012 5069 5018
rect 5011 4978 5023 5012
rect 5057 5009 5069 5012
rect 5296 5009 5302 5021
rect 5057 4981 5302 5009
rect 5057 4978 5069 4981
rect 5011 4972 5069 4978
rect 5296 4969 5302 4981
rect 5354 4969 5360 5021
rect 5584 4969 5590 5021
rect 5642 4969 5648 5021
rect 5698 5018 5726 5129
rect 8755 5126 8767 5160
rect 8801 5157 8813 5160
rect 11728 5157 11734 5169
rect 8801 5129 11734 5157
rect 8801 5126 8813 5129
rect 8755 5120 8813 5126
rect 11728 5117 11734 5129
rect 11786 5117 11792 5169
rect 5875 5086 5933 5092
rect 5875 5052 5887 5086
rect 5921 5083 5933 5086
rect 5921 5055 7262 5083
rect 5921 5052 5933 5055
rect 5875 5046 5933 5052
rect 7234 5021 7262 5055
rect 10576 5043 10582 5095
rect 10634 5083 10640 5095
rect 12211 5086 12269 5092
rect 12211 5083 12223 5086
rect 10634 5055 12223 5083
rect 10634 5043 10640 5055
rect 12211 5052 12223 5055
rect 12257 5052 12269 5086
rect 12211 5046 12269 5052
rect 5683 5012 5741 5018
rect 5683 4978 5695 5012
rect 5729 4978 5741 5012
rect 5683 4972 5741 4978
rect 7120 4969 7126 5021
rect 7178 4969 7184 5021
rect 7216 4969 7222 5021
rect 7274 4969 7280 5021
rect 10384 4969 10390 5021
rect 10442 5009 10448 5021
rect 10675 5012 10733 5018
rect 10675 5009 10687 5012
rect 10442 4981 10687 5009
rect 10442 4969 10448 4981
rect 10675 4978 10687 4981
rect 10721 4978 10733 5012
rect 10675 4972 10733 4978
rect 9526 4947 9578 4953
rect 4528 4895 4534 4947
rect 4586 4935 4592 4947
rect 4627 4938 4685 4944
rect 4627 4935 4639 4938
rect 4586 4907 4639 4935
rect 4586 4895 4592 4907
rect 4627 4904 4639 4907
rect 4673 4904 4685 4938
rect 4627 4898 4685 4904
rect 6736 4895 6742 4947
rect 6794 4895 6800 4947
rect 8656 4935 8662 4947
rect 8304 4907 8662 4935
rect 8656 4895 8662 4907
rect 8714 4935 8720 4947
rect 8714 4907 9526 4935
rect 8714 4895 8720 4907
rect 11059 4938 11117 4944
rect 11059 4904 11071 4938
rect 11105 4904 11117 4938
rect 11059 4898 11117 4904
rect 9526 4889 9578 4895
rect 11074 4861 11102 4898
rect 10594 4833 11102 4861
rect 10594 4799 10622 4833
rect 10576 4747 10582 4799
rect 10634 4747 10640 4799
rect 1152 4688 13056 4710
rect 1152 4636 1966 4688
rect 2018 4636 2030 4688
rect 2082 4636 2094 4688
rect 2146 4636 2158 4688
rect 2210 4636 2222 4688
rect 2274 4636 2286 4688
rect 2338 4636 7966 4688
rect 8018 4636 8030 4688
rect 8082 4636 8094 4688
rect 8146 4636 8158 4688
rect 8210 4636 8222 4688
rect 8274 4636 8286 4688
rect 8338 4636 13056 4688
rect 1152 4614 13056 4636
rect 8656 4565 8662 4577
rect 6082 4537 8662 4565
rect 6082 4403 6110 4537
rect 8656 4525 8662 4537
rect 8714 4525 8720 4577
rect 8560 4451 8566 4503
rect 8618 4451 8624 4503
rect 7216 4377 7222 4429
rect 7274 4377 7280 4429
rect 5971 4346 6029 4352
rect 5971 4312 5983 4346
rect 6017 4343 6029 4346
rect 8179 4346 8237 4352
rect 6017 4315 6302 4343
rect 6017 4312 6029 4315
rect 5971 4306 6029 4312
rect 4051 4272 4109 4278
rect 4051 4238 4063 4272
rect 4097 4269 4109 4272
rect 4528 4269 4534 4281
rect 4097 4241 4534 4269
rect 4097 4238 4109 4241
rect 4051 4232 4109 4238
rect 4528 4229 4534 4241
rect 4586 4229 4592 4281
rect 3955 4124 4013 4130
rect 3955 4090 3967 4124
rect 4001 4121 4013 4124
rect 4240 4121 4246 4133
rect 4001 4093 4246 4121
rect 4001 4090 4013 4093
rect 3955 4084 4013 4090
rect 4240 4081 4246 4093
rect 4298 4081 4304 4133
rect 4339 4124 4397 4130
rect 4339 4090 4351 4124
rect 4385 4121 4397 4124
rect 4432 4121 4438 4133
rect 4385 4093 4438 4121
rect 4385 4090 4397 4093
rect 4339 4084 4397 4090
rect 4432 4081 4438 4093
rect 4490 4081 4496 4133
rect 6274 4121 6302 4315
rect 8179 4312 8191 4346
rect 8225 4343 8237 4346
rect 8464 4343 8470 4355
rect 8225 4315 8470 4343
rect 8225 4312 8237 4315
rect 8179 4306 8237 4312
rect 8464 4303 8470 4315
rect 8522 4303 8528 4355
rect 6355 4272 6413 4278
rect 6355 4238 6367 4272
rect 6401 4238 6413 4272
rect 6355 4232 6413 4238
rect 6370 4195 6398 4232
rect 7120 4229 7126 4281
rect 7178 4269 7184 4281
rect 7888 4269 7894 4281
rect 7178 4241 7894 4269
rect 7178 4229 7184 4241
rect 7888 4229 7894 4241
rect 7946 4269 7952 4281
rect 8578 4278 8606 4451
rect 10480 4417 10486 4429
rect 10114 4389 10486 4417
rect 10114 4343 10142 4389
rect 10480 4377 10486 4389
rect 10538 4377 10544 4429
rect 10768 4377 10774 4429
rect 10826 4377 10832 4429
rect 9538 4315 10142 4343
rect 8563 4272 8621 4278
rect 8563 4269 8575 4272
rect 7946 4241 8575 4269
rect 7946 4229 7952 4241
rect 8563 4238 8575 4241
rect 8609 4238 8621 4272
rect 8563 4232 8621 4238
rect 9424 4229 9430 4281
rect 9482 4229 9488 4281
rect 6736 4195 6742 4207
rect 6370 4167 6742 4195
rect 6736 4155 6742 4167
rect 6794 4195 6800 4207
rect 9538 4195 9566 4315
rect 10384 4303 10390 4355
rect 10442 4343 10448 4355
rect 10867 4346 10925 4352
rect 10867 4343 10879 4346
rect 10442 4315 10879 4343
rect 10442 4303 10448 4315
rect 10867 4312 10879 4315
rect 10913 4312 10925 4346
rect 10867 4306 10925 4312
rect 9616 4229 9622 4281
rect 9674 4269 9680 4281
rect 10003 4272 10061 4278
rect 10003 4269 10015 4272
rect 9674 4241 10015 4269
rect 9674 4229 9680 4241
rect 10003 4238 10015 4241
rect 10049 4238 10061 4272
rect 10003 4232 10061 4238
rect 12499 4272 12557 4278
rect 12499 4238 12511 4272
rect 12545 4269 12557 4272
rect 12784 4269 12790 4281
rect 12545 4241 12790 4269
rect 12545 4238 12557 4241
rect 12499 4232 12557 4238
rect 12784 4229 12790 4241
rect 12842 4229 12848 4281
rect 12688 4195 12694 4207
rect 6794 4167 9566 4195
rect 9730 4167 12694 4195
rect 6794 4155 6800 4167
rect 6547 4124 6605 4130
rect 6547 4121 6559 4124
rect 6274 4093 6559 4121
rect 6547 4090 6559 4093
rect 6593 4121 6605 4124
rect 6640 4121 6646 4133
rect 6593 4093 6646 4121
rect 6593 4090 6605 4093
rect 6547 4084 6605 4090
rect 6640 4081 6646 4093
rect 6698 4081 6704 4133
rect 7024 4081 7030 4133
rect 7082 4121 7088 4133
rect 8752 4121 8758 4133
rect 7082 4093 8758 4121
rect 7082 4081 7088 4093
rect 8752 4081 8758 4093
rect 8810 4081 8816 4133
rect 9730 4130 9758 4167
rect 12688 4155 12694 4167
rect 12746 4155 12752 4207
rect 9715 4124 9773 4130
rect 9715 4090 9727 4124
rect 9761 4090 9773 4124
rect 9715 4084 9773 4090
rect 10291 4124 10349 4130
rect 10291 4090 10303 4124
rect 10337 4121 10349 4124
rect 11440 4121 11446 4133
rect 10337 4093 11446 4121
rect 10337 4090 10349 4093
rect 10291 4084 10349 4090
rect 11440 4081 11446 4093
rect 11498 4081 11504 4133
rect 1152 4022 13056 4044
rect 1152 3970 4966 4022
rect 5018 3970 5030 4022
rect 5082 3970 5094 4022
rect 5146 3970 5158 4022
rect 5210 3970 5222 4022
rect 5274 3970 5286 4022
rect 5338 3970 10966 4022
rect 11018 3970 11030 4022
rect 11082 3970 11094 4022
rect 11146 3970 11158 4022
rect 11210 3970 11222 4022
rect 11274 3970 11286 4022
rect 11338 3970 13056 4022
rect 1152 3948 13056 3970
rect 6451 3902 6509 3908
rect 6451 3868 6463 3902
rect 6497 3899 6509 3902
rect 6736 3899 6742 3911
rect 6497 3871 6742 3899
rect 6497 3868 6509 3871
rect 6451 3862 6509 3868
rect 6736 3859 6742 3871
rect 6794 3859 6800 3911
rect 7120 3859 7126 3911
rect 7178 3859 7184 3911
rect 7696 3859 7702 3911
rect 7754 3899 7760 3911
rect 10291 3902 10349 3908
rect 7754 3871 9470 3899
rect 7754 3859 7760 3871
rect 6163 3828 6221 3834
rect 6163 3794 6175 3828
rect 6209 3825 6221 3828
rect 7138 3825 7166 3859
rect 6209 3797 7166 3825
rect 7234 3797 8414 3825
rect 6209 3794 6221 3797
rect 6163 3788 6221 3794
rect 4144 3711 4150 3763
rect 4202 3751 4208 3763
rect 7024 3751 7030 3763
rect 4202 3723 5726 3751
rect 4202 3711 4208 3723
rect 4240 3637 4246 3689
rect 4298 3677 4304 3689
rect 4531 3680 4589 3686
rect 4531 3677 4543 3680
rect 4298 3649 4543 3677
rect 4298 3637 4304 3649
rect 4531 3646 4543 3649
rect 4577 3646 4589 3680
rect 4531 3640 4589 3646
rect 4258 3529 4286 3637
rect 5698 3603 5726 3723
rect 6754 3723 7030 3751
rect 6256 3637 6262 3689
rect 6314 3677 6320 3689
rect 6754 3686 6782 3723
rect 7024 3711 7030 3723
rect 7082 3711 7088 3763
rect 7120 3711 7126 3763
rect 7178 3711 7184 3763
rect 7234 3760 7262 3797
rect 8386 3763 8414 3797
rect 8656 3785 8662 3837
rect 8714 3785 8720 3837
rect 9442 3825 9470 3871
rect 10291 3868 10303 3902
rect 10337 3899 10349 3902
rect 10384 3899 10390 3911
rect 10337 3871 10390 3899
rect 10337 3868 10349 3871
rect 10291 3862 10349 3868
rect 10384 3859 10390 3871
rect 10442 3859 10448 3911
rect 12499 3902 12557 3908
rect 12499 3868 12511 3902
rect 12545 3899 12557 3902
rect 12880 3899 12886 3911
rect 12545 3871 12886 3899
rect 12545 3868 12557 3871
rect 12499 3862 12557 3868
rect 12880 3859 12886 3871
rect 12938 3859 12944 3911
rect 10483 3828 10541 3834
rect 10483 3825 10495 3828
rect 9442 3797 10495 3825
rect 10483 3794 10495 3797
rect 10529 3825 10541 3828
rect 10576 3825 10582 3837
rect 10529 3797 10582 3825
rect 10529 3794 10541 3797
rect 10483 3788 10541 3794
rect 10576 3785 10582 3797
rect 10634 3785 10640 3837
rect 10690 3797 12254 3825
rect 7219 3754 7277 3760
rect 7219 3720 7231 3754
rect 7265 3720 7277 3754
rect 7795 3754 7853 3760
rect 7795 3751 7807 3754
rect 7219 3714 7277 3720
rect 7330 3723 7807 3751
rect 6739 3680 6797 3686
rect 6739 3677 6751 3680
rect 6314 3649 6751 3677
rect 6314 3637 6320 3649
rect 6739 3646 6751 3649
rect 6785 3646 6797 3680
rect 7138 3677 7166 3711
rect 7330 3677 7358 3723
rect 7795 3720 7807 3723
rect 7841 3720 7853 3754
rect 7795 3714 7853 3720
rect 8368 3711 8374 3763
rect 8426 3711 8432 3763
rect 8674 3686 8702 3785
rect 9040 3711 9046 3763
rect 9098 3751 9104 3763
rect 10690 3751 10718 3797
rect 9098 3723 10718 3751
rect 9098 3711 9104 3723
rect 10768 3711 10774 3763
rect 10826 3751 10832 3763
rect 12226 3760 12254 3797
rect 11059 3754 11117 3760
rect 11059 3751 11071 3754
rect 10826 3723 11071 3751
rect 10826 3711 10832 3723
rect 11059 3720 11071 3723
rect 11105 3720 11117 3754
rect 11059 3714 11117 3720
rect 12211 3754 12269 3760
rect 12211 3720 12223 3754
rect 12257 3720 12269 3754
rect 12211 3714 12269 3720
rect 8659 3680 8717 3686
rect 8659 3677 8671 3680
rect 7138 3649 7358 3677
rect 7522 3649 8671 3677
rect 6739 3640 6797 3646
rect 7216 3603 7222 3615
rect 5698 3589 7222 3603
rect 5712 3575 7222 3589
rect 7216 3563 7222 3575
rect 7274 3563 7280 3615
rect 7522 3603 7550 3649
rect 8659 3646 8671 3649
rect 8705 3646 8717 3680
rect 8659 3640 8717 3646
rect 10192 3637 10198 3689
rect 10250 3677 10256 3689
rect 10675 3680 10733 3686
rect 10675 3677 10687 3680
rect 10250 3649 10687 3677
rect 10250 3637 10256 3649
rect 10675 3646 10687 3649
rect 10721 3677 10733 3680
rect 11248 3677 11254 3689
rect 10721 3649 11254 3677
rect 10721 3646 10733 3649
rect 10675 3640 10733 3646
rect 11248 3637 11254 3649
rect 11306 3637 11312 3689
rect 7426 3575 7550 3603
rect 8275 3606 8333 3612
rect 7426 3529 7454 3575
rect 8275 3572 8287 3606
rect 8321 3603 8333 3606
rect 8368 3603 8374 3615
rect 8321 3575 8374 3603
rect 8321 3572 8333 3575
rect 8275 3566 8333 3572
rect 8368 3563 8374 3575
rect 8426 3563 8432 3615
rect 9616 3563 9622 3615
rect 9674 3563 9680 3615
rect 11347 3606 11405 3612
rect 11347 3572 11359 3606
rect 11393 3603 11405 3606
rect 12304 3603 12310 3615
rect 11393 3575 12310 3603
rect 11393 3572 11405 3575
rect 11347 3566 11405 3572
rect 12304 3563 12310 3575
rect 12362 3563 12368 3615
rect 10000 3529 10006 3541
rect 4258 3501 7454 3529
rect 7522 3501 10006 3529
rect 6544 3415 6550 3467
rect 6602 3455 6608 3467
rect 7120 3455 7126 3467
rect 6602 3427 7126 3455
rect 6602 3415 6608 3427
rect 7120 3415 7126 3427
rect 7178 3415 7184 3467
rect 7522 3464 7550 3501
rect 10000 3489 10006 3501
rect 10058 3489 10064 3541
rect 10192 3489 10198 3541
rect 10250 3529 10256 3541
rect 12112 3529 12118 3541
rect 10250 3501 12118 3529
rect 10250 3489 10256 3501
rect 12112 3489 12118 3501
rect 12170 3489 12176 3541
rect 7507 3458 7565 3464
rect 7507 3424 7519 3458
rect 7553 3424 7565 3458
rect 7507 3418 7565 3424
rect 8083 3458 8141 3464
rect 8083 3424 8095 3458
rect 8129 3455 8141 3458
rect 9808 3455 9814 3467
rect 8129 3427 9814 3455
rect 8129 3424 8141 3427
rect 8083 3418 8141 3424
rect 9808 3415 9814 3427
rect 9866 3415 9872 3467
rect 1152 3356 13056 3378
rect 1152 3304 1966 3356
rect 2018 3304 2030 3356
rect 2082 3304 2094 3356
rect 2146 3304 2158 3356
rect 2210 3304 2222 3356
rect 2274 3304 2286 3356
rect 2338 3304 7966 3356
rect 8018 3304 8030 3356
rect 8082 3304 8094 3356
rect 8146 3304 8158 3356
rect 8210 3304 8222 3356
rect 8274 3304 8286 3356
rect 8338 3304 13056 3356
rect 1152 3282 13056 3304
rect 4720 3193 4726 3245
rect 4778 3193 4784 3245
rect 6256 3193 6262 3245
rect 6314 3193 6320 3245
rect 6544 3193 6550 3245
rect 6602 3193 6608 3245
rect 6640 3193 6646 3245
rect 6698 3233 6704 3245
rect 8464 3233 8470 3245
rect 6698 3205 8470 3233
rect 6698 3193 6704 3205
rect 8464 3193 8470 3205
rect 8522 3193 8528 3245
rect 9235 3236 9293 3242
rect 9235 3202 9247 3236
rect 9281 3233 9293 3236
rect 9904 3233 9910 3245
rect 9281 3205 9910 3233
rect 9281 3202 9293 3205
rect 9235 3196 9293 3202
rect 9904 3193 9910 3205
rect 9962 3193 9968 3245
rect 10192 3193 10198 3245
rect 10250 3193 10256 3245
rect 10576 3193 10582 3245
rect 10634 3193 10640 3245
rect 10768 3193 10774 3245
rect 10826 3233 10832 3245
rect 11632 3233 11638 3245
rect 10826 3205 11638 3233
rect 10826 3193 10832 3205
rect 11632 3193 11638 3205
rect 11690 3193 11696 3245
rect 12496 3193 12502 3245
rect 12554 3193 12560 3245
rect 4432 3119 4438 3171
rect 4490 3159 4496 3171
rect 10210 3159 10238 3193
rect 4490 3131 10238 3159
rect 10594 3159 10622 3193
rect 10594 3131 11198 3159
rect 4490 3119 4496 3131
rect 9622 3097 9674 3103
rect 7216 3045 7222 3097
rect 7274 3045 7280 3097
rect 11170 3094 11198 3131
rect 11248 3119 11254 3171
rect 11306 3119 11312 3171
rect 11155 3088 11213 3094
rect 11155 3054 11167 3088
rect 11201 3054 11213 3088
rect 11266 3085 11294 3119
rect 11635 3088 11693 3094
rect 11635 3085 11647 3088
rect 11266 3057 11647 3085
rect 11155 3048 11213 3054
rect 11635 3054 11647 3057
rect 11681 3054 11693 3088
rect 11635 3048 11693 3054
rect 9622 3039 9674 3045
rect 4432 2971 4438 3023
rect 4490 2971 4496 3023
rect 6067 3014 6125 3020
rect 6067 2980 6079 3014
rect 6113 3011 6125 3014
rect 7120 3011 7126 3023
rect 6113 2983 7126 3011
rect 6113 2980 6125 2983
rect 6067 2974 6125 2980
rect 7120 2971 7126 2983
rect 7178 2971 7184 3023
rect 7696 2971 7702 3023
rect 7754 2971 7760 3023
rect 7888 2971 7894 3023
rect 7946 3011 7952 3023
rect 8179 3014 8237 3020
rect 8179 3011 8191 3014
rect 7946 2983 8191 3011
rect 7946 2971 7952 2983
rect 8179 2980 8191 2983
rect 8225 2980 8237 3014
rect 8179 2974 8237 2980
rect 8464 2971 8470 3023
rect 8522 3011 8528 3023
rect 10768 3011 10774 3023
rect 8522 2983 10774 3011
rect 8522 2971 8528 2983
rect 10768 2971 10774 2983
rect 10826 2971 10832 3023
rect 11827 3014 11885 3020
rect 11827 3011 11839 3014
rect 10882 2983 11839 3011
rect 2035 2940 2093 2946
rect 2035 2906 2047 2940
rect 2081 2937 2093 2940
rect 3376 2937 3382 2949
rect 2081 2909 3382 2937
rect 2081 2906 2093 2909
rect 2035 2900 2093 2906
rect 3376 2897 3382 2909
rect 3434 2897 3440 2949
rect 7714 2937 7742 2971
rect 8563 2940 8621 2946
rect 8563 2937 8575 2940
rect 7714 2909 8575 2937
rect 8563 2906 8575 2909
rect 8609 2906 8621 2940
rect 8563 2900 8621 2906
rect 9904 2897 9910 2949
rect 9962 2937 9968 2949
rect 10882 2937 10910 2983
rect 11827 2980 11839 2983
rect 11873 2980 11885 3014
rect 11827 2974 11885 2980
rect 9962 2909 10910 2937
rect 9962 2897 9968 2909
rect 12208 2897 12214 2949
rect 12266 2897 12272 2949
rect 1744 2749 1750 2801
rect 1802 2749 1808 2801
rect 1152 2690 13056 2712
rect 1152 2638 4966 2690
rect 5018 2638 5030 2690
rect 5082 2638 5094 2690
rect 5146 2638 5158 2690
rect 5210 2638 5222 2690
rect 5274 2638 5286 2690
rect 5338 2638 10966 2690
rect 11018 2638 11030 2690
rect 11082 2638 11094 2690
rect 11146 2638 11158 2690
rect 11210 2638 11222 2690
rect 11274 2638 11286 2690
rect 11338 2638 13056 2690
rect 1152 2616 13056 2638
<< via1 >>
rect 4966 14626 5018 14678
rect 5030 14626 5082 14678
rect 5094 14626 5146 14678
rect 5158 14626 5210 14678
rect 5222 14626 5274 14678
rect 5286 14626 5338 14678
rect 10966 14626 11018 14678
rect 11030 14626 11082 14678
rect 11094 14626 11146 14678
rect 11158 14626 11210 14678
rect 11222 14626 11274 14678
rect 11286 14626 11338 14678
rect 1846 14367 1898 14419
rect 3286 14410 3338 14419
rect 3286 14376 3295 14410
rect 3295 14376 3329 14410
rect 3329 14376 3338 14410
rect 3286 14367 3338 14376
rect 6166 14367 6218 14419
rect 7894 14410 7946 14419
rect 7894 14376 7903 14410
rect 7903 14376 7937 14410
rect 7937 14376 7946 14410
rect 7894 14367 7946 14376
rect 11542 14515 11594 14567
rect 9142 14410 9194 14419
rect 9142 14376 9151 14410
rect 9151 14376 9185 14410
rect 9185 14376 9194 14410
rect 9142 14367 9194 14376
rect 9334 14367 9386 14419
rect 1750 14262 1802 14271
rect 1750 14228 1759 14262
rect 1759 14228 1793 14262
rect 1793 14228 1802 14262
rect 1750 14219 1802 14228
rect 5590 14336 5642 14345
rect 5590 14302 5599 14336
rect 5599 14302 5633 14336
rect 5633 14302 5642 14336
rect 5590 14293 5642 14302
rect 5686 14293 5738 14345
rect 1942 14145 1994 14197
rect 3382 14262 3434 14271
rect 3382 14228 3391 14262
rect 3391 14228 3425 14262
rect 3425 14228 3434 14262
rect 3382 14219 3434 14228
rect 3958 14219 4010 14271
rect 4054 14219 4106 14271
rect 11062 14293 11114 14345
rect 6550 14145 6602 14197
rect 5686 14071 5738 14123
rect 7990 14262 8042 14271
rect 7990 14228 7999 14262
rect 7999 14228 8033 14262
rect 8033 14228 8042 14262
rect 7990 14219 8042 14228
rect 12310 14367 12362 14419
rect 12022 14293 12074 14345
rect 8662 14145 8714 14197
rect 8854 14145 8906 14197
rect 10006 14145 10058 14197
rect 11446 14145 11498 14197
rect 9622 14071 9674 14123
rect 1966 13960 2018 14012
rect 2030 13960 2082 14012
rect 2094 13960 2146 14012
rect 2158 13960 2210 14012
rect 2222 13960 2274 14012
rect 2286 13960 2338 14012
rect 7966 13960 8018 14012
rect 8030 13960 8082 14012
rect 8094 13960 8146 14012
rect 8158 13960 8210 14012
rect 8222 13960 8274 14012
rect 8286 13960 8338 14012
rect 3286 13849 3338 13901
rect 4246 13849 4298 13901
rect 7894 13849 7946 13901
rect 8566 13849 8618 13901
rect 11062 13892 11114 13901
rect 11062 13858 11071 13892
rect 11071 13858 11105 13892
rect 11105 13858 11114 13892
rect 11062 13849 11114 13858
rect 4054 13744 4106 13753
rect 4054 13710 4063 13744
rect 4063 13710 4097 13744
rect 4097 13710 4106 13744
rect 4054 13701 4106 13710
rect 3574 13627 3626 13679
rect 4246 13670 4298 13679
rect 4246 13636 4255 13670
rect 4255 13636 4289 13670
rect 4289 13636 4298 13670
rect 4246 13627 4298 13636
rect 3958 13553 4010 13605
rect 4438 13596 4490 13605
rect 4438 13562 4447 13596
rect 4447 13562 4481 13596
rect 4481 13562 4490 13596
rect 4438 13553 4490 13562
rect 5590 13775 5642 13827
rect 5686 13701 5738 13753
rect 5494 13670 5546 13679
rect 5494 13636 5519 13670
rect 5519 13636 5546 13670
rect 5494 13627 5546 13636
rect 9238 13701 9290 13753
rect 5782 13596 5834 13605
rect 5782 13562 5791 13596
rect 5791 13562 5825 13596
rect 5825 13562 5834 13596
rect 5782 13553 5834 13562
rect 7798 13553 7850 13605
rect 8662 13479 8714 13531
rect 8950 13553 9002 13605
rect 12406 13553 12458 13605
rect 12790 13553 12842 13605
rect 9430 13405 9482 13457
rect 9814 13405 9866 13457
rect 11830 13405 11882 13457
rect 12406 13405 12458 13457
rect 4966 13294 5018 13346
rect 5030 13294 5082 13346
rect 5094 13294 5146 13346
rect 5158 13294 5210 13346
rect 5222 13294 5274 13346
rect 5286 13294 5338 13346
rect 10966 13294 11018 13346
rect 11030 13294 11082 13346
rect 11094 13294 11146 13346
rect 11158 13294 11210 13346
rect 11222 13294 11274 13346
rect 11286 13294 11338 13346
rect 1750 13183 1802 13235
rect 4438 13183 4490 13235
rect 6166 13226 6218 13235
rect 6166 13192 6175 13226
rect 6175 13192 6209 13226
rect 6209 13192 6218 13226
rect 6166 13183 6218 13192
rect 9334 13183 9386 13235
rect 10678 13183 10730 13235
rect 8470 13109 8522 13161
rect 8662 13109 8714 13161
rect 10006 13109 10058 13161
rect 12022 13226 12074 13235
rect 12022 13192 12031 13226
rect 12031 13192 12065 13226
rect 12065 13192 12074 13226
rect 12022 13183 12074 13192
rect 12310 13183 12362 13235
rect 790 12961 842 13013
rect 3574 12961 3626 13013
rect 4438 12961 4490 13013
rect 5494 13035 5546 13087
rect 9814 13035 9866 13087
rect 10198 12961 10250 13013
rect 10678 13035 10730 13087
rect 10774 13078 10826 13087
rect 10774 13044 10783 13078
rect 10783 13044 10817 13078
rect 10817 13044 10826 13078
rect 10774 13035 10826 13044
rect 11446 13035 11498 13087
rect 12214 13078 12266 13087
rect 12214 13044 12223 13078
rect 12223 13044 12257 13078
rect 12257 13044 12266 13078
rect 12214 13035 12266 13044
rect 4054 12813 4106 12865
rect 8758 12887 8810 12939
rect 9238 12813 9290 12865
rect 12502 12782 12554 12791
rect 12502 12748 12511 12782
rect 12511 12748 12545 12782
rect 12545 12748 12554 12782
rect 12502 12739 12554 12748
rect 1966 12628 2018 12680
rect 2030 12628 2082 12680
rect 2094 12628 2146 12680
rect 2158 12628 2210 12680
rect 2222 12628 2274 12680
rect 2286 12628 2338 12680
rect 7966 12628 8018 12680
rect 8030 12628 8082 12680
rect 8094 12628 8146 12680
rect 8158 12628 8210 12680
rect 8222 12628 8274 12680
rect 8286 12628 8338 12680
rect 1846 12517 1898 12569
rect 9142 12517 9194 12569
rect 9910 12517 9962 12569
rect 4246 12369 4298 12421
rect 8758 12443 8810 12495
rect 10678 12369 10730 12421
rect 3574 12295 3626 12347
rect 7222 12295 7274 12347
rect 7798 12295 7850 12347
rect 10870 12338 10922 12347
rect 10870 12304 10879 12338
rect 10879 12304 10913 12338
rect 10913 12304 10922 12338
rect 10870 12295 10922 12304
rect 6550 12221 6602 12273
rect 8950 12221 9002 12273
rect 10486 12264 10538 12273
rect 10486 12230 10495 12264
rect 10495 12230 10529 12264
rect 10529 12230 10538 12264
rect 10486 12221 10538 12230
rect 4966 11962 5018 12014
rect 5030 11962 5082 12014
rect 5094 11962 5146 12014
rect 5158 11962 5210 12014
rect 5222 11962 5274 12014
rect 5286 11962 5338 12014
rect 10966 11962 11018 12014
rect 11030 11962 11082 12014
rect 11094 11962 11146 12014
rect 11158 11962 11210 12014
rect 11222 11962 11274 12014
rect 11286 11962 11338 12014
rect 9430 11894 9482 11903
rect 9430 11860 9439 11894
rect 9439 11860 9473 11894
rect 9473 11860 9482 11894
rect 9430 11851 9482 11860
rect 10486 11703 10538 11755
rect 2614 11672 2666 11681
rect 2614 11638 2623 11672
rect 2623 11638 2657 11672
rect 2657 11638 2666 11672
rect 2614 11629 2666 11638
rect 2806 11629 2858 11681
rect 10966 11629 11018 11681
rect 1750 11555 1802 11607
rect 4630 11555 4682 11607
rect 12502 11598 12554 11607
rect 12502 11564 12511 11598
rect 12511 11564 12545 11598
rect 12545 11564 12554 11598
rect 12502 11555 12554 11564
rect 2710 11407 2762 11459
rect 8470 11407 8522 11459
rect 10678 11481 10730 11533
rect 1966 11296 2018 11348
rect 2030 11296 2082 11348
rect 2094 11296 2146 11348
rect 2158 11296 2210 11348
rect 2222 11296 2274 11348
rect 2286 11296 2338 11348
rect 7966 11296 8018 11348
rect 8030 11296 8082 11348
rect 8094 11296 8146 11348
rect 8158 11296 8210 11348
rect 8222 11296 8274 11348
rect 8286 11296 8338 11348
rect 2614 11185 2666 11237
rect 4630 11228 4682 11237
rect 4630 11194 4639 11228
rect 4639 11194 4673 11228
rect 4673 11194 4682 11228
rect 4630 11185 4682 11194
rect 7222 11228 7274 11237
rect 7222 11194 7231 11228
rect 7231 11194 7265 11228
rect 7265 11194 7274 11228
rect 7222 11185 7274 11194
rect 12982 11185 13034 11237
rect 10966 11154 11018 11163
rect 4150 11037 4202 11089
rect 7222 11037 7274 11089
rect 2710 10963 2762 11015
rect 3382 10963 3434 11015
rect 4822 11006 4874 11015
rect 4822 10972 4831 11006
rect 4831 10972 4865 11006
rect 4865 10972 4874 11006
rect 4822 10963 4874 10972
rect 5494 10963 5546 11015
rect 10966 11120 10975 11154
rect 10975 11120 11009 11154
rect 11009 11120 11018 11154
rect 10966 11111 11018 11120
rect 8470 11037 8522 11089
rect 8662 11006 8714 11015
rect 8662 10972 8671 11006
rect 8671 10972 8705 11006
rect 8705 10972 8714 11006
rect 8662 10963 8714 10972
rect 5782 10889 5834 10941
rect 8470 10932 8522 10941
rect 8470 10898 8479 10932
rect 8479 10898 8513 10932
rect 8513 10898 8522 10932
rect 8470 10889 8522 10898
rect 3574 10741 3626 10793
rect 3862 10741 3914 10793
rect 7510 10741 7562 10793
rect 9046 10932 9098 10941
rect 9046 10898 9055 10932
rect 9055 10898 9089 10932
rect 9089 10898 9098 10932
rect 9046 10889 9098 10898
rect 10870 10889 10922 10941
rect 11734 10889 11786 10941
rect 11926 10784 11978 10793
rect 11926 10750 11935 10784
rect 11935 10750 11969 10784
rect 11969 10750 11978 10784
rect 11926 10741 11978 10750
rect 4966 10630 5018 10682
rect 5030 10630 5082 10682
rect 5094 10630 5146 10682
rect 5158 10630 5210 10682
rect 5222 10630 5274 10682
rect 5286 10630 5338 10682
rect 10966 10630 11018 10682
rect 11030 10630 11082 10682
rect 11094 10630 11146 10682
rect 11158 10630 11210 10682
rect 11222 10630 11274 10682
rect 11286 10630 11338 10682
rect 4054 10519 4106 10571
rect 4822 10519 4874 10571
rect 5782 10519 5834 10571
rect 2806 10297 2858 10349
rect 3766 10340 3818 10349
rect 3766 10306 3775 10340
rect 3775 10306 3809 10340
rect 3809 10306 3818 10340
rect 3766 10297 3818 10306
rect 3862 10340 3914 10349
rect 3862 10306 3871 10340
rect 3871 10306 3905 10340
rect 3905 10306 3914 10340
rect 3862 10297 3914 10306
rect 7126 10445 7178 10497
rect 9142 10445 9194 10497
rect 2422 10223 2474 10275
rect 5686 10149 5738 10201
rect 10102 10371 10154 10423
rect 10966 10371 11018 10423
rect 9046 10297 9098 10349
rect 7222 10223 7274 10275
rect 3382 10075 3434 10127
rect 7126 10075 7178 10127
rect 7318 10075 7370 10127
rect 9526 10223 9578 10275
rect 9142 10149 9194 10201
rect 10294 10149 10346 10201
rect 10198 10075 10250 10127
rect 10582 10075 10634 10127
rect 12502 10118 12554 10127
rect 12502 10084 12511 10118
rect 12511 10084 12545 10118
rect 12545 10084 12554 10118
rect 12502 10075 12554 10084
rect 1966 9964 2018 10016
rect 2030 9964 2082 10016
rect 2094 9964 2146 10016
rect 2158 9964 2210 10016
rect 2222 9964 2274 10016
rect 2286 9964 2338 10016
rect 7966 9964 8018 10016
rect 8030 9964 8082 10016
rect 8094 9964 8146 10016
rect 8158 9964 8210 10016
rect 8222 9964 8274 10016
rect 8286 9964 8338 10016
rect 3766 9853 3818 9905
rect 9046 9853 9098 9905
rect 11542 9853 11594 9905
rect 2806 9705 2858 9757
rect 7222 9779 7274 9831
rect 8470 9705 8522 9757
rect 8662 9705 8714 9757
rect 9526 9748 9578 9757
rect 9526 9714 9535 9748
rect 9535 9714 9569 9748
rect 9569 9714 9578 9748
rect 9526 9705 9578 9714
rect 10678 9705 10730 9757
rect 3478 9631 3530 9683
rect 3574 9631 3626 9683
rect 4534 9631 4586 9683
rect 7510 9631 7562 9683
rect 8566 9631 8618 9683
rect 4150 9557 4202 9609
rect 5782 9557 5834 9609
rect 6646 9600 6698 9609
rect 6646 9566 6655 9600
rect 6655 9566 6689 9600
rect 6689 9566 6698 9600
rect 6646 9557 6698 9566
rect 8758 9557 8810 9609
rect 10966 9631 11018 9683
rect 10486 9600 10538 9609
rect 10486 9566 10495 9600
rect 10495 9566 10529 9600
rect 10529 9566 10538 9600
rect 10486 9557 10538 9566
rect 7414 9409 7466 9461
rect 10102 9452 10154 9461
rect 10102 9418 10111 9452
rect 10111 9418 10145 9452
rect 10145 9418 10154 9452
rect 10102 9409 10154 9418
rect 4966 9298 5018 9350
rect 5030 9298 5082 9350
rect 5094 9298 5146 9350
rect 5158 9298 5210 9350
rect 5222 9298 5274 9350
rect 5286 9298 5338 9350
rect 10966 9298 11018 9350
rect 11030 9298 11082 9350
rect 11094 9298 11146 9350
rect 11158 9298 11210 9350
rect 11222 9298 11274 9350
rect 11286 9298 11338 9350
rect 4630 9187 4682 9239
rect 10870 9187 10922 9239
rect 11350 9230 11402 9239
rect 11350 9196 11359 9230
rect 11359 9196 11393 9230
rect 11393 9196 11402 9230
rect 11350 9187 11402 9196
rect 12502 9230 12554 9239
rect 12502 9196 12511 9230
rect 12511 9196 12545 9230
rect 12545 9196 12554 9230
rect 12502 9187 12554 9196
rect 2710 9113 2762 9165
rect 1846 8743 1898 8795
rect 2998 9008 3050 9017
rect 2998 8974 3007 9008
rect 3007 8974 3041 9008
rect 3041 8974 3050 9008
rect 2998 8965 3050 8974
rect 5398 9039 5450 9091
rect 5782 9039 5834 9091
rect 7414 9113 7466 9165
rect 5206 9008 5258 9017
rect 5206 8974 5215 9008
rect 5215 8974 5249 9008
rect 5249 8974 5258 9008
rect 5206 8965 5258 8974
rect 5302 9008 5354 9017
rect 5302 8974 5311 9008
rect 5311 8974 5345 9008
rect 5345 8974 5354 9008
rect 5302 8965 5354 8974
rect 3478 8891 3530 8943
rect 10102 9039 10154 9091
rect 10966 9039 11018 9091
rect 9814 8965 9866 9017
rect 3382 8817 3434 8869
rect 7126 8891 7178 8943
rect 8566 8891 8618 8943
rect 10678 8891 10730 8943
rect 5590 8817 5642 8869
rect 4342 8743 4394 8795
rect 5782 8743 5834 8795
rect 9046 8786 9098 8795
rect 9046 8752 9055 8786
rect 9055 8752 9089 8786
rect 9089 8752 9098 8786
rect 9046 8743 9098 8752
rect 1966 8632 2018 8684
rect 2030 8632 2082 8684
rect 2094 8632 2146 8684
rect 2158 8632 2210 8684
rect 2222 8632 2274 8684
rect 2286 8632 2338 8684
rect 7966 8632 8018 8684
rect 8030 8632 8082 8684
rect 8094 8632 8146 8684
rect 8158 8632 8210 8684
rect 8222 8632 8274 8684
rect 8286 8632 8338 8684
rect 1846 8521 1898 8573
rect 5398 8564 5450 8573
rect 5398 8530 5407 8564
rect 5407 8530 5441 8564
rect 5441 8530 5450 8564
rect 5398 8521 5450 8530
rect 10774 8521 10826 8573
rect 6646 8447 6698 8499
rect 1750 8342 1802 8351
rect 1750 8308 1759 8342
rect 1759 8308 1793 8342
rect 1793 8308 1802 8342
rect 1750 8299 1802 8308
rect 6742 8373 6794 8425
rect 2422 8299 2474 8351
rect 2806 8299 2858 8351
rect 7798 8299 7850 8351
rect 9814 8299 9866 8351
rect 10678 8373 10730 8425
rect 10966 8299 11018 8351
rect 2518 8268 2570 8277
rect 2518 8234 2527 8268
rect 2527 8234 2561 8268
rect 2561 8234 2570 8268
rect 2518 8225 2570 8234
rect 4246 8268 4298 8277
rect 4246 8234 4255 8268
rect 4255 8234 4289 8268
rect 4289 8234 4298 8268
rect 4246 8225 4298 8234
rect 7702 8268 7754 8277
rect 7702 8234 7711 8268
rect 7711 8234 7745 8268
rect 7745 8234 7754 8268
rect 7702 8225 7754 8234
rect 10486 8268 10538 8277
rect 10486 8234 10495 8268
rect 10495 8234 10529 8268
rect 10529 8234 10538 8268
rect 10486 8225 10538 8234
rect 5302 8151 5354 8203
rect 1654 8120 1706 8129
rect 1654 8086 1663 8120
rect 1663 8086 1697 8120
rect 1697 8086 1706 8120
rect 1654 8077 1706 8086
rect 1942 8120 1994 8129
rect 1942 8086 1951 8120
rect 1951 8086 1985 8120
rect 1985 8086 1994 8120
rect 1942 8077 1994 8086
rect 3670 8120 3722 8129
rect 3670 8086 3679 8120
rect 3679 8086 3713 8120
rect 3713 8086 3722 8120
rect 3670 8077 3722 8086
rect 4438 8077 4490 8129
rect 10678 8077 10730 8129
rect 4966 7966 5018 8018
rect 5030 7966 5082 8018
rect 5094 7966 5146 8018
rect 5158 7966 5210 8018
rect 5222 7966 5274 8018
rect 5286 7966 5338 8018
rect 10966 7966 11018 8018
rect 11030 7966 11082 8018
rect 11094 7966 11146 8018
rect 11158 7966 11210 8018
rect 11222 7966 11274 8018
rect 11286 7966 11338 8018
rect 1654 7855 1706 7907
rect 1942 7855 1994 7907
rect 2326 7855 2378 7907
rect 2518 7855 2570 7907
rect 3670 7855 3722 7907
rect 4246 7855 4298 7907
rect 12886 7855 12938 7907
rect 4822 7781 4874 7833
rect 5398 7781 5450 7833
rect 9814 7781 9866 7833
rect 4630 7676 4682 7685
rect 4630 7642 4639 7676
rect 4639 7642 4673 7676
rect 4673 7642 4682 7676
rect 4630 7633 4682 7642
rect 6742 7750 6794 7759
rect 6742 7716 6751 7750
rect 6751 7716 6785 7750
rect 6785 7716 6794 7750
rect 6742 7707 6794 7716
rect 10390 7707 10442 7759
rect 5014 7633 5066 7685
rect 5782 7676 5834 7685
rect 5782 7642 5791 7676
rect 5791 7642 5825 7676
rect 5825 7642 5834 7676
rect 5782 7633 5834 7642
rect 7126 7633 7178 7685
rect 7510 7633 7562 7685
rect 2998 7559 3050 7611
rect 3862 7602 3914 7611
rect 3862 7568 3871 7602
rect 3871 7568 3905 7602
rect 3905 7568 3914 7602
rect 3862 7559 3914 7568
rect 7894 7559 7946 7611
rect 9430 7559 9482 7611
rect 12310 7559 12362 7611
rect 1966 7300 2018 7352
rect 2030 7300 2082 7352
rect 2094 7300 2146 7352
rect 2158 7300 2210 7352
rect 2222 7300 2274 7352
rect 2286 7300 2338 7352
rect 7966 7300 8018 7352
rect 8030 7300 8082 7352
rect 8094 7300 8146 7352
rect 8158 7300 8210 7352
rect 8222 7300 8274 7352
rect 8286 7300 8338 7352
rect 4342 7115 4394 7167
rect 6646 7189 6698 7241
rect 2422 7041 2474 7093
rect 3478 6967 3530 7019
rect 6742 7041 6794 7093
rect 7798 7084 7850 7093
rect 7798 7050 7807 7084
rect 7807 7050 7841 7084
rect 7841 7050 7850 7084
rect 7798 7041 7850 7050
rect 9430 7115 9482 7167
rect 4438 6967 4490 7019
rect 3862 6936 3914 6945
rect 3862 6902 3871 6936
rect 3871 6902 3905 6936
rect 3905 6902 3914 6936
rect 3862 6893 3914 6902
rect 3958 6893 4010 6945
rect 5590 6967 5642 7019
rect 12502 7084 12554 7093
rect 12502 7050 12511 7084
rect 12511 7050 12545 7084
rect 12545 7050 12554 7084
rect 12502 7041 12554 7050
rect 5014 6893 5066 6945
rect 7126 6893 7178 6945
rect 8566 6967 8618 7019
rect 4342 6819 4394 6871
rect 10390 6893 10442 6945
rect 11638 6936 11690 6945
rect 11638 6902 11647 6936
rect 11647 6902 11681 6936
rect 11681 6902 11690 6936
rect 11638 6893 11690 6902
rect 8566 6819 8618 6871
rect 11926 6862 11978 6871
rect 11926 6828 11935 6862
rect 11935 6828 11969 6862
rect 11969 6828 11978 6862
rect 11926 6819 11978 6828
rect 4630 6788 4682 6797
rect 4630 6754 4639 6788
rect 4639 6754 4673 6788
rect 4673 6754 4682 6788
rect 4630 6745 4682 6754
rect 4822 6745 4874 6797
rect 7894 6745 7946 6797
rect 10870 6745 10922 6797
rect 4966 6634 5018 6686
rect 5030 6634 5082 6686
rect 5094 6634 5146 6686
rect 5158 6634 5210 6686
rect 5222 6634 5274 6686
rect 5286 6634 5338 6686
rect 10966 6634 11018 6686
rect 11030 6634 11082 6686
rect 11094 6634 11146 6686
rect 11158 6634 11210 6686
rect 11222 6634 11274 6686
rect 11286 6634 11338 6686
rect 3958 6566 4010 6575
rect 3958 6532 3967 6566
rect 3967 6532 4001 6566
rect 4001 6532 4010 6566
rect 3958 6523 4010 6532
rect 4342 6523 4394 6575
rect 4342 6375 4394 6427
rect 4822 6523 4874 6575
rect 9622 6523 9674 6575
rect 7702 6375 7754 6427
rect 10294 6375 10346 6427
rect 2422 6301 2474 6353
rect 7894 6301 7946 6353
rect 8566 6301 8618 6353
rect 9430 6227 9482 6279
rect 2422 6153 2474 6205
rect 8566 6153 8618 6205
rect 12502 6270 12554 6279
rect 12502 6236 12511 6270
rect 12511 6236 12545 6270
rect 12545 6236 12554 6270
rect 12502 6227 12554 6236
rect 3382 6122 3434 6131
rect 3382 6088 3391 6122
rect 3391 6088 3425 6122
rect 3425 6088 3434 6122
rect 3382 6079 3434 6088
rect 5590 6122 5642 6131
rect 5590 6088 5599 6122
rect 5599 6088 5633 6122
rect 5633 6088 5642 6122
rect 5590 6079 5642 6088
rect 10774 6079 10826 6131
rect 11350 6122 11402 6131
rect 11350 6088 11359 6122
rect 11359 6088 11393 6122
rect 11393 6088 11402 6122
rect 11350 6079 11402 6088
rect 1966 5968 2018 6020
rect 2030 5968 2082 6020
rect 2094 5968 2146 6020
rect 2158 5968 2210 6020
rect 2222 5968 2274 6020
rect 2286 5968 2338 6020
rect 7966 5968 8018 6020
rect 8030 5968 8082 6020
rect 8094 5968 8146 6020
rect 8158 5968 8210 6020
rect 8222 5968 8274 6020
rect 8286 5968 8338 6020
rect 2422 5857 2474 5909
rect 4342 5857 4394 5909
rect 4630 5709 4682 5761
rect 6742 5709 6794 5761
rect 10486 5752 10538 5761
rect 10486 5718 10495 5752
rect 10495 5718 10529 5752
rect 10529 5718 10538 5752
rect 10486 5709 10538 5718
rect 10774 5709 10826 5761
rect 12598 5709 12650 5761
rect 3382 5635 3434 5687
rect 4726 5635 4778 5687
rect 3286 5413 3338 5465
rect 4438 5487 4490 5539
rect 6646 5487 6698 5539
rect 7318 5635 7370 5687
rect 10870 5678 10922 5687
rect 10870 5644 10879 5678
rect 10879 5644 10913 5678
rect 10913 5644 10922 5678
rect 10870 5635 10922 5644
rect 9430 5561 9482 5613
rect 10006 5604 10058 5613
rect 10006 5570 10015 5604
rect 10015 5570 10049 5604
rect 10049 5570 10058 5604
rect 10006 5561 10058 5570
rect 4150 5413 4202 5465
rect 5782 5413 5834 5465
rect 9526 5456 9578 5465
rect 9526 5422 9535 5456
rect 9535 5422 9569 5456
rect 9569 5422 9578 5456
rect 9526 5413 9578 5422
rect 10294 5456 10346 5465
rect 10294 5422 10303 5456
rect 10303 5422 10337 5456
rect 10337 5422 10346 5456
rect 10294 5413 10346 5422
rect 12214 5413 12266 5465
rect 4966 5302 5018 5354
rect 5030 5302 5082 5354
rect 5094 5302 5146 5354
rect 5158 5302 5210 5354
rect 5222 5302 5274 5354
rect 5286 5302 5338 5354
rect 10966 5302 11018 5354
rect 11030 5302 11082 5354
rect 11094 5302 11146 5354
rect 11158 5302 11210 5354
rect 11222 5302 11274 5354
rect 11286 5302 11338 5354
rect 3286 5191 3338 5243
rect 4726 5191 4778 5243
rect 5302 5234 5354 5243
rect 5302 5200 5311 5234
rect 5311 5200 5345 5234
rect 5345 5200 5354 5234
rect 5302 5191 5354 5200
rect 5686 5191 5738 5243
rect 7126 5191 7178 5243
rect 8374 5191 8426 5243
rect 12502 5234 12554 5243
rect 12502 5200 12511 5234
rect 12511 5200 12545 5234
rect 12545 5200 12554 5234
rect 12502 5191 12554 5200
rect 4726 5086 4778 5095
rect 4726 5052 4735 5086
rect 4735 5052 4769 5086
rect 4769 5052 4778 5086
rect 4726 5043 4778 5052
rect 5494 5043 5546 5095
rect 5302 4969 5354 5021
rect 5590 5012 5642 5021
rect 5590 4978 5599 5012
rect 5599 4978 5633 5012
rect 5633 4978 5642 5012
rect 5590 4969 5642 4978
rect 11734 5117 11786 5169
rect 10582 5043 10634 5095
rect 7126 5012 7178 5021
rect 7126 4978 7135 5012
rect 7135 4978 7169 5012
rect 7169 4978 7178 5012
rect 7126 4969 7178 4978
rect 7222 4969 7274 5021
rect 10390 4969 10442 5021
rect 4534 4895 4586 4947
rect 6742 4938 6794 4947
rect 6742 4904 6751 4938
rect 6751 4904 6785 4938
rect 6785 4904 6794 4938
rect 6742 4895 6794 4904
rect 8662 4895 8714 4947
rect 9526 4895 9578 4947
rect 10582 4747 10634 4799
rect 1966 4636 2018 4688
rect 2030 4636 2082 4688
rect 2094 4636 2146 4688
rect 2158 4636 2210 4688
rect 2222 4636 2274 4688
rect 2286 4636 2338 4688
rect 7966 4636 8018 4688
rect 8030 4636 8082 4688
rect 8094 4636 8146 4688
rect 8158 4636 8210 4688
rect 8222 4636 8274 4688
rect 8286 4636 8338 4688
rect 8662 4525 8714 4577
rect 8566 4451 8618 4503
rect 7222 4377 7274 4429
rect 4534 4229 4586 4281
rect 4246 4081 4298 4133
rect 4438 4081 4490 4133
rect 8470 4303 8522 4355
rect 7126 4229 7178 4281
rect 7894 4229 7946 4281
rect 10486 4420 10538 4429
rect 10486 4386 10495 4420
rect 10495 4386 10529 4420
rect 10529 4386 10538 4420
rect 10486 4377 10538 4386
rect 10774 4377 10826 4429
rect 9430 4272 9482 4281
rect 9430 4238 9439 4272
rect 9439 4238 9473 4272
rect 9473 4238 9482 4272
rect 9430 4229 9482 4238
rect 6742 4155 6794 4207
rect 10390 4303 10442 4355
rect 9622 4229 9674 4281
rect 12790 4229 12842 4281
rect 6646 4081 6698 4133
rect 7030 4081 7082 4133
rect 8758 4081 8810 4133
rect 12694 4155 12746 4207
rect 11446 4081 11498 4133
rect 4966 3970 5018 4022
rect 5030 3970 5082 4022
rect 5094 3970 5146 4022
rect 5158 3970 5210 4022
rect 5222 3970 5274 4022
rect 5286 3970 5338 4022
rect 10966 3970 11018 4022
rect 11030 3970 11082 4022
rect 11094 3970 11146 4022
rect 11158 3970 11210 4022
rect 11222 3970 11274 4022
rect 11286 3970 11338 4022
rect 6742 3859 6794 3911
rect 7126 3859 7178 3911
rect 7702 3859 7754 3911
rect 4150 3754 4202 3763
rect 4150 3720 4159 3754
rect 4159 3720 4193 3754
rect 4193 3720 4202 3754
rect 4150 3711 4202 3720
rect 4246 3637 4298 3689
rect 6262 3637 6314 3689
rect 7030 3711 7082 3763
rect 7126 3711 7178 3763
rect 8662 3785 8714 3837
rect 10390 3859 10442 3911
rect 12886 3859 12938 3911
rect 10582 3785 10634 3837
rect 8374 3711 8426 3763
rect 9046 3711 9098 3763
rect 10774 3711 10826 3763
rect 7222 3563 7274 3615
rect 10198 3637 10250 3689
rect 11254 3637 11306 3689
rect 8374 3563 8426 3615
rect 9622 3563 9674 3615
rect 12310 3563 12362 3615
rect 6550 3415 6602 3467
rect 7126 3415 7178 3467
rect 10006 3489 10058 3541
rect 10198 3489 10250 3541
rect 12118 3489 12170 3541
rect 9814 3415 9866 3467
rect 1966 3304 2018 3356
rect 2030 3304 2082 3356
rect 2094 3304 2146 3356
rect 2158 3304 2210 3356
rect 2222 3304 2274 3356
rect 2286 3304 2338 3356
rect 7966 3304 8018 3356
rect 8030 3304 8082 3356
rect 8094 3304 8146 3356
rect 8158 3304 8210 3356
rect 8222 3304 8274 3356
rect 8286 3304 8338 3356
rect 4726 3236 4778 3245
rect 4726 3202 4735 3236
rect 4735 3202 4769 3236
rect 4769 3202 4778 3236
rect 4726 3193 4778 3202
rect 6262 3236 6314 3245
rect 6262 3202 6271 3236
rect 6271 3202 6305 3236
rect 6305 3202 6314 3236
rect 6262 3193 6314 3202
rect 6550 3236 6602 3245
rect 6550 3202 6559 3236
rect 6559 3202 6593 3236
rect 6593 3202 6602 3236
rect 6550 3193 6602 3202
rect 6646 3193 6698 3245
rect 8470 3193 8522 3245
rect 9910 3193 9962 3245
rect 10198 3193 10250 3245
rect 10582 3193 10634 3245
rect 10774 3193 10826 3245
rect 11638 3193 11690 3245
rect 12502 3236 12554 3245
rect 12502 3202 12511 3236
rect 12511 3202 12545 3236
rect 12545 3202 12554 3236
rect 12502 3193 12554 3202
rect 4438 3119 4490 3171
rect 7222 3045 7274 3097
rect 9622 3045 9674 3097
rect 11254 3119 11306 3171
rect 4438 3014 4490 3023
rect 4438 2980 4447 3014
rect 4447 2980 4481 3014
rect 4481 2980 4490 3014
rect 4438 2971 4490 2980
rect 7126 2971 7178 3023
rect 7702 2971 7754 3023
rect 7894 2971 7946 3023
rect 8470 2971 8522 3023
rect 10774 3014 10826 3023
rect 10774 2980 10783 3014
rect 10783 2980 10817 3014
rect 10817 2980 10826 3014
rect 10774 2971 10826 2980
rect 3382 2897 3434 2949
rect 9910 2897 9962 2949
rect 12214 2940 12266 2949
rect 12214 2906 12223 2940
rect 12223 2906 12257 2940
rect 12257 2906 12266 2940
rect 12214 2897 12266 2906
rect 1750 2792 1802 2801
rect 1750 2758 1759 2792
rect 1759 2758 1793 2792
rect 1793 2758 1802 2792
rect 1750 2749 1802 2758
rect 4966 2638 5018 2690
rect 5030 2638 5082 2690
rect 5094 2638 5146 2690
rect 5158 2638 5210 2690
rect 5222 2638 5274 2690
rect 5286 2638 5338 2690
rect 10966 2638 11018 2690
rect 11030 2638 11082 2690
rect 11094 2638 11146 2690
rect 11158 2638 11210 2690
rect 11222 2638 11274 2690
rect 11286 2638 11338 2690
<< metal2 >>
rect 788 16522 844 17322
rect 1940 16522 1996 17322
rect 3092 16664 3148 17322
rect 3092 16636 3422 16664
rect 3092 16522 3148 16636
rect 802 13019 830 16522
rect 1846 14419 1898 14425
rect 1846 14361 1898 14367
rect 1750 14271 1802 14277
rect 1750 14213 1802 14219
rect 1762 13241 1790 14213
rect 1750 13235 1802 13241
rect 1750 13177 1802 13183
rect 790 13013 842 13019
rect 790 12955 842 12961
rect 1858 12575 1886 14361
rect 1954 14203 1982 16522
rect 3286 14419 3338 14425
rect 3286 14361 3338 14367
rect 1942 14197 1994 14203
rect 1942 14139 1994 14145
rect 1964 14014 2340 14023
rect 2020 14012 2044 14014
rect 2100 14012 2124 14014
rect 2180 14012 2204 14014
rect 2260 14012 2284 14014
rect 2020 13960 2030 14012
rect 2274 13960 2284 14012
rect 2020 13958 2044 13960
rect 2100 13958 2124 13960
rect 2180 13958 2204 13960
rect 2260 13958 2284 13960
rect 1964 13949 2340 13958
rect 3298 13907 3326 14361
rect 3394 14277 3422 16636
rect 4244 16522 4300 17322
rect 5396 16664 5452 17322
rect 5396 16636 5726 16664
rect 5396 16522 5452 16636
rect 3382 14271 3434 14277
rect 3382 14213 3434 14219
rect 3958 14271 4010 14277
rect 3958 14213 4010 14219
rect 4054 14271 4106 14277
rect 4054 14213 4106 14219
rect 3286 13901 3338 13907
rect 3286 13843 3338 13849
rect 3574 13679 3626 13685
rect 3574 13621 3626 13627
rect 3586 13019 3614 13621
rect 3970 13611 3998 14213
rect 4066 13759 4094 14213
rect 4258 13907 4286 16522
rect 4964 14680 5340 14689
rect 5020 14678 5044 14680
rect 5100 14678 5124 14680
rect 5180 14678 5204 14680
rect 5260 14678 5284 14680
rect 5020 14626 5030 14678
rect 5274 14626 5284 14678
rect 5020 14624 5044 14626
rect 5100 14624 5124 14626
rect 5180 14624 5204 14626
rect 5260 14624 5284 14626
rect 4964 14615 5340 14624
rect 5698 14351 5726 16636
rect 6548 16522 6604 17322
rect 7700 16664 7756 17322
rect 7700 16636 8030 16664
rect 7700 16522 7756 16636
rect 6166 14419 6218 14425
rect 6166 14361 6218 14367
rect 5590 14345 5642 14351
rect 5590 14287 5642 14293
rect 5686 14345 5738 14351
rect 5686 14287 5738 14293
rect 4246 13901 4298 13907
rect 4246 13843 4298 13849
rect 5602 13833 5630 14287
rect 5686 14123 5738 14129
rect 5686 14065 5738 14071
rect 5590 13827 5642 13833
rect 5590 13769 5642 13775
rect 5698 13759 5726 14065
rect 4054 13753 4106 13759
rect 5686 13753 5738 13759
rect 4054 13695 4106 13701
rect 5602 13701 5686 13704
rect 5602 13695 5738 13701
rect 3958 13605 4010 13611
rect 3958 13547 4010 13553
rect 3574 13013 3626 13019
rect 3574 12955 3626 12961
rect 1964 12682 2340 12691
rect 2020 12680 2044 12682
rect 2100 12680 2124 12682
rect 2180 12680 2204 12682
rect 2260 12680 2284 12682
rect 2020 12628 2030 12680
rect 2274 12628 2284 12680
rect 2020 12626 2044 12628
rect 2100 12626 2124 12628
rect 2180 12626 2204 12628
rect 2260 12626 2284 12628
rect 1964 12617 2340 12626
rect 1846 12569 1898 12575
rect 1846 12511 1898 12517
rect 3586 12353 3614 12955
rect 4066 12871 4094 13695
rect 4246 13679 4298 13685
rect 4246 13621 4298 13627
rect 5494 13679 5546 13685
rect 5494 13621 5546 13627
rect 5602 13676 5726 13695
rect 4054 12865 4106 12871
rect 4054 12807 4106 12813
rect 3574 12347 3626 12353
rect 3574 12289 3626 12295
rect 2614 11681 2666 11687
rect 2614 11623 2666 11629
rect 2806 11681 2858 11687
rect 2806 11623 2858 11629
rect 1750 11607 1802 11613
rect 1750 11549 1802 11555
rect 1762 8357 1790 11549
rect 1964 11350 2340 11359
rect 2020 11348 2044 11350
rect 2100 11348 2124 11350
rect 2180 11348 2204 11350
rect 2260 11348 2284 11350
rect 2020 11296 2030 11348
rect 2274 11296 2284 11348
rect 2020 11294 2044 11296
rect 2100 11294 2124 11296
rect 2180 11294 2204 11296
rect 2260 11294 2284 11296
rect 1964 11285 2340 11294
rect 2626 11243 2654 11623
rect 2710 11459 2762 11465
rect 2710 11401 2762 11407
rect 2614 11237 2666 11243
rect 2614 11179 2666 11185
rect 2722 11021 2750 11401
rect 2710 11015 2762 11021
rect 2710 10957 2762 10963
rect 2422 10275 2474 10281
rect 2422 10217 2474 10223
rect 1964 10018 2340 10027
rect 2020 10016 2044 10018
rect 2100 10016 2124 10018
rect 2180 10016 2204 10018
rect 2260 10016 2284 10018
rect 2020 9964 2030 10016
rect 2274 9964 2284 10016
rect 2020 9962 2044 9964
rect 2100 9962 2124 9964
rect 2180 9962 2204 9964
rect 2260 9962 2284 9964
rect 1964 9953 2340 9962
rect 1846 8795 1898 8801
rect 1846 8737 1898 8743
rect 1858 8579 1886 8737
rect 1964 8686 2340 8695
rect 2020 8684 2044 8686
rect 2100 8684 2124 8686
rect 2180 8684 2204 8686
rect 2260 8684 2284 8686
rect 2020 8632 2030 8684
rect 2274 8632 2284 8684
rect 2020 8630 2044 8632
rect 2100 8630 2124 8632
rect 2180 8630 2204 8632
rect 2260 8630 2284 8632
rect 1964 8621 2340 8630
rect 1846 8573 1898 8579
rect 2434 8524 2462 10217
rect 2722 9171 2750 10957
rect 2818 10355 2846 11623
rect 3382 11015 3434 11021
rect 3382 10957 3434 10963
rect 2806 10349 2858 10355
rect 2806 10291 2858 10297
rect 2818 9763 2846 10291
rect 3394 10133 3422 10957
rect 3574 10793 3626 10799
rect 3574 10735 3626 10741
rect 3862 10793 3914 10799
rect 3862 10735 3914 10741
rect 3382 10127 3434 10133
rect 3382 10069 3434 10075
rect 2806 9757 2858 9763
rect 2806 9699 2858 9705
rect 2710 9165 2762 9171
rect 2710 9107 2762 9113
rect 1846 8515 1898 8521
rect 2338 8496 2462 8524
rect 1750 8351 1802 8357
rect 1750 8293 1802 8299
rect 1654 8129 1706 8135
rect 1654 8071 1706 8077
rect 1942 8129 1994 8135
rect 1942 8071 1994 8077
rect 1666 7913 1694 8071
rect 1954 7913 1982 8071
rect 2338 7913 2366 8496
rect 2818 8357 2846 9699
rect 2998 9017 3050 9023
rect 2998 8959 3050 8965
rect 2422 8351 2474 8357
rect 2422 8293 2474 8299
rect 2806 8351 2858 8357
rect 2806 8293 2858 8299
rect 1654 7907 1706 7913
rect 1654 7849 1706 7855
rect 1942 7907 1994 7913
rect 1942 7849 1994 7855
rect 2326 7907 2378 7913
rect 2326 7849 2378 7855
rect 1964 7354 2340 7363
rect 2020 7352 2044 7354
rect 2100 7352 2124 7354
rect 2180 7352 2204 7354
rect 2260 7352 2284 7354
rect 2020 7300 2030 7352
rect 2274 7300 2284 7352
rect 2020 7298 2044 7300
rect 2100 7298 2124 7300
rect 2180 7298 2204 7300
rect 2260 7298 2284 7300
rect 1964 7289 2340 7298
rect 2434 7099 2462 8293
rect 2518 8277 2570 8283
rect 2518 8219 2570 8225
rect 2530 7913 2558 8219
rect 2518 7907 2570 7913
rect 2518 7849 2570 7855
rect 3010 7617 3038 8959
rect 3394 8875 3422 10069
rect 3586 9689 3614 10735
rect 3874 10355 3902 10735
rect 4066 10577 4094 12807
rect 4258 12427 4286 13621
rect 4438 13605 4490 13611
rect 4438 13547 4490 13553
rect 4450 13241 4478 13547
rect 4964 13348 5340 13357
rect 5020 13346 5044 13348
rect 5100 13346 5124 13348
rect 5180 13346 5204 13348
rect 5260 13346 5284 13348
rect 5020 13294 5030 13346
rect 5274 13294 5284 13346
rect 5020 13292 5044 13294
rect 5100 13292 5124 13294
rect 5180 13292 5204 13294
rect 5260 13292 5284 13294
rect 4964 13283 5340 13292
rect 4438 13235 4490 13241
rect 4438 13177 4490 13183
rect 5506 13093 5534 13621
rect 5494 13087 5546 13093
rect 5494 13029 5546 13035
rect 4438 13013 4490 13019
rect 5602 12974 5630 13676
rect 5782 13605 5834 13611
rect 5782 13547 5834 13553
rect 4438 12955 4490 12961
rect 4246 12421 4298 12427
rect 4246 12363 4298 12369
rect 4150 11089 4202 11095
rect 4150 11031 4202 11037
rect 4054 10571 4106 10577
rect 4054 10513 4106 10519
rect 3766 10349 3818 10355
rect 3766 10291 3818 10297
rect 3862 10349 3914 10355
rect 3862 10291 3914 10297
rect 3778 9911 3806 10291
rect 3766 9905 3818 9911
rect 3766 9847 3818 9853
rect 3478 9683 3530 9689
rect 3478 9625 3530 9631
rect 3574 9683 3626 9689
rect 3574 9625 3626 9631
rect 3490 8949 3518 9625
rect 4162 9615 4190 11031
rect 4150 9609 4202 9615
rect 4150 9551 4202 9557
rect 3478 8943 3530 8949
rect 3478 8885 3530 8891
rect 3382 8869 3434 8875
rect 3382 8811 3434 8817
rect 2998 7611 3050 7617
rect 2998 7553 3050 7559
rect 2422 7093 2474 7099
rect 2422 7035 2474 7041
rect 2434 6359 2462 7035
rect 3490 7025 3518 8885
rect 4342 8795 4394 8801
rect 4342 8737 4394 8743
rect 4246 8277 4298 8283
rect 4246 8219 4298 8225
rect 3670 8129 3722 8135
rect 3670 8071 3722 8077
rect 3682 7913 3710 8071
rect 4258 7913 4286 8219
rect 3670 7907 3722 7913
rect 3670 7849 3722 7855
rect 4246 7907 4298 7913
rect 4246 7849 4298 7855
rect 3862 7611 3914 7617
rect 3862 7553 3914 7559
rect 3478 7019 3530 7025
rect 3478 6961 3530 6967
rect 3874 6951 3902 7553
rect 4354 7173 4382 8737
rect 4450 8135 4478 12955
rect 5410 12946 5630 12974
rect 5794 12974 5822 13547
rect 6178 13241 6206 14361
rect 6562 14203 6590 16522
rect 7894 14419 7946 14425
rect 7894 14361 7946 14367
rect 6550 14197 6602 14203
rect 6550 14139 6602 14145
rect 7906 13907 7934 14361
rect 8002 14277 8030 16636
rect 8852 16522 8908 17322
rect 10004 16522 10060 17322
rect 11156 16664 11212 17322
rect 11156 16636 11486 16664
rect 11156 16522 11212 16636
rect 8660 16382 8716 16391
rect 8578 16340 8660 16368
rect 7990 14271 8042 14277
rect 7990 14213 8042 14219
rect 7964 14014 8340 14023
rect 8020 14012 8044 14014
rect 8100 14012 8124 14014
rect 8180 14012 8204 14014
rect 8260 14012 8284 14014
rect 8020 13960 8030 14012
rect 8274 13960 8284 14012
rect 8020 13958 8044 13960
rect 8100 13958 8124 13960
rect 8180 13958 8204 13960
rect 8260 13958 8284 13960
rect 7964 13949 8340 13958
rect 8578 13907 8606 16340
rect 8660 16317 8716 16326
rect 8660 15198 8716 15207
rect 8660 15133 8716 15142
rect 8674 14203 8702 15133
rect 8866 14203 8894 16522
rect 9908 15790 9964 15799
rect 9908 15725 9964 15734
rect 9142 14419 9194 14425
rect 9142 14361 9194 14367
rect 9334 14419 9386 14425
rect 9334 14361 9386 14367
rect 8662 14197 8714 14203
rect 8662 14139 8714 14145
rect 8854 14197 8906 14203
rect 8854 14139 8906 14145
rect 7894 13901 7946 13907
rect 7894 13843 7946 13849
rect 8566 13901 8618 13907
rect 8566 13843 8618 13849
rect 7798 13605 7850 13611
rect 7798 13547 7850 13553
rect 8950 13605 9002 13611
rect 8950 13547 9002 13553
rect 6166 13235 6218 13241
rect 6166 13177 6218 13183
rect 5794 12946 5918 12974
rect 4964 12016 5340 12025
rect 5020 12014 5044 12016
rect 5100 12014 5124 12016
rect 5180 12014 5204 12016
rect 5260 12014 5284 12016
rect 5020 11962 5030 12014
rect 5274 11962 5284 12014
rect 5020 11960 5044 11962
rect 5100 11960 5124 11962
rect 5180 11960 5204 11962
rect 5260 11960 5284 11962
rect 4964 11951 5340 11960
rect 4630 11607 4682 11613
rect 4630 11549 4682 11555
rect 4642 11243 4670 11549
rect 4630 11237 4682 11243
rect 4630 11179 4682 11185
rect 4822 11015 4874 11021
rect 4822 10957 4874 10963
rect 4834 10577 4862 10957
rect 4964 10684 5340 10693
rect 5020 10682 5044 10684
rect 5100 10682 5124 10684
rect 5180 10682 5204 10684
rect 5260 10682 5284 10684
rect 5020 10630 5030 10682
rect 5274 10630 5284 10682
rect 5020 10628 5044 10630
rect 5100 10628 5124 10630
rect 5180 10628 5204 10630
rect 5260 10628 5284 10630
rect 4964 10619 5340 10628
rect 4822 10571 4874 10577
rect 4822 10513 4874 10519
rect 4534 9683 4586 9689
rect 4534 9625 4586 9631
rect 4438 8129 4490 8135
rect 4438 8071 4490 8077
rect 4342 7167 4394 7173
rect 4342 7109 4394 7115
rect 4438 7019 4490 7025
rect 4438 6961 4490 6967
rect 3862 6945 3914 6951
rect 3862 6887 3914 6893
rect 3958 6945 4010 6951
rect 3958 6887 4010 6893
rect 3970 6581 3998 6887
rect 4342 6871 4394 6877
rect 4342 6813 4394 6819
rect 4354 6581 4382 6813
rect 3958 6575 4010 6581
rect 3958 6517 4010 6523
rect 4342 6575 4394 6581
rect 4342 6517 4394 6523
rect 4342 6427 4394 6433
rect 4342 6369 4394 6375
rect 2422 6353 2474 6359
rect 2422 6295 2474 6301
rect 2422 6205 2474 6211
rect 2422 6147 2474 6153
rect 1964 6022 2340 6031
rect 2020 6020 2044 6022
rect 2100 6020 2124 6022
rect 2180 6020 2204 6022
rect 2260 6020 2284 6022
rect 2020 5968 2030 6020
rect 2274 5968 2284 6020
rect 2020 5966 2044 5968
rect 2100 5966 2124 5968
rect 2180 5966 2204 5968
rect 2260 5966 2284 5968
rect 1964 5957 2340 5966
rect 2434 5915 2462 6147
rect 3382 6131 3434 6137
rect 3382 6073 3434 6079
rect 2422 5909 2474 5915
rect 2422 5851 2474 5857
rect 3394 5693 3422 6073
rect 4354 5915 4382 6369
rect 4342 5909 4394 5915
rect 4342 5851 4394 5857
rect 3382 5687 3434 5693
rect 3382 5629 3434 5635
rect 3286 5465 3338 5471
rect 3286 5407 3338 5413
rect 3298 5249 3326 5407
rect 3286 5243 3338 5249
rect 3286 5185 3338 5191
rect 1964 4690 2340 4699
rect 2020 4688 2044 4690
rect 2100 4688 2124 4690
rect 2180 4688 2204 4690
rect 2260 4688 2284 4690
rect 2020 4636 2030 4688
rect 2274 4636 2284 4688
rect 2020 4634 2044 4636
rect 2100 4634 2124 4636
rect 2180 4634 2204 4636
rect 2260 4634 2284 4636
rect 1964 4625 2340 4634
rect 1964 3358 2340 3367
rect 2020 3356 2044 3358
rect 2100 3356 2124 3358
rect 2180 3356 2204 3358
rect 2260 3356 2284 3358
rect 2020 3304 2030 3356
rect 2274 3304 2284 3356
rect 2020 3302 2044 3304
rect 2100 3302 2124 3304
rect 2180 3302 2204 3304
rect 2260 3302 2284 3304
rect 1964 3293 2340 3302
rect 3394 2955 3422 5629
rect 4450 5545 4478 6961
rect 4438 5539 4490 5545
rect 4438 5481 4490 5487
rect 4150 5465 4202 5471
rect 4150 5407 4202 5413
rect 4162 3769 4190 5407
rect 4546 4953 4574 9625
rect 5410 9560 5438 12946
rect 5494 11015 5546 11021
rect 5494 10957 5546 10963
rect 4834 9532 5438 9560
rect 4630 9239 4682 9245
rect 4630 9181 4682 9187
rect 4642 7691 4670 9181
rect 4834 7839 4862 9532
rect 4964 9352 5340 9361
rect 5020 9350 5044 9352
rect 5100 9350 5124 9352
rect 5180 9350 5204 9352
rect 5260 9350 5284 9352
rect 5020 9298 5030 9350
rect 5274 9298 5284 9350
rect 5020 9296 5044 9298
rect 5100 9296 5124 9298
rect 5180 9296 5204 9298
rect 5260 9296 5284 9298
rect 4964 9287 5340 9296
rect 5204 9130 5260 9139
rect 5204 9065 5260 9074
rect 5398 9091 5450 9097
rect 5218 9023 5246 9065
rect 5398 9033 5450 9039
rect 5206 9017 5258 9023
rect 5206 8959 5258 8965
rect 5302 9017 5354 9023
rect 5302 8959 5354 8965
rect 5314 8228 5342 8959
rect 5410 8579 5438 9033
rect 5398 8573 5450 8579
rect 5398 8515 5450 8521
rect 5314 8209 5438 8228
rect 5302 8203 5438 8209
rect 5354 8200 5438 8203
rect 5302 8145 5354 8151
rect 4964 8020 5340 8029
rect 5020 8018 5044 8020
rect 5100 8018 5124 8020
rect 5180 8018 5204 8020
rect 5260 8018 5284 8020
rect 5020 7966 5030 8018
rect 5274 7966 5284 8018
rect 5020 7964 5044 7966
rect 5100 7964 5124 7966
rect 5180 7964 5204 7966
rect 5260 7964 5284 7966
rect 4964 7955 5340 7964
rect 5410 7839 5438 8200
rect 4822 7833 4874 7839
rect 4822 7775 4874 7781
rect 5398 7833 5450 7839
rect 5398 7775 5450 7781
rect 4630 7685 4682 7691
rect 4630 7627 4682 7633
rect 5014 7685 5066 7691
rect 5014 7627 5066 7633
rect 4642 6896 4670 7627
rect 5026 6951 5054 7627
rect 5014 6945 5066 6951
rect 4642 6868 4766 6896
rect 5014 6887 5066 6893
rect 4630 6797 4682 6803
rect 4630 6739 4682 6745
rect 4642 5767 4670 6739
rect 4630 5761 4682 5767
rect 4630 5703 4682 5709
rect 4738 5693 4766 6868
rect 4822 6797 4874 6803
rect 4822 6739 4874 6745
rect 4834 6581 4862 6739
rect 4964 6688 5340 6697
rect 5020 6686 5044 6688
rect 5100 6686 5124 6688
rect 5180 6686 5204 6688
rect 5260 6686 5284 6688
rect 5020 6634 5030 6686
rect 5274 6634 5284 6686
rect 5020 6632 5044 6634
rect 5100 6632 5124 6634
rect 5180 6632 5204 6634
rect 5260 6632 5284 6634
rect 4964 6623 5340 6632
rect 4822 6575 4874 6581
rect 4822 6517 4874 6523
rect 4726 5687 4778 5693
rect 4726 5629 4778 5635
rect 4738 5249 4766 5629
rect 4964 5356 5340 5365
rect 5020 5354 5044 5356
rect 5100 5354 5124 5356
rect 5180 5354 5204 5356
rect 5260 5354 5284 5356
rect 5020 5302 5030 5354
rect 5274 5302 5284 5354
rect 5020 5300 5044 5302
rect 5100 5300 5124 5302
rect 5180 5300 5204 5302
rect 5260 5300 5284 5302
rect 4964 5291 5340 5300
rect 4726 5243 4778 5249
rect 4726 5185 4778 5191
rect 5302 5243 5354 5249
rect 5302 5185 5354 5191
rect 4726 5095 4778 5101
rect 4726 5037 4778 5043
rect 4534 4947 4586 4953
rect 4534 4889 4586 4895
rect 4546 4287 4574 4889
rect 4534 4281 4586 4287
rect 4534 4223 4586 4229
rect 4246 4133 4298 4139
rect 4246 4075 4298 4081
rect 4438 4133 4490 4139
rect 4438 4075 4490 4081
rect 4150 3763 4202 3769
rect 4150 3705 4202 3711
rect 4258 3695 4286 4075
rect 4246 3689 4298 3695
rect 4246 3631 4298 3637
rect 4450 3177 4478 4075
rect 4738 3251 4766 5037
rect 5314 5027 5342 5185
rect 5506 5101 5534 10957
rect 5782 10941 5834 10947
rect 5782 10883 5834 10889
rect 5794 10577 5822 10883
rect 5782 10571 5834 10577
rect 5782 10513 5834 10519
rect 5686 10201 5738 10207
rect 5686 10143 5738 10149
rect 5590 8869 5642 8875
rect 5590 8811 5642 8817
rect 5602 7025 5630 8811
rect 5590 7019 5642 7025
rect 5590 6961 5642 6967
rect 5590 6131 5642 6137
rect 5590 6073 5642 6079
rect 5494 5095 5546 5101
rect 5494 5037 5546 5043
rect 5602 5027 5630 6073
rect 5698 5249 5726 10143
rect 5782 9609 5834 9615
rect 5782 9551 5834 9557
rect 5794 9097 5822 9551
rect 5782 9091 5834 9097
rect 5782 9033 5834 9039
rect 5782 8795 5834 8801
rect 5782 8737 5834 8743
rect 5794 7691 5822 8737
rect 5782 7685 5834 7691
rect 5782 7627 5834 7633
rect 5890 7488 5918 12946
rect 7810 12353 7838 13547
rect 8662 13531 8714 13537
rect 8662 13473 8714 13479
rect 8674 13167 8702 13473
rect 8470 13161 8522 13167
rect 8470 13103 8522 13109
rect 8662 13161 8714 13167
rect 8662 13103 8714 13109
rect 8482 12974 8510 13103
rect 8386 12946 8510 12974
rect 7964 12682 8340 12691
rect 8020 12680 8044 12682
rect 8100 12680 8124 12682
rect 8180 12680 8204 12682
rect 8260 12680 8284 12682
rect 8020 12628 8030 12680
rect 8274 12628 8284 12680
rect 8020 12626 8044 12628
rect 8100 12626 8124 12628
rect 8180 12626 8204 12628
rect 8260 12626 8284 12628
rect 7964 12617 8340 12626
rect 7222 12347 7274 12353
rect 7222 12289 7274 12295
rect 7798 12347 7850 12353
rect 7798 12289 7850 12295
rect 6550 12273 6602 12279
rect 6550 12215 6602 12221
rect 5794 7460 5918 7488
rect 5794 5471 5822 7460
rect 5782 5465 5834 5471
rect 5782 5407 5834 5413
rect 5686 5243 5738 5249
rect 5686 5185 5738 5191
rect 5302 5021 5354 5027
rect 5302 4963 5354 4969
rect 5590 5021 5642 5027
rect 5590 4963 5642 4969
rect 4964 4024 5340 4033
rect 5020 4022 5044 4024
rect 5100 4022 5124 4024
rect 5180 4022 5204 4024
rect 5260 4022 5284 4024
rect 5020 3970 5030 4022
rect 5274 3970 5284 4022
rect 5020 3968 5044 3970
rect 5100 3968 5124 3970
rect 5180 3968 5204 3970
rect 5260 3968 5284 3970
rect 4964 3959 5340 3968
rect 6262 3689 6314 3695
rect 6262 3631 6314 3637
rect 6274 3251 6302 3631
rect 6562 3473 6590 12215
rect 7234 11243 7262 12289
rect 7964 11350 8340 11359
rect 8020 11348 8044 11350
rect 8100 11348 8124 11350
rect 8180 11348 8204 11350
rect 8260 11348 8284 11350
rect 8020 11296 8030 11348
rect 8274 11296 8284 11348
rect 8020 11294 8044 11296
rect 8100 11294 8124 11296
rect 8180 11294 8204 11296
rect 8260 11294 8284 11296
rect 7964 11285 8340 11294
rect 7222 11237 7274 11243
rect 7222 11179 7274 11185
rect 7222 11089 7274 11095
rect 7222 11031 7274 11037
rect 7126 10497 7178 10503
rect 7126 10439 7178 10445
rect 7138 10133 7166 10439
rect 7234 10281 7262 11031
rect 7510 10793 7562 10799
rect 7510 10735 7562 10741
rect 7222 10275 7274 10281
rect 7222 10217 7274 10223
rect 7126 10127 7178 10133
rect 7126 10069 7178 10075
rect 7234 9837 7262 10217
rect 7318 10127 7370 10133
rect 7318 10069 7370 10075
rect 7222 9831 7274 9837
rect 7222 9773 7274 9779
rect 6646 9609 6698 9615
rect 6646 9551 6698 9557
rect 6658 8505 6686 9551
rect 7126 8943 7178 8949
rect 7126 8885 7178 8891
rect 7138 8820 7166 8885
rect 7330 8820 7358 10069
rect 7522 9689 7550 10735
rect 7964 10018 8340 10027
rect 8020 10016 8044 10018
rect 8100 10016 8124 10018
rect 8180 10016 8204 10018
rect 8260 10016 8284 10018
rect 8020 9964 8030 10016
rect 8274 9964 8284 10016
rect 8020 9962 8044 9964
rect 8100 9962 8124 9964
rect 8180 9962 8204 9964
rect 8260 9962 8284 9964
rect 7964 9953 8340 9962
rect 7510 9683 7562 9689
rect 7510 9625 7562 9631
rect 7414 9461 7466 9467
rect 7414 9403 7466 9409
rect 7426 9171 7454 9403
rect 7414 9165 7466 9171
rect 7414 9107 7466 9113
rect 7138 8792 7358 8820
rect 6646 8499 6698 8505
rect 6646 8441 6698 8447
rect 6658 7247 6686 8441
rect 6742 8425 6794 8431
rect 6742 8367 6794 8373
rect 6754 7765 6782 8367
rect 6742 7759 6794 7765
rect 6742 7701 6794 7707
rect 6646 7241 6698 7247
rect 6646 7183 6698 7189
rect 6658 5545 6686 7183
rect 6754 7099 6782 7701
rect 7126 7685 7178 7691
rect 7126 7627 7178 7633
rect 6742 7093 6794 7099
rect 6742 7035 6794 7041
rect 6754 5767 6782 7035
rect 7138 6951 7166 7627
rect 7126 6945 7178 6951
rect 7126 6887 7178 6893
rect 6742 5761 6794 5767
rect 6742 5703 6794 5709
rect 6646 5539 6698 5545
rect 6646 5481 6698 5487
rect 7138 5249 7166 6887
rect 7330 5693 7358 8792
rect 7522 7691 7550 9625
rect 7964 8686 8340 8695
rect 8020 8684 8044 8686
rect 8100 8684 8124 8686
rect 8180 8684 8204 8686
rect 8260 8684 8284 8686
rect 8020 8632 8030 8684
rect 8274 8632 8284 8684
rect 8020 8630 8044 8632
rect 8100 8630 8124 8632
rect 8180 8630 8204 8632
rect 8260 8630 8284 8632
rect 7964 8621 8340 8630
rect 7798 8351 7850 8357
rect 7798 8293 7850 8299
rect 7702 8277 7754 8283
rect 7702 8219 7754 8225
rect 7510 7685 7562 7691
rect 7510 7627 7562 7633
rect 7714 6433 7742 8219
rect 7810 7099 7838 8293
rect 7894 7611 7946 7617
rect 7894 7553 7946 7559
rect 7798 7093 7850 7099
rect 7798 7035 7850 7041
rect 7906 6803 7934 7553
rect 7964 7354 8340 7363
rect 8020 7352 8044 7354
rect 8100 7352 8124 7354
rect 8180 7352 8204 7354
rect 8260 7352 8284 7354
rect 8020 7300 8030 7352
rect 8274 7300 8284 7352
rect 8020 7298 8044 7300
rect 8100 7298 8124 7300
rect 8180 7298 8204 7300
rect 8260 7298 8284 7300
rect 7964 7289 8340 7298
rect 7894 6797 7946 6803
rect 7894 6739 7946 6745
rect 7702 6427 7754 6433
rect 7702 6369 7754 6375
rect 7318 5687 7370 5693
rect 7318 5629 7370 5635
rect 7126 5243 7178 5249
rect 7126 5185 7178 5191
rect 7126 5021 7178 5027
rect 7126 4963 7178 4969
rect 7222 5021 7274 5027
rect 7222 4963 7274 4969
rect 6742 4947 6794 4953
rect 6742 4889 6794 4895
rect 6754 4213 6782 4889
rect 7138 4287 7166 4963
rect 7234 4435 7262 4963
rect 7222 4429 7274 4435
rect 7222 4371 7274 4377
rect 7126 4281 7178 4287
rect 7126 4223 7178 4229
rect 6742 4207 6794 4213
rect 6742 4149 6794 4155
rect 6646 4133 6698 4139
rect 6646 4075 6698 4081
rect 6550 3467 6602 3473
rect 6550 3409 6602 3415
rect 6562 3251 6590 3409
rect 6658 3251 6686 4075
rect 6754 3917 6782 4149
rect 7030 4133 7082 4139
rect 7030 4075 7082 4081
rect 6742 3911 6794 3917
rect 6742 3853 6794 3859
rect 7042 3769 7070 4075
rect 7138 3917 7166 4223
rect 7126 3911 7178 3917
rect 7126 3853 7178 3859
rect 7030 3763 7082 3769
rect 7030 3705 7082 3711
rect 7126 3763 7178 3769
rect 7126 3705 7178 3711
rect 7138 3473 7166 3705
rect 7234 3621 7262 4371
rect 7714 3917 7742 6369
rect 7906 6359 7934 6739
rect 7894 6353 7946 6359
rect 7894 6295 7946 6301
rect 7964 6022 8340 6031
rect 8020 6020 8044 6022
rect 8100 6020 8124 6022
rect 8180 6020 8204 6022
rect 8260 6020 8284 6022
rect 8020 5968 8030 6020
rect 8274 5968 8284 6020
rect 8020 5966 8044 5968
rect 8100 5966 8124 5968
rect 8180 5966 8204 5968
rect 8260 5966 8284 5968
rect 7964 5957 8340 5966
rect 8386 5249 8414 12946
rect 8758 12939 8810 12945
rect 8758 12881 8810 12887
rect 8770 12501 8798 12881
rect 8758 12495 8810 12501
rect 8758 12437 8810 12443
rect 8962 12372 8990 13547
rect 9154 12575 9182 14361
rect 9238 13753 9290 13759
rect 9238 13695 9290 13701
rect 9250 12871 9278 13695
rect 9346 13241 9374 14361
rect 9622 14123 9674 14129
rect 9622 14065 9674 14071
rect 9430 13457 9482 13463
rect 9430 13399 9482 13405
rect 9334 13235 9386 13241
rect 9334 13177 9386 13183
rect 9238 12865 9290 12871
rect 9238 12807 9290 12813
rect 9142 12569 9194 12575
rect 9142 12511 9194 12517
rect 8962 12344 9182 12372
rect 8950 12273 9002 12279
rect 8950 12215 9002 12221
rect 8470 11459 8522 11465
rect 8470 11401 8522 11407
rect 8482 11095 8510 11401
rect 8470 11089 8522 11095
rect 8470 11031 8522 11037
rect 8482 10947 8510 11031
rect 8662 11015 8714 11021
rect 8662 10957 8714 10963
rect 8470 10941 8522 10947
rect 8470 10883 8522 10889
rect 8482 9763 8510 10883
rect 8674 9763 8702 10957
rect 8470 9757 8522 9763
rect 8470 9699 8522 9705
rect 8662 9757 8714 9763
rect 8962 9745 8990 12215
rect 9046 10941 9098 10947
rect 9046 10883 9098 10889
rect 9058 10355 9086 10883
rect 9154 10503 9182 12344
rect 9442 11909 9470 13399
rect 9430 11903 9482 11909
rect 9430 11845 9482 11851
rect 9142 10497 9194 10503
rect 9142 10439 9194 10445
rect 9046 10349 9098 10355
rect 9046 10291 9098 10297
rect 9058 9911 9086 10291
rect 9154 10207 9182 10439
rect 9526 10275 9578 10281
rect 9526 10217 9578 10223
rect 9142 10201 9194 10207
rect 9142 10143 9194 10149
rect 9046 9905 9098 9911
rect 9046 9847 9098 9853
rect 9538 9763 9566 10217
rect 9526 9757 9578 9763
rect 8962 9717 9086 9745
rect 8662 9699 8714 9705
rect 8566 9683 8618 9689
rect 8566 9625 8618 9631
rect 8578 8949 8606 9625
rect 8758 9609 8810 9615
rect 8758 9551 8810 9557
rect 8566 8943 8618 8949
rect 8566 8885 8618 8891
rect 8482 7025 8606 7044
rect 8482 7019 8618 7025
rect 8482 7016 8566 7019
rect 8374 5243 8426 5249
rect 8374 5185 8426 5191
rect 7964 4690 8340 4699
rect 8020 4688 8044 4690
rect 8100 4688 8124 4690
rect 8180 4688 8204 4690
rect 8260 4688 8284 4690
rect 8020 4636 8030 4688
rect 8274 4636 8284 4688
rect 8020 4634 8044 4636
rect 8100 4634 8124 4636
rect 8180 4634 8204 4636
rect 8260 4634 8284 4636
rect 7964 4625 8340 4634
rect 7894 4281 7946 4287
rect 7894 4223 7946 4229
rect 7702 3911 7754 3917
rect 7702 3853 7754 3859
rect 7222 3615 7274 3621
rect 7222 3557 7274 3563
rect 7126 3467 7178 3473
rect 7126 3409 7178 3415
rect 4726 3245 4778 3251
rect 4726 3187 4778 3193
rect 6262 3245 6314 3251
rect 6262 3187 6314 3193
rect 6550 3245 6602 3251
rect 6550 3187 6602 3193
rect 6646 3245 6698 3251
rect 6646 3187 6698 3193
rect 4438 3171 4490 3177
rect 4438 3113 4490 3119
rect 7234 3103 7262 3557
rect 7222 3097 7274 3103
rect 7222 3039 7274 3045
rect 7714 3029 7742 3853
rect 7906 3029 7934 4223
rect 8386 3769 8414 5185
rect 8482 4380 8510 7016
rect 8566 6961 8618 6967
rect 8566 6871 8618 6877
rect 8566 6813 8618 6819
rect 8578 6359 8606 6813
rect 8566 6353 8618 6359
rect 8566 6295 8618 6301
rect 8566 6205 8618 6211
rect 8566 6147 8618 6153
rect 8578 4509 8606 6147
rect 8662 4947 8714 4953
rect 8662 4889 8714 4895
rect 8674 4583 8702 4889
rect 8662 4577 8714 4583
rect 8662 4519 8714 4525
rect 8566 4503 8618 4509
rect 8566 4445 8618 4451
rect 8482 4361 8702 4380
rect 8470 4355 8702 4361
rect 8522 4352 8702 4355
rect 8470 4297 8522 4303
rect 8674 3843 8702 4352
rect 8770 4139 8798 9551
rect 9058 8801 9086 9717
rect 9526 9699 9578 9705
rect 9046 8795 9098 8801
rect 9046 8737 9098 8743
rect 8758 4133 8810 4139
rect 8758 4075 8810 4081
rect 8662 3837 8714 3843
rect 8662 3779 8714 3785
rect 9058 3769 9086 8737
rect 9430 7611 9482 7617
rect 9430 7553 9482 7559
rect 9442 7173 9470 7553
rect 9430 7167 9482 7173
rect 9430 7109 9482 7115
rect 9442 6285 9470 7109
rect 9634 6581 9662 14065
rect 9814 13457 9866 13463
rect 9814 13399 9866 13405
rect 9826 13093 9854 13399
rect 9814 13087 9866 13093
rect 9814 13029 9866 13035
rect 9922 12575 9950 15725
rect 10018 14203 10046 16522
rect 10964 14680 11340 14689
rect 11020 14678 11044 14680
rect 11100 14678 11124 14680
rect 11180 14678 11204 14680
rect 11260 14678 11284 14680
rect 11020 14626 11030 14678
rect 11274 14626 11284 14678
rect 11020 14624 11044 14626
rect 11100 14624 11124 14626
rect 11180 14624 11204 14626
rect 11260 14624 11284 14626
rect 10964 14615 11340 14624
rect 10676 14458 10732 14467
rect 10676 14393 10732 14402
rect 10006 14197 10058 14203
rect 10006 14139 10058 14145
rect 10690 13241 10718 14393
rect 11062 14345 11114 14351
rect 11062 14287 11114 14293
rect 11074 13907 11102 14287
rect 11458 14203 11486 16636
rect 12308 16522 12364 17322
rect 13460 16664 13516 17322
rect 13186 16636 13516 16664
rect 11542 14567 11594 14573
rect 11542 14509 11594 14515
rect 11446 14197 11498 14203
rect 11446 14139 11498 14145
rect 11062 13901 11114 13907
rect 11062 13843 11114 13849
rect 10964 13348 11340 13357
rect 11020 13346 11044 13348
rect 11100 13346 11124 13348
rect 11180 13346 11204 13348
rect 11260 13346 11284 13348
rect 11020 13294 11030 13346
rect 11274 13294 11284 13346
rect 11020 13292 11044 13294
rect 11100 13292 11124 13294
rect 11180 13292 11204 13294
rect 11260 13292 11284 13294
rect 10964 13283 11340 13292
rect 10678 13235 10730 13241
rect 10678 13177 10730 13183
rect 10006 13161 10058 13167
rect 10006 13103 10058 13109
rect 9910 12569 9962 12575
rect 9910 12511 9962 12517
rect 9814 9017 9866 9023
rect 9814 8959 9866 8965
rect 9826 8357 9854 8959
rect 9814 8351 9866 8357
rect 9814 8293 9866 8299
rect 9826 7839 9854 8293
rect 9814 7833 9866 7839
rect 9814 7775 9866 7781
rect 9622 6575 9674 6581
rect 9622 6517 9674 6523
rect 9430 6279 9482 6285
rect 9430 6221 9482 6227
rect 9442 5619 9470 6221
rect 9430 5613 9482 5619
rect 9430 5555 9482 5561
rect 9442 4287 9470 5555
rect 9526 5465 9578 5471
rect 9526 5407 9578 5413
rect 9538 4953 9566 5407
rect 9526 4947 9578 4953
rect 9526 4889 9578 4895
rect 9430 4281 9482 4287
rect 9430 4223 9482 4229
rect 9538 4084 9566 4889
rect 9634 4287 9662 6517
rect 10018 5619 10046 13103
rect 10678 13087 10730 13093
rect 10678 13029 10730 13035
rect 10774 13087 10826 13093
rect 10774 13029 10826 13035
rect 11446 13087 11498 13093
rect 11446 13029 11498 13035
rect 10198 13013 10250 13019
rect 10198 12955 10250 12961
rect 10102 10423 10154 10429
rect 10102 10365 10154 10371
rect 10114 9560 10142 10365
rect 10210 10133 10238 12955
rect 10690 12427 10718 13029
rect 10678 12421 10730 12427
rect 10678 12363 10730 12369
rect 10486 12273 10538 12279
rect 10486 12215 10538 12221
rect 10498 11761 10526 12215
rect 10486 11755 10538 11761
rect 10486 11697 10538 11703
rect 10294 10201 10346 10207
rect 10294 10143 10346 10149
rect 10198 10127 10250 10133
rect 10198 10069 10250 10075
rect 10114 9532 10238 9560
rect 10102 9461 10154 9467
rect 10102 9403 10154 9409
rect 10114 9097 10142 9403
rect 10102 9091 10154 9097
rect 10102 9033 10154 9039
rect 10006 5613 10058 5619
rect 10006 5555 10058 5561
rect 9622 4281 9674 4287
rect 9622 4223 9674 4229
rect 9538 4056 9662 4084
rect 8374 3763 8426 3769
rect 8374 3705 8426 3711
rect 9046 3763 9098 3769
rect 9046 3705 9098 3711
rect 9634 3621 9662 4056
rect 10018 3640 10046 5555
rect 10210 3695 10238 9532
rect 10306 6433 10334 10143
rect 10498 9615 10526 11697
rect 10690 11539 10718 12363
rect 10678 11533 10730 11539
rect 10678 11475 10730 11481
rect 10582 10127 10634 10133
rect 10582 10069 10634 10075
rect 10486 9609 10538 9615
rect 10486 9551 10538 9557
rect 10486 8277 10538 8283
rect 10486 8219 10538 8225
rect 10390 7759 10442 7765
rect 10390 7701 10442 7707
rect 10402 6951 10430 7701
rect 10390 6945 10442 6951
rect 10390 6887 10442 6893
rect 10294 6427 10346 6433
rect 10294 6369 10346 6375
rect 10294 5465 10346 5471
rect 10294 5407 10346 5413
rect 8374 3615 8426 3621
rect 8374 3557 8426 3563
rect 9622 3615 9674 3621
rect 9622 3557 9674 3563
rect 9922 3612 10046 3640
rect 10198 3689 10250 3695
rect 10198 3631 10250 3637
rect 8386 3492 8414 3557
rect 8386 3464 8510 3492
rect 7964 3358 8340 3367
rect 8020 3356 8044 3358
rect 8100 3356 8124 3358
rect 8180 3356 8204 3358
rect 8260 3356 8284 3358
rect 8020 3304 8030 3356
rect 8274 3304 8284 3356
rect 8020 3302 8044 3304
rect 8100 3302 8124 3304
rect 8180 3302 8204 3304
rect 8260 3302 8284 3304
rect 7964 3293 8340 3302
rect 8482 3251 8510 3464
rect 8470 3245 8522 3251
rect 8470 3187 8522 3193
rect 8482 3029 8510 3187
rect 9634 3103 9662 3557
rect 9814 3467 9866 3473
rect 9814 3409 9866 3415
rect 9622 3097 9674 3103
rect 9622 3039 9674 3045
rect 4438 3023 4490 3029
rect 4438 2965 4490 2971
rect 7126 3023 7178 3029
rect 7126 2965 7178 2971
rect 7702 3023 7754 3029
rect 7702 2965 7754 2971
rect 7894 3023 7946 3029
rect 7894 2965 7946 2971
rect 8470 3023 8522 3029
rect 8470 2965 8522 2971
rect 3382 2949 3434 2955
rect 3382 2891 3434 2897
rect 1750 2801 1802 2807
rect 1750 2743 1802 2749
rect 1556 680 1612 800
rect 1762 680 1790 2743
rect 1556 652 1790 680
rect 4340 680 4396 800
rect 4450 680 4478 2965
rect 4964 2692 5340 2701
rect 5020 2690 5044 2692
rect 5100 2690 5124 2692
rect 5180 2690 5204 2692
rect 5260 2690 5284 2692
rect 5020 2638 5030 2690
rect 5274 2638 5284 2690
rect 5020 2636 5044 2638
rect 5100 2636 5124 2638
rect 5180 2636 5204 2638
rect 5260 2636 5284 2638
rect 4964 2627 5340 2636
rect 7138 800 7166 2965
rect 9826 999 9854 3409
rect 9922 3251 9950 3612
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10198 3541 10250 3547
rect 10198 3483 10250 3489
rect 9910 3245 9962 3251
rect 9910 3187 9962 3193
rect 9910 2949 9962 2955
rect 9910 2891 9962 2897
rect 9812 990 9868 999
rect 9812 925 9868 934
rect 9922 800 9950 2891
rect 10018 2183 10046 3483
rect 10210 3251 10238 3483
rect 10198 3245 10250 3251
rect 10198 3187 10250 3193
rect 10004 2174 10060 2183
rect 10004 2109 10060 2118
rect 10306 1591 10334 5407
rect 10402 5027 10430 6887
rect 10498 5767 10526 8219
rect 10486 5761 10538 5767
rect 10486 5703 10538 5709
rect 10390 5021 10442 5027
rect 10390 4963 10442 4969
rect 10402 4361 10430 4963
rect 10498 4435 10526 5703
rect 10594 5101 10622 10069
rect 10678 9757 10730 9763
rect 10678 9699 10730 9705
rect 10690 8949 10718 9699
rect 10678 8943 10730 8949
rect 10678 8885 10730 8891
rect 10690 8431 10718 8885
rect 10786 8579 10814 13029
rect 10870 12347 10922 12353
rect 10870 12289 10922 12295
rect 10882 10947 10910 12289
rect 10964 12016 11340 12025
rect 11020 12014 11044 12016
rect 11100 12014 11124 12016
rect 11180 12014 11204 12016
rect 11260 12014 11284 12016
rect 11020 11962 11030 12014
rect 11274 11962 11284 12014
rect 11020 11960 11044 11962
rect 11100 11960 11124 11962
rect 11180 11960 11204 11962
rect 11260 11960 11284 11962
rect 10964 11951 11340 11960
rect 10966 11681 11018 11687
rect 10966 11623 11018 11629
rect 10978 11169 11006 11623
rect 10966 11163 11018 11169
rect 10966 11105 11018 11111
rect 10870 10941 10922 10947
rect 10870 10883 10922 10889
rect 10964 10684 11340 10693
rect 11020 10682 11044 10684
rect 11100 10682 11124 10684
rect 11180 10682 11204 10684
rect 11260 10682 11284 10684
rect 11020 10630 11030 10682
rect 11274 10630 11284 10682
rect 11020 10628 11044 10630
rect 11100 10628 11124 10630
rect 11180 10628 11204 10630
rect 11260 10628 11284 10630
rect 10964 10619 11340 10628
rect 10966 10423 11018 10429
rect 10966 10365 11018 10371
rect 10978 9689 11006 10365
rect 10966 9683 11018 9689
rect 10966 9625 11018 9631
rect 10978 9560 11006 9625
rect 10882 9532 11006 9560
rect 10882 9245 10910 9532
rect 10964 9352 11340 9361
rect 11020 9350 11044 9352
rect 11100 9350 11124 9352
rect 11180 9350 11204 9352
rect 11260 9350 11284 9352
rect 11020 9298 11030 9350
rect 11274 9298 11284 9350
rect 11020 9296 11044 9298
rect 11100 9296 11124 9298
rect 11180 9296 11204 9298
rect 11260 9296 11284 9298
rect 10964 9287 11340 9296
rect 11458 9264 11486 13029
rect 11554 9911 11582 14509
rect 12322 14425 12350 16522
rect 12310 14419 12362 14425
rect 12310 14361 12362 14367
rect 12022 14345 12074 14351
rect 12022 14287 12074 14293
rect 11830 13457 11882 13463
rect 11828 13422 11830 13431
rect 11882 13422 11884 13431
rect 11828 13357 11884 13366
rect 12034 13241 12062 14287
rect 12308 14014 12364 14023
rect 12308 13949 12364 13958
rect 12322 13241 12350 13949
rect 12406 13605 12458 13611
rect 12790 13605 12842 13611
rect 12458 13553 12638 13556
rect 12406 13547 12638 13553
rect 12790 13547 12842 13553
rect 12418 13528 12638 13547
rect 12406 13457 12458 13463
rect 12406 13399 12458 13405
rect 12022 13235 12074 13241
rect 12022 13177 12074 13183
rect 12310 13235 12362 13241
rect 12310 13177 12362 13183
rect 12214 13087 12266 13093
rect 12214 13029 12266 13035
rect 12226 12974 12254 13029
rect 12130 12946 12254 12974
rect 11734 10941 11786 10947
rect 11734 10883 11786 10889
rect 11542 9905 11594 9911
rect 11542 9847 11594 9853
rect 11362 9245 11486 9264
rect 10870 9239 10922 9245
rect 10870 9181 10922 9187
rect 11350 9239 11486 9245
rect 11402 9236 11486 9239
rect 11350 9181 11402 9187
rect 10966 9091 11018 9097
rect 10966 9033 11018 9039
rect 10774 8573 10826 8579
rect 10774 8515 10826 8521
rect 10678 8425 10730 8431
rect 10678 8367 10730 8373
rect 10978 8357 11006 9033
rect 10966 8351 11018 8357
rect 10966 8293 11018 8299
rect 10678 8129 10730 8135
rect 10678 8071 10730 8077
rect 10582 5095 10634 5101
rect 10582 5037 10634 5043
rect 10582 4799 10634 4805
rect 10582 4741 10634 4747
rect 10486 4429 10538 4435
rect 10486 4371 10538 4377
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10402 3917 10430 4297
rect 10390 3911 10442 3917
rect 10390 3853 10442 3859
rect 10594 3843 10622 4741
rect 10690 4232 10718 8071
rect 10964 8020 11340 8029
rect 11020 8018 11044 8020
rect 11100 8018 11124 8020
rect 11180 8018 11204 8020
rect 11260 8018 11284 8020
rect 11020 7966 11030 8018
rect 11274 7966 11284 8018
rect 11020 7964 11044 7966
rect 11100 7964 11124 7966
rect 11180 7964 11204 7966
rect 11260 7964 11284 7966
rect 10964 7955 11340 7964
rect 11638 6945 11690 6951
rect 11638 6887 11690 6893
rect 10870 6797 10922 6803
rect 10870 6739 10922 6745
rect 10774 6131 10826 6137
rect 10774 6073 10826 6079
rect 10786 5767 10814 6073
rect 10774 5761 10826 5767
rect 10774 5703 10826 5709
rect 10786 4435 10814 5703
rect 10882 5693 10910 6739
rect 10964 6688 11340 6697
rect 11020 6686 11044 6688
rect 11100 6686 11124 6688
rect 11180 6686 11204 6688
rect 11260 6686 11284 6688
rect 11020 6634 11030 6686
rect 11274 6634 11284 6686
rect 11020 6632 11044 6634
rect 11100 6632 11124 6634
rect 11180 6632 11204 6634
rect 11260 6632 11284 6634
rect 10964 6623 11340 6632
rect 11350 6131 11402 6137
rect 11350 6073 11402 6079
rect 11362 5735 11390 6073
rect 11348 5726 11404 5735
rect 10870 5687 10922 5693
rect 11348 5661 11404 5670
rect 10870 5629 10922 5635
rect 10964 5356 11340 5365
rect 11020 5354 11044 5356
rect 11100 5354 11124 5356
rect 11180 5354 11204 5356
rect 11260 5354 11284 5356
rect 11020 5302 11030 5354
rect 11274 5302 11284 5354
rect 11020 5300 11044 5302
rect 11100 5300 11124 5302
rect 11180 5300 11204 5302
rect 11260 5300 11284 5302
rect 10964 5291 11340 5300
rect 10774 4429 10826 4435
rect 10774 4371 10826 4377
rect 10690 4204 10814 4232
rect 10582 3837 10634 3843
rect 10582 3779 10634 3785
rect 10594 3251 10622 3779
rect 10786 3769 10814 4204
rect 11446 4133 11498 4139
rect 11446 4075 11498 4081
rect 10964 4024 11340 4033
rect 11020 4022 11044 4024
rect 11100 4022 11124 4024
rect 11180 4022 11204 4024
rect 11260 4022 11284 4024
rect 11020 3970 11030 4022
rect 11274 3970 11284 4022
rect 11020 3968 11044 3970
rect 11100 3968 11124 3970
rect 11180 3968 11204 3970
rect 11260 3968 11284 3970
rect 10964 3959 11340 3968
rect 10774 3763 10826 3769
rect 10774 3705 10826 3711
rect 11254 3689 11306 3695
rect 11254 3631 11306 3637
rect 10582 3245 10634 3251
rect 10582 3187 10634 3193
rect 10774 3245 10826 3251
rect 10774 3187 10826 3193
rect 10786 3029 10814 3187
rect 11266 3177 11294 3631
rect 11254 3171 11306 3177
rect 11254 3113 11306 3119
rect 10774 3023 10826 3029
rect 10774 2965 10826 2971
rect 11458 2775 11486 4075
rect 11650 3251 11678 6887
rect 11746 5175 11774 10883
rect 11926 10793 11978 10799
rect 11926 10735 11978 10741
rect 11938 10471 11966 10735
rect 11924 10462 11980 10471
rect 11924 10397 11980 10406
rect 11924 6910 11980 6919
rect 11924 6845 11926 6854
rect 11978 6845 11980 6854
rect 11926 6813 11978 6819
rect 11734 5169 11786 5175
rect 11734 5111 11786 5117
rect 12130 3547 12158 12946
rect 12418 12839 12446 13399
rect 12404 12830 12460 12839
rect 12404 12765 12460 12774
rect 12502 12791 12554 12797
rect 12502 12733 12554 12739
rect 12514 12247 12542 12733
rect 12500 12238 12556 12247
rect 12500 12173 12556 12182
rect 12502 11607 12554 11613
rect 12502 11549 12554 11555
rect 12514 11063 12542 11549
rect 12500 11054 12556 11063
rect 12500 10989 12556 10998
rect 12502 10127 12554 10133
rect 12502 10069 12554 10075
rect 12514 9879 12542 10069
rect 12500 9870 12556 9879
rect 12500 9805 12556 9814
rect 12500 9278 12556 9287
rect 12500 9213 12502 9222
rect 12554 9213 12556 9222
rect 12502 9181 12554 9187
rect 12500 8094 12556 8103
rect 12500 8029 12556 8038
rect 12310 7611 12362 7617
rect 12310 7553 12362 7559
rect 12322 7511 12350 7553
rect 12308 7502 12364 7511
rect 12308 7437 12364 7446
rect 12514 7099 12542 8029
rect 12502 7093 12554 7099
rect 12502 7035 12554 7041
rect 12500 6318 12556 6327
rect 12500 6253 12502 6262
rect 12554 6253 12556 6262
rect 12502 6221 12554 6227
rect 12610 5767 12638 13528
rect 12598 5761 12650 5767
rect 12598 5703 12650 5709
rect 12214 5465 12266 5471
rect 12214 5407 12266 5413
rect 12118 3541 12170 3547
rect 12118 3483 12170 3489
rect 11638 3245 11690 3251
rect 11638 3187 11690 3193
rect 12226 2955 12254 5407
rect 12502 5243 12554 5249
rect 12502 5185 12554 5191
rect 12514 5143 12542 5185
rect 12500 5134 12556 5143
rect 12500 5069 12556 5078
rect 12802 4287 12830 13547
rect 12980 11646 13036 11655
rect 12980 11581 13036 11590
rect 12994 11243 13022 11581
rect 12982 11237 13034 11243
rect 12982 11179 13034 11185
rect 13186 9139 13214 16636
rect 13460 16522 13516 16636
rect 13172 9130 13228 9139
rect 13172 9065 13228 9074
rect 12884 8686 12940 8695
rect 12884 8621 12940 8630
rect 12898 7913 12926 8621
rect 12886 7907 12938 7913
rect 12886 7849 12938 7855
rect 12884 4542 12940 4551
rect 12884 4477 12940 4486
rect 12790 4281 12842 4287
rect 12790 4223 12842 4229
rect 12694 4207 12746 4213
rect 12694 4149 12746 4155
rect 12500 3950 12556 3959
rect 12500 3885 12556 3894
rect 12310 3615 12362 3621
rect 12310 3557 12362 3563
rect 12322 3367 12350 3557
rect 12308 3358 12364 3367
rect 12308 3293 12364 3302
rect 12514 3251 12542 3885
rect 12502 3245 12554 3251
rect 12502 3187 12554 3193
rect 12214 2949 12266 2955
rect 12214 2891 12266 2897
rect 11444 2766 11500 2775
rect 11444 2701 11500 2710
rect 10964 2692 11340 2701
rect 11020 2690 11044 2692
rect 11100 2690 11124 2692
rect 11180 2690 11204 2692
rect 11260 2690 11284 2692
rect 11020 2638 11030 2690
rect 11274 2638 11284 2690
rect 11020 2636 11044 2638
rect 11100 2636 11124 2638
rect 11180 2636 11204 2638
rect 11260 2636 11284 2638
rect 10964 2627 11340 2636
rect 10292 1582 10348 1591
rect 10292 1517 10348 1526
rect 12706 800 12734 4149
rect 12898 3917 12926 4477
rect 12886 3911 12938 3917
rect 12886 3853 12938 3859
rect 4340 652 4478 680
rect 1556 0 1612 652
rect 4340 0 4396 652
rect 7124 0 7180 800
rect 9908 0 9964 800
rect 12692 0 12748 800
<< via2 >>
rect 1964 14012 2020 14014
rect 2044 14012 2100 14014
rect 2124 14012 2180 14014
rect 2204 14012 2260 14014
rect 2284 14012 2340 14014
rect 1964 13960 1966 14012
rect 1966 13960 2018 14012
rect 2018 13960 2020 14012
rect 2044 13960 2082 14012
rect 2082 13960 2094 14012
rect 2094 13960 2100 14012
rect 2124 13960 2146 14012
rect 2146 13960 2158 14012
rect 2158 13960 2180 14012
rect 2204 13960 2210 14012
rect 2210 13960 2222 14012
rect 2222 13960 2260 14012
rect 2284 13960 2286 14012
rect 2286 13960 2338 14012
rect 2338 13960 2340 14012
rect 1964 13958 2020 13960
rect 2044 13958 2100 13960
rect 2124 13958 2180 13960
rect 2204 13958 2260 13960
rect 2284 13958 2340 13960
rect 4964 14678 5020 14680
rect 5044 14678 5100 14680
rect 5124 14678 5180 14680
rect 5204 14678 5260 14680
rect 5284 14678 5340 14680
rect 4964 14626 4966 14678
rect 4966 14626 5018 14678
rect 5018 14626 5020 14678
rect 5044 14626 5082 14678
rect 5082 14626 5094 14678
rect 5094 14626 5100 14678
rect 5124 14626 5146 14678
rect 5146 14626 5158 14678
rect 5158 14626 5180 14678
rect 5204 14626 5210 14678
rect 5210 14626 5222 14678
rect 5222 14626 5260 14678
rect 5284 14626 5286 14678
rect 5286 14626 5338 14678
rect 5338 14626 5340 14678
rect 4964 14624 5020 14626
rect 5044 14624 5100 14626
rect 5124 14624 5180 14626
rect 5204 14624 5260 14626
rect 5284 14624 5340 14626
rect 1964 12680 2020 12682
rect 2044 12680 2100 12682
rect 2124 12680 2180 12682
rect 2204 12680 2260 12682
rect 2284 12680 2340 12682
rect 1964 12628 1966 12680
rect 1966 12628 2018 12680
rect 2018 12628 2020 12680
rect 2044 12628 2082 12680
rect 2082 12628 2094 12680
rect 2094 12628 2100 12680
rect 2124 12628 2146 12680
rect 2146 12628 2158 12680
rect 2158 12628 2180 12680
rect 2204 12628 2210 12680
rect 2210 12628 2222 12680
rect 2222 12628 2260 12680
rect 2284 12628 2286 12680
rect 2286 12628 2338 12680
rect 2338 12628 2340 12680
rect 1964 12626 2020 12628
rect 2044 12626 2100 12628
rect 2124 12626 2180 12628
rect 2204 12626 2260 12628
rect 2284 12626 2340 12628
rect 1964 11348 2020 11350
rect 2044 11348 2100 11350
rect 2124 11348 2180 11350
rect 2204 11348 2260 11350
rect 2284 11348 2340 11350
rect 1964 11296 1966 11348
rect 1966 11296 2018 11348
rect 2018 11296 2020 11348
rect 2044 11296 2082 11348
rect 2082 11296 2094 11348
rect 2094 11296 2100 11348
rect 2124 11296 2146 11348
rect 2146 11296 2158 11348
rect 2158 11296 2180 11348
rect 2204 11296 2210 11348
rect 2210 11296 2222 11348
rect 2222 11296 2260 11348
rect 2284 11296 2286 11348
rect 2286 11296 2338 11348
rect 2338 11296 2340 11348
rect 1964 11294 2020 11296
rect 2044 11294 2100 11296
rect 2124 11294 2180 11296
rect 2204 11294 2260 11296
rect 2284 11294 2340 11296
rect 1964 10016 2020 10018
rect 2044 10016 2100 10018
rect 2124 10016 2180 10018
rect 2204 10016 2260 10018
rect 2284 10016 2340 10018
rect 1964 9964 1966 10016
rect 1966 9964 2018 10016
rect 2018 9964 2020 10016
rect 2044 9964 2082 10016
rect 2082 9964 2094 10016
rect 2094 9964 2100 10016
rect 2124 9964 2146 10016
rect 2146 9964 2158 10016
rect 2158 9964 2180 10016
rect 2204 9964 2210 10016
rect 2210 9964 2222 10016
rect 2222 9964 2260 10016
rect 2284 9964 2286 10016
rect 2286 9964 2338 10016
rect 2338 9964 2340 10016
rect 1964 9962 2020 9964
rect 2044 9962 2100 9964
rect 2124 9962 2180 9964
rect 2204 9962 2260 9964
rect 2284 9962 2340 9964
rect 1964 8684 2020 8686
rect 2044 8684 2100 8686
rect 2124 8684 2180 8686
rect 2204 8684 2260 8686
rect 2284 8684 2340 8686
rect 1964 8632 1966 8684
rect 1966 8632 2018 8684
rect 2018 8632 2020 8684
rect 2044 8632 2082 8684
rect 2082 8632 2094 8684
rect 2094 8632 2100 8684
rect 2124 8632 2146 8684
rect 2146 8632 2158 8684
rect 2158 8632 2180 8684
rect 2204 8632 2210 8684
rect 2210 8632 2222 8684
rect 2222 8632 2260 8684
rect 2284 8632 2286 8684
rect 2286 8632 2338 8684
rect 2338 8632 2340 8684
rect 1964 8630 2020 8632
rect 2044 8630 2100 8632
rect 2124 8630 2180 8632
rect 2204 8630 2260 8632
rect 2284 8630 2340 8632
rect 1964 7352 2020 7354
rect 2044 7352 2100 7354
rect 2124 7352 2180 7354
rect 2204 7352 2260 7354
rect 2284 7352 2340 7354
rect 1964 7300 1966 7352
rect 1966 7300 2018 7352
rect 2018 7300 2020 7352
rect 2044 7300 2082 7352
rect 2082 7300 2094 7352
rect 2094 7300 2100 7352
rect 2124 7300 2146 7352
rect 2146 7300 2158 7352
rect 2158 7300 2180 7352
rect 2204 7300 2210 7352
rect 2210 7300 2222 7352
rect 2222 7300 2260 7352
rect 2284 7300 2286 7352
rect 2286 7300 2338 7352
rect 2338 7300 2340 7352
rect 1964 7298 2020 7300
rect 2044 7298 2100 7300
rect 2124 7298 2180 7300
rect 2204 7298 2260 7300
rect 2284 7298 2340 7300
rect 4964 13346 5020 13348
rect 5044 13346 5100 13348
rect 5124 13346 5180 13348
rect 5204 13346 5260 13348
rect 5284 13346 5340 13348
rect 4964 13294 4966 13346
rect 4966 13294 5018 13346
rect 5018 13294 5020 13346
rect 5044 13294 5082 13346
rect 5082 13294 5094 13346
rect 5094 13294 5100 13346
rect 5124 13294 5146 13346
rect 5146 13294 5158 13346
rect 5158 13294 5180 13346
rect 5204 13294 5210 13346
rect 5210 13294 5222 13346
rect 5222 13294 5260 13346
rect 5284 13294 5286 13346
rect 5286 13294 5338 13346
rect 5338 13294 5340 13346
rect 4964 13292 5020 13294
rect 5044 13292 5100 13294
rect 5124 13292 5180 13294
rect 5204 13292 5260 13294
rect 5284 13292 5340 13294
rect 7964 14012 8020 14014
rect 8044 14012 8100 14014
rect 8124 14012 8180 14014
rect 8204 14012 8260 14014
rect 8284 14012 8340 14014
rect 7964 13960 7966 14012
rect 7966 13960 8018 14012
rect 8018 13960 8020 14012
rect 8044 13960 8082 14012
rect 8082 13960 8094 14012
rect 8094 13960 8100 14012
rect 8124 13960 8146 14012
rect 8146 13960 8158 14012
rect 8158 13960 8180 14012
rect 8204 13960 8210 14012
rect 8210 13960 8222 14012
rect 8222 13960 8260 14012
rect 8284 13960 8286 14012
rect 8286 13960 8338 14012
rect 8338 13960 8340 14012
rect 7964 13958 8020 13960
rect 8044 13958 8100 13960
rect 8124 13958 8180 13960
rect 8204 13958 8260 13960
rect 8284 13958 8340 13960
rect 8660 16326 8716 16382
rect 8660 15142 8716 15198
rect 9908 15734 9964 15790
rect 4964 12014 5020 12016
rect 5044 12014 5100 12016
rect 5124 12014 5180 12016
rect 5204 12014 5260 12016
rect 5284 12014 5340 12016
rect 4964 11962 4966 12014
rect 4966 11962 5018 12014
rect 5018 11962 5020 12014
rect 5044 11962 5082 12014
rect 5082 11962 5094 12014
rect 5094 11962 5100 12014
rect 5124 11962 5146 12014
rect 5146 11962 5158 12014
rect 5158 11962 5180 12014
rect 5204 11962 5210 12014
rect 5210 11962 5222 12014
rect 5222 11962 5260 12014
rect 5284 11962 5286 12014
rect 5286 11962 5338 12014
rect 5338 11962 5340 12014
rect 4964 11960 5020 11962
rect 5044 11960 5100 11962
rect 5124 11960 5180 11962
rect 5204 11960 5260 11962
rect 5284 11960 5340 11962
rect 4964 10682 5020 10684
rect 5044 10682 5100 10684
rect 5124 10682 5180 10684
rect 5204 10682 5260 10684
rect 5284 10682 5340 10684
rect 4964 10630 4966 10682
rect 4966 10630 5018 10682
rect 5018 10630 5020 10682
rect 5044 10630 5082 10682
rect 5082 10630 5094 10682
rect 5094 10630 5100 10682
rect 5124 10630 5146 10682
rect 5146 10630 5158 10682
rect 5158 10630 5180 10682
rect 5204 10630 5210 10682
rect 5210 10630 5222 10682
rect 5222 10630 5260 10682
rect 5284 10630 5286 10682
rect 5286 10630 5338 10682
rect 5338 10630 5340 10682
rect 4964 10628 5020 10630
rect 5044 10628 5100 10630
rect 5124 10628 5180 10630
rect 5204 10628 5260 10630
rect 5284 10628 5340 10630
rect 1964 6020 2020 6022
rect 2044 6020 2100 6022
rect 2124 6020 2180 6022
rect 2204 6020 2260 6022
rect 2284 6020 2340 6022
rect 1964 5968 1966 6020
rect 1966 5968 2018 6020
rect 2018 5968 2020 6020
rect 2044 5968 2082 6020
rect 2082 5968 2094 6020
rect 2094 5968 2100 6020
rect 2124 5968 2146 6020
rect 2146 5968 2158 6020
rect 2158 5968 2180 6020
rect 2204 5968 2210 6020
rect 2210 5968 2222 6020
rect 2222 5968 2260 6020
rect 2284 5968 2286 6020
rect 2286 5968 2338 6020
rect 2338 5968 2340 6020
rect 1964 5966 2020 5968
rect 2044 5966 2100 5968
rect 2124 5966 2180 5968
rect 2204 5966 2260 5968
rect 2284 5966 2340 5968
rect 1964 4688 2020 4690
rect 2044 4688 2100 4690
rect 2124 4688 2180 4690
rect 2204 4688 2260 4690
rect 2284 4688 2340 4690
rect 1964 4636 1966 4688
rect 1966 4636 2018 4688
rect 2018 4636 2020 4688
rect 2044 4636 2082 4688
rect 2082 4636 2094 4688
rect 2094 4636 2100 4688
rect 2124 4636 2146 4688
rect 2146 4636 2158 4688
rect 2158 4636 2180 4688
rect 2204 4636 2210 4688
rect 2210 4636 2222 4688
rect 2222 4636 2260 4688
rect 2284 4636 2286 4688
rect 2286 4636 2338 4688
rect 2338 4636 2340 4688
rect 1964 4634 2020 4636
rect 2044 4634 2100 4636
rect 2124 4634 2180 4636
rect 2204 4634 2260 4636
rect 2284 4634 2340 4636
rect 1964 3356 2020 3358
rect 2044 3356 2100 3358
rect 2124 3356 2180 3358
rect 2204 3356 2260 3358
rect 2284 3356 2340 3358
rect 1964 3304 1966 3356
rect 1966 3304 2018 3356
rect 2018 3304 2020 3356
rect 2044 3304 2082 3356
rect 2082 3304 2094 3356
rect 2094 3304 2100 3356
rect 2124 3304 2146 3356
rect 2146 3304 2158 3356
rect 2158 3304 2180 3356
rect 2204 3304 2210 3356
rect 2210 3304 2222 3356
rect 2222 3304 2260 3356
rect 2284 3304 2286 3356
rect 2286 3304 2338 3356
rect 2338 3304 2340 3356
rect 1964 3302 2020 3304
rect 2044 3302 2100 3304
rect 2124 3302 2180 3304
rect 2204 3302 2260 3304
rect 2284 3302 2340 3304
rect 4964 9350 5020 9352
rect 5044 9350 5100 9352
rect 5124 9350 5180 9352
rect 5204 9350 5260 9352
rect 5284 9350 5340 9352
rect 4964 9298 4966 9350
rect 4966 9298 5018 9350
rect 5018 9298 5020 9350
rect 5044 9298 5082 9350
rect 5082 9298 5094 9350
rect 5094 9298 5100 9350
rect 5124 9298 5146 9350
rect 5146 9298 5158 9350
rect 5158 9298 5180 9350
rect 5204 9298 5210 9350
rect 5210 9298 5222 9350
rect 5222 9298 5260 9350
rect 5284 9298 5286 9350
rect 5286 9298 5338 9350
rect 5338 9298 5340 9350
rect 4964 9296 5020 9298
rect 5044 9296 5100 9298
rect 5124 9296 5180 9298
rect 5204 9296 5260 9298
rect 5284 9296 5340 9298
rect 5204 9074 5260 9130
rect 4964 8018 5020 8020
rect 5044 8018 5100 8020
rect 5124 8018 5180 8020
rect 5204 8018 5260 8020
rect 5284 8018 5340 8020
rect 4964 7966 4966 8018
rect 4966 7966 5018 8018
rect 5018 7966 5020 8018
rect 5044 7966 5082 8018
rect 5082 7966 5094 8018
rect 5094 7966 5100 8018
rect 5124 7966 5146 8018
rect 5146 7966 5158 8018
rect 5158 7966 5180 8018
rect 5204 7966 5210 8018
rect 5210 7966 5222 8018
rect 5222 7966 5260 8018
rect 5284 7966 5286 8018
rect 5286 7966 5338 8018
rect 5338 7966 5340 8018
rect 4964 7964 5020 7966
rect 5044 7964 5100 7966
rect 5124 7964 5180 7966
rect 5204 7964 5260 7966
rect 5284 7964 5340 7966
rect 4964 6686 5020 6688
rect 5044 6686 5100 6688
rect 5124 6686 5180 6688
rect 5204 6686 5260 6688
rect 5284 6686 5340 6688
rect 4964 6634 4966 6686
rect 4966 6634 5018 6686
rect 5018 6634 5020 6686
rect 5044 6634 5082 6686
rect 5082 6634 5094 6686
rect 5094 6634 5100 6686
rect 5124 6634 5146 6686
rect 5146 6634 5158 6686
rect 5158 6634 5180 6686
rect 5204 6634 5210 6686
rect 5210 6634 5222 6686
rect 5222 6634 5260 6686
rect 5284 6634 5286 6686
rect 5286 6634 5338 6686
rect 5338 6634 5340 6686
rect 4964 6632 5020 6634
rect 5044 6632 5100 6634
rect 5124 6632 5180 6634
rect 5204 6632 5260 6634
rect 5284 6632 5340 6634
rect 4964 5354 5020 5356
rect 5044 5354 5100 5356
rect 5124 5354 5180 5356
rect 5204 5354 5260 5356
rect 5284 5354 5340 5356
rect 4964 5302 4966 5354
rect 4966 5302 5018 5354
rect 5018 5302 5020 5354
rect 5044 5302 5082 5354
rect 5082 5302 5094 5354
rect 5094 5302 5100 5354
rect 5124 5302 5146 5354
rect 5146 5302 5158 5354
rect 5158 5302 5180 5354
rect 5204 5302 5210 5354
rect 5210 5302 5222 5354
rect 5222 5302 5260 5354
rect 5284 5302 5286 5354
rect 5286 5302 5338 5354
rect 5338 5302 5340 5354
rect 4964 5300 5020 5302
rect 5044 5300 5100 5302
rect 5124 5300 5180 5302
rect 5204 5300 5260 5302
rect 5284 5300 5340 5302
rect 7964 12680 8020 12682
rect 8044 12680 8100 12682
rect 8124 12680 8180 12682
rect 8204 12680 8260 12682
rect 8284 12680 8340 12682
rect 7964 12628 7966 12680
rect 7966 12628 8018 12680
rect 8018 12628 8020 12680
rect 8044 12628 8082 12680
rect 8082 12628 8094 12680
rect 8094 12628 8100 12680
rect 8124 12628 8146 12680
rect 8146 12628 8158 12680
rect 8158 12628 8180 12680
rect 8204 12628 8210 12680
rect 8210 12628 8222 12680
rect 8222 12628 8260 12680
rect 8284 12628 8286 12680
rect 8286 12628 8338 12680
rect 8338 12628 8340 12680
rect 7964 12626 8020 12628
rect 8044 12626 8100 12628
rect 8124 12626 8180 12628
rect 8204 12626 8260 12628
rect 8284 12626 8340 12628
rect 4964 4022 5020 4024
rect 5044 4022 5100 4024
rect 5124 4022 5180 4024
rect 5204 4022 5260 4024
rect 5284 4022 5340 4024
rect 4964 3970 4966 4022
rect 4966 3970 5018 4022
rect 5018 3970 5020 4022
rect 5044 3970 5082 4022
rect 5082 3970 5094 4022
rect 5094 3970 5100 4022
rect 5124 3970 5146 4022
rect 5146 3970 5158 4022
rect 5158 3970 5180 4022
rect 5204 3970 5210 4022
rect 5210 3970 5222 4022
rect 5222 3970 5260 4022
rect 5284 3970 5286 4022
rect 5286 3970 5338 4022
rect 5338 3970 5340 4022
rect 4964 3968 5020 3970
rect 5044 3968 5100 3970
rect 5124 3968 5180 3970
rect 5204 3968 5260 3970
rect 5284 3968 5340 3970
rect 7964 11348 8020 11350
rect 8044 11348 8100 11350
rect 8124 11348 8180 11350
rect 8204 11348 8260 11350
rect 8284 11348 8340 11350
rect 7964 11296 7966 11348
rect 7966 11296 8018 11348
rect 8018 11296 8020 11348
rect 8044 11296 8082 11348
rect 8082 11296 8094 11348
rect 8094 11296 8100 11348
rect 8124 11296 8146 11348
rect 8146 11296 8158 11348
rect 8158 11296 8180 11348
rect 8204 11296 8210 11348
rect 8210 11296 8222 11348
rect 8222 11296 8260 11348
rect 8284 11296 8286 11348
rect 8286 11296 8338 11348
rect 8338 11296 8340 11348
rect 7964 11294 8020 11296
rect 8044 11294 8100 11296
rect 8124 11294 8180 11296
rect 8204 11294 8260 11296
rect 8284 11294 8340 11296
rect 7964 10016 8020 10018
rect 8044 10016 8100 10018
rect 8124 10016 8180 10018
rect 8204 10016 8260 10018
rect 8284 10016 8340 10018
rect 7964 9964 7966 10016
rect 7966 9964 8018 10016
rect 8018 9964 8020 10016
rect 8044 9964 8082 10016
rect 8082 9964 8094 10016
rect 8094 9964 8100 10016
rect 8124 9964 8146 10016
rect 8146 9964 8158 10016
rect 8158 9964 8180 10016
rect 8204 9964 8210 10016
rect 8210 9964 8222 10016
rect 8222 9964 8260 10016
rect 8284 9964 8286 10016
rect 8286 9964 8338 10016
rect 8338 9964 8340 10016
rect 7964 9962 8020 9964
rect 8044 9962 8100 9964
rect 8124 9962 8180 9964
rect 8204 9962 8260 9964
rect 8284 9962 8340 9964
rect 7964 8684 8020 8686
rect 8044 8684 8100 8686
rect 8124 8684 8180 8686
rect 8204 8684 8260 8686
rect 8284 8684 8340 8686
rect 7964 8632 7966 8684
rect 7966 8632 8018 8684
rect 8018 8632 8020 8684
rect 8044 8632 8082 8684
rect 8082 8632 8094 8684
rect 8094 8632 8100 8684
rect 8124 8632 8146 8684
rect 8146 8632 8158 8684
rect 8158 8632 8180 8684
rect 8204 8632 8210 8684
rect 8210 8632 8222 8684
rect 8222 8632 8260 8684
rect 8284 8632 8286 8684
rect 8286 8632 8338 8684
rect 8338 8632 8340 8684
rect 7964 8630 8020 8632
rect 8044 8630 8100 8632
rect 8124 8630 8180 8632
rect 8204 8630 8260 8632
rect 8284 8630 8340 8632
rect 7964 7352 8020 7354
rect 8044 7352 8100 7354
rect 8124 7352 8180 7354
rect 8204 7352 8260 7354
rect 8284 7352 8340 7354
rect 7964 7300 7966 7352
rect 7966 7300 8018 7352
rect 8018 7300 8020 7352
rect 8044 7300 8082 7352
rect 8082 7300 8094 7352
rect 8094 7300 8100 7352
rect 8124 7300 8146 7352
rect 8146 7300 8158 7352
rect 8158 7300 8180 7352
rect 8204 7300 8210 7352
rect 8210 7300 8222 7352
rect 8222 7300 8260 7352
rect 8284 7300 8286 7352
rect 8286 7300 8338 7352
rect 8338 7300 8340 7352
rect 7964 7298 8020 7300
rect 8044 7298 8100 7300
rect 8124 7298 8180 7300
rect 8204 7298 8260 7300
rect 8284 7298 8340 7300
rect 7964 6020 8020 6022
rect 8044 6020 8100 6022
rect 8124 6020 8180 6022
rect 8204 6020 8260 6022
rect 8284 6020 8340 6022
rect 7964 5968 7966 6020
rect 7966 5968 8018 6020
rect 8018 5968 8020 6020
rect 8044 5968 8082 6020
rect 8082 5968 8094 6020
rect 8094 5968 8100 6020
rect 8124 5968 8146 6020
rect 8146 5968 8158 6020
rect 8158 5968 8180 6020
rect 8204 5968 8210 6020
rect 8210 5968 8222 6020
rect 8222 5968 8260 6020
rect 8284 5968 8286 6020
rect 8286 5968 8338 6020
rect 8338 5968 8340 6020
rect 7964 5966 8020 5968
rect 8044 5966 8100 5968
rect 8124 5966 8180 5968
rect 8204 5966 8260 5968
rect 8284 5966 8340 5968
rect 7964 4688 8020 4690
rect 8044 4688 8100 4690
rect 8124 4688 8180 4690
rect 8204 4688 8260 4690
rect 8284 4688 8340 4690
rect 7964 4636 7966 4688
rect 7966 4636 8018 4688
rect 8018 4636 8020 4688
rect 8044 4636 8082 4688
rect 8082 4636 8094 4688
rect 8094 4636 8100 4688
rect 8124 4636 8146 4688
rect 8146 4636 8158 4688
rect 8158 4636 8180 4688
rect 8204 4636 8210 4688
rect 8210 4636 8222 4688
rect 8222 4636 8260 4688
rect 8284 4636 8286 4688
rect 8286 4636 8338 4688
rect 8338 4636 8340 4688
rect 7964 4634 8020 4636
rect 8044 4634 8100 4636
rect 8124 4634 8180 4636
rect 8204 4634 8260 4636
rect 8284 4634 8340 4636
rect 10964 14678 11020 14680
rect 11044 14678 11100 14680
rect 11124 14678 11180 14680
rect 11204 14678 11260 14680
rect 11284 14678 11340 14680
rect 10964 14626 10966 14678
rect 10966 14626 11018 14678
rect 11018 14626 11020 14678
rect 11044 14626 11082 14678
rect 11082 14626 11094 14678
rect 11094 14626 11100 14678
rect 11124 14626 11146 14678
rect 11146 14626 11158 14678
rect 11158 14626 11180 14678
rect 11204 14626 11210 14678
rect 11210 14626 11222 14678
rect 11222 14626 11260 14678
rect 11284 14626 11286 14678
rect 11286 14626 11338 14678
rect 11338 14626 11340 14678
rect 10964 14624 11020 14626
rect 11044 14624 11100 14626
rect 11124 14624 11180 14626
rect 11204 14624 11260 14626
rect 11284 14624 11340 14626
rect 10676 14402 10732 14458
rect 10964 13346 11020 13348
rect 11044 13346 11100 13348
rect 11124 13346 11180 13348
rect 11204 13346 11260 13348
rect 11284 13346 11340 13348
rect 10964 13294 10966 13346
rect 10966 13294 11018 13346
rect 11018 13294 11020 13346
rect 11044 13294 11082 13346
rect 11082 13294 11094 13346
rect 11094 13294 11100 13346
rect 11124 13294 11146 13346
rect 11146 13294 11158 13346
rect 11158 13294 11180 13346
rect 11204 13294 11210 13346
rect 11210 13294 11222 13346
rect 11222 13294 11260 13346
rect 11284 13294 11286 13346
rect 11286 13294 11338 13346
rect 11338 13294 11340 13346
rect 10964 13292 11020 13294
rect 11044 13292 11100 13294
rect 11124 13292 11180 13294
rect 11204 13292 11260 13294
rect 11284 13292 11340 13294
rect 7964 3356 8020 3358
rect 8044 3356 8100 3358
rect 8124 3356 8180 3358
rect 8204 3356 8260 3358
rect 8284 3356 8340 3358
rect 7964 3304 7966 3356
rect 7966 3304 8018 3356
rect 8018 3304 8020 3356
rect 8044 3304 8082 3356
rect 8082 3304 8094 3356
rect 8094 3304 8100 3356
rect 8124 3304 8146 3356
rect 8146 3304 8158 3356
rect 8158 3304 8180 3356
rect 8204 3304 8210 3356
rect 8210 3304 8222 3356
rect 8222 3304 8260 3356
rect 8284 3304 8286 3356
rect 8286 3304 8338 3356
rect 8338 3304 8340 3356
rect 7964 3302 8020 3304
rect 8044 3302 8100 3304
rect 8124 3302 8180 3304
rect 8204 3302 8260 3304
rect 8284 3302 8340 3304
rect 4964 2690 5020 2692
rect 5044 2690 5100 2692
rect 5124 2690 5180 2692
rect 5204 2690 5260 2692
rect 5284 2690 5340 2692
rect 4964 2638 4966 2690
rect 4966 2638 5018 2690
rect 5018 2638 5020 2690
rect 5044 2638 5082 2690
rect 5082 2638 5094 2690
rect 5094 2638 5100 2690
rect 5124 2638 5146 2690
rect 5146 2638 5158 2690
rect 5158 2638 5180 2690
rect 5204 2638 5210 2690
rect 5210 2638 5222 2690
rect 5222 2638 5260 2690
rect 5284 2638 5286 2690
rect 5286 2638 5338 2690
rect 5338 2638 5340 2690
rect 4964 2636 5020 2638
rect 5044 2636 5100 2638
rect 5124 2636 5180 2638
rect 5204 2636 5260 2638
rect 5284 2636 5340 2638
rect 9812 934 9868 990
rect 10004 2118 10060 2174
rect 10964 12014 11020 12016
rect 11044 12014 11100 12016
rect 11124 12014 11180 12016
rect 11204 12014 11260 12016
rect 11284 12014 11340 12016
rect 10964 11962 10966 12014
rect 10966 11962 11018 12014
rect 11018 11962 11020 12014
rect 11044 11962 11082 12014
rect 11082 11962 11094 12014
rect 11094 11962 11100 12014
rect 11124 11962 11146 12014
rect 11146 11962 11158 12014
rect 11158 11962 11180 12014
rect 11204 11962 11210 12014
rect 11210 11962 11222 12014
rect 11222 11962 11260 12014
rect 11284 11962 11286 12014
rect 11286 11962 11338 12014
rect 11338 11962 11340 12014
rect 10964 11960 11020 11962
rect 11044 11960 11100 11962
rect 11124 11960 11180 11962
rect 11204 11960 11260 11962
rect 11284 11960 11340 11962
rect 10964 10682 11020 10684
rect 11044 10682 11100 10684
rect 11124 10682 11180 10684
rect 11204 10682 11260 10684
rect 11284 10682 11340 10684
rect 10964 10630 10966 10682
rect 10966 10630 11018 10682
rect 11018 10630 11020 10682
rect 11044 10630 11082 10682
rect 11082 10630 11094 10682
rect 11094 10630 11100 10682
rect 11124 10630 11146 10682
rect 11146 10630 11158 10682
rect 11158 10630 11180 10682
rect 11204 10630 11210 10682
rect 11210 10630 11222 10682
rect 11222 10630 11260 10682
rect 11284 10630 11286 10682
rect 11286 10630 11338 10682
rect 11338 10630 11340 10682
rect 10964 10628 11020 10630
rect 11044 10628 11100 10630
rect 11124 10628 11180 10630
rect 11204 10628 11260 10630
rect 11284 10628 11340 10630
rect 10964 9350 11020 9352
rect 11044 9350 11100 9352
rect 11124 9350 11180 9352
rect 11204 9350 11260 9352
rect 11284 9350 11340 9352
rect 10964 9298 10966 9350
rect 10966 9298 11018 9350
rect 11018 9298 11020 9350
rect 11044 9298 11082 9350
rect 11082 9298 11094 9350
rect 11094 9298 11100 9350
rect 11124 9298 11146 9350
rect 11146 9298 11158 9350
rect 11158 9298 11180 9350
rect 11204 9298 11210 9350
rect 11210 9298 11222 9350
rect 11222 9298 11260 9350
rect 11284 9298 11286 9350
rect 11286 9298 11338 9350
rect 11338 9298 11340 9350
rect 10964 9296 11020 9298
rect 11044 9296 11100 9298
rect 11124 9296 11180 9298
rect 11204 9296 11260 9298
rect 11284 9296 11340 9298
rect 11828 13405 11830 13422
rect 11830 13405 11882 13422
rect 11882 13405 11884 13422
rect 11828 13366 11884 13405
rect 12308 13958 12364 14014
rect 10964 8018 11020 8020
rect 11044 8018 11100 8020
rect 11124 8018 11180 8020
rect 11204 8018 11260 8020
rect 11284 8018 11340 8020
rect 10964 7966 10966 8018
rect 10966 7966 11018 8018
rect 11018 7966 11020 8018
rect 11044 7966 11082 8018
rect 11082 7966 11094 8018
rect 11094 7966 11100 8018
rect 11124 7966 11146 8018
rect 11146 7966 11158 8018
rect 11158 7966 11180 8018
rect 11204 7966 11210 8018
rect 11210 7966 11222 8018
rect 11222 7966 11260 8018
rect 11284 7966 11286 8018
rect 11286 7966 11338 8018
rect 11338 7966 11340 8018
rect 10964 7964 11020 7966
rect 11044 7964 11100 7966
rect 11124 7964 11180 7966
rect 11204 7964 11260 7966
rect 11284 7964 11340 7966
rect 10964 6686 11020 6688
rect 11044 6686 11100 6688
rect 11124 6686 11180 6688
rect 11204 6686 11260 6688
rect 11284 6686 11340 6688
rect 10964 6634 10966 6686
rect 10966 6634 11018 6686
rect 11018 6634 11020 6686
rect 11044 6634 11082 6686
rect 11082 6634 11094 6686
rect 11094 6634 11100 6686
rect 11124 6634 11146 6686
rect 11146 6634 11158 6686
rect 11158 6634 11180 6686
rect 11204 6634 11210 6686
rect 11210 6634 11222 6686
rect 11222 6634 11260 6686
rect 11284 6634 11286 6686
rect 11286 6634 11338 6686
rect 11338 6634 11340 6686
rect 10964 6632 11020 6634
rect 11044 6632 11100 6634
rect 11124 6632 11180 6634
rect 11204 6632 11260 6634
rect 11284 6632 11340 6634
rect 11348 5670 11404 5726
rect 10964 5354 11020 5356
rect 11044 5354 11100 5356
rect 11124 5354 11180 5356
rect 11204 5354 11260 5356
rect 11284 5354 11340 5356
rect 10964 5302 10966 5354
rect 10966 5302 11018 5354
rect 11018 5302 11020 5354
rect 11044 5302 11082 5354
rect 11082 5302 11094 5354
rect 11094 5302 11100 5354
rect 11124 5302 11146 5354
rect 11146 5302 11158 5354
rect 11158 5302 11180 5354
rect 11204 5302 11210 5354
rect 11210 5302 11222 5354
rect 11222 5302 11260 5354
rect 11284 5302 11286 5354
rect 11286 5302 11338 5354
rect 11338 5302 11340 5354
rect 10964 5300 11020 5302
rect 11044 5300 11100 5302
rect 11124 5300 11180 5302
rect 11204 5300 11260 5302
rect 11284 5300 11340 5302
rect 10964 4022 11020 4024
rect 11044 4022 11100 4024
rect 11124 4022 11180 4024
rect 11204 4022 11260 4024
rect 11284 4022 11340 4024
rect 10964 3970 10966 4022
rect 10966 3970 11018 4022
rect 11018 3970 11020 4022
rect 11044 3970 11082 4022
rect 11082 3970 11094 4022
rect 11094 3970 11100 4022
rect 11124 3970 11146 4022
rect 11146 3970 11158 4022
rect 11158 3970 11180 4022
rect 11204 3970 11210 4022
rect 11210 3970 11222 4022
rect 11222 3970 11260 4022
rect 11284 3970 11286 4022
rect 11286 3970 11338 4022
rect 11338 3970 11340 4022
rect 10964 3968 11020 3970
rect 11044 3968 11100 3970
rect 11124 3968 11180 3970
rect 11204 3968 11260 3970
rect 11284 3968 11340 3970
rect 11924 10406 11980 10462
rect 11924 6871 11980 6910
rect 11924 6854 11926 6871
rect 11926 6854 11978 6871
rect 11978 6854 11980 6871
rect 12404 12774 12460 12830
rect 12500 12182 12556 12238
rect 12500 10998 12556 11054
rect 12500 9814 12556 9870
rect 12500 9239 12556 9278
rect 12500 9222 12502 9239
rect 12502 9222 12554 9239
rect 12554 9222 12556 9239
rect 12500 8038 12556 8094
rect 12308 7446 12364 7502
rect 12500 6279 12556 6318
rect 12500 6262 12502 6279
rect 12502 6262 12554 6279
rect 12554 6262 12556 6279
rect 12500 5078 12556 5134
rect 12980 11590 13036 11646
rect 13172 9074 13228 9130
rect 12884 8630 12940 8686
rect 12884 4486 12940 4542
rect 12500 3894 12556 3950
rect 12308 3302 12364 3358
rect 11444 2710 11500 2766
rect 10964 2690 11020 2692
rect 11044 2690 11100 2692
rect 11124 2690 11180 2692
rect 11204 2690 11260 2692
rect 11284 2690 11340 2692
rect 10964 2638 10966 2690
rect 10966 2638 11018 2690
rect 11018 2638 11020 2690
rect 11044 2638 11082 2690
rect 11082 2638 11094 2690
rect 11094 2638 11100 2690
rect 11124 2638 11146 2690
rect 11146 2638 11158 2690
rect 11158 2638 11180 2690
rect 11204 2638 11210 2690
rect 11210 2638 11222 2690
rect 11222 2638 11260 2690
rect 11284 2638 11286 2690
rect 11286 2638 11338 2690
rect 11338 2638 11340 2690
rect 10964 2636 11020 2638
rect 11044 2636 11100 2638
rect 11124 2636 11180 2638
rect 11204 2636 11260 2638
rect 11284 2636 11340 2638
rect 10292 1526 10348 1582
<< metal3 >>
rect 8655 16384 8721 16387
rect 13498 16384 14298 16414
rect 8655 16382 14298 16384
rect 8655 16326 8660 16382
rect 8716 16326 14298 16382
rect 8655 16324 14298 16326
rect 8655 16321 8721 16324
rect 13498 16294 14298 16324
rect 9903 15792 9969 15795
rect 13498 15792 14298 15822
rect 9903 15790 14298 15792
rect 9903 15734 9908 15790
rect 9964 15734 14298 15790
rect 9903 15732 14298 15734
rect 9903 15729 9969 15732
rect 13498 15702 14298 15732
rect 8655 15200 8721 15203
rect 13498 15200 14298 15230
rect 8655 15198 14298 15200
rect 8655 15142 8660 15198
rect 8716 15142 14298 15198
rect 8655 15140 14298 15142
rect 8655 15137 8721 15140
rect 13498 15110 14298 15140
rect 4954 14684 5350 14685
rect 4954 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5350 14684
rect 4954 14619 5350 14620
rect 10954 14684 11350 14685
rect 10954 14620 10960 14684
rect 11024 14620 11040 14684
rect 11104 14620 11120 14684
rect 11184 14620 11200 14684
rect 11264 14620 11280 14684
rect 11344 14620 11350 14684
rect 10954 14619 11350 14620
rect 13498 14608 14298 14638
rect 11586 14548 14298 14608
rect 10671 14460 10737 14463
rect 11586 14460 11646 14548
rect 13498 14518 14298 14548
rect 10671 14458 11646 14460
rect 10671 14402 10676 14458
rect 10732 14402 11646 14458
rect 10671 14400 11646 14402
rect 10671 14397 10737 14400
rect 1954 14018 2350 14019
rect 1954 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2350 14018
rect 1954 13953 2350 13954
rect 7954 14018 8350 14019
rect 7954 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8350 14018
rect 7954 13953 8350 13954
rect 12303 14016 12369 14019
rect 13498 14016 14298 14046
rect 12303 14014 14298 14016
rect 12303 13958 12308 14014
rect 12364 13958 14298 14014
rect 12303 13956 14298 13958
rect 12303 13953 12369 13956
rect 13498 13926 14298 13956
rect 11823 13424 11889 13427
rect 13498 13424 14298 13454
rect 11823 13422 14298 13424
rect 11823 13366 11828 13422
rect 11884 13366 14298 13422
rect 11823 13364 14298 13366
rect 11823 13361 11889 13364
rect 4954 13352 5350 13353
rect 4954 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5350 13352
rect 4954 13287 5350 13288
rect 10954 13352 11350 13353
rect 10954 13288 10960 13352
rect 11024 13288 11040 13352
rect 11104 13288 11120 13352
rect 11184 13288 11200 13352
rect 11264 13288 11280 13352
rect 11344 13288 11350 13352
rect 13498 13334 14298 13364
rect 10954 13287 11350 13288
rect 12399 12832 12465 12835
rect 13498 12832 14298 12862
rect 12399 12830 14298 12832
rect 12399 12774 12404 12830
rect 12460 12774 14298 12830
rect 12399 12772 14298 12774
rect 12399 12769 12465 12772
rect 13498 12742 14298 12772
rect 1954 12686 2350 12687
rect 1954 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2350 12686
rect 1954 12621 2350 12622
rect 7954 12686 8350 12687
rect 7954 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8350 12686
rect 7954 12621 8350 12622
rect 12495 12240 12561 12243
rect 13498 12240 14298 12270
rect 12495 12238 14298 12240
rect 12495 12182 12500 12238
rect 12556 12182 14298 12238
rect 12495 12180 14298 12182
rect 12495 12177 12561 12180
rect 13498 12150 14298 12180
rect 4954 12020 5350 12021
rect 4954 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5350 12020
rect 4954 11955 5350 11956
rect 10954 12020 11350 12021
rect 10954 11956 10960 12020
rect 11024 11956 11040 12020
rect 11104 11956 11120 12020
rect 11184 11956 11200 12020
rect 11264 11956 11280 12020
rect 11344 11956 11350 12020
rect 10954 11955 11350 11956
rect 12975 11648 13041 11651
rect 13498 11648 14298 11678
rect 12975 11646 14298 11648
rect 12975 11590 12980 11646
rect 13036 11590 14298 11646
rect 12975 11588 14298 11590
rect 12975 11585 13041 11588
rect 13498 11558 14298 11588
rect 1954 11354 2350 11355
rect 1954 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2350 11354
rect 1954 11289 2350 11290
rect 7954 11354 8350 11355
rect 7954 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8350 11354
rect 7954 11289 8350 11290
rect 12495 11056 12561 11059
rect 13498 11056 14298 11086
rect 12495 11054 14298 11056
rect 12495 10998 12500 11054
rect 12556 10998 14298 11054
rect 12495 10996 14298 10998
rect 12495 10993 12561 10996
rect 13498 10966 14298 10996
rect 4954 10688 5350 10689
rect 4954 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5350 10688
rect 4954 10623 5350 10624
rect 10954 10688 11350 10689
rect 10954 10624 10960 10688
rect 11024 10624 11040 10688
rect 11104 10624 11120 10688
rect 11184 10624 11200 10688
rect 11264 10624 11280 10688
rect 11344 10624 11350 10688
rect 10954 10623 11350 10624
rect 11919 10464 11985 10467
rect 13498 10464 14298 10494
rect 11919 10462 14298 10464
rect 11919 10406 11924 10462
rect 11980 10406 14298 10462
rect 11919 10404 14298 10406
rect 11919 10401 11985 10404
rect 13498 10374 14298 10404
rect 1954 10022 2350 10023
rect 1954 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2350 10022
rect 1954 9957 2350 9958
rect 7954 10022 8350 10023
rect 7954 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8350 10022
rect 7954 9957 8350 9958
rect 12495 9872 12561 9875
rect 13498 9872 14298 9902
rect 12495 9870 14298 9872
rect 12495 9814 12500 9870
rect 12556 9814 14298 9870
rect 12495 9812 14298 9814
rect 12495 9809 12561 9812
rect 13498 9782 14298 9812
rect 4954 9356 5350 9357
rect 4954 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5350 9356
rect 4954 9291 5350 9292
rect 10954 9356 11350 9357
rect 10954 9292 10960 9356
rect 11024 9292 11040 9356
rect 11104 9292 11120 9356
rect 11184 9292 11200 9356
rect 11264 9292 11280 9356
rect 11344 9292 11350 9356
rect 10954 9291 11350 9292
rect 12495 9280 12561 9283
rect 13498 9280 14298 9310
rect 12495 9278 14298 9280
rect 12495 9222 12500 9278
rect 12556 9222 14298 9278
rect 12495 9220 14298 9222
rect 12495 9217 12561 9220
rect 13498 9190 14298 9220
rect 5199 9132 5265 9135
rect 13167 9132 13233 9135
rect 5199 9130 13233 9132
rect 5199 9074 5204 9130
rect 5260 9074 13172 9130
rect 13228 9074 13233 9130
rect 5199 9072 13233 9074
rect 5199 9069 5265 9072
rect 13167 9069 13233 9072
rect 1954 8690 2350 8691
rect 1954 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2350 8690
rect 1954 8625 2350 8626
rect 7954 8690 8350 8691
rect 7954 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8350 8690
rect 7954 8625 8350 8626
rect 12879 8688 12945 8691
rect 13498 8688 14298 8718
rect 12879 8686 14298 8688
rect 12879 8630 12884 8686
rect 12940 8630 14298 8686
rect 12879 8628 14298 8630
rect 12879 8625 12945 8628
rect 13498 8598 14298 8628
rect 12495 8096 12561 8099
rect 13498 8096 14298 8126
rect 12495 8094 14298 8096
rect 12495 8038 12500 8094
rect 12556 8038 14298 8094
rect 12495 8036 14298 8038
rect 12495 8033 12561 8036
rect 4954 8024 5350 8025
rect 4954 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5350 8024
rect 4954 7959 5350 7960
rect 10954 8024 11350 8025
rect 10954 7960 10960 8024
rect 11024 7960 11040 8024
rect 11104 7960 11120 8024
rect 11184 7960 11200 8024
rect 11264 7960 11280 8024
rect 11344 7960 11350 8024
rect 13498 8006 14298 8036
rect 10954 7959 11350 7960
rect 12303 7504 12369 7507
rect 13498 7504 14298 7534
rect 12303 7502 14298 7504
rect 12303 7446 12308 7502
rect 12364 7446 14298 7502
rect 12303 7444 14298 7446
rect 12303 7441 12369 7444
rect 13498 7414 14298 7444
rect 1954 7358 2350 7359
rect 1954 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2350 7358
rect 1954 7293 2350 7294
rect 7954 7358 8350 7359
rect 7954 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8350 7358
rect 7954 7293 8350 7294
rect 11919 6912 11985 6915
rect 13498 6912 14298 6942
rect 11919 6910 14298 6912
rect 11919 6854 11924 6910
rect 11980 6854 14298 6910
rect 11919 6852 14298 6854
rect 11919 6849 11985 6852
rect 13498 6822 14298 6852
rect 4954 6692 5350 6693
rect 4954 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5350 6692
rect 4954 6627 5350 6628
rect 10954 6692 11350 6693
rect 10954 6628 10960 6692
rect 11024 6628 11040 6692
rect 11104 6628 11120 6692
rect 11184 6628 11200 6692
rect 11264 6628 11280 6692
rect 11344 6628 11350 6692
rect 10954 6627 11350 6628
rect 12495 6320 12561 6323
rect 13498 6320 14298 6350
rect 12495 6318 14298 6320
rect 12495 6262 12500 6318
rect 12556 6262 14298 6318
rect 12495 6260 14298 6262
rect 12495 6257 12561 6260
rect 13498 6230 14298 6260
rect 1954 6026 2350 6027
rect 1954 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2350 6026
rect 1954 5961 2350 5962
rect 7954 6026 8350 6027
rect 7954 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8350 6026
rect 7954 5961 8350 5962
rect 11343 5728 11409 5731
rect 13498 5728 14298 5758
rect 11343 5726 14298 5728
rect 11343 5670 11348 5726
rect 11404 5670 14298 5726
rect 11343 5668 14298 5670
rect 11343 5665 11409 5668
rect 13498 5638 14298 5668
rect 4954 5360 5350 5361
rect 4954 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5350 5360
rect 4954 5295 5350 5296
rect 10954 5360 11350 5361
rect 10954 5296 10960 5360
rect 11024 5296 11040 5360
rect 11104 5296 11120 5360
rect 11184 5296 11200 5360
rect 11264 5296 11280 5360
rect 11344 5296 11350 5360
rect 10954 5295 11350 5296
rect 12495 5136 12561 5139
rect 13498 5136 14298 5166
rect 12495 5134 14298 5136
rect 12495 5078 12500 5134
rect 12556 5078 14298 5134
rect 12495 5076 14298 5078
rect 12495 5073 12561 5076
rect 13498 5046 14298 5076
rect 1954 4694 2350 4695
rect 1954 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2350 4694
rect 1954 4629 2350 4630
rect 7954 4694 8350 4695
rect 7954 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8350 4694
rect 7954 4629 8350 4630
rect 12879 4544 12945 4547
rect 13498 4544 14298 4574
rect 12879 4542 14298 4544
rect 12879 4486 12884 4542
rect 12940 4486 14298 4542
rect 12879 4484 14298 4486
rect 12879 4481 12945 4484
rect 13498 4454 14298 4484
rect 4954 4028 5350 4029
rect 4954 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5350 4028
rect 4954 3963 5350 3964
rect 10954 4028 11350 4029
rect 10954 3964 10960 4028
rect 11024 3964 11040 4028
rect 11104 3964 11120 4028
rect 11184 3964 11200 4028
rect 11264 3964 11280 4028
rect 11344 3964 11350 4028
rect 10954 3963 11350 3964
rect 12495 3952 12561 3955
rect 13498 3952 14298 3982
rect 12495 3950 14298 3952
rect 12495 3894 12500 3950
rect 12556 3894 14298 3950
rect 12495 3892 14298 3894
rect 12495 3889 12561 3892
rect 13498 3862 14298 3892
rect 1954 3362 2350 3363
rect 1954 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2350 3362
rect 1954 3297 2350 3298
rect 7954 3362 8350 3363
rect 7954 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8350 3362
rect 7954 3297 8350 3298
rect 12303 3360 12369 3363
rect 13498 3360 14298 3390
rect 12303 3358 14298 3360
rect 12303 3302 12308 3358
rect 12364 3302 14298 3358
rect 12303 3300 14298 3302
rect 12303 3297 12369 3300
rect 13498 3270 14298 3300
rect 11439 2768 11505 2771
rect 13498 2768 14298 2798
rect 11439 2766 14298 2768
rect 11439 2710 11444 2766
rect 11500 2710 14298 2766
rect 11439 2708 14298 2710
rect 11439 2705 11505 2708
rect 4954 2696 5350 2697
rect 4954 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5350 2696
rect 4954 2631 5350 2632
rect 10954 2696 11350 2697
rect 10954 2632 10960 2696
rect 11024 2632 11040 2696
rect 11104 2632 11120 2696
rect 11184 2632 11200 2696
rect 11264 2632 11280 2696
rect 11344 2632 11350 2696
rect 13498 2678 14298 2708
rect 10954 2631 11350 2632
rect 9999 2176 10065 2179
rect 13498 2176 14298 2206
rect 9999 2174 14298 2176
rect 9999 2118 10004 2174
rect 10060 2118 14298 2174
rect 9999 2116 14298 2118
rect 9999 2113 10065 2116
rect 13498 2086 14298 2116
rect 10287 1584 10353 1587
rect 13498 1584 14298 1614
rect 10287 1582 14298 1584
rect 10287 1526 10292 1582
rect 10348 1526 14298 1582
rect 10287 1524 14298 1526
rect 10287 1521 10353 1524
rect 13498 1494 14298 1524
rect 9807 992 9873 995
rect 13498 992 14298 1022
rect 9807 990 14298 992
rect 9807 934 9812 990
rect 9868 934 14298 990
rect 9807 932 14298 934
rect 9807 929 9873 932
rect 13498 902 14298 932
<< via3 >>
rect 4960 14680 5024 14684
rect 4960 14624 4964 14680
rect 4964 14624 5020 14680
rect 5020 14624 5024 14680
rect 4960 14620 5024 14624
rect 5040 14680 5104 14684
rect 5040 14624 5044 14680
rect 5044 14624 5100 14680
rect 5100 14624 5104 14680
rect 5040 14620 5104 14624
rect 5120 14680 5184 14684
rect 5120 14624 5124 14680
rect 5124 14624 5180 14680
rect 5180 14624 5184 14680
rect 5120 14620 5184 14624
rect 5200 14680 5264 14684
rect 5200 14624 5204 14680
rect 5204 14624 5260 14680
rect 5260 14624 5264 14680
rect 5200 14620 5264 14624
rect 5280 14680 5344 14684
rect 5280 14624 5284 14680
rect 5284 14624 5340 14680
rect 5340 14624 5344 14680
rect 5280 14620 5344 14624
rect 10960 14680 11024 14684
rect 10960 14624 10964 14680
rect 10964 14624 11020 14680
rect 11020 14624 11024 14680
rect 10960 14620 11024 14624
rect 11040 14680 11104 14684
rect 11040 14624 11044 14680
rect 11044 14624 11100 14680
rect 11100 14624 11104 14680
rect 11040 14620 11104 14624
rect 11120 14680 11184 14684
rect 11120 14624 11124 14680
rect 11124 14624 11180 14680
rect 11180 14624 11184 14680
rect 11120 14620 11184 14624
rect 11200 14680 11264 14684
rect 11200 14624 11204 14680
rect 11204 14624 11260 14680
rect 11260 14624 11264 14680
rect 11200 14620 11264 14624
rect 11280 14680 11344 14684
rect 11280 14624 11284 14680
rect 11284 14624 11340 14680
rect 11340 14624 11344 14680
rect 11280 14620 11344 14624
rect 1960 14014 2024 14018
rect 1960 13958 1964 14014
rect 1964 13958 2020 14014
rect 2020 13958 2024 14014
rect 1960 13954 2024 13958
rect 2040 14014 2104 14018
rect 2040 13958 2044 14014
rect 2044 13958 2100 14014
rect 2100 13958 2104 14014
rect 2040 13954 2104 13958
rect 2120 14014 2184 14018
rect 2120 13958 2124 14014
rect 2124 13958 2180 14014
rect 2180 13958 2184 14014
rect 2120 13954 2184 13958
rect 2200 14014 2264 14018
rect 2200 13958 2204 14014
rect 2204 13958 2260 14014
rect 2260 13958 2264 14014
rect 2200 13954 2264 13958
rect 2280 14014 2344 14018
rect 2280 13958 2284 14014
rect 2284 13958 2340 14014
rect 2340 13958 2344 14014
rect 2280 13954 2344 13958
rect 7960 14014 8024 14018
rect 7960 13958 7964 14014
rect 7964 13958 8020 14014
rect 8020 13958 8024 14014
rect 7960 13954 8024 13958
rect 8040 14014 8104 14018
rect 8040 13958 8044 14014
rect 8044 13958 8100 14014
rect 8100 13958 8104 14014
rect 8040 13954 8104 13958
rect 8120 14014 8184 14018
rect 8120 13958 8124 14014
rect 8124 13958 8180 14014
rect 8180 13958 8184 14014
rect 8120 13954 8184 13958
rect 8200 14014 8264 14018
rect 8200 13958 8204 14014
rect 8204 13958 8260 14014
rect 8260 13958 8264 14014
rect 8200 13954 8264 13958
rect 8280 14014 8344 14018
rect 8280 13958 8284 14014
rect 8284 13958 8340 14014
rect 8340 13958 8344 14014
rect 8280 13954 8344 13958
rect 4960 13348 5024 13352
rect 4960 13292 4964 13348
rect 4964 13292 5020 13348
rect 5020 13292 5024 13348
rect 4960 13288 5024 13292
rect 5040 13348 5104 13352
rect 5040 13292 5044 13348
rect 5044 13292 5100 13348
rect 5100 13292 5104 13348
rect 5040 13288 5104 13292
rect 5120 13348 5184 13352
rect 5120 13292 5124 13348
rect 5124 13292 5180 13348
rect 5180 13292 5184 13348
rect 5120 13288 5184 13292
rect 5200 13348 5264 13352
rect 5200 13292 5204 13348
rect 5204 13292 5260 13348
rect 5260 13292 5264 13348
rect 5200 13288 5264 13292
rect 5280 13348 5344 13352
rect 5280 13292 5284 13348
rect 5284 13292 5340 13348
rect 5340 13292 5344 13348
rect 5280 13288 5344 13292
rect 10960 13348 11024 13352
rect 10960 13292 10964 13348
rect 10964 13292 11020 13348
rect 11020 13292 11024 13348
rect 10960 13288 11024 13292
rect 11040 13348 11104 13352
rect 11040 13292 11044 13348
rect 11044 13292 11100 13348
rect 11100 13292 11104 13348
rect 11040 13288 11104 13292
rect 11120 13348 11184 13352
rect 11120 13292 11124 13348
rect 11124 13292 11180 13348
rect 11180 13292 11184 13348
rect 11120 13288 11184 13292
rect 11200 13348 11264 13352
rect 11200 13292 11204 13348
rect 11204 13292 11260 13348
rect 11260 13292 11264 13348
rect 11200 13288 11264 13292
rect 11280 13348 11344 13352
rect 11280 13292 11284 13348
rect 11284 13292 11340 13348
rect 11340 13292 11344 13348
rect 11280 13288 11344 13292
rect 1960 12682 2024 12686
rect 1960 12626 1964 12682
rect 1964 12626 2020 12682
rect 2020 12626 2024 12682
rect 1960 12622 2024 12626
rect 2040 12682 2104 12686
rect 2040 12626 2044 12682
rect 2044 12626 2100 12682
rect 2100 12626 2104 12682
rect 2040 12622 2104 12626
rect 2120 12682 2184 12686
rect 2120 12626 2124 12682
rect 2124 12626 2180 12682
rect 2180 12626 2184 12682
rect 2120 12622 2184 12626
rect 2200 12682 2264 12686
rect 2200 12626 2204 12682
rect 2204 12626 2260 12682
rect 2260 12626 2264 12682
rect 2200 12622 2264 12626
rect 2280 12682 2344 12686
rect 2280 12626 2284 12682
rect 2284 12626 2340 12682
rect 2340 12626 2344 12682
rect 2280 12622 2344 12626
rect 7960 12682 8024 12686
rect 7960 12626 7964 12682
rect 7964 12626 8020 12682
rect 8020 12626 8024 12682
rect 7960 12622 8024 12626
rect 8040 12682 8104 12686
rect 8040 12626 8044 12682
rect 8044 12626 8100 12682
rect 8100 12626 8104 12682
rect 8040 12622 8104 12626
rect 8120 12682 8184 12686
rect 8120 12626 8124 12682
rect 8124 12626 8180 12682
rect 8180 12626 8184 12682
rect 8120 12622 8184 12626
rect 8200 12682 8264 12686
rect 8200 12626 8204 12682
rect 8204 12626 8260 12682
rect 8260 12626 8264 12682
rect 8200 12622 8264 12626
rect 8280 12682 8344 12686
rect 8280 12626 8284 12682
rect 8284 12626 8340 12682
rect 8340 12626 8344 12682
rect 8280 12622 8344 12626
rect 4960 12016 5024 12020
rect 4960 11960 4964 12016
rect 4964 11960 5020 12016
rect 5020 11960 5024 12016
rect 4960 11956 5024 11960
rect 5040 12016 5104 12020
rect 5040 11960 5044 12016
rect 5044 11960 5100 12016
rect 5100 11960 5104 12016
rect 5040 11956 5104 11960
rect 5120 12016 5184 12020
rect 5120 11960 5124 12016
rect 5124 11960 5180 12016
rect 5180 11960 5184 12016
rect 5120 11956 5184 11960
rect 5200 12016 5264 12020
rect 5200 11960 5204 12016
rect 5204 11960 5260 12016
rect 5260 11960 5264 12016
rect 5200 11956 5264 11960
rect 5280 12016 5344 12020
rect 5280 11960 5284 12016
rect 5284 11960 5340 12016
rect 5340 11960 5344 12016
rect 5280 11956 5344 11960
rect 10960 12016 11024 12020
rect 10960 11960 10964 12016
rect 10964 11960 11020 12016
rect 11020 11960 11024 12016
rect 10960 11956 11024 11960
rect 11040 12016 11104 12020
rect 11040 11960 11044 12016
rect 11044 11960 11100 12016
rect 11100 11960 11104 12016
rect 11040 11956 11104 11960
rect 11120 12016 11184 12020
rect 11120 11960 11124 12016
rect 11124 11960 11180 12016
rect 11180 11960 11184 12016
rect 11120 11956 11184 11960
rect 11200 12016 11264 12020
rect 11200 11960 11204 12016
rect 11204 11960 11260 12016
rect 11260 11960 11264 12016
rect 11200 11956 11264 11960
rect 11280 12016 11344 12020
rect 11280 11960 11284 12016
rect 11284 11960 11340 12016
rect 11340 11960 11344 12016
rect 11280 11956 11344 11960
rect 1960 11350 2024 11354
rect 1960 11294 1964 11350
rect 1964 11294 2020 11350
rect 2020 11294 2024 11350
rect 1960 11290 2024 11294
rect 2040 11350 2104 11354
rect 2040 11294 2044 11350
rect 2044 11294 2100 11350
rect 2100 11294 2104 11350
rect 2040 11290 2104 11294
rect 2120 11350 2184 11354
rect 2120 11294 2124 11350
rect 2124 11294 2180 11350
rect 2180 11294 2184 11350
rect 2120 11290 2184 11294
rect 2200 11350 2264 11354
rect 2200 11294 2204 11350
rect 2204 11294 2260 11350
rect 2260 11294 2264 11350
rect 2200 11290 2264 11294
rect 2280 11350 2344 11354
rect 2280 11294 2284 11350
rect 2284 11294 2340 11350
rect 2340 11294 2344 11350
rect 2280 11290 2344 11294
rect 7960 11350 8024 11354
rect 7960 11294 7964 11350
rect 7964 11294 8020 11350
rect 8020 11294 8024 11350
rect 7960 11290 8024 11294
rect 8040 11350 8104 11354
rect 8040 11294 8044 11350
rect 8044 11294 8100 11350
rect 8100 11294 8104 11350
rect 8040 11290 8104 11294
rect 8120 11350 8184 11354
rect 8120 11294 8124 11350
rect 8124 11294 8180 11350
rect 8180 11294 8184 11350
rect 8120 11290 8184 11294
rect 8200 11350 8264 11354
rect 8200 11294 8204 11350
rect 8204 11294 8260 11350
rect 8260 11294 8264 11350
rect 8200 11290 8264 11294
rect 8280 11350 8344 11354
rect 8280 11294 8284 11350
rect 8284 11294 8340 11350
rect 8340 11294 8344 11350
rect 8280 11290 8344 11294
rect 4960 10684 5024 10688
rect 4960 10628 4964 10684
rect 4964 10628 5020 10684
rect 5020 10628 5024 10684
rect 4960 10624 5024 10628
rect 5040 10684 5104 10688
rect 5040 10628 5044 10684
rect 5044 10628 5100 10684
rect 5100 10628 5104 10684
rect 5040 10624 5104 10628
rect 5120 10684 5184 10688
rect 5120 10628 5124 10684
rect 5124 10628 5180 10684
rect 5180 10628 5184 10684
rect 5120 10624 5184 10628
rect 5200 10684 5264 10688
rect 5200 10628 5204 10684
rect 5204 10628 5260 10684
rect 5260 10628 5264 10684
rect 5200 10624 5264 10628
rect 5280 10684 5344 10688
rect 5280 10628 5284 10684
rect 5284 10628 5340 10684
rect 5340 10628 5344 10684
rect 5280 10624 5344 10628
rect 10960 10684 11024 10688
rect 10960 10628 10964 10684
rect 10964 10628 11020 10684
rect 11020 10628 11024 10684
rect 10960 10624 11024 10628
rect 11040 10684 11104 10688
rect 11040 10628 11044 10684
rect 11044 10628 11100 10684
rect 11100 10628 11104 10684
rect 11040 10624 11104 10628
rect 11120 10684 11184 10688
rect 11120 10628 11124 10684
rect 11124 10628 11180 10684
rect 11180 10628 11184 10684
rect 11120 10624 11184 10628
rect 11200 10684 11264 10688
rect 11200 10628 11204 10684
rect 11204 10628 11260 10684
rect 11260 10628 11264 10684
rect 11200 10624 11264 10628
rect 11280 10684 11344 10688
rect 11280 10628 11284 10684
rect 11284 10628 11340 10684
rect 11340 10628 11344 10684
rect 11280 10624 11344 10628
rect 1960 10018 2024 10022
rect 1960 9962 1964 10018
rect 1964 9962 2020 10018
rect 2020 9962 2024 10018
rect 1960 9958 2024 9962
rect 2040 10018 2104 10022
rect 2040 9962 2044 10018
rect 2044 9962 2100 10018
rect 2100 9962 2104 10018
rect 2040 9958 2104 9962
rect 2120 10018 2184 10022
rect 2120 9962 2124 10018
rect 2124 9962 2180 10018
rect 2180 9962 2184 10018
rect 2120 9958 2184 9962
rect 2200 10018 2264 10022
rect 2200 9962 2204 10018
rect 2204 9962 2260 10018
rect 2260 9962 2264 10018
rect 2200 9958 2264 9962
rect 2280 10018 2344 10022
rect 2280 9962 2284 10018
rect 2284 9962 2340 10018
rect 2340 9962 2344 10018
rect 2280 9958 2344 9962
rect 7960 10018 8024 10022
rect 7960 9962 7964 10018
rect 7964 9962 8020 10018
rect 8020 9962 8024 10018
rect 7960 9958 8024 9962
rect 8040 10018 8104 10022
rect 8040 9962 8044 10018
rect 8044 9962 8100 10018
rect 8100 9962 8104 10018
rect 8040 9958 8104 9962
rect 8120 10018 8184 10022
rect 8120 9962 8124 10018
rect 8124 9962 8180 10018
rect 8180 9962 8184 10018
rect 8120 9958 8184 9962
rect 8200 10018 8264 10022
rect 8200 9962 8204 10018
rect 8204 9962 8260 10018
rect 8260 9962 8264 10018
rect 8200 9958 8264 9962
rect 8280 10018 8344 10022
rect 8280 9962 8284 10018
rect 8284 9962 8340 10018
rect 8340 9962 8344 10018
rect 8280 9958 8344 9962
rect 4960 9352 5024 9356
rect 4960 9296 4964 9352
rect 4964 9296 5020 9352
rect 5020 9296 5024 9352
rect 4960 9292 5024 9296
rect 5040 9352 5104 9356
rect 5040 9296 5044 9352
rect 5044 9296 5100 9352
rect 5100 9296 5104 9352
rect 5040 9292 5104 9296
rect 5120 9352 5184 9356
rect 5120 9296 5124 9352
rect 5124 9296 5180 9352
rect 5180 9296 5184 9352
rect 5120 9292 5184 9296
rect 5200 9352 5264 9356
rect 5200 9296 5204 9352
rect 5204 9296 5260 9352
rect 5260 9296 5264 9352
rect 5200 9292 5264 9296
rect 5280 9352 5344 9356
rect 5280 9296 5284 9352
rect 5284 9296 5340 9352
rect 5340 9296 5344 9352
rect 5280 9292 5344 9296
rect 10960 9352 11024 9356
rect 10960 9296 10964 9352
rect 10964 9296 11020 9352
rect 11020 9296 11024 9352
rect 10960 9292 11024 9296
rect 11040 9352 11104 9356
rect 11040 9296 11044 9352
rect 11044 9296 11100 9352
rect 11100 9296 11104 9352
rect 11040 9292 11104 9296
rect 11120 9352 11184 9356
rect 11120 9296 11124 9352
rect 11124 9296 11180 9352
rect 11180 9296 11184 9352
rect 11120 9292 11184 9296
rect 11200 9352 11264 9356
rect 11200 9296 11204 9352
rect 11204 9296 11260 9352
rect 11260 9296 11264 9352
rect 11200 9292 11264 9296
rect 11280 9352 11344 9356
rect 11280 9296 11284 9352
rect 11284 9296 11340 9352
rect 11340 9296 11344 9352
rect 11280 9292 11344 9296
rect 1960 8686 2024 8690
rect 1960 8630 1964 8686
rect 1964 8630 2020 8686
rect 2020 8630 2024 8686
rect 1960 8626 2024 8630
rect 2040 8686 2104 8690
rect 2040 8630 2044 8686
rect 2044 8630 2100 8686
rect 2100 8630 2104 8686
rect 2040 8626 2104 8630
rect 2120 8686 2184 8690
rect 2120 8630 2124 8686
rect 2124 8630 2180 8686
rect 2180 8630 2184 8686
rect 2120 8626 2184 8630
rect 2200 8686 2264 8690
rect 2200 8630 2204 8686
rect 2204 8630 2260 8686
rect 2260 8630 2264 8686
rect 2200 8626 2264 8630
rect 2280 8686 2344 8690
rect 2280 8630 2284 8686
rect 2284 8630 2340 8686
rect 2340 8630 2344 8686
rect 2280 8626 2344 8630
rect 7960 8686 8024 8690
rect 7960 8630 7964 8686
rect 7964 8630 8020 8686
rect 8020 8630 8024 8686
rect 7960 8626 8024 8630
rect 8040 8686 8104 8690
rect 8040 8630 8044 8686
rect 8044 8630 8100 8686
rect 8100 8630 8104 8686
rect 8040 8626 8104 8630
rect 8120 8686 8184 8690
rect 8120 8630 8124 8686
rect 8124 8630 8180 8686
rect 8180 8630 8184 8686
rect 8120 8626 8184 8630
rect 8200 8686 8264 8690
rect 8200 8630 8204 8686
rect 8204 8630 8260 8686
rect 8260 8630 8264 8686
rect 8200 8626 8264 8630
rect 8280 8686 8344 8690
rect 8280 8630 8284 8686
rect 8284 8630 8340 8686
rect 8340 8630 8344 8686
rect 8280 8626 8344 8630
rect 4960 8020 5024 8024
rect 4960 7964 4964 8020
rect 4964 7964 5020 8020
rect 5020 7964 5024 8020
rect 4960 7960 5024 7964
rect 5040 8020 5104 8024
rect 5040 7964 5044 8020
rect 5044 7964 5100 8020
rect 5100 7964 5104 8020
rect 5040 7960 5104 7964
rect 5120 8020 5184 8024
rect 5120 7964 5124 8020
rect 5124 7964 5180 8020
rect 5180 7964 5184 8020
rect 5120 7960 5184 7964
rect 5200 8020 5264 8024
rect 5200 7964 5204 8020
rect 5204 7964 5260 8020
rect 5260 7964 5264 8020
rect 5200 7960 5264 7964
rect 5280 8020 5344 8024
rect 5280 7964 5284 8020
rect 5284 7964 5340 8020
rect 5340 7964 5344 8020
rect 5280 7960 5344 7964
rect 10960 8020 11024 8024
rect 10960 7964 10964 8020
rect 10964 7964 11020 8020
rect 11020 7964 11024 8020
rect 10960 7960 11024 7964
rect 11040 8020 11104 8024
rect 11040 7964 11044 8020
rect 11044 7964 11100 8020
rect 11100 7964 11104 8020
rect 11040 7960 11104 7964
rect 11120 8020 11184 8024
rect 11120 7964 11124 8020
rect 11124 7964 11180 8020
rect 11180 7964 11184 8020
rect 11120 7960 11184 7964
rect 11200 8020 11264 8024
rect 11200 7964 11204 8020
rect 11204 7964 11260 8020
rect 11260 7964 11264 8020
rect 11200 7960 11264 7964
rect 11280 8020 11344 8024
rect 11280 7964 11284 8020
rect 11284 7964 11340 8020
rect 11340 7964 11344 8020
rect 11280 7960 11344 7964
rect 1960 7354 2024 7358
rect 1960 7298 1964 7354
rect 1964 7298 2020 7354
rect 2020 7298 2024 7354
rect 1960 7294 2024 7298
rect 2040 7354 2104 7358
rect 2040 7298 2044 7354
rect 2044 7298 2100 7354
rect 2100 7298 2104 7354
rect 2040 7294 2104 7298
rect 2120 7354 2184 7358
rect 2120 7298 2124 7354
rect 2124 7298 2180 7354
rect 2180 7298 2184 7354
rect 2120 7294 2184 7298
rect 2200 7354 2264 7358
rect 2200 7298 2204 7354
rect 2204 7298 2260 7354
rect 2260 7298 2264 7354
rect 2200 7294 2264 7298
rect 2280 7354 2344 7358
rect 2280 7298 2284 7354
rect 2284 7298 2340 7354
rect 2340 7298 2344 7354
rect 2280 7294 2344 7298
rect 7960 7354 8024 7358
rect 7960 7298 7964 7354
rect 7964 7298 8020 7354
rect 8020 7298 8024 7354
rect 7960 7294 8024 7298
rect 8040 7354 8104 7358
rect 8040 7298 8044 7354
rect 8044 7298 8100 7354
rect 8100 7298 8104 7354
rect 8040 7294 8104 7298
rect 8120 7354 8184 7358
rect 8120 7298 8124 7354
rect 8124 7298 8180 7354
rect 8180 7298 8184 7354
rect 8120 7294 8184 7298
rect 8200 7354 8264 7358
rect 8200 7298 8204 7354
rect 8204 7298 8260 7354
rect 8260 7298 8264 7354
rect 8200 7294 8264 7298
rect 8280 7354 8344 7358
rect 8280 7298 8284 7354
rect 8284 7298 8340 7354
rect 8340 7298 8344 7354
rect 8280 7294 8344 7298
rect 4960 6688 5024 6692
rect 4960 6632 4964 6688
rect 4964 6632 5020 6688
rect 5020 6632 5024 6688
rect 4960 6628 5024 6632
rect 5040 6688 5104 6692
rect 5040 6632 5044 6688
rect 5044 6632 5100 6688
rect 5100 6632 5104 6688
rect 5040 6628 5104 6632
rect 5120 6688 5184 6692
rect 5120 6632 5124 6688
rect 5124 6632 5180 6688
rect 5180 6632 5184 6688
rect 5120 6628 5184 6632
rect 5200 6688 5264 6692
rect 5200 6632 5204 6688
rect 5204 6632 5260 6688
rect 5260 6632 5264 6688
rect 5200 6628 5264 6632
rect 5280 6688 5344 6692
rect 5280 6632 5284 6688
rect 5284 6632 5340 6688
rect 5340 6632 5344 6688
rect 5280 6628 5344 6632
rect 10960 6688 11024 6692
rect 10960 6632 10964 6688
rect 10964 6632 11020 6688
rect 11020 6632 11024 6688
rect 10960 6628 11024 6632
rect 11040 6688 11104 6692
rect 11040 6632 11044 6688
rect 11044 6632 11100 6688
rect 11100 6632 11104 6688
rect 11040 6628 11104 6632
rect 11120 6688 11184 6692
rect 11120 6632 11124 6688
rect 11124 6632 11180 6688
rect 11180 6632 11184 6688
rect 11120 6628 11184 6632
rect 11200 6688 11264 6692
rect 11200 6632 11204 6688
rect 11204 6632 11260 6688
rect 11260 6632 11264 6688
rect 11200 6628 11264 6632
rect 11280 6688 11344 6692
rect 11280 6632 11284 6688
rect 11284 6632 11340 6688
rect 11340 6632 11344 6688
rect 11280 6628 11344 6632
rect 1960 6022 2024 6026
rect 1960 5966 1964 6022
rect 1964 5966 2020 6022
rect 2020 5966 2024 6022
rect 1960 5962 2024 5966
rect 2040 6022 2104 6026
rect 2040 5966 2044 6022
rect 2044 5966 2100 6022
rect 2100 5966 2104 6022
rect 2040 5962 2104 5966
rect 2120 6022 2184 6026
rect 2120 5966 2124 6022
rect 2124 5966 2180 6022
rect 2180 5966 2184 6022
rect 2120 5962 2184 5966
rect 2200 6022 2264 6026
rect 2200 5966 2204 6022
rect 2204 5966 2260 6022
rect 2260 5966 2264 6022
rect 2200 5962 2264 5966
rect 2280 6022 2344 6026
rect 2280 5966 2284 6022
rect 2284 5966 2340 6022
rect 2340 5966 2344 6022
rect 2280 5962 2344 5966
rect 7960 6022 8024 6026
rect 7960 5966 7964 6022
rect 7964 5966 8020 6022
rect 8020 5966 8024 6022
rect 7960 5962 8024 5966
rect 8040 6022 8104 6026
rect 8040 5966 8044 6022
rect 8044 5966 8100 6022
rect 8100 5966 8104 6022
rect 8040 5962 8104 5966
rect 8120 6022 8184 6026
rect 8120 5966 8124 6022
rect 8124 5966 8180 6022
rect 8180 5966 8184 6022
rect 8120 5962 8184 5966
rect 8200 6022 8264 6026
rect 8200 5966 8204 6022
rect 8204 5966 8260 6022
rect 8260 5966 8264 6022
rect 8200 5962 8264 5966
rect 8280 6022 8344 6026
rect 8280 5966 8284 6022
rect 8284 5966 8340 6022
rect 8340 5966 8344 6022
rect 8280 5962 8344 5966
rect 4960 5356 5024 5360
rect 4960 5300 4964 5356
rect 4964 5300 5020 5356
rect 5020 5300 5024 5356
rect 4960 5296 5024 5300
rect 5040 5356 5104 5360
rect 5040 5300 5044 5356
rect 5044 5300 5100 5356
rect 5100 5300 5104 5356
rect 5040 5296 5104 5300
rect 5120 5356 5184 5360
rect 5120 5300 5124 5356
rect 5124 5300 5180 5356
rect 5180 5300 5184 5356
rect 5120 5296 5184 5300
rect 5200 5356 5264 5360
rect 5200 5300 5204 5356
rect 5204 5300 5260 5356
rect 5260 5300 5264 5356
rect 5200 5296 5264 5300
rect 5280 5356 5344 5360
rect 5280 5300 5284 5356
rect 5284 5300 5340 5356
rect 5340 5300 5344 5356
rect 5280 5296 5344 5300
rect 10960 5356 11024 5360
rect 10960 5300 10964 5356
rect 10964 5300 11020 5356
rect 11020 5300 11024 5356
rect 10960 5296 11024 5300
rect 11040 5356 11104 5360
rect 11040 5300 11044 5356
rect 11044 5300 11100 5356
rect 11100 5300 11104 5356
rect 11040 5296 11104 5300
rect 11120 5356 11184 5360
rect 11120 5300 11124 5356
rect 11124 5300 11180 5356
rect 11180 5300 11184 5356
rect 11120 5296 11184 5300
rect 11200 5356 11264 5360
rect 11200 5300 11204 5356
rect 11204 5300 11260 5356
rect 11260 5300 11264 5356
rect 11200 5296 11264 5300
rect 11280 5356 11344 5360
rect 11280 5300 11284 5356
rect 11284 5300 11340 5356
rect 11340 5300 11344 5356
rect 11280 5296 11344 5300
rect 1960 4690 2024 4694
rect 1960 4634 1964 4690
rect 1964 4634 2020 4690
rect 2020 4634 2024 4690
rect 1960 4630 2024 4634
rect 2040 4690 2104 4694
rect 2040 4634 2044 4690
rect 2044 4634 2100 4690
rect 2100 4634 2104 4690
rect 2040 4630 2104 4634
rect 2120 4690 2184 4694
rect 2120 4634 2124 4690
rect 2124 4634 2180 4690
rect 2180 4634 2184 4690
rect 2120 4630 2184 4634
rect 2200 4690 2264 4694
rect 2200 4634 2204 4690
rect 2204 4634 2260 4690
rect 2260 4634 2264 4690
rect 2200 4630 2264 4634
rect 2280 4690 2344 4694
rect 2280 4634 2284 4690
rect 2284 4634 2340 4690
rect 2340 4634 2344 4690
rect 2280 4630 2344 4634
rect 7960 4690 8024 4694
rect 7960 4634 7964 4690
rect 7964 4634 8020 4690
rect 8020 4634 8024 4690
rect 7960 4630 8024 4634
rect 8040 4690 8104 4694
rect 8040 4634 8044 4690
rect 8044 4634 8100 4690
rect 8100 4634 8104 4690
rect 8040 4630 8104 4634
rect 8120 4690 8184 4694
rect 8120 4634 8124 4690
rect 8124 4634 8180 4690
rect 8180 4634 8184 4690
rect 8120 4630 8184 4634
rect 8200 4690 8264 4694
rect 8200 4634 8204 4690
rect 8204 4634 8260 4690
rect 8260 4634 8264 4690
rect 8200 4630 8264 4634
rect 8280 4690 8344 4694
rect 8280 4634 8284 4690
rect 8284 4634 8340 4690
rect 8340 4634 8344 4690
rect 8280 4630 8344 4634
rect 4960 4024 5024 4028
rect 4960 3968 4964 4024
rect 4964 3968 5020 4024
rect 5020 3968 5024 4024
rect 4960 3964 5024 3968
rect 5040 4024 5104 4028
rect 5040 3968 5044 4024
rect 5044 3968 5100 4024
rect 5100 3968 5104 4024
rect 5040 3964 5104 3968
rect 5120 4024 5184 4028
rect 5120 3968 5124 4024
rect 5124 3968 5180 4024
rect 5180 3968 5184 4024
rect 5120 3964 5184 3968
rect 5200 4024 5264 4028
rect 5200 3968 5204 4024
rect 5204 3968 5260 4024
rect 5260 3968 5264 4024
rect 5200 3964 5264 3968
rect 5280 4024 5344 4028
rect 5280 3968 5284 4024
rect 5284 3968 5340 4024
rect 5340 3968 5344 4024
rect 5280 3964 5344 3968
rect 10960 4024 11024 4028
rect 10960 3968 10964 4024
rect 10964 3968 11020 4024
rect 11020 3968 11024 4024
rect 10960 3964 11024 3968
rect 11040 4024 11104 4028
rect 11040 3968 11044 4024
rect 11044 3968 11100 4024
rect 11100 3968 11104 4024
rect 11040 3964 11104 3968
rect 11120 4024 11184 4028
rect 11120 3968 11124 4024
rect 11124 3968 11180 4024
rect 11180 3968 11184 4024
rect 11120 3964 11184 3968
rect 11200 4024 11264 4028
rect 11200 3968 11204 4024
rect 11204 3968 11260 4024
rect 11260 3968 11264 4024
rect 11200 3964 11264 3968
rect 11280 4024 11344 4028
rect 11280 3968 11284 4024
rect 11284 3968 11340 4024
rect 11340 3968 11344 4024
rect 11280 3964 11344 3968
rect 1960 3358 2024 3362
rect 1960 3302 1964 3358
rect 1964 3302 2020 3358
rect 2020 3302 2024 3358
rect 1960 3298 2024 3302
rect 2040 3358 2104 3362
rect 2040 3302 2044 3358
rect 2044 3302 2100 3358
rect 2100 3302 2104 3358
rect 2040 3298 2104 3302
rect 2120 3358 2184 3362
rect 2120 3302 2124 3358
rect 2124 3302 2180 3358
rect 2180 3302 2184 3358
rect 2120 3298 2184 3302
rect 2200 3358 2264 3362
rect 2200 3302 2204 3358
rect 2204 3302 2260 3358
rect 2260 3302 2264 3358
rect 2200 3298 2264 3302
rect 2280 3358 2344 3362
rect 2280 3302 2284 3358
rect 2284 3302 2340 3358
rect 2340 3302 2344 3358
rect 2280 3298 2344 3302
rect 7960 3358 8024 3362
rect 7960 3302 7964 3358
rect 7964 3302 8020 3358
rect 8020 3302 8024 3358
rect 7960 3298 8024 3302
rect 8040 3358 8104 3362
rect 8040 3302 8044 3358
rect 8044 3302 8100 3358
rect 8100 3302 8104 3358
rect 8040 3298 8104 3302
rect 8120 3358 8184 3362
rect 8120 3302 8124 3358
rect 8124 3302 8180 3358
rect 8180 3302 8184 3358
rect 8120 3298 8184 3302
rect 8200 3358 8264 3362
rect 8200 3302 8204 3358
rect 8204 3302 8260 3358
rect 8260 3302 8264 3358
rect 8200 3298 8264 3302
rect 8280 3358 8344 3362
rect 8280 3302 8284 3358
rect 8284 3302 8340 3358
rect 8340 3302 8344 3358
rect 8280 3298 8344 3302
rect 4960 2692 5024 2696
rect 4960 2636 4964 2692
rect 4964 2636 5020 2692
rect 5020 2636 5024 2692
rect 4960 2632 5024 2636
rect 5040 2692 5104 2696
rect 5040 2636 5044 2692
rect 5044 2636 5100 2692
rect 5100 2636 5104 2692
rect 5040 2632 5104 2636
rect 5120 2692 5184 2696
rect 5120 2636 5124 2692
rect 5124 2636 5180 2692
rect 5180 2636 5184 2692
rect 5120 2632 5184 2636
rect 5200 2692 5264 2696
rect 5200 2636 5204 2692
rect 5204 2636 5260 2692
rect 5260 2636 5264 2692
rect 5200 2632 5264 2636
rect 5280 2692 5344 2696
rect 5280 2636 5284 2692
rect 5284 2636 5340 2692
rect 5340 2636 5344 2692
rect 5280 2632 5344 2636
rect 10960 2692 11024 2696
rect 10960 2636 10964 2692
rect 10964 2636 11020 2692
rect 11020 2636 11024 2692
rect 10960 2632 11024 2636
rect 11040 2692 11104 2696
rect 11040 2636 11044 2692
rect 11044 2636 11100 2692
rect 11100 2636 11104 2692
rect 11040 2632 11104 2636
rect 11120 2692 11184 2696
rect 11120 2636 11124 2692
rect 11124 2636 11180 2692
rect 11180 2636 11184 2692
rect 11120 2632 11184 2636
rect 11200 2692 11264 2696
rect 11200 2636 11204 2692
rect 11204 2636 11260 2692
rect 11260 2636 11264 2692
rect 11200 2632 11264 2636
rect 11280 2692 11344 2696
rect 11280 2636 11284 2692
rect 11284 2636 11340 2692
rect 11340 2636 11344 2692
rect 11280 2632 11344 2636
<< metal4 >>
rect 1952 14018 2352 14700
rect 1952 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2352 14018
rect 1952 12686 2352 13954
rect 1952 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2352 12686
rect 1952 11354 2352 12622
rect 1952 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2352 11354
rect 1952 10022 2352 11290
rect 1952 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2352 10022
rect 1952 8690 2352 9958
rect 1952 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2352 8690
rect 1952 7358 2352 8626
rect 1952 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2352 7358
rect 1952 6026 2352 7294
rect 1952 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2352 6026
rect 1952 4694 2352 5962
rect 1952 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2352 4694
rect 1952 3362 2352 4630
rect 1952 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2352 3362
rect 1952 2616 2352 3298
rect 4952 14684 5352 14700
rect 4952 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5352 14684
rect 4952 13352 5352 14620
rect 4952 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5352 13352
rect 4952 12020 5352 13288
rect 4952 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5352 12020
rect 4952 10688 5352 11956
rect 4952 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5352 10688
rect 4952 9356 5352 10624
rect 4952 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5352 9356
rect 4952 8024 5352 9292
rect 4952 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5352 8024
rect 4952 6692 5352 7960
rect 4952 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5352 6692
rect 4952 5360 5352 6628
rect 4952 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5352 5360
rect 4952 4028 5352 5296
rect 4952 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5352 4028
rect 4952 2696 5352 3964
rect 4952 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5352 2696
rect 4952 2616 5352 2632
rect 7952 14018 8352 14700
rect 7952 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8352 14018
rect 7952 12686 8352 13954
rect 7952 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8352 12686
rect 7952 11354 8352 12622
rect 7952 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8352 11354
rect 7952 10022 8352 11290
rect 7952 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8352 10022
rect 7952 8690 8352 9958
rect 7952 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8352 8690
rect 7952 7358 8352 8626
rect 7952 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8352 7358
rect 7952 6026 8352 7294
rect 7952 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8352 6026
rect 7952 4694 8352 5962
rect 7952 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8352 4694
rect 7952 3362 8352 4630
rect 7952 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8352 3362
rect 7952 2616 8352 3298
rect 10952 14684 11352 14700
rect 10952 14620 10960 14684
rect 11024 14620 11040 14684
rect 11104 14620 11120 14684
rect 11184 14620 11200 14684
rect 11264 14620 11280 14684
rect 11344 14620 11352 14684
rect 10952 13352 11352 14620
rect 10952 13288 10960 13352
rect 11024 13288 11040 13352
rect 11104 13288 11120 13352
rect 11184 13288 11200 13352
rect 11264 13288 11280 13352
rect 11344 13288 11352 13352
rect 10952 12020 11352 13288
rect 10952 11956 10960 12020
rect 11024 11956 11040 12020
rect 11104 11956 11120 12020
rect 11184 11956 11200 12020
rect 11264 11956 11280 12020
rect 11344 11956 11352 12020
rect 10952 10688 11352 11956
rect 10952 10624 10960 10688
rect 11024 10624 11040 10688
rect 11104 10624 11120 10688
rect 11184 10624 11200 10688
rect 11264 10624 11280 10688
rect 11344 10624 11352 10688
rect 10952 9356 11352 10624
rect 10952 9292 10960 9356
rect 11024 9292 11040 9356
rect 11104 9292 11120 9356
rect 11184 9292 11200 9356
rect 11264 9292 11280 9356
rect 11344 9292 11352 9356
rect 10952 8024 11352 9292
rect 10952 7960 10960 8024
rect 11024 7960 11040 8024
rect 11104 7960 11120 8024
rect 11184 7960 11200 8024
rect 11264 7960 11280 8024
rect 11344 7960 11352 8024
rect 10952 6692 11352 7960
rect 10952 6628 10960 6692
rect 11024 6628 11040 6692
rect 11104 6628 11120 6692
rect 11184 6628 11200 6692
rect 11264 6628 11280 6692
rect 11344 6628 11352 6692
rect 10952 5360 11352 6628
rect 10952 5296 10960 5360
rect 11024 5296 11040 5360
rect 11104 5296 11120 5360
rect 11184 5296 11200 5360
rect 11264 5296 11280 5360
rect 11344 5296 11352 5360
rect 10952 4028 11352 5296
rect 10952 3964 10960 4028
rect 11024 3964 11040 4028
rect 11104 3964 11120 4028
rect 11184 3964 11200 4028
rect 11264 3964 11280 4028
rect 11344 3964 11352 4028
rect 10952 2696 11352 3964
rect 10952 2632 10960 2696
rect 11024 2632 11040 2696
rect 11104 2632 11120 2696
rect 11184 2632 11200 2696
rect 11264 2632 11280 2696
rect 11344 2632 11352 2696
rect 10952 2616 11352 2632
use sky130_fd_sc_hs__and2_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 11616 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 12576 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__and4bb_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 2304 0 -1 9324
box -38 -49 998 715
use sky130_fd_sc_hs__mux2_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 2880 0 1 5328
box -38 -49 902 715
use sky130_fd_sc_hs__or2b_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 5280 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__clkbuf_1  _24_
timestamp 1723858470
transform -1 0 2592 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 5376 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  _26_
timestamp 1723858470
transform 1 0 3552 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _27_
timestamp 1723858470
transform -1 0 5664 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nand2b_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 4608 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_1  _29_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 5568 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__or2_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 4320 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 1632 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__and3_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 3552 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_1  _33_
timestamp 1723858470
transform -1 0 4992 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  _34_
timestamp 1723858470
transform -1 0 2688 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__nor2_1  _35_
timestamp 1723858470
transform 1 0 1536 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand3_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 6912 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__xor2_1  _37_
timestamp 1723858470
transform 1 0 3840 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__nor2_1  _38_
timestamp 1723858470
transform 1 0 1824 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__dfxtp_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 1824 0 -1 6660
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _40_
timestamp 1723858470
transform 1 0 4032 0 -1 6660
box -38 -49 1670 715
use sky130_fd_sc_hs__dfrtp_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 4128 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _42_
timestamp 1723858470
transform -1 0 8640 0 1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _43_
timestamp 1723858470
transform 1 0 8256 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _44_
timestamp 1723858470
transform 1 0 9024 0 1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _45_
timestamp 1723858470
transform 1 0 8064 0 -1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _46_
timestamp 1723858470
transform -1 0 7872 0 1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _47_
timestamp 1723858470
transform -1 0 6720 0 1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _48_
timestamp 1723858470
transform 1 0 6720 0 1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _49_
timestamp 1723858470
transform 1 0 9024 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _50_
timestamp 1723858470
transform 1 0 5184 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfxtp_1  _51_
timestamp 1723858470
transform 1 0 3840 0 1 7992
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _52_
timestamp 1723858470
transform -1 0 4416 0 -1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _53_
timestamp 1723858470
transform 1 0 1920 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _54_
timestamp 1723858470
transform 1 0 2112 0 1 7992
box -38 -49 1670 715
use sky130_fd_sc_hs__dfrtp_1  _55_
timestamp 1723858470
transform -1 0 6336 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _56_
timestamp 1723858470
transform 1 0 8352 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _57_
timestamp 1723858470
transform 1 0 7008 0 -1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _58_
timestamp 1723858470
transform -1 0 7680 0 1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _59_
timestamp 1723858470
transform -1 0 7776 0 1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _60_
timestamp 1723858470
transform 1 0 7776 0 -1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _61_
timestamp 1723858470
transform -1 0 11136 0 -1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _62_
timestamp 1723858470
transform -1 0 11232 0 1 2664
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _63_
timestamp 1723858470
transform -1 0 8640 0 1 2664
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _64_
timestamp 1723858470
transform -1 0 11520 0 -1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _65_
timestamp 1723858470
transform 1 0 10464 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _66_
timestamp 1723858470
transform 1 0 10464 0 1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _67_
timestamp 1723858470
transform 1 0 10464 0 1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _68_
timestamp 1723858470
transform 1 0 9312 0 -1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _69_
timestamp 1723858470
transform 1 0 10464 0 1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _70_
timestamp 1723858470
transform 1 0 10464 0 1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _71_
timestamp 1723858470
transform -1 0 6432 0 1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _72_
timestamp 1723858470
transform 1 0 6720 0 -1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _73_
timestamp 1723858470
transform 1 0 9024 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _74_
timestamp 1723858470
transform -1 0 10176 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _75_
timestamp 1723858470
transform -1 0 8928 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _76_
timestamp 1723858470
transform 1 0 5760 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _77_
timestamp 1723858470
transform 1 0 4128 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _78_
timestamp 1723858470
transform -1 0 6048 0 -1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _79_
timestamp 1723858470
transform -1 0 4128 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _80_
timestamp 1723858470
transform -1 0 3744 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _81_
timestamp 1723858470
transform -1 0 3744 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_0_CLK $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 5280 0 -1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1723858470
transform -1 0 3456 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1723858470
transform -1 0 3456 0 1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__buf_1  fanout1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 6816 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  fanout2
timestamp 1723858470
transform 1 0 9792 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  fanout44 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 5376 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  fanout45
timestamp 1723858470
transform -1 0 8352 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__buf_2  fanout46 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 6144 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  fanout47
timestamp 1723858470
transform -1 0 7008 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_4  fanout48 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform -1 0 9696 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__buf_2  fanout49
timestamp 1723858470
transform -1 0 8928 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__buf_1  fanout50
timestamp 1723858470
transform -1 0 12096 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__buf_1  fanout51
timestamp 1723858470
transform 1 0 4896 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__buf_2  fanout52
timestamp 1723858470
transform 1 0 8256 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  fanout53
timestamp 1723858470
transform -1 0 9792 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  fanout54
timestamp 1723858470
transform -1 0 6912 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  fanout55
timestamp 1723858470
transform -1 0 5664 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  fanout56
timestamp 1723858470
transform 1 0 3840 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  fanout57
timestamp 1723858470
transform 1 0 4512 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__buf_2  fanout58
timestamp 1723858470
transform 1 0 3840 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  fanout59
timestamp 1723858470
transform -1 0 3168 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_2  fanout60
timestamp 1723858470
transform -1 0 2016 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  fanout61
timestamp 1723858470
transform -1 0 10848 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  fanout62
timestamp 1723858470
transform -1 0 8352 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_4 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 1536 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 2208 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_19
timestamp 1723858470
transform 1 0 2976 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 3840 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 4224 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_38
timestamp 1723858470
transform 1 0 4800 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_46
timestamp 1723858470
transform 1 0 5568 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_78
timestamp 1723858470
transform 1 0 8640 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_80
timestamp 1723858470
transform 1 0 8832 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_105
timestamp 1723858470
transform 1 0 11232 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_107
timestamp 1723858470
transform 1 0 11424 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_113
timestamp 1723858470
transform 1 0 12000 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_4
timestamp 1723858470
transform 1 0 1536 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_12
timestamp 1723858470
transform 1 0 2304 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_20
timestamp 1723858470
transform 1 0 3072 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_1_28
timestamp 1723858470
transform 1 0 3840 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_30
timestamp 1723858470
transform 1 0 4032 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_1_59
timestamp 1723858470
transform 1 0 6816 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_61
timestamp 1723858470
transform 1 0 7008 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_101
timestamp 1723858470
transform 1 0 10848 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_1_109
timestamp 1723858470
transform 1 0 11616 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_113
timestamp 1723858470
transform 1 0 12000 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_4
timestamp 1723858470
transform 1 0 1536 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_12
timestamp 1723858470
transform 1 0 2304 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_2_20
timestamp 1723858470
transform 1 0 3072 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_24
timestamp 1723858470
transform 1 0 3456 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_26
timestamp 1723858470
transform 1 0 3648 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_78
timestamp 1723858470
transform 1 0 8640 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_80
timestamp 1723858470
transform 1 0 8832 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_82
timestamp 1723858470
transform 1 0 9024 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_84
timestamp 1723858470
transform 1 0 9216 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_4
timestamp 1723858470
transform 1 0 1536 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_12
timestamp 1723858470
transform 1 0 2304 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_20
timestamp 1723858470
transform 1 0 3072 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_3_28
timestamp 1723858470
transform 1 0 3840 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_32
timestamp 1723858470
transform 1 0 4224 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_34
timestamp 1723858470
transform 1 0 4416 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_52
timestamp 1723858470
transform 1 0 6144 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_55
timestamp 1723858470
transform 1 0 6432 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6624 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_3_104
timestamp 1723858470
transform 1 0 11136 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_3_109
timestamp 1723858470
transform 1 0 11616 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_113
timestamp 1723858470
transform 1 0 12000 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_4
timestamp 1723858470
transform 1 0 1536 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_8
timestamp 1723858470
transform 1 0 1920 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_10
timestamp 1723858470
transform 1 0 2112 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_15
timestamp 1723858470
transform 1 0 2592 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_17
timestamp 1723858470
transform 1 0 2784 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_28
timestamp 1723858470
transform 1 0 3840 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_44
timestamp 1723858470
transform 1 0 5376 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_4_68
timestamp 1723858470
transform 1 0 7680 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_76
timestamp 1723858470
transform 1 0 8448 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_80
timestamp 1723858470
transform 1 0 8832 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_82
timestamp 1723858470
transform 1 0 9024 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_89
timestamp 1723858470
transform 1 0 9696 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_4
timestamp 1723858470
transform 1 0 1536 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_6
timestamp 1723858470
transform 1 0 1728 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_24
timestamp 1723858470
transform 1 0 3456 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_5_47
timestamp 1723858470
transform 1 0 5664 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_51
timestamp 1723858470
transform 1 0 6048 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_53
timestamp 1723858470
transform 1 0 6240 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_55
timestamp 1723858470
transform 1 0 6432 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_5_63
timestamp 1723858470
transform 1 0 7200 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_67
timestamp 1723858470
transform 1 0 7584 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_92
timestamp 1723858470
transform 1 0 9984 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_100
timestamp 1723858470
transform 1 0 10752 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_109
timestamp 1723858470
transform 1 0 11616 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_6_24
timestamp 1723858470
transform 1 0 3456 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_6_26
timestamp 1723858470
transform 1 0 3648 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_6_70
timestamp 1723858470
transform 1 0 7872 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_6_74
timestamp 1723858470
transform 1 0 8256 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_6_105
timestamp 1723858470
transform 1 0 11232 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_6_107
timestamp 1723858470
transform 1 0 11424 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_4
timestamp 1723858470
transform 1 0 1536 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_8
timestamp 1723858470
transform 1 0 1920 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_14
timestamp 1723858470
transform 1 0 2496 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_26
timestamp 1723858470
transform 1 0 3648 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_32
timestamp 1723858470
transform 1 0 4224 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_41
timestamp 1723858470
transform 1 0 5088 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_49
timestamp 1723858470
transform 1 0 5856 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_53
timestamp 1723858470
transform 1 0 6240 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 6432 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_61
timestamp 1723858470
transform 1 0 7008 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_69
timestamp 1723858470
transform 1 0 7776 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_71
timestamp 1723858470
transform 1 0 7968 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_95
timestamp 1723858470
transform 1 0 10272 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_99
timestamp 1723858470
transform 1 0 10656 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_101
timestamp 1723858470
transform 1 0 10848 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_109
timestamp 1723858470
transform 1 0 11616 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_113
timestamp 1723858470
transform 1 0 12000 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_8_45
timestamp 1723858470
transform 1 0 5472 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_69
timestamp 1723858470
transform 1 0 7776 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_8_77
timestamp 1723858470
transform 1 0 8544 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_82
timestamp 1723858470
transform 1 0 9024 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_8_90
timestamp 1723858470
transform 1 0 9792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_8_94
timestamp 1723858470
transform 1 0 10176 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_8_96
timestamp 1723858470
transform 1 0 10368 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_9_4
timestamp 1723858470
transform 1 0 1536 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_9_22
timestamp 1723858470
transform 1 0 3264 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_9_60
timestamp 1723858470
transform 1 0 6912 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_9_84
timestamp 1723858470
transform 1 0 9216 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_9_109
timestamp 1723858470
transform 1 0 11616 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_9_113
timestamp 1723858470
transform 1 0 12000 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_24
timestamp 1723858470
transform 1 0 3456 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_26
timestamp 1723858470
transform 1 0 3648 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_33
timestamp 1723858470
transform 1 0 4320 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_82
timestamp 1723858470
transform 1 0 9024 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_84
timestamp 1723858470
transform 1 0 9216 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_94
timestamp 1723858470
transform 1 0 10176 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_96
timestamp 1723858470
transform 1 0 10368 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_4
timestamp 1723858470
transform 1 0 1536 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_60
timestamp 1723858470
transform 1 0 6912 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_68
timestamp 1723858470
transform 1 0 7680 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_70
timestamp 1723858470
transform 1 0 7872 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_98
timestamp 1723858470
transform 1 0 10560 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_106
timestamp 1723858470
transform 1 0 11328 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_109
timestamp 1723858470
transform 1 0 11616 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_113
timestamp 1723858470
transform 1 0 12000 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_4
timestamp 1723858470
transform 1 0 1536 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_12_16
timestamp 1723858470
transform 1 0 2688 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_24
timestamp 1723858470
transform 1 0 3456 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_26
timestamp 1723858470
transform 1 0 3648 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_12_28
timestamp 1723858470
transform 1 0 3840 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_40
timestamp 1723858470
transform 1 0 4992 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_12_65
timestamp 1723858470
transform 1 0 7392 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_73
timestamp 1723858470
transform 1 0 8160 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_79
timestamp 1723858470
transform 1 0 8736 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_105
timestamp 1723858470
transform 1 0 11232 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_107
timestamp 1723858470
transform 1 0 11424 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_4
timestamp 1723858470
transform 1 0 1536 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_13_12
timestamp 1723858470
transform 1 0 2304 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_34
timestamp 1723858470
transform 1 0 4416 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_42
timestamp 1723858470
transform 1 0 5184 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_13_50
timestamp 1723858470
transform 1 0 5952 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_55
timestamp 1723858470
transform 1 0 6432 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_63
timestamp 1723858470
transform 1 0 7200 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_71
timestamp 1723858470
transform 1 0 7968 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_13_79
timestamp 1723858470
transform 1 0 8736 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_13_83
timestamp 1723858470
transform 1 0 9120 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_13_109
timestamp 1723858470
transform 1 0 11616 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_13_113
timestamp 1723858470
transform 1 0 12000 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_28
timestamp 1723858470
transform 1 0 3840 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_36
timestamp 1723858470
transform 1 0 4608 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_44
timestamp 1723858470
transform 1 0 5376 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_14_52
timestamp 1723858470
transform 1 0 6144 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_14_56
timestamp 1723858470
transform 1 0 6528 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_82
timestamp 1723858470
transform 1 0 9024 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_14_90
timestamp 1723858470
transform 1 0 9792 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_55
timestamp 1723858470
transform 1 0 6432 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_63
timestamp 1723858470
transform 1 0 7200 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_94
timestamp 1723858470
transform 1 0 10176 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_16_39
timestamp 1723858470
transform 1 0 4896 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_43
timestamp 1723858470
transform 1 0 5280 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_16_105
timestamp 1723858470
transform 1 0 11232 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_107
timestamp 1723858470
transform 1 0 11424 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_4
timestamp 1723858470
transform 1 0 1536 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_15
timestamp 1723858470
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_51
timestamp 1723858470
transform 1 0 6048 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_53
timestamp 1723858470
transform 1 0 6240 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_55
timestamp 1723858470
transform 1 0 6432 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_17_88
timestamp 1723858470
transform 1 0 9600 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_92
timestamp 1723858470
transform 1 0 9984 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_99
timestamp 1723858470
transform 1 0 10656 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_101
timestamp 1723858470
transform 1 0 10848 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_119
timestamp 1723858470
transform 1 0 12576 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd2_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 5568 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__clkbuf_1  hold2
timestamp 1723858470
transform -1 0 5856 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold3
timestamp 1723858470
transform -1 0 4224 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold4
timestamp 1723858470
transform -1 0 2304 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold5
timestamp 1723858470
transform -1 0 3648 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold6
timestamp 1723858470
transform -1 0 4608 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold7
timestamp 1723858470
transform -1 0 2784 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold8
timestamp 1723858470
transform 1 0 2112 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold9
timestamp 1723858470
transform -1 0 4608 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  hold10
timestamp 1723858470
transform -1 0 3456 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  input1
timestamp 1723858470
transform 1 0 5952 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  input2
timestamp 1723858470
transform -1 0 12000 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  input3
timestamp 1723858470
transform 1 0 1536 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  input4
timestamp 1723858470
transform 1 0 4416 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_4  output5
timestamp 1723858470
transform -1 0 12672 0 -1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output6
timestamp 1723858470
transform -1 0 12096 0 1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output7
timestamp 1723858470
transform -1 0 11520 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output8
timestamp 1723858470
transform -1 0 12672 0 1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output9
timestamp 1723858470
transform -1 0 12672 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output10
timestamp 1723858470
transform -1 0 12672 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output11
timestamp 1723858470
transform -1 0 12672 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output12
timestamp 1723858470
transform -1 0 12096 0 1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output13
timestamp 1723858470
transform -1 0 12672 0 -1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output14
timestamp 1723858470
transform 1 0 10944 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output15
timestamp 1723858470
transform -1 0 9888 0 1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output16
timestamp 1723858470
transform 1 0 1632 0 1 2664
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output17
timestamp 1723858470
transform -1 0 2592 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output18
timestamp 1723858470
transform -1 0 3744 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output19
timestamp 1723858470
transform -1 0 4896 0 1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output20
timestamp 1723858470
transform -1 0 7776 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output21
timestamp 1723858470
transform -1 0 7200 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output22
timestamp 1723858470
transform -1 0 8352 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output23
timestamp 1723858470
transform -1 0 9600 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output24
timestamp 1723858470
transform -1 0 10656 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output25
timestamp 1723858470
transform -1 0 12192 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output26
timestamp 1723858470
transform -1 0 12672 0 1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output27
timestamp 1723858470
transform -1 0 12672 0 -1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output28
timestamp 1723858470
transform 1 0 12096 0 1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output29
timestamp 1723858470
transform 1 0 11520 0 1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output30
timestamp 1723858470
transform 1 0 10944 0 -1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output31
timestamp 1723858470
transform 1 0 10368 0 -1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output32
timestamp 1723858470
transform 1 0 8352 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output33
timestamp 1723858470
transform 1 0 9888 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output34
timestamp 1723858470
transform 1 0 8352 0 1 13320
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output35
timestamp 1723858470
transform -1 0 8256 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output36
timestamp 1723858470
transform -1 0 10464 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output37
timestamp 1723858470
transform -1 0 7680 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output38
timestamp 1723858470
transform -1 0 10464 0 1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output39
timestamp 1723858470
transform -1 0 11520 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output40
timestamp 1723858470
transform -1 0 12672 0 1 2664
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output41
timestamp 1723858470
transform -1 0 12672 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output42
timestamp 1723858470
transform -1 0 12672 0 -1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  output43
timestamp 1723858470
transform -1 0 11520 0 -1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__decap_4  PHY_0
timestamp 1723858470
transform 1 0 1152 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_1
timestamp 1723858470
transform -1 0 13056 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_2
timestamp 1723858470
transform 1 0 1152 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_3
timestamp 1723858470
transform -1 0 13056 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_4
timestamp 1723858470
transform 1 0 1152 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_5
timestamp 1723858470
transform -1 0 13056 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_6
timestamp 1723858470
transform 1 0 1152 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_7
timestamp 1723858470
transform -1 0 13056 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_8
timestamp 1723858470
transform 1 0 1152 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_9
timestamp 1723858470
transform -1 0 13056 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_10
timestamp 1723858470
transform 1 0 1152 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_11
timestamp 1723858470
transform -1 0 13056 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_12
timestamp 1723858470
transform 1 0 1152 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_13
timestamp 1723858470
transform -1 0 13056 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_14
timestamp 1723858470
transform 1 0 1152 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_15
timestamp 1723858470
transform -1 0 13056 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_16
timestamp 1723858470
transform 1 0 1152 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_17
timestamp 1723858470
transform -1 0 13056 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_18
timestamp 1723858470
transform 1 0 1152 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_19
timestamp 1723858470
transform -1 0 13056 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_20
timestamp 1723858470
transform 1 0 1152 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_21
timestamp 1723858470
transform -1 0 13056 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_22
timestamp 1723858470
transform 1 0 1152 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_23
timestamp 1723858470
transform -1 0 13056 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_24
timestamp 1723858470
transform 1 0 1152 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_25
timestamp 1723858470
transform -1 0 13056 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_26
timestamp 1723858470
transform 1 0 1152 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_27
timestamp 1723858470
transform -1 0 13056 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_28
timestamp 1723858470
transform 1 0 1152 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_29
timestamp 1723858470
transform -1 0 13056 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_30
timestamp 1723858470
transform 1 0 1152 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_31
timestamp 1723858470
transform -1 0 13056 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_32
timestamp 1723858470
transform 1 0 1152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_33
timestamp 1723858470
transform -1 0 13056 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_34
timestamp 1723858470
transform 1 0 1152 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_35
timestamp 1723858470
transform -1 0 13056 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_36 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1723858470
transform 1 0 3744 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_37
timestamp 1723858470
transform 1 0 6336 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_38
timestamp 1723858470
transform 1 0 8928 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_39
timestamp 1723858470
transform 1 0 11520 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_40
timestamp 1723858470
transform 1 0 6336 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_41
timestamp 1723858470
transform 1 0 11520 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_42
timestamp 1723858470
transform 1 0 3744 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_43
timestamp 1723858470
transform 1 0 8928 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_44
timestamp 1723858470
transform 1 0 6336 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_45
timestamp 1723858470
transform 1 0 11520 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_46
timestamp 1723858470
transform 1 0 3744 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_47
timestamp 1723858470
transform 1 0 8928 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_48
timestamp 1723858470
transform 1 0 6336 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_49
timestamp 1723858470
transform 1 0 11520 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_50
timestamp 1723858470
transform 1 0 3744 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_51
timestamp 1723858470
transform 1 0 8928 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_52
timestamp 1723858470
transform 1 0 6336 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_53
timestamp 1723858470
transform 1 0 11520 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_54
timestamp 1723858470
transform 1 0 3744 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_55
timestamp 1723858470
transform 1 0 8928 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_56
timestamp 1723858470
transform 1 0 6336 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_57
timestamp 1723858470
transform 1 0 11520 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_58
timestamp 1723858470
transform 1 0 3744 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_59
timestamp 1723858470
transform 1 0 8928 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_60
timestamp 1723858470
transform 1 0 6336 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_61
timestamp 1723858470
transform 1 0 11520 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_62
timestamp 1723858470
transform 1 0 3744 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_63
timestamp 1723858470
transform 1 0 8928 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_64
timestamp 1723858470
transform 1 0 6336 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_65
timestamp 1723858470
transform 1 0 11520 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_66
timestamp 1723858470
transform 1 0 3744 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_67
timestamp 1723858470
transform 1 0 8928 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_68
timestamp 1723858470
transform 1 0 6336 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_69
timestamp 1723858470
transform 1 0 11520 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_70
timestamp 1723858470
transform 1 0 3744 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_71
timestamp 1723858470
transform 1 0 8928 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_72
timestamp 1723858470
transform 1 0 3744 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_73
timestamp 1723858470
transform 1 0 6336 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_74
timestamp 1723858470
transform 1 0 8928 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_75
timestamp 1723858470
transform 1 0 11520 0 -1 14652
box -38 -49 134 715
<< labels >>
flabel metal3 s 13498 6230 14298 6350 0 FreeSans 480 0 0 0 CF[0]
port 0 nsew signal tristate
flabel metal3 s 13498 6822 14298 6942 0 FreeSans 480 0 0 0 CF[1]
port 1 nsew signal tristate
flabel metal3 s 13498 7414 14298 7534 0 FreeSans 480 0 0 0 CF[2]
port 2 nsew signal tristate
flabel metal3 s 13498 8006 14298 8126 0 FreeSans 480 0 0 0 CF[3]
port 3 nsew signal tristate
flabel metal3 s 13498 8598 14298 8718 0 FreeSans 480 0 0 0 CF[4]
port 4 nsew signal tristate
flabel metal3 s 13498 9190 14298 9310 0 FreeSans 480 0 0 0 CF[5]
port 5 nsew signal tristate
flabel metal3 s 13498 9782 14298 9902 0 FreeSans 480 0 0 0 CF[6]
port 6 nsew signal tristate
flabel metal3 s 13498 10374 14298 10494 0 FreeSans 480 0 0 0 CF[7]
port 7 nsew signal tristate
flabel metal3 s 13498 10966 14298 11086 0 FreeSans 480 0 0 0 CF[8]
port 8 nsew signal tristate
flabel metal2 s 12308 16522 12364 17322 0 FreeSans 224 90 0 0 CKO
port 9 nsew signal tristate
flabel metal2 s 12692 0 12748 800 0 FreeSans 224 90 0 0 CKS
port 10 nsew signal tristate
flabel metal2 s 1556 0 1612 800 0 FreeSans 224 90 0 0 CKSB
port 11 nsew signal tristate
flabel metal2 s 13460 16522 13516 17322 0 FreeSans 224 90 0 0 CLK
port 12 nsew signal input
flabel metal2 s 7124 0 7180 800 0 FreeSans 224 90 0 0 CMP_N
port 13 nsew signal input
flabel metal2 s 9908 0 9964 800 0 FreeSans 224 90 0 0 CMP_P
port 14 nsew signal input
flabel metal2 s 1940 16522 1996 17322 0 FreeSans 224 90 0 0 DATA[0]
port 15 nsew signal tristate
flabel metal2 s 3092 16522 3148 17322 0 FreeSans 224 90 0 0 DATA[1]
port 16 nsew signal tristate
flabel metal2 s 4244 16522 4300 17322 0 FreeSans 224 90 0 0 DATA[2]
port 17 nsew signal tristate
flabel metal2 s 5396 16522 5452 17322 0 FreeSans 224 90 0 0 DATA[3]
port 18 nsew signal tristate
flabel metal2 s 6548 16522 6604 17322 0 FreeSans 224 90 0 0 DATA[4]
port 19 nsew signal tristate
flabel metal2 s 7700 16522 7756 17322 0 FreeSans 224 90 0 0 DATA[5]
port 20 nsew signal tristate
flabel metal2 s 8852 16522 8908 17322 0 FreeSans 224 90 0 0 DATA[6]
port 21 nsew signal tristate
flabel metal2 s 10004 16522 10060 17322 0 FreeSans 224 90 0 0 DATA[7]
port 22 nsew signal tristate
flabel metal2 s 11156 16522 11212 17322 0 FreeSans 224 90 0 0 DATA[8]
port 23 nsew signal tristate
flabel metal2 s 788 16522 844 17322 0 FreeSans 224 90 0 0 EN
port 24 nsew signal input
flabel metal2 s 4340 0 4396 800 0 FreeSans 224 90 0 0 RDY
port 25 nsew signal input
flabel metal3 s 13498 11558 14298 11678 0 FreeSans 480 0 0 0 SWN[0]
port 26 nsew signal tristate
flabel metal3 s 13498 12150 14298 12270 0 FreeSans 480 0 0 0 SWN[1]
port 27 nsew signal tristate
flabel metal3 s 13498 12742 14298 12862 0 FreeSans 480 0 0 0 SWN[2]
port 28 nsew signal tristate
flabel metal3 s 13498 13334 14298 13454 0 FreeSans 480 0 0 0 SWN[3]
port 29 nsew signal tristate
flabel metal3 s 13498 13926 14298 14046 0 FreeSans 480 0 0 0 SWN[4]
port 30 nsew signal tristate
flabel metal3 s 13498 14518 14298 14638 0 FreeSans 480 0 0 0 SWN[5]
port 31 nsew signal tristate
flabel metal3 s 13498 15110 14298 15230 0 FreeSans 480 0 0 0 SWN[6]
port 32 nsew signal tristate
flabel metal3 s 13498 15702 14298 15822 0 FreeSans 480 0 0 0 SWN[7]
port 33 nsew signal tristate
flabel metal3 s 13498 16294 14298 16414 0 FreeSans 480 0 0 0 SWN[8]
port 34 nsew signal tristate
flabel metal3 s 13498 902 14298 1022 0 FreeSans 480 0 0 0 SWP[0]
port 35 nsew signal tristate
flabel metal3 s 13498 1494 14298 1614 0 FreeSans 480 0 0 0 SWP[1]
port 36 nsew signal tristate
flabel metal3 s 13498 2086 14298 2206 0 FreeSans 480 0 0 0 SWP[2]
port 37 nsew signal tristate
flabel metal3 s 13498 2678 14298 2798 0 FreeSans 480 0 0 0 SWP[3]
port 38 nsew signal tristate
flabel metal3 s 13498 3270 14298 3390 0 FreeSans 480 0 0 0 SWP[4]
port 39 nsew signal tristate
flabel metal3 s 13498 3862 14298 3982 0 FreeSans 480 0 0 0 SWP[5]
port 40 nsew signal tristate
flabel metal3 s 13498 4454 14298 4574 0 FreeSans 480 0 0 0 SWP[6]
port 41 nsew signal tristate
flabel metal3 s 13498 5046 14298 5166 0 FreeSans 480 0 0 0 SWP[7]
port 42 nsew signal tristate
flabel metal3 s 13498 5638 14298 5758 0 FreeSans 480 0 0 0 SWP[8]
port 43 nsew signal tristate
flabel metal4 s 4952 2616 5352 14700 0 FreeSans 1920 90 0 0 VGND
port 44 nsew ground bidirectional
flabel metal4 s 10952 2616 11352 14700 0 FreeSans 1920 90 0 0 VGND
port 44 nsew ground bidirectional
flabel metal4 s 1952 2616 2352 14700 0 FreeSans 1920 90 0 0 VPWR
port 45 nsew power bidirectional
flabel metal4 s 7952 2616 8352 14700 0 FreeSans 1920 90 0 0 VPWR
port 45 nsew power bidirectional
rlabel metal1 7104 14652 7104 14652 0 VGND
rlabel metal1 7104 13986 7104 13986 0 VPWR
rlabel via2 12528 6271 12528 6271 0 CF[0]
rlabel via2 11952 6863 11952 6863 0 CF[1]
rlabel metal1 11856 7585 11856 7585 0 CF[2]
rlabel metal2 12528 7566 12528 7566 0 CF[3]
rlabel metal1 12720 7881 12720 7881 0 CF[4]
rlabel via2 12528 9231 12528 9231 0 CF[5]
rlabel metal2 12528 9971 12528 9971 0 CF[6]
rlabel metal3 12729 10434 12729 10434 0 CF[7]
rlabel metal2 12528 11303 12528 11303 0 CF[8]
rlabel metal1 11568 14245 11568 14245 0 CKO
rlabel metal1 11232 4181 11232 4181 0 CKS
rlabel metal2 1687 666 1687 666 0 CKSB
rlabel metal2 13337 16650 13337 16650 0 CLK
rlabel metal1 6624 2997 6624 2997 0 CMP_N
rlabel metal1 10416 2923 10416 2923 0 CMP_P
rlabel metal1 2112 14171 2112 14171 0 DATA[0]
rlabel metal2 3408 15447 3408 15447 0 DATA[1]
rlabel metal1 4416 13875 4416 13875 0 DATA[2]
rlabel metal2 5712 15484 5712 15484 0 DATA[3]
rlabel metal1 6720 14171 6720 14171 0 DATA[4]
rlabel metal2 8016 15447 8016 15447 0 DATA[5]
rlabel metal1 9072 14171 9072 14171 0 DATA[6]
rlabel metal1 10176 14171 10176 14171 0 DATA[7]
rlabel metal1 11664 14171 11664 14171 0 DATA[8]
rlabel metal1 1200 12987 1200 12987 0 EN
rlabel metal2 4423 666 4423 666 0 RDY
rlabel metal1 12768 11211 12768 11211 0 SWN[0]
rlabel metal2 12528 12487 12528 12487 0 SWN[1]
rlabel metal1 12336 13431 12336 13431 0 SWN[2]
rlabel metal1 11760 13431 11760 13431 0 SWN[3]
rlabel metal1 11712 13135 11712 13135 0 SWN[4]
rlabel metal1 10608 13209 10608 13209 0 SWN[5]
rlabel metal1 8592 14171 8592 14171 0 SWN[6]
rlabel metal3 11721 15762 11721 15762 0 SWN[7]
rlabel metal1 8544 13875 8544 13875 0 SWN[8]
rlabel metal3 11673 962 11673 962 0 SWP[0]
rlabel metal3 11913 1554 11913 1554 0 SWP[1]
rlabel metal3 11769 2146 11769 2146 0 SWP[2]
rlabel metal3 12489 2738 12489 2738 0 SWP[3]
rlabel metal1 11856 3589 11856 3589 0 SWP[4]
rlabel metal2 12528 3570 12528 3570 0 SWP[5]
rlabel metal1 12720 3885 12720 3885 0 SWP[6]
rlabel metal2 12528 5161 12528 5161 0 SWP[7]
rlabel metal2 11376 5901 11376 5901 0 SWP[8]
rlabel metal1 2352 5883 2352 5883 0 _00_
rlabel metal1 4464 6475 4464 6475 0 _01_
rlabel metal2 5808 8214 5808 8214 0 _02_
rlabel metal2 4656 11396 4656 11396 0 _03_
rlabel metal1 1920 7659 1920 7659 0 _04_
rlabel metal1 1968 7807 1968 7807 0 _05_
rlabel metal2 12048 13764 12048 13764 0 _06_
rlabel metal2 4656 8436 4656 8436 0 _07_
rlabel metal1 4080 5513 4080 5513 0 _08_
rlabel metal1 2544 5698 2544 5698 0 _09_
rlabel metal1 4512 5883 4512 5883 0 _10_
rlabel metal2 3984 6734 3984 6734 0 _11_
rlabel metal1 1872 8251 1872 8251 0 _12_
rlabel metal1 3840 9879 3840 9879 0 _13_
rlabel metal1 2352 10915 2352 10915 0 _14_
rlabel metal1 4080 10286 4080 10286 0 _15_
rlabel metal1 2304 11211 2304 11211 0 _16_
rlabel metal1 4368 7030 4368 7030 0 _17_
rlabel metal1 2256 8880 2256 8880 0 _18_
rlabel metal1 5280 9065 5280 9065 0 clk_div_0.COUNT\[0\]
rlabel metal1 2784 11433 2784 11433 0 clk_div_0.COUNT\[1\]
rlabel metal1 3456 10101 3456 10101 0 clk_div_0.COUNT\[2\]
rlabel metal1 3888 7659 3888 7659 0 clk_div_0.COUNT\[3\]
rlabel metal1 3456 9657 3456 9657 0 clknet_0_CLK
rlabel metal1 2304 8325 2304 8325 0 clknet_1_0__leaf_CLK
rlabel metal2 2832 10693 2832 10693 0 clknet_1_1__leaf_CLK
rlabel metal1 7968 13579 7968 13579 0 cyclic_flag_0.FINAL
rlabel metal1 6768 3700 6768 3700 0 net1
rlabel metal1 10944 8325 10944 8325 0 net10
rlabel metal1 10944 9657 10944 9657 0 net11
rlabel metal1 11280 10915 11280 10915 0 net12
rlabel metal1 5856 10323 5856 10323 0 net13
rlabel metal1 11376 14430 11376 14430 0 net14
rlabel metal2 5616 5550 5616 5550 0 net15
rlabel metal2 3408 4514 3408 4514 0 net16
rlabel metal1 1824 12543 1824 12543 0 net17
rlabel metal1 2544 13875 2544 13875 0 net18
rlabel metal1 3264 13209 3264 13209 0 net19
rlabel metal1 10464 3663 10464 3663 0 net2
rlabel metal1 5616 14430 5616 14430 0 net20
rlabel metal1 6480 14393 6480 14393 0 net21
rlabel metal1 7872 13875 7872 13875 0 net22
rlabel metal1 8064 12543 8064 12543 0 net23
rlabel metal1 8736 13209 8736 13209 0 net24
rlabel metal2 11088 14097 11088 14097 0 net25
rlabel metal1 12000 10915 12000 10915 0 net26
rlabel metal2 12240 13010 12240 13010 0 net27
rlabel metal1 12672 13579 12672 13579 0 net28
rlabel metal2 12528 13542 12528 13542 0 net29
rlabel metal1 1824 13209 1824 13209 0 net3
rlabel metal1 11424 13061 11424 13061 0 net30
rlabel metal1 11616 8547 11616 8547 0 net31
rlabel metal1 10176 14541 10176 14541 0 net32
rlabel metal1 10320 12210 10320 12210 0 net33
rlabel metal1 8784 13542 8784 13542 0 net34
rlabel metal2 6576 7733 6576 7733 0 net35
rlabel metal1 3696 13542 3696 13542 0 net36
rlabel metal1 4080 13098 4080 13098 0 net37
rlabel metal1 6600 14245 6600 14245 0 net38
rlabel metal1 4368 12987 4368 12987 0 net39
rlabel metal1 5136 5069 5136 5069 0 net4
rlabel metal2 5808 13269 5808 13269 0 net40
rlabel metal2 9072 6253 9072 6253 0 net41
rlabel metal1 10176 12987 10176 12987 0 net42
rlabel metal1 9024 13579 9024 13579 0 net43
rlabel metal1 5864 13653 5864 13653 0 net44
rlabel metal1 5520 13579 5520 13579 0 net45
rlabel metal2 7248 3737 7248 3737 0 net46
rlabel metal2 6768 8066 6768 8066 0 net47
rlabel metal2 9648 3330 9648 3330 0 net48
rlabel metal1 9360 5587 9360 5587 0 net49
rlabel metal1 8592 4366 8592 4366 0 net5
rlabel metal2 10800 5069 10800 5069 0 net50
rlabel metal1 8496 6956 8496 6956 0 net51
rlabel metal1 11232 13209 11232 13209 0 net52
rlabel metal2 10704 8658 10704 8658 0 net53
rlabel metal2 8592 9287 8592 9287 0 net54
rlabel metal1 5520 5217 5520 5217 0 net55
rlabel metal1 7680 6993 7680 6993 0 net56
rlabel metal1 4608 4921 4608 4921 0 net57
rlabel metal2 4080 13986 4080 13986 0 net58
rlabel metal1 3456 14319 3456 14319 0 net59
rlabel metal2 10800 3108 10800 3108 0 net6
rlabel metal1 5849 13727 5849 13727 0 net60
rlabel metal1 7776 6401 7776 6401 0 net61
rlabel metal1 7104 8917 7104 8917 0 net62
rlabel metal1 1680 10989 1680 10989 0 net63
rlabel metal1 4896 7881 4896 7881 0 net64
rlabel metal1 3456 7585 3456 7585 0 net65
rlabel metal1 2064 8362 2064 8362 0 net66
rlabel metal2 2544 8066 2544 8066 0 net67
rlabel metal1 3456 10915 3456 10915 0 net68
rlabel metal2 1776 9953 1776 9953 0 net69
rlabel metal1 10752 7733 10752 7733 0 net7
rlabel metal1 2400 7881 2400 7881 0 net70
rlabel metal1 3792 5587 3792 5587 0 net71
rlabel metal1 1824 10915 1824 10915 0 net72
rlabel metal2 10512 6993 10512 6993 0 net73
rlabel metal2 10128 9250 10128 9250 0 net74
rlabel metal1 8064 6327 8064 6327 0 net8
rlabel metal1 11184 7807 11184 7807 0 net9
<< properties >>
string FIXED_BBOX 0 0 14298 17322
<< end >>
