magic
tech sky130A
magscale 1 2
timestamp 1757383169
<< metal3 >>
rect -32264 5612 -31492 5640
rect -32264 5188 -31576 5612
rect -31512 5188 -31492 5612
rect -32264 5160 -31492 5188
rect -31252 5612 -30480 5640
rect -31252 5188 -30564 5612
rect -30500 5188 -30480 5612
rect -31252 5160 -30480 5188
rect -30240 5612 -29468 5640
rect -30240 5188 -29552 5612
rect -29488 5188 -29468 5612
rect -30240 5160 -29468 5188
rect -29228 5612 -28456 5640
rect -29228 5188 -28540 5612
rect -28476 5188 -28456 5612
rect -29228 5160 -28456 5188
rect -28216 5612 -27444 5640
rect -28216 5188 -27528 5612
rect -27464 5188 -27444 5612
rect -28216 5160 -27444 5188
rect -27204 5612 -26432 5640
rect -27204 5188 -26516 5612
rect -26452 5188 -26432 5612
rect -27204 5160 -26432 5188
rect -26192 5612 -25420 5640
rect -26192 5188 -25504 5612
rect -25440 5188 -25420 5612
rect -26192 5160 -25420 5188
rect -25180 5612 -24408 5640
rect -25180 5188 -24492 5612
rect -24428 5188 -24408 5612
rect -25180 5160 -24408 5188
rect -24168 5612 -23396 5640
rect -24168 5188 -23480 5612
rect -23416 5188 -23396 5612
rect -24168 5160 -23396 5188
rect -23156 5612 -22384 5640
rect -23156 5188 -22468 5612
rect -22404 5188 -22384 5612
rect -23156 5160 -22384 5188
rect -22144 5612 -21372 5640
rect -22144 5188 -21456 5612
rect -21392 5188 -21372 5612
rect -22144 5160 -21372 5188
rect -21132 5612 -20360 5640
rect -21132 5188 -20444 5612
rect -20380 5188 -20360 5612
rect -21132 5160 -20360 5188
rect -20120 5612 -19348 5640
rect -20120 5188 -19432 5612
rect -19368 5188 -19348 5612
rect -20120 5160 -19348 5188
rect -19108 5612 -18336 5640
rect -19108 5188 -18420 5612
rect -18356 5188 -18336 5612
rect -19108 5160 -18336 5188
rect -18096 5612 -17324 5640
rect -18096 5188 -17408 5612
rect -17344 5188 -17324 5612
rect -18096 5160 -17324 5188
rect -17084 5612 -16312 5640
rect -17084 5188 -16396 5612
rect -16332 5188 -16312 5612
rect -17084 5160 -16312 5188
rect -16072 5612 -15300 5640
rect -16072 5188 -15384 5612
rect -15320 5188 -15300 5612
rect -16072 5160 -15300 5188
rect -15060 5612 -14288 5640
rect -15060 5188 -14372 5612
rect -14308 5188 -14288 5612
rect -15060 5160 -14288 5188
rect -14048 5612 -13276 5640
rect -14048 5188 -13360 5612
rect -13296 5188 -13276 5612
rect -14048 5160 -13276 5188
rect -13036 5612 -12264 5640
rect -13036 5188 -12348 5612
rect -12284 5188 -12264 5612
rect -13036 5160 -12264 5188
rect -12024 5612 -11252 5640
rect -12024 5188 -11336 5612
rect -11272 5188 -11252 5612
rect -12024 5160 -11252 5188
rect -11012 5612 -10240 5640
rect -11012 5188 -10324 5612
rect -10260 5188 -10240 5612
rect -11012 5160 -10240 5188
rect -10000 5612 -9228 5640
rect -10000 5188 -9312 5612
rect -9248 5188 -9228 5612
rect -10000 5160 -9228 5188
rect -8988 5612 -8216 5640
rect -8988 5188 -8300 5612
rect -8236 5188 -8216 5612
rect -8988 5160 -8216 5188
rect -7976 5612 -7204 5640
rect -7976 5188 -7288 5612
rect -7224 5188 -7204 5612
rect -7976 5160 -7204 5188
rect -6964 5612 -6192 5640
rect -6964 5188 -6276 5612
rect -6212 5188 -6192 5612
rect -6964 5160 -6192 5188
rect -5952 5612 -5180 5640
rect -5952 5188 -5264 5612
rect -5200 5188 -5180 5612
rect -5952 5160 -5180 5188
rect -4940 5612 -4168 5640
rect -4940 5188 -4252 5612
rect -4188 5188 -4168 5612
rect -4940 5160 -4168 5188
rect -3928 5612 -3156 5640
rect -3928 5188 -3240 5612
rect -3176 5188 -3156 5612
rect -3928 5160 -3156 5188
rect -2916 5612 -2144 5640
rect -2916 5188 -2228 5612
rect -2164 5188 -2144 5612
rect -2916 5160 -2144 5188
rect -1904 5612 -1132 5640
rect -1904 5188 -1216 5612
rect -1152 5188 -1132 5612
rect -1904 5160 -1132 5188
rect -892 5612 -120 5640
rect -892 5188 -204 5612
rect -140 5188 -120 5612
rect -892 5160 -120 5188
rect 120 5612 892 5640
rect 120 5188 808 5612
rect 872 5188 892 5612
rect 120 5160 892 5188
rect 1132 5612 1904 5640
rect 1132 5188 1820 5612
rect 1884 5188 1904 5612
rect 1132 5160 1904 5188
rect 2144 5612 2916 5640
rect 2144 5188 2832 5612
rect 2896 5188 2916 5612
rect 2144 5160 2916 5188
rect 3156 5612 3928 5640
rect 3156 5188 3844 5612
rect 3908 5188 3928 5612
rect 3156 5160 3928 5188
rect 4168 5612 4940 5640
rect 4168 5188 4856 5612
rect 4920 5188 4940 5612
rect 4168 5160 4940 5188
rect 5180 5612 5952 5640
rect 5180 5188 5868 5612
rect 5932 5188 5952 5612
rect 5180 5160 5952 5188
rect 6192 5612 6964 5640
rect 6192 5188 6880 5612
rect 6944 5188 6964 5612
rect 6192 5160 6964 5188
rect 7204 5612 7976 5640
rect 7204 5188 7892 5612
rect 7956 5188 7976 5612
rect 7204 5160 7976 5188
rect 8216 5612 8988 5640
rect 8216 5188 8904 5612
rect 8968 5188 8988 5612
rect 8216 5160 8988 5188
rect 9228 5612 10000 5640
rect 9228 5188 9916 5612
rect 9980 5188 10000 5612
rect 9228 5160 10000 5188
rect 10240 5612 11012 5640
rect 10240 5188 10928 5612
rect 10992 5188 11012 5612
rect 10240 5160 11012 5188
rect 11252 5612 12024 5640
rect 11252 5188 11940 5612
rect 12004 5188 12024 5612
rect 11252 5160 12024 5188
rect 12264 5612 13036 5640
rect 12264 5188 12952 5612
rect 13016 5188 13036 5612
rect 12264 5160 13036 5188
rect 13276 5612 14048 5640
rect 13276 5188 13964 5612
rect 14028 5188 14048 5612
rect 13276 5160 14048 5188
rect 14288 5612 15060 5640
rect 14288 5188 14976 5612
rect 15040 5188 15060 5612
rect 14288 5160 15060 5188
rect 15300 5612 16072 5640
rect 15300 5188 15988 5612
rect 16052 5188 16072 5612
rect 15300 5160 16072 5188
rect 16312 5612 17084 5640
rect 16312 5188 17000 5612
rect 17064 5188 17084 5612
rect 16312 5160 17084 5188
rect 17324 5612 18096 5640
rect 17324 5188 18012 5612
rect 18076 5188 18096 5612
rect 17324 5160 18096 5188
rect 18336 5612 19108 5640
rect 18336 5188 19024 5612
rect 19088 5188 19108 5612
rect 18336 5160 19108 5188
rect 19348 5612 20120 5640
rect 19348 5188 20036 5612
rect 20100 5188 20120 5612
rect 19348 5160 20120 5188
rect 20360 5612 21132 5640
rect 20360 5188 21048 5612
rect 21112 5188 21132 5612
rect 20360 5160 21132 5188
rect 21372 5612 22144 5640
rect 21372 5188 22060 5612
rect 22124 5188 22144 5612
rect 21372 5160 22144 5188
rect 22384 5612 23156 5640
rect 22384 5188 23072 5612
rect 23136 5188 23156 5612
rect 22384 5160 23156 5188
rect 23396 5612 24168 5640
rect 23396 5188 24084 5612
rect 24148 5188 24168 5612
rect 23396 5160 24168 5188
rect 24408 5612 25180 5640
rect 24408 5188 25096 5612
rect 25160 5188 25180 5612
rect 24408 5160 25180 5188
rect 25420 5612 26192 5640
rect 25420 5188 26108 5612
rect 26172 5188 26192 5612
rect 25420 5160 26192 5188
rect 26432 5612 27204 5640
rect 26432 5188 27120 5612
rect 27184 5188 27204 5612
rect 26432 5160 27204 5188
rect 27444 5612 28216 5640
rect 27444 5188 28132 5612
rect 28196 5188 28216 5612
rect 27444 5160 28216 5188
rect 28456 5612 29228 5640
rect 28456 5188 29144 5612
rect 29208 5188 29228 5612
rect 28456 5160 29228 5188
rect 29468 5612 30240 5640
rect 29468 5188 30156 5612
rect 30220 5188 30240 5612
rect 29468 5160 30240 5188
rect 30480 5612 31252 5640
rect 30480 5188 31168 5612
rect 31232 5188 31252 5612
rect 30480 5160 31252 5188
rect 31492 5612 32264 5640
rect 31492 5188 32180 5612
rect 32244 5188 32264 5612
rect 31492 5160 32264 5188
rect -32264 4892 -31492 4920
rect -32264 4468 -31576 4892
rect -31512 4468 -31492 4892
rect -32264 4440 -31492 4468
rect -31252 4892 -30480 4920
rect -31252 4468 -30564 4892
rect -30500 4468 -30480 4892
rect -31252 4440 -30480 4468
rect -30240 4892 -29468 4920
rect -30240 4468 -29552 4892
rect -29488 4468 -29468 4892
rect -30240 4440 -29468 4468
rect -29228 4892 -28456 4920
rect -29228 4468 -28540 4892
rect -28476 4468 -28456 4892
rect -29228 4440 -28456 4468
rect -28216 4892 -27444 4920
rect -28216 4468 -27528 4892
rect -27464 4468 -27444 4892
rect -28216 4440 -27444 4468
rect -27204 4892 -26432 4920
rect -27204 4468 -26516 4892
rect -26452 4468 -26432 4892
rect -27204 4440 -26432 4468
rect -26192 4892 -25420 4920
rect -26192 4468 -25504 4892
rect -25440 4468 -25420 4892
rect -26192 4440 -25420 4468
rect -25180 4892 -24408 4920
rect -25180 4468 -24492 4892
rect -24428 4468 -24408 4892
rect -25180 4440 -24408 4468
rect -24168 4892 -23396 4920
rect -24168 4468 -23480 4892
rect -23416 4468 -23396 4892
rect -24168 4440 -23396 4468
rect -23156 4892 -22384 4920
rect -23156 4468 -22468 4892
rect -22404 4468 -22384 4892
rect -23156 4440 -22384 4468
rect -22144 4892 -21372 4920
rect -22144 4468 -21456 4892
rect -21392 4468 -21372 4892
rect -22144 4440 -21372 4468
rect -21132 4892 -20360 4920
rect -21132 4468 -20444 4892
rect -20380 4468 -20360 4892
rect -21132 4440 -20360 4468
rect -20120 4892 -19348 4920
rect -20120 4468 -19432 4892
rect -19368 4468 -19348 4892
rect -20120 4440 -19348 4468
rect -19108 4892 -18336 4920
rect -19108 4468 -18420 4892
rect -18356 4468 -18336 4892
rect -19108 4440 -18336 4468
rect -18096 4892 -17324 4920
rect -18096 4468 -17408 4892
rect -17344 4468 -17324 4892
rect -18096 4440 -17324 4468
rect -17084 4892 -16312 4920
rect -17084 4468 -16396 4892
rect -16332 4468 -16312 4892
rect -17084 4440 -16312 4468
rect -16072 4892 -15300 4920
rect -16072 4468 -15384 4892
rect -15320 4468 -15300 4892
rect -16072 4440 -15300 4468
rect -15060 4892 -14288 4920
rect -15060 4468 -14372 4892
rect -14308 4468 -14288 4892
rect -15060 4440 -14288 4468
rect -14048 4892 -13276 4920
rect -14048 4468 -13360 4892
rect -13296 4468 -13276 4892
rect -14048 4440 -13276 4468
rect -13036 4892 -12264 4920
rect -13036 4468 -12348 4892
rect -12284 4468 -12264 4892
rect -13036 4440 -12264 4468
rect -12024 4892 -11252 4920
rect -12024 4468 -11336 4892
rect -11272 4468 -11252 4892
rect -12024 4440 -11252 4468
rect -11012 4892 -10240 4920
rect -11012 4468 -10324 4892
rect -10260 4468 -10240 4892
rect -11012 4440 -10240 4468
rect -10000 4892 -9228 4920
rect -10000 4468 -9312 4892
rect -9248 4468 -9228 4892
rect -10000 4440 -9228 4468
rect -8988 4892 -8216 4920
rect -8988 4468 -8300 4892
rect -8236 4468 -8216 4892
rect -8988 4440 -8216 4468
rect -7976 4892 -7204 4920
rect -7976 4468 -7288 4892
rect -7224 4468 -7204 4892
rect -7976 4440 -7204 4468
rect -6964 4892 -6192 4920
rect -6964 4468 -6276 4892
rect -6212 4468 -6192 4892
rect -6964 4440 -6192 4468
rect -5952 4892 -5180 4920
rect -5952 4468 -5264 4892
rect -5200 4468 -5180 4892
rect -5952 4440 -5180 4468
rect -4940 4892 -4168 4920
rect -4940 4468 -4252 4892
rect -4188 4468 -4168 4892
rect -4940 4440 -4168 4468
rect -3928 4892 -3156 4920
rect -3928 4468 -3240 4892
rect -3176 4468 -3156 4892
rect -3928 4440 -3156 4468
rect -2916 4892 -2144 4920
rect -2916 4468 -2228 4892
rect -2164 4468 -2144 4892
rect -2916 4440 -2144 4468
rect -1904 4892 -1132 4920
rect -1904 4468 -1216 4892
rect -1152 4468 -1132 4892
rect -1904 4440 -1132 4468
rect -892 4892 -120 4920
rect -892 4468 -204 4892
rect -140 4468 -120 4892
rect -892 4440 -120 4468
rect 120 4892 892 4920
rect 120 4468 808 4892
rect 872 4468 892 4892
rect 120 4440 892 4468
rect 1132 4892 1904 4920
rect 1132 4468 1820 4892
rect 1884 4468 1904 4892
rect 1132 4440 1904 4468
rect 2144 4892 2916 4920
rect 2144 4468 2832 4892
rect 2896 4468 2916 4892
rect 2144 4440 2916 4468
rect 3156 4892 3928 4920
rect 3156 4468 3844 4892
rect 3908 4468 3928 4892
rect 3156 4440 3928 4468
rect 4168 4892 4940 4920
rect 4168 4468 4856 4892
rect 4920 4468 4940 4892
rect 4168 4440 4940 4468
rect 5180 4892 5952 4920
rect 5180 4468 5868 4892
rect 5932 4468 5952 4892
rect 5180 4440 5952 4468
rect 6192 4892 6964 4920
rect 6192 4468 6880 4892
rect 6944 4468 6964 4892
rect 6192 4440 6964 4468
rect 7204 4892 7976 4920
rect 7204 4468 7892 4892
rect 7956 4468 7976 4892
rect 7204 4440 7976 4468
rect 8216 4892 8988 4920
rect 8216 4468 8904 4892
rect 8968 4468 8988 4892
rect 8216 4440 8988 4468
rect 9228 4892 10000 4920
rect 9228 4468 9916 4892
rect 9980 4468 10000 4892
rect 9228 4440 10000 4468
rect 10240 4892 11012 4920
rect 10240 4468 10928 4892
rect 10992 4468 11012 4892
rect 10240 4440 11012 4468
rect 11252 4892 12024 4920
rect 11252 4468 11940 4892
rect 12004 4468 12024 4892
rect 11252 4440 12024 4468
rect 12264 4892 13036 4920
rect 12264 4468 12952 4892
rect 13016 4468 13036 4892
rect 12264 4440 13036 4468
rect 13276 4892 14048 4920
rect 13276 4468 13964 4892
rect 14028 4468 14048 4892
rect 13276 4440 14048 4468
rect 14288 4892 15060 4920
rect 14288 4468 14976 4892
rect 15040 4468 15060 4892
rect 14288 4440 15060 4468
rect 15300 4892 16072 4920
rect 15300 4468 15988 4892
rect 16052 4468 16072 4892
rect 15300 4440 16072 4468
rect 16312 4892 17084 4920
rect 16312 4468 17000 4892
rect 17064 4468 17084 4892
rect 16312 4440 17084 4468
rect 17324 4892 18096 4920
rect 17324 4468 18012 4892
rect 18076 4468 18096 4892
rect 17324 4440 18096 4468
rect 18336 4892 19108 4920
rect 18336 4468 19024 4892
rect 19088 4468 19108 4892
rect 18336 4440 19108 4468
rect 19348 4892 20120 4920
rect 19348 4468 20036 4892
rect 20100 4468 20120 4892
rect 19348 4440 20120 4468
rect 20360 4892 21132 4920
rect 20360 4468 21048 4892
rect 21112 4468 21132 4892
rect 20360 4440 21132 4468
rect 21372 4892 22144 4920
rect 21372 4468 22060 4892
rect 22124 4468 22144 4892
rect 21372 4440 22144 4468
rect 22384 4892 23156 4920
rect 22384 4468 23072 4892
rect 23136 4468 23156 4892
rect 22384 4440 23156 4468
rect 23396 4892 24168 4920
rect 23396 4468 24084 4892
rect 24148 4468 24168 4892
rect 23396 4440 24168 4468
rect 24408 4892 25180 4920
rect 24408 4468 25096 4892
rect 25160 4468 25180 4892
rect 24408 4440 25180 4468
rect 25420 4892 26192 4920
rect 25420 4468 26108 4892
rect 26172 4468 26192 4892
rect 25420 4440 26192 4468
rect 26432 4892 27204 4920
rect 26432 4468 27120 4892
rect 27184 4468 27204 4892
rect 26432 4440 27204 4468
rect 27444 4892 28216 4920
rect 27444 4468 28132 4892
rect 28196 4468 28216 4892
rect 27444 4440 28216 4468
rect 28456 4892 29228 4920
rect 28456 4468 29144 4892
rect 29208 4468 29228 4892
rect 28456 4440 29228 4468
rect 29468 4892 30240 4920
rect 29468 4468 30156 4892
rect 30220 4468 30240 4892
rect 29468 4440 30240 4468
rect 30480 4892 31252 4920
rect 30480 4468 31168 4892
rect 31232 4468 31252 4892
rect 30480 4440 31252 4468
rect 31492 4892 32264 4920
rect 31492 4468 32180 4892
rect 32244 4468 32264 4892
rect 31492 4440 32264 4468
rect -32264 4172 -31492 4200
rect -32264 3748 -31576 4172
rect -31512 3748 -31492 4172
rect -32264 3720 -31492 3748
rect -31252 4172 -30480 4200
rect -31252 3748 -30564 4172
rect -30500 3748 -30480 4172
rect -31252 3720 -30480 3748
rect -30240 4172 -29468 4200
rect -30240 3748 -29552 4172
rect -29488 3748 -29468 4172
rect -30240 3720 -29468 3748
rect -29228 4172 -28456 4200
rect -29228 3748 -28540 4172
rect -28476 3748 -28456 4172
rect -29228 3720 -28456 3748
rect -28216 4172 -27444 4200
rect -28216 3748 -27528 4172
rect -27464 3748 -27444 4172
rect -28216 3720 -27444 3748
rect -27204 4172 -26432 4200
rect -27204 3748 -26516 4172
rect -26452 3748 -26432 4172
rect -27204 3720 -26432 3748
rect -26192 4172 -25420 4200
rect -26192 3748 -25504 4172
rect -25440 3748 -25420 4172
rect -26192 3720 -25420 3748
rect -25180 4172 -24408 4200
rect -25180 3748 -24492 4172
rect -24428 3748 -24408 4172
rect -25180 3720 -24408 3748
rect -24168 4172 -23396 4200
rect -24168 3748 -23480 4172
rect -23416 3748 -23396 4172
rect -24168 3720 -23396 3748
rect -23156 4172 -22384 4200
rect -23156 3748 -22468 4172
rect -22404 3748 -22384 4172
rect -23156 3720 -22384 3748
rect -22144 4172 -21372 4200
rect -22144 3748 -21456 4172
rect -21392 3748 -21372 4172
rect -22144 3720 -21372 3748
rect -21132 4172 -20360 4200
rect -21132 3748 -20444 4172
rect -20380 3748 -20360 4172
rect -21132 3720 -20360 3748
rect -20120 4172 -19348 4200
rect -20120 3748 -19432 4172
rect -19368 3748 -19348 4172
rect -20120 3720 -19348 3748
rect -19108 4172 -18336 4200
rect -19108 3748 -18420 4172
rect -18356 3748 -18336 4172
rect -19108 3720 -18336 3748
rect -18096 4172 -17324 4200
rect -18096 3748 -17408 4172
rect -17344 3748 -17324 4172
rect -18096 3720 -17324 3748
rect -17084 4172 -16312 4200
rect -17084 3748 -16396 4172
rect -16332 3748 -16312 4172
rect -17084 3720 -16312 3748
rect -16072 4172 -15300 4200
rect -16072 3748 -15384 4172
rect -15320 3748 -15300 4172
rect -16072 3720 -15300 3748
rect -15060 4172 -14288 4200
rect -15060 3748 -14372 4172
rect -14308 3748 -14288 4172
rect -15060 3720 -14288 3748
rect -14048 4172 -13276 4200
rect -14048 3748 -13360 4172
rect -13296 3748 -13276 4172
rect -14048 3720 -13276 3748
rect -13036 4172 -12264 4200
rect -13036 3748 -12348 4172
rect -12284 3748 -12264 4172
rect -13036 3720 -12264 3748
rect -12024 4172 -11252 4200
rect -12024 3748 -11336 4172
rect -11272 3748 -11252 4172
rect -12024 3720 -11252 3748
rect -11012 4172 -10240 4200
rect -11012 3748 -10324 4172
rect -10260 3748 -10240 4172
rect -11012 3720 -10240 3748
rect -10000 4172 -9228 4200
rect -10000 3748 -9312 4172
rect -9248 3748 -9228 4172
rect -10000 3720 -9228 3748
rect -8988 4172 -8216 4200
rect -8988 3748 -8300 4172
rect -8236 3748 -8216 4172
rect -8988 3720 -8216 3748
rect -7976 4172 -7204 4200
rect -7976 3748 -7288 4172
rect -7224 3748 -7204 4172
rect -7976 3720 -7204 3748
rect -6964 4172 -6192 4200
rect -6964 3748 -6276 4172
rect -6212 3748 -6192 4172
rect -6964 3720 -6192 3748
rect -5952 4172 -5180 4200
rect -5952 3748 -5264 4172
rect -5200 3748 -5180 4172
rect -5952 3720 -5180 3748
rect -4940 4172 -4168 4200
rect -4940 3748 -4252 4172
rect -4188 3748 -4168 4172
rect -4940 3720 -4168 3748
rect -3928 4172 -3156 4200
rect -3928 3748 -3240 4172
rect -3176 3748 -3156 4172
rect -3928 3720 -3156 3748
rect -2916 4172 -2144 4200
rect -2916 3748 -2228 4172
rect -2164 3748 -2144 4172
rect -2916 3720 -2144 3748
rect -1904 4172 -1132 4200
rect -1904 3748 -1216 4172
rect -1152 3748 -1132 4172
rect -1904 3720 -1132 3748
rect -892 4172 -120 4200
rect -892 3748 -204 4172
rect -140 3748 -120 4172
rect -892 3720 -120 3748
rect 120 4172 892 4200
rect 120 3748 808 4172
rect 872 3748 892 4172
rect 120 3720 892 3748
rect 1132 4172 1904 4200
rect 1132 3748 1820 4172
rect 1884 3748 1904 4172
rect 1132 3720 1904 3748
rect 2144 4172 2916 4200
rect 2144 3748 2832 4172
rect 2896 3748 2916 4172
rect 2144 3720 2916 3748
rect 3156 4172 3928 4200
rect 3156 3748 3844 4172
rect 3908 3748 3928 4172
rect 3156 3720 3928 3748
rect 4168 4172 4940 4200
rect 4168 3748 4856 4172
rect 4920 3748 4940 4172
rect 4168 3720 4940 3748
rect 5180 4172 5952 4200
rect 5180 3748 5868 4172
rect 5932 3748 5952 4172
rect 5180 3720 5952 3748
rect 6192 4172 6964 4200
rect 6192 3748 6880 4172
rect 6944 3748 6964 4172
rect 6192 3720 6964 3748
rect 7204 4172 7976 4200
rect 7204 3748 7892 4172
rect 7956 3748 7976 4172
rect 7204 3720 7976 3748
rect 8216 4172 8988 4200
rect 8216 3748 8904 4172
rect 8968 3748 8988 4172
rect 8216 3720 8988 3748
rect 9228 4172 10000 4200
rect 9228 3748 9916 4172
rect 9980 3748 10000 4172
rect 9228 3720 10000 3748
rect 10240 4172 11012 4200
rect 10240 3748 10928 4172
rect 10992 3748 11012 4172
rect 10240 3720 11012 3748
rect 11252 4172 12024 4200
rect 11252 3748 11940 4172
rect 12004 3748 12024 4172
rect 11252 3720 12024 3748
rect 12264 4172 13036 4200
rect 12264 3748 12952 4172
rect 13016 3748 13036 4172
rect 12264 3720 13036 3748
rect 13276 4172 14048 4200
rect 13276 3748 13964 4172
rect 14028 3748 14048 4172
rect 13276 3720 14048 3748
rect 14288 4172 15060 4200
rect 14288 3748 14976 4172
rect 15040 3748 15060 4172
rect 14288 3720 15060 3748
rect 15300 4172 16072 4200
rect 15300 3748 15988 4172
rect 16052 3748 16072 4172
rect 15300 3720 16072 3748
rect 16312 4172 17084 4200
rect 16312 3748 17000 4172
rect 17064 3748 17084 4172
rect 16312 3720 17084 3748
rect 17324 4172 18096 4200
rect 17324 3748 18012 4172
rect 18076 3748 18096 4172
rect 17324 3720 18096 3748
rect 18336 4172 19108 4200
rect 18336 3748 19024 4172
rect 19088 3748 19108 4172
rect 18336 3720 19108 3748
rect 19348 4172 20120 4200
rect 19348 3748 20036 4172
rect 20100 3748 20120 4172
rect 19348 3720 20120 3748
rect 20360 4172 21132 4200
rect 20360 3748 21048 4172
rect 21112 3748 21132 4172
rect 20360 3720 21132 3748
rect 21372 4172 22144 4200
rect 21372 3748 22060 4172
rect 22124 3748 22144 4172
rect 21372 3720 22144 3748
rect 22384 4172 23156 4200
rect 22384 3748 23072 4172
rect 23136 3748 23156 4172
rect 22384 3720 23156 3748
rect 23396 4172 24168 4200
rect 23396 3748 24084 4172
rect 24148 3748 24168 4172
rect 23396 3720 24168 3748
rect 24408 4172 25180 4200
rect 24408 3748 25096 4172
rect 25160 3748 25180 4172
rect 24408 3720 25180 3748
rect 25420 4172 26192 4200
rect 25420 3748 26108 4172
rect 26172 3748 26192 4172
rect 25420 3720 26192 3748
rect 26432 4172 27204 4200
rect 26432 3748 27120 4172
rect 27184 3748 27204 4172
rect 26432 3720 27204 3748
rect 27444 4172 28216 4200
rect 27444 3748 28132 4172
rect 28196 3748 28216 4172
rect 27444 3720 28216 3748
rect 28456 4172 29228 4200
rect 28456 3748 29144 4172
rect 29208 3748 29228 4172
rect 28456 3720 29228 3748
rect 29468 4172 30240 4200
rect 29468 3748 30156 4172
rect 30220 3748 30240 4172
rect 29468 3720 30240 3748
rect 30480 4172 31252 4200
rect 30480 3748 31168 4172
rect 31232 3748 31252 4172
rect 30480 3720 31252 3748
rect 31492 4172 32264 4200
rect 31492 3748 32180 4172
rect 32244 3748 32264 4172
rect 31492 3720 32264 3748
rect -32264 3452 -31492 3480
rect -32264 3028 -31576 3452
rect -31512 3028 -31492 3452
rect -32264 3000 -31492 3028
rect -31252 3452 -30480 3480
rect -31252 3028 -30564 3452
rect -30500 3028 -30480 3452
rect -31252 3000 -30480 3028
rect -30240 3452 -29468 3480
rect -30240 3028 -29552 3452
rect -29488 3028 -29468 3452
rect -30240 3000 -29468 3028
rect -29228 3452 -28456 3480
rect -29228 3028 -28540 3452
rect -28476 3028 -28456 3452
rect -29228 3000 -28456 3028
rect -28216 3452 -27444 3480
rect -28216 3028 -27528 3452
rect -27464 3028 -27444 3452
rect -28216 3000 -27444 3028
rect -27204 3452 -26432 3480
rect -27204 3028 -26516 3452
rect -26452 3028 -26432 3452
rect -27204 3000 -26432 3028
rect -26192 3452 -25420 3480
rect -26192 3028 -25504 3452
rect -25440 3028 -25420 3452
rect -26192 3000 -25420 3028
rect -25180 3452 -24408 3480
rect -25180 3028 -24492 3452
rect -24428 3028 -24408 3452
rect -25180 3000 -24408 3028
rect -24168 3452 -23396 3480
rect -24168 3028 -23480 3452
rect -23416 3028 -23396 3452
rect -24168 3000 -23396 3028
rect -23156 3452 -22384 3480
rect -23156 3028 -22468 3452
rect -22404 3028 -22384 3452
rect -23156 3000 -22384 3028
rect -22144 3452 -21372 3480
rect -22144 3028 -21456 3452
rect -21392 3028 -21372 3452
rect -22144 3000 -21372 3028
rect -21132 3452 -20360 3480
rect -21132 3028 -20444 3452
rect -20380 3028 -20360 3452
rect -21132 3000 -20360 3028
rect -20120 3452 -19348 3480
rect -20120 3028 -19432 3452
rect -19368 3028 -19348 3452
rect -20120 3000 -19348 3028
rect -19108 3452 -18336 3480
rect -19108 3028 -18420 3452
rect -18356 3028 -18336 3452
rect -19108 3000 -18336 3028
rect -18096 3452 -17324 3480
rect -18096 3028 -17408 3452
rect -17344 3028 -17324 3452
rect -18096 3000 -17324 3028
rect -17084 3452 -16312 3480
rect -17084 3028 -16396 3452
rect -16332 3028 -16312 3452
rect -17084 3000 -16312 3028
rect -16072 3452 -15300 3480
rect -16072 3028 -15384 3452
rect -15320 3028 -15300 3452
rect -16072 3000 -15300 3028
rect -15060 3452 -14288 3480
rect -15060 3028 -14372 3452
rect -14308 3028 -14288 3452
rect -15060 3000 -14288 3028
rect -14048 3452 -13276 3480
rect -14048 3028 -13360 3452
rect -13296 3028 -13276 3452
rect -14048 3000 -13276 3028
rect -13036 3452 -12264 3480
rect -13036 3028 -12348 3452
rect -12284 3028 -12264 3452
rect -13036 3000 -12264 3028
rect -12024 3452 -11252 3480
rect -12024 3028 -11336 3452
rect -11272 3028 -11252 3452
rect -12024 3000 -11252 3028
rect -11012 3452 -10240 3480
rect -11012 3028 -10324 3452
rect -10260 3028 -10240 3452
rect -11012 3000 -10240 3028
rect -10000 3452 -9228 3480
rect -10000 3028 -9312 3452
rect -9248 3028 -9228 3452
rect -10000 3000 -9228 3028
rect -8988 3452 -8216 3480
rect -8988 3028 -8300 3452
rect -8236 3028 -8216 3452
rect -8988 3000 -8216 3028
rect -7976 3452 -7204 3480
rect -7976 3028 -7288 3452
rect -7224 3028 -7204 3452
rect -7976 3000 -7204 3028
rect -6964 3452 -6192 3480
rect -6964 3028 -6276 3452
rect -6212 3028 -6192 3452
rect -6964 3000 -6192 3028
rect -5952 3452 -5180 3480
rect -5952 3028 -5264 3452
rect -5200 3028 -5180 3452
rect -5952 3000 -5180 3028
rect -4940 3452 -4168 3480
rect -4940 3028 -4252 3452
rect -4188 3028 -4168 3452
rect -4940 3000 -4168 3028
rect -3928 3452 -3156 3480
rect -3928 3028 -3240 3452
rect -3176 3028 -3156 3452
rect -3928 3000 -3156 3028
rect -2916 3452 -2144 3480
rect -2916 3028 -2228 3452
rect -2164 3028 -2144 3452
rect -2916 3000 -2144 3028
rect -1904 3452 -1132 3480
rect -1904 3028 -1216 3452
rect -1152 3028 -1132 3452
rect -1904 3000 -1132 3028
rect -892 3452 -120 3480
rect -892 3028 -204 3452
rect -140 3028 -120 3452
rect -892 3000 -120 3028
rect 120 3452 892 3480
rect 120 3028 808 3452
rect 872 3028 892 3452
rect 120 3000 892 3028
rect 1132 3452 1904 3480
rect 1132 3028 1820 3452
rect 1884 3028 1904 3452
rect 1132 3000 1904 3028
rect 2144 3452 2916 3480
rect 2144 3028 2832 3452
rect 2896 3028 2916 3452
rect 2144 3000 2916 3028
rect 3156 3452 3928 3480
rect 3156 3028 3844 3452
rect 3908 3028 3928 3452
rect 3156 3000 3928 3028
rect 4168 3452 4940 3480
rect 4168 3028 4856 3452
rect 4920 3028 4940 3452
rect 4168 3000 4940 3028
rect 5180 3452 5952 3480
rect 5180 3028 5868 3452
rect 5932 3028 5952 3452
rect 5180 3000 5952 3028
rect 6192 3452 6964 3480
rect 6192 3028 6880 3452
rect 6944 3028 6964 3452
rect 6192 3000 6964 3028
rect 7204 3452 7976 3480
rect 7204 3028 7892 3452
rect 7956 3028 7976 3452
rect 7204 3000 7976 3028
rect 8216 3452 8988 3480
rect 8216 3028 8904 3452
rect 8968 3028 8988 3452
rect 8216 3000 8988 3028
rect 9228 3452 10000 3480
rect 9228 3028 9916 3452
rect 9980 3028 10000 3452
rect 9228 3000 10000 3028
rect 10240 3452 11012 3480
rect 10240 3028 10928 3452
rect 10992 3028 11012 3452
rect 10240 3000 11012 3028
rect 11252 3452 12024 3480
rect 11252 3028 11940 3452
rect 12004 3028 12024 3452
rect 11252 3000 12024 3028
rect 12264 3452 13036 3480
rect 12264 3028 12952 3452
rect 13016 3028 13036 3452
rect 12264 3000 13036 3028
rect 13276 3452 14048 3480
rect 13276 3028 13964 3452
rect 14028 3028 14048 3452
rect 13276 3000 14048 3028
rect 14288 3452 15060 3480
rect 14288 3028 14976 3452
rect 15040 3028 15060 3452
rect 14288 3000 15060 3028
rect 15300 3452 16072 3480
rect 15300 3028 15988 3452
rect 16052 3028 16072 3452
rect 15300 3000 16072 3028
rect 16312 3452 17084 3480
rect 16312 3028 17000 3452
rect 17064 3028 17084 3452
rect 16312 3000 17084 3028
rect 17324 3452 18096 3480
rect 17324 3028 18012 3452
rect 18076 3028 18096 3452
rect 17324 3000 18096 3028
rect 18336 3452 19108 3480
rect 18336 3028 19024 3452
rect 19088 3028 19108 3452
rect 18336 3000 19108 3028
rect 19348 3452 20120 3480
rect 19348 3028 20036 3452
rect 20100 3028 20120 3452
rect 19348 3000 20120 3028
rect 20360 3452 21132 3480
rect 20360 3028 21048 3452
rect 21112 3028 21132 3452
rect 20360 3000 21132 3028
rect 21372 3452 22144 3480
rect 21372 3028 22060 3452
rect 22124 3028 22144 3452
rect 21372 3000 22144 3028
rect 22384 3452 23156 3480
rect 22384 3028 23072 3452
rect 23136 3028 23156 3452
rect 22384 3000 23156 3028
rect 23396 3452 24168 3480
rect 23396 3028 24084 3452
rect 24148 3028 24168 3452
rect 23396 3000 24168 3028
rect 24408 3452 25180 3480
rect 24408 3028 25096 3452
rect 25160 3028 25180 3452
rect 24408 3000 25180 3028
rect 25420 3452 26192 3480
rect 25420 3028 26108 3452
rect 26172 3028 26192 3452
rect 25420 3000 26192 3028
rect 26432 3452 27204 3480
rect 26432 3028 27120 3452
rect 27184 3028 27204 3452
rect 26432 3000 27204 3028
rect 27444 3452 28216 3480
rect 27444 3028 28132 3452
rect 28196 3028 28216 3452
rect 27444 3000 28216 3028
rect 28456 3452 29228 3480
rect 28456 3028 29144 3452
rect 29208 3028 29228 3452
rect 28456 3000 29228 3028
rect 29468 3452 30240 3480
rect 29468 3028 30156 3452
rect 30220 3028 30240 3452
rect 29468 3000 30240 3028
rect 30480 3452 31252 3480
rect 30480 3028 31168 3452
rect 31232 3028 31252 3452
rect 30480 3000 31252 3028
rect 31492 3452 32264 3480
rect 31492 3028 32180 3452
rect 32244 3028 32264 3452
rect 31492 3000 32264 3028
rect -32264 2732 -31492 2760
rect -32264 2308 -31576 2732
rect -31512 2308 -31492 2732
rect -32264 2280 -31492 2308
rect -31252 2732 -30480 2760
rect -31252 2308 -30564 2732
rect -30500 2308 -30480 2732
rect -31252 2280 -30480 2308
rect -30240 2732 -29468 2760
rect -30240 2308 -29552 2732
rect -29488 2308 -29468 2732
rect -30240 2280 -29468 2308
rect -29228 2732 -28456 2760
rect -29228 2308 -28540 2732
rect -28476 2308 -28456 2732
rect -29228 2280 -28456 2308
rect -28216 2732 -27444 2760
rect -28216 2308 -27528 2732
rect -27464 2308 -27444 2732
rect -28216 2280 -27444 2308
rect -27204 2732 -26432 2760
rect -27204 2308 -26516 2732
rect -26452 2308 -26432 2732
rect -27204 2280 -26432 2308
rect -26192 2732 -25420 2760
rect -26192 2308 -25504 2732
rect -25440 2308 -25420 2732
rect -26192 2280 -25420 2308
rect -25180 2732 -24408 2760
rect -25180 2308 -24492 2732
rect -24428 2308 -24408 2732
rect -25180 2280 -24408 2308
rect -24168 2732 -23396 2760
rect -24168 2308 -23480 2732
rect -23416 2308 -23396 2732
rect -24168 2280 -23396 2308
rect -23156 2732 -22384 2760
rect -23156 2308 -22468 2732
rect -22404 2308 -22384 2732
rect -23156 2280 -22384 2308
rect -22144 2732 -21372 2760
rect -22144 2308 -21456 2732
rect -21392 2308 -21372 2732
rect -22144 2280 -21372 2308
rect -21132 2732 -20360 2760
rect -21132 2308 -20444 2732
rect -20380 2308 -20360 2732
rect -21132 2280 -20360 2308
rect -20120 2732 -19348 2760
rect -20120 2308 -19432 2732
rect -19368 2308 -19348 2732
rect -20120 2280 -19348 2308
rect -19108 2732 -18336 2760
rect -19108 2308 -18420 2732
rect -18356 2308 -18336 2732
rect -19108 2280 -18336 2308
rect -18096 2732 -17324 2760
rect -18096 2308 -17408 2732
rect -17344 2308 -17324 2732
rect -18096 2280 -17324 2308
rect -17084 2732 -16312 2760
rect -17084 2308 -16396 2732
rect -16332 2308 -16312 2732
rect -17084 2280 -16312 2308
rect -16072 2732 -15300 2760
rect -16072 2308 -15384 2732
rect -15320 2308 -15300 2732
rect -16072 2280 -15300 2308
rect -15060 2732 -14288 2760
rect -15060 2308 -14372 2732
rect -14308 2308 -14288 2732
rect -15060 2280 -14288 2308
rect -14048 2732 -13276 2760
rect -14048 2308 -13360 2732
rect -13296 2308 -13276 2732
rect -14048 2280 -13276 2308
rect -13036 2732 -12264 2760
rect -13036 2308 -12348 2732
rect -12284 2308 -12264 2732
rect -13036 2280 -12264 2308
rect -12024 2732 -11252 2760
rect -12024 2308 -11336 2732
rect -11272 2308 -11252 2732
rect -12024 2280 -11252 2308
rect -11012 2732 -10240 2760
rect -11012 2308 -10324 2732
rect -10260 2308 -10240 2732
rect -11012 2280 -10240 2308
rect -10000 2732 -9228 2760
rect -10000 2308 -9312 2732
rect -9248 2308 -9228 2732
rect -10000 2280 -9228 2308
rect -8988 2732 -8216 2760
rect -8988 2308 -8300 2732
rect -8236 2308 -8216 2732
rect -8988 2280 -8216 2308
rect -7976 2732 -7204 2760
rect -7976 2308 -7288 2732
rect -7224 2308 -7204 2732
rect -7976 2280 -7204 2308
rect -6964 2732 -6192 2760
rect -6964 2308 -6276 2732
rect -6212 2308 -6192 2732
rect -6964 2280 -6192 2308
rect -5952 2732 -5180 2760
rect -5952 2308 -5264 2732
rect -5200 2308 -5180 2732
rect -5952 2280 -5180 2308
rect -4940 2732 -4168 2760
rect -4940 2308 -4252 2732
rect -4188 2308 -4168 2732
rect -4940 2280 -4168 2308
rect -3928 2732 -3156 2760
rect -3928 2308 -3240 2732
rect -3176 2308 -3156 2732
rect -3928 2280 -3156 2308
rect -2916 2732 -2144 2760
rect -2916 2308 -2228 2732
rect -2164 2308 -2144 2732
rect -2916 2280 -2144 2308
rect -1904 2732 -1132 2760
rect -1904 2308 -1216 2732
rect -1152 2308 -1132 2732
rect -1904 2280 -1132 2308
rect -892 2732 -120 2760
rect -892 2308 -204 2732
rect -140 2308 -120 2732
rect -892 2280 -120 2308
rect 120 2732 892 2760
rect 120 2308 808 2732
rect 872 2308 892 2732
rect 120 2280 892 2308
rect 1132 2732 1904 2760
rect 1132 2308 1820 2732
rect 1884 2308 1904 2732
rect 1132 2280 1904 2308
rect 2144 2732 2916 2760
rect 2144 2308 2832 2732
rect 2896 2308 2916 2732
rect 2144 2280 2916 2308
rect 3156 2732 3928 2760
rect 3156 2308 3844 2732
rect 3908 2308 3928 2732
rect 3156 2280 3928 2308
rect 4168 2732 4940 2760
rect 4168 2308 4856 2732
rect 4920 2308 4940 2732
rect 4168 2280 4940 2308
rect 5180 2732 5952 2760
rect 5180 2308 5868 2732
rect 5932 2308 5952 2732
rect 5180 2280 5952 2308
rect 6192 2732 6964 2760
rect 6192 2308 6880 2732
rect 6944 2308 6964 2732
rect 6192 2280 6964 2308
rect 7204 2732 7976 2760
rect 7204 2308 7892 2732
rect 7956 2308 7976 2732
rect 7204 2280 7976 2308
rect 8216 2732 8988 2760
rect 8216 2308 8904 2732
rect 8968 2308 8988 2732
rect 8216 2280 8988 2308
rect 9228 2732 10000 2760
rect 9228 2308 9916 2732
rect 9980 2308 10000 2732
rect 9228 2280 10000 2308
rect 10240 2732 11012 2760
rect 10240 2308 10928 2732
rect 10992 2308 11012 2732
rect 10240 2280 11012 2308
rect 11252 2732 12024 2760
rect 11252 2308 11940 2732
rect 12004 2308 12024 2732
rect 11252 2280 12024 2308
rect 12264 2732 13036 2760
rect 12264 2308 12952 2732
rect 13016 2308 13036 2732
rect 12264 2280 13036 2308
rect 13276 2732 14048 2760
rect 13276 2308 13964 2732
rect 14028 2308 14048 2732
rect 13276 2280 14048 2308
rect 14288 2732 15060 2760
rect 14288 2308 14976 2732
rect 15040 2308 15060 2732
rect 14288 2280 15060 2308
rect 15300 2732 16072 2760
rect 15300 2308 15988 2732
rect 16052 2308 16072 2732
rect 15300 2280 16072 2308
rect 16312 2732 17084 2760
rect 16312 2308 17000 2732
rect 17064 2308 17084 2732
rect 16312 2280 17084 2308
rect 17324 2732 18096 2760
rect 17324 2308 18012 2732
rect 18076 2308 18096 2732
rect 17324 2280 18096 2308
rect 18336 2732 19108 2760
rect 18336 2308 19024 2732
rect 19088 2308 19108 2732
rect 18336 2280 19108 2308
rect 19348 2732 20120 2760
rect 19348 2308 20036 2732
rect 20100 2308 20120 2732
rect 19348 2280 20120 2308
rect 20360 2732 21132 2760
rect 20360 2308 21048 2732
rect 21112 2308 21132 2732
rect 20360 2280 21132 2308
rect 21372 2732 22144 2760
rect 21372 2308 22060 2732
rect 22124 2308 22144 2732
rect 21372 2280 22144 2308
rect 22384 2732 23156 2760
rect 22384 2308 23072 2732
rect 23136 2308 23156 2732
rect 22384 2280 23156 2308
rect 23396 2732 24168 2760
rect 23396 2308 24084 2732
rect 24148 2308 24168 2732
rect 23396 2280 24168 2308
rect 24408 2732 25180 2760
rect 24408 2308 25096 2732
rect 25160 2308 25180 2732
rect 24408 2280 25180 2308
rect 25420 2732 26192 2760
rect 25420 2308 26108 2732
rect 26172 2308 26192 2732
rect 25420 2280 26192 2308
rect 26432 2732 27204 2760
rect 26432 2308 27120 2732
rect 27184 2308 27204 2732
rect 26432 2280 27204 2308
rect 27444 2732 28216 2760
rect 27444 2308 28132 2732
rect 28196 2308 28216 2732
rect 27444 2280 28216 2308
rect 28456 2732 29228 2760
rect 28456 2308 29144 2732
rect 29208 2308 29228 2732
rect 28456 2280 29228 2308
rect 29468 2732 30240 2760
rect 29468 2308 30156 2732
rect 30220 2308 30240 2732
rect 29468 2280 30240 2308
rect 30480 2732 31252 2760
rect 30480 2308 31168 2732
rect 31232 2308 31252 2732
rect 30480 2280 31252 2308
rect 31492 2732 32264 2760
rect 31492 2308 32180 2732
rect 32244 2308 32264 2732
rect 31492 2280 32264 2308
rect -32264 2012 -31492 2040
rect -32264 1588 -31576 2012
rect -31512 1588 -31492 2012
rect -32264 1560 -31492 1588
rect -31252 2012 -30480 2040
rect -31252 1588 -30564 2012
rect -30500 1588 -30480 2012
rect -31252 1560 -30480 1588
rect -30240 2012 -29468 2040
rect -30240 1588 -29552 2012
rect -29488 1588 -29468 2012
rect -30240 1560 -29468 1588
rect -29228 2012 -28456 2040
rect -29228 1588 -28540 2012
rect -28476 1588 -28456 2012
rect -29228 1560 -28456 1588
rect -28216 2012 -27444 2040
rect -28216 1588 -27528 2012
rect -27464 1588 -27444 2012
rect -28216 1560 -27444 1588
rect -27204 2012 -26432 2040
rect -27204 1588 -26516 2012
rect -26452 1588 -26432 2012
rect -27204 1560 -26432 1588
rect -26192 2012 -25420 2040
rect -26192 1588 -25504 2012
rect -25440 1588 -25420 2012
rect -26192 1560 -25420 1588
rect -25180 2012 -24408 2040
rect -25180 1588 -24492 2012
rect -24428 1588 -24408 2012
rect -25180 1560 -24408 1588
rect -24168 2012 -23396 2040
rect -24168 1588 -23480 2012
rect -23416 1588 -23396 2012
rect -24168 1560 -23396 1588
rect -23156 2012 -22384 2040
rect -23156 1588 -22468 2012
rect -22404 1588 -22384 2012
rect -23156 1560 -22384 1588
rect -22144 2012 -21372 2040
rect -22144 1588 -21456 2012
rect -21392 1588 -21372 2012
rect -22144 1560 -21372 1588
rect -21132 2012 -20360 2040
rect -21132 1588 -20444 2012
rect -20380 1588 -20360 2012
rect -21132 1560 -20360 1588
rect -20120 2012 -19348 2040
rect -20120 1588 -19432 2012
rect -19368 1588 -19348 2012
rect -20120 1560 -19348 1588
rect -19108 2012 -18336 2040
rect -19108 1588 -18420 2012
rect -18356 1588 -18336 2012
rect -19108 1560 -18336 1588
rect -18096 2012 -17324 2040
rect -18096 1588 -17408 2012
rect -17344 1588 -17324 2012
rect -18096 1560 -17324 1588
rect -17084 2012 -16312 2040
rect -17084 1588 -16396 2012
rect -16332 1588 -16312 2012
rect -17084 1560 -16312 1588
rect -16072 2012 -15300 2040
rect -16072 1588 -15384 2012
rect -15320 1588 -15300 2012
rect -16072 1560 -15300 1588
rect -15060 2012 -14288 2040
rect -15060 1588 -14372 2012
rect -14308 1588 -14288 2012
rect -15060 1560 -14288 1588
rect -14048 2012 -13276 2040
rect -14048 1588 -13360 2012
rect -13296 1588 -13276 2012
rect -14048 1560 -13276 1588
rect -13036 2012 -12264 2040
rect -13036 1588 -12348 2012
rect -12284 1588 -12264 2012
rect -13036 1560 -12264 1588
rect -12024 2012 -11252 2040
rect -12024 1588 -11336 2012
rect -11272 1588 -11252 2012
rect -12024 1560 -11252 1588
rect -11012 2012 -10240 2040
rect -11012 1588 -10324 2012
rect -10260 1588 -10240 2012
rect -11012 1560 -10240 1588
rect -10000 2012 -9228 2040
rect -10000 1588 -9312 2012
rect -9248 1588 -9228 2012
rect -10000 1560 -9228 1588
rect -8988 2012 -8216 2040
rect -8988 1588 -8300 2012
rect -8236 1588 -8216 2012
rect -8988 1560 -8216 1588
rect -7976 2012 -7204 2040
rect -7976 1588 -7288 2012
rect -7224 1588 -7204 2012
rect -7976 1560 -7204 1588
rect -6964 2012 -6192 2040
rect -6964 1588 -6276 2012
rect -6212 1588 -6192 2012
rect -6964 1560 -6192 1588
rect -5952 2012 -5180 2040
rect -5952 1588 -5264 2012
rect -5200 1588 -5180 2012
rect -5952 1560 -5180 1588
rect -4940 2012 -4168 2040
rect -4940 1588 -4252 2012
rect -4188 1588 -4168 2012
rect -4940 1560 -4168 1588
rect -3928 2012 -3156 2040
rect -3928 1588 -3240 2012
rect -3176 1588 -3156 2012
rect -3928 1560 -3156 1588
rect -2916 2012 -2144 2040
rect -2916 1588 -2228 2012
rect -2164 1588 -2144 2012
rect -2916 1560 -2144 1588
rect -1904 2012 -1132 2040
rect -1904 1588 -1216 2012
rect -1152 1588 -1132 2012
rect -1904 1560 -1132 1588
rect -892 2012 -120 2040
rect -892 1588 -204 2012
rect -140 1588 -120 2012
rect -892 1560 -120 1588
rect 120 2012 892 2040
rect 120 1588 808 2012
rect 872 1588 892 2012
rect 120 1560 892 1588
rect 1132 2012 1904 2040
rect 1132 1588 1820 2012
rect 1884 1588 1904 2012
rect 1132 1560 1904 1588
rect 2144 2012 2916 2040
rect 2144 1588 2832 2012
rect 2896 1588 2916 2012
rect 2144 1560 2916 1588
rect 3156 2012 3928 2040
rect 3156 1588 3844 2012
rect 3908 1588 3928 2012
rect 3156 1560 3928 1588
rect 4168 2012 4940 2040
rect 4168 1588 4856 2012
rect 4920 1588 4940 2012
rect 4168 1560 4940 1588
rect 5180 2012 5952 2040
rect 5180 1588 5868 2012
rect 5932 1588 5952 2012
rect 5180 1560 5952 1588
rect 6192 2012 6964 2040
rect 6192 1588 6880 2012
rect 6944 1588 6964 2012
rect 6192 1560 6964 1588
rect 7204 2012 7976 2040
rect 7204 1588 7892 2012
rect 7956 1588 7976 2012
rect 7204 1560 7976 1588
rect 8216 2012 8988 2040
rect 8216 1588 8904 2012
rect 8968 1588 8988 2012
rect 8216 1560 8988 1588
rect 9228 2012 10000 2040
rect 9228 1588 9916 2012
rect 9980 1588 10000 2012
rect 9228 1560 10000 1588
rect 10240 2012 11012 2040
rect 10240 1588 10928 2012
rect 10992 1588 11012 2012
rect 10240 1560 11012 1588
rect 11252 2012 12024 2040
rect 11252 1588 11940 2012
rect 12004 1588 12024 2012
rect 11252 1560 12024 1588
rect 12264 2012 13036 2040
rect 12264 1588 12952 2012
rect 13016 1588 13036 2012
rect 12264 1560 13036 1588
rect 13276 2012 14048 2040
rect 13276 1588 13964 2012
rect 14028 1588 14048 2012
rect 13276 1560 14048 1588
rect 14288 2012 15060 2040
rect 14288 1588 14976 2012
rect 15040 1588 15060 2012
rect 14288 1560 15060 1588
rect 15300 2012 16072 2040
rect 15300 1588 15988 2012
rect 16052 1588 16072 2012
rect 15300 1560 16072 1588
rect 16312 2012 17084 2040
rect 16312 1588 17000 2012
rect 17064 1588 17084 2012
rect 16312 1560 17084 1588
rect 17324 2012 18096 2040
rect 17324 1588 18012 2012
rect 18076 1588 18096 2012
rect 17324 1560 18096 1588
rect 18336 2012 19108 2040
rect 18336 1588 19024 2012
rect 19088 1588 19108 2012
rect 18336 1560 19108 1588
rect 19348 2012 20120 2040
rect 19348 1588 20036 2012
rect 20100 1588 20120 2012
rect 19348 1560 20120 1588
rect 20360 2012 21132 2040
rect 20360 1588 21048 2012
rect 21112 1588 21132 2012
rect 20360 1560 21132 1588
rect 21372 2012 22144 2040
rect 21372 1588 22060 2012
rect 22124 1588 22144 2012
rect 21372 1560 22144 1588
rect 22384 2012 23156 2040
rect 22384 1588 23072 2012
rect 23136 1588 23156 2012
rect 22384 1560 23156 1588
rect 23396 2012 24168 2040
rect 23396 1588 24084 2012
rect 24148 1588 24168 2012
rect 23396 1560 24168 1588
rect 24408 2012 25180 2040
rect 24408 1588 25096 2012
rect 25160 1588 25180 2012
rect 24408 1560 25180 1588
rect 25420 2012 26192 2040
rect 25420 1588 26108 2012
rect 26172 1588 26192 2012
rect 25420 1560 26192 1588
rect 26432 2012 27204 2040
rect 26432 1588 27120 2012
rect 27184 1588 27204 2012
rect 26432 1560 27204 1588
rect 27444 2012 28216 2040
rect 27444 1588 28132 2012
rect 28196 1588 28216 2012
rect 27444 1560 28216 1588
rect 28456 2012 29228 2040
rect 28456 1588 29144 2012
rect 29208 1588 29228 2012
rect 28456 1560 29228 1588
rect 29468 2012 30240 2040
rect 29468 1588 30156 2012
rect 30220 1588 30240 2012
rect 29468 1560 30240 1588
rect 30480 2012 31252 2040
rect 30480 1588 31168 2012
rect 31232 1588 31252 2012
rect 30480 1560 31252 1588
rect 31492 2012 32264 2040
rect 31492 1588 32180 2012
rect 32244 1588 32264 2012
rect 31492 1560 32264 1588
rect -32264 1292 -31492 1320
rect -32264 868 -31576 1292
rect -31512 868 -31492 1292
rect -32264 840 -31492 868
rect -31252 1292 -30480 1320
rect -31252 868 -30564 1292
rect -30500 868 -30480 1292
rect -31252 840 -30480 868
rect -30240 1292 -29468 1320
rect -30240 868 -29552 1292
rect -29488 868 -29468 1292
rect -30240 840 -29468 868
rect -29228 1292 -28456 1320
rect -29228 868 -28540 1292
rect -28476 868 -28456 1292
rect -29228 840 -28456 868
rect -28216 1292 -27444 1320
rect -28216 868 -27528 1292
rect -27464 868 -27444 1292
rect -28216 840 -27444 868
rect -27204 1292 -26432 1320
rect -27204 868 -26516 1292
rect -26452 868 -26432 1292
rect -27204 840 -26432 868
rect -26192 1292 -25420 1320
rect -26192 868 -25504 1292
rect -25440 868 -25420 1292
rect -26192 840 -25420 868
rect -25180 1292 -24408 1320
rect -25180 868 -24492 1292
rect -24428 868 -24408 1292
rect -25180 840 -24408 868
rect -24168 1292 -23396 1320
rect -24168 868 -23480 1292
rect -23416 868 -23396 1292
rect -24168 840 -23396 868
rect -23156 1292 -22384 1320
rect -23156 868 -22468 1292
rect -22404 868 -22384 1292
rect -23156 840 -22384 868
rect -22144 1292 -21372 1320
rect -22144 868 -21456 1292
rect -21392 868 -21372 1292
rect -22144 840 -21372 868
rect -21132 1292 -20360 1320
rect -21132 868 -20444 1292
rect -20380 868 -20360 1292
rect -21132 840 -20360 868
rect -20120 1292 -19348 1320
rect -20120 868 -19432 1292
rect -19368 868 -19348 1292
rect -20120 840 -19348 868
rect -19108 1292 -18336 1320
rect -19108 868 -18420 1292
rect -18356 868 -18336 1292
rect -19108 840 -18336 868
rect -18096 1292 -17324 1320
rect -18096 868 -17408 1292
rect -17344 868 -17324 1292
rect -18096 840 -17324 868
rect -17084 1292 -16312 1320
rect -17084 868 -16396 1292
rect -16332 868 -16312 1292
rect -17084 840 -16312 868
rect -16072 1292 -15300 1320
rect -16072 868 -15384 1292
rect -15320 868 -15300 1292
rect -16072 840 -15300 868
rect -15060 1292 -14288 1320
rect -15060 868 -14372 1292
rect -14308 868 -14288 1292
rect -15060 840 -14288 868
rect -14048 1292 -13276 1320
rect -14048 868 -13360 1292
rect -13296 868 -13276 1292
rect -14048 840 -13276 868
rect -13036 1292 -12264 1320
rect -13036 868 -12348 1292
rect -12284 868 -12264 1292
rect -13036 840 -12264 868
rect -12024 1292 -11252 1320
rect -12024 868 -11336 1292
rect -11272 868 -11252 1292
rect -12024 840 -11252 868
rect -11012 1292 -10240 1320
rect -11012 868 -10324 1292
rect -10260 868 -10240 1292
rect -11012 840 -10240 868
rect -10000 1292 -9228 1320
rect -10000 868 -9312 1292
rect -9248 868 -9228 1292
rect -10000 840 -9228 868
rect -8988 1292 -8216 1320
rect -8988 868 -8300 1292
rect -8236 868 -8216 1292
rect -8988 840 -8216 868
rect -7976 1292 -7204 1320
rect -7976 868 -7288 1292
rect -7224 868 -7204 1292
rect -7976 840 -7204 868
rect -6964 1292 -6192 1320
rect -6964 868 -6276 1292
rect -6212 868 -6192 1292
rect -6964 840 -6192 868
rect -5952 1292 -5180 1320
rect -5952 868 -5264 1292
rect -5200 868 -5180 1292
rect -5952 840 -5180 868
rect -4940 1292 -4168 1320
rect -4940 868 -4252 1292
rect -4188 868 -4168 1292
rect -4940 840 -4168 868
rect -3928 1292 -3156 1320
rect -3928 868 -3240 1292
rect -3176 868 -3156 1292
rect -3928 840 -3156 868
rect -2916 1292 -2144 1320
rect -2916 868 -2228 1292
rect -2164 868 -2144 1292
rect -2916 840 -2144 868
rect -1904 1292 -1132 1320
rect -1904 868 -1216 1292
rect -1152 868 -1132 1292
rect -1904 840 -1132 868
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect 1132 1292 1904 1320
rect 1132 868 1820 1292
rect 1884 868 1904 1292
rect 1132 840 1904 868
rect 2144 1292 2916 1320
rect 2144 868 2832 1292
rect 2896 868 2916 1292
rect 2144 840 2916 868
rect 3156 1292 3928 1320
rect 3156 868 3844 1292
rect 3908 868 3928 1292
rect 3156 840 3928 868
rect 4168 1292 4940 1320
rect 4168 868 4856 1292
rect 4920 868 4940 1292
rect 4168 840 4940 868
rect 5180 1292 5952 1320
rect 5180 868 5868 1292
rect 5932 868 5952 1292
rect 5180 840 5952 868
rect 6192 1292 6964 1320
rect 6192 868 6880 1292
rect 6944 868 6964 1292
rect 6192 840 6964 868
rect 7204 1292 7976 1320
rect 7204 868 7892 1292
rect 7956 868 7976 1292
rect 7204 840 7976 868
rect 8216 1292 8988 1320
rect 8216 868 8904 1292
rect 8968 868 8988 1292
rect 8216 840 8988 868
rect 9228 1292 10000 1320
rect 9228 868 9916 1292
rect 9980 868 10000 1292
rect 9228 840 10000 868
rect 10240 1292 11012 1320
rect 10240 868 10928 1292
rect 10992 868 11012 1292
rect 10240 840 11012 868
rect 11252 1292 12024 1320
rect 11252 868 11940 1292
rect 12004 868 12024 1292
rect 11252 840 12024 868
rect 12264 1292 13036 1320
rect 12264 868 12952 1292
rect 13016 868 13036 1292
rect 12264 840 13036 868
rect 13276 1292 14048 1320
rect 13276 868 13964 1292
rect 14028 868 14048 1292
rect 13276 840 14048 868
rect 14288 1292 15060 1320
rect 14288 868 14976 1292
rect 15040 868 15060 1292
rect 14288 840 15060 868
rect 15300 1292 16072 1320
rect 15300 868 15988 1292
rect 16052 868 16072 1292
rect 15300 840 16072 868
rect 16312 1292 17084 1320
rect 16312 868 17000 1292
rect 17064 868 17084 1292
rect 16312 840 17084 868
rect 17324 1292 18096 1320
rect 17324 868 18012 1292
rect 18076 868 18096 1292
rect 17324 840 18096 868
rect 18336 1292 19108 1320
rect 18336 868 19024 1292
rect 19088 868 19108 1292
rect 18336 840 19108 868
rect 19348 1292 20120 1320
rect 19348 868 20036 1292
rect 20100 868 20120 1292
rect 19348 840 20120 868
rect 20360 1292 21132 1320
rect 20360 868 21048 1292
rect 21112 868 21132 1292
rect 20360 840 21132 868
rect 21372 1292 22144 1320
rect 21372 868 22060 1292
rect 22124 868 22144 1292
rect 21372 840 22144 868
rect 22384 1292 23156 1320
rect 22384 868 23072 1292
rect 23136 868 23156 1292
rect 22384 840 23156 868
rect 23396 1292 24168 1320
rect 23396 868 24084 1292
rect 24148 868 24168 1292
rect 23396 840 24168 868
rect 24408 1292 25180 1320
rect 24408 868 25096 1292
rect 25160 868 25180 1292
rect 24408 840 25180 868
rect 25420 1292 26192 1320
rect 25420 868 26108 1292
rect 26172 868 26192 1292
rect 25420 840 26192 868
rect 26432 1292 27204 1320
rect 26432 868 27120 1292
rect 27184 868 27204 1292
rect 26432 840 27204 868
rect 27444 1292 28216 1320
rect 27444 868 28132 1292
rect 28196 868 28216 1292
rect 27444 840 28216 868
rect 28456 1292 29228 1320
rect 28456 868 29144 1292
rect 29208 868 29228 1292
rect 28456 840 29228 868
rect 29468 1292 30240 1320
rect 29468 868 30156 1292
rect 30220 868 30240 1292
rect 29468 840 30240 868
rect 30480 1292 31252 1320
rect 30480 868 31168 1292
rect 31232 868 31252 1292
rect 30480 840 31252 868
rect 31492 1292 32264 1320
rect 31492 868 32180 1292
rect 32244 868 32264 1292
rect 31492 840 32264 868
rect -32264 572 -31492 600
rect -32264 148 -31576 572
rect -31512 148 -31492 572
rect -32264 120 -31492 148
rect -31252 572 -30480 600
rect -31252 148 -30564 572
rect -30500 148 -30480 572
rect -31252 120 -30480 148
rect -30240 572 -29468 600
rect -30240 148 -29552 572
rect -29488 148 -29468 572
rect -30240 120 -29468 148
rect -29228 572 -28456 600
rect -29228 148 -28540 572
rect -28476 148 -28456 572
rect -29228 120 -28456 148
rect -28216 572 -27444 600
rect -28216 148 -27528 572
rect -27464 148 -27444 572
rect -28216 120 -27444 148
rect -27204 572 -26432 600
rect -27204 148 -26516 572
rect -26452 148 -26432 572
rect -27204 120 -26432 148
rect -26192 572 -25420 600
rect -26192 148 -25504 572
rect -25440 148 -25420 572
rect -26192 120 -25420 148
rect -25180 572 -24408 600
rect -25180 148 -24492 572
rect -24428 148 -24408 572
rect -25180 120 -24408 148
rect -24168 572 -23396 600
rect -24168 148 -23480 572
rect -23416 148 -23396 572
rect -24168 120 -23396 148
rect -23156 572 -22384 600
rect -23156 148 -22468 572
rect -22404 148 -22384 572
rect -23156 120 -22384 148
rect -22144 572 -21372 600
rect -22144 148 -21456 572
rect -21392 148 -21372 572
rect -22144 120 -21372 148
rect -21132 572 -20360 600
rect -21132 148 -20444 572
rect -20380 148 -20360 572
rect -21132 120 -20360 148
rect -20120 572 -19348 600
rect -20120 148 -19432 572
rect -19368 148 -19348 572
rect -20120 120 -19348 148
rect -19108 572 -18336 600
rect -19108 148 -18420 572
rect -18356 148 -18336 572
rect -19108 120 -18336 148
rect -18096 572 -17324 600
rect -18096 148 -17408 572
rect -17344 148 -17324 572
rect -18096 120 -17324 148
rect -17084 572 -16312 600
rect -17084 148 -16396 572
rect -16332 148 -16312 572
rect -17084 120 -16312 148
rect -16072 572 -15300 600
rect -16072 148 -15384 572
rect -15320 148 -15300 572
rect -16072 120 -15300 148
rect -15060 572 -14288 600
rect -15060 148 -14372 572
rect -14308 148 -14288 572
rect -15060 120 -14288 148
rect -14048 572 -13276 600
rect -14048 148 -13360 572
rect -13296 148 -13276 572
rect -14048 120 -13276 148
rect -13036 572 -12264 600
rect -13036 148 -12348 572
rect -12284 148 -12264 572
rect -13036 120 -12264 148
rect -12024 572 -11252 600
rect -12024 148 -11336 572
rect -11272 148 -11252 572
rect -12024 120 -11252 148
rect -11012 572 -10240 600
rect -11012 148 -10324 572
rect -10260 148 -10240 572
rect -11012 120 -10240 148
rect -10000 572 -9228 600
rect -10000 148 -9312 572
rect -9248 148 -9228 572
rect -10000 120 -9228 148
rect -8988 572 -8216 600
rect -8988 148 -8300 572
rect -8236 148 -8216 572
rect -8988 120 -8216 148
rect -7976 572 -7204 600
rect -7976 148 -7288 572
rect -7224 148 -7204 572
rect -7976 120 -7204 148
rect -6964 572 -6192 600
rect -6964 148 -6276 572
rect -6212 148 -6192 572
rect -6964 120 -6192 148
rect -5952 572 -5180 600
rect -5952 148 -5264 572
rect -5200 148 -5180 572
rect -5952 120 -5180 148
rect -4940 572 -4168 600
rect -4940 148 -4252 572
rect -4188 148 -4168 572
rect -4940 120 -4168 148
rect -3928 572 -3156 600
rect -3928 148 -3240 572
rect -3176 148 -3156 572
rect -3928 120 -3156 148
rect -2916 572 -2144 600
rect -2916 148 -2228 572
rect -2164 148 -2144 572
rect -2916 120 -2144 148
rect -1904 572 -1132 600
rect -1904 148 -1216 572
rect -1152 148 -1132 572
rect -1904 120 -1132 148
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect 1132 572 1904 600
rect 1132 148 1820 572
rect 1884 148 1904 572
rect 1132 120 1904 148
rect 2144 572 2916 600
rect 2144 148 2832 572
rect 2896 148 2916 572
rect 2144 120 2916 148
rect 3156 572 3928 600
rect 3156 148 3844 572
rect 3908 148 3928 572
rect 3156 120 3928 148
rect 4168 572 4940 600
rect 4168 148 4856 572
rect 4920 148 4940 572
rect 4168 120 4940 148
rect 5180 572 5952 600
rect 5180 148 5868 572
rect 5932 148 5952 572
rect 5180 120 5952 148
rect 6192 572 6964 600
rect 6192 148 6880 572
rect 6944 148 6964 572
rect 6192 120 6964 148
rect 7204 572 7976 600
rect 7204 148 7892 572
rect 7956 148 7976 572
rect 7204 120 7976 148
rect 8216 572 8988 600
rect 8216 148 8904 572
rect 8968 148 8988 572
rect 8216 120 8988 148
rect 9228 572 10000 600
rect 9228 148 9916 572
rect 9980 148 10000 572
rect 9228 120 10000 148
rect 10240 572 11012 600
rect 10240 148 10928 572
rect 10992 148 11012 572
rect 10240 120 11012 148
rect 11252 572 12024 600
rect 11252 148 11940 572
rect 12004 148 12024 572
rect 11252 120 12024 148
rect 12264 572 13036 600
rect 12264 148 12952 572
rect 13016 148 13036 572
rect 12264 120 13036 148
rect 13276 572 14048 600
rect 13276 148 13964 572
rect 14028 148 14048 572
rect 13276 120 14048 148
rect 14288 572 15060 600
rect 14288 148 14976 572
rect 15040 148 15060 572
rect 14288 120 15060 148
rect 15300 572 16072 600
rect 15300 148 15988 572
rect 16052 148 16072 572
rect 15300 120 16072 148
rect 16312 572 17084 600
rect 16312 148 17000 572
rect 17064 148 17084 572
rect 16312 120 17084 148
rect 17324 572 18096 600
rect 17324 148 18012 572
rect 18076 148 18096 572
rect 17324 120 18096 148
rect 18336 572 19108 600
rect 18336 148 19024 572
rect 19088 148 19108 572
rect 18336 120 19108 148
rect 19348 572 20120 600
rect 19348 148 20036 572
rect 20100 148 20120 572
rect 19348 120 20120 148
rect 20360 572 21132 600
rect 20360 148 21048 572
rect 21112 148 21132 572
rect 20360 120 21132 148
rect 21372 572 22144 600
rect 21372 148 22060 572
rect 22124 148 22144 572
rect 21372 120 22144 148
rect 22384 572 23156 600
rect 22384 148 23072 572
rect 23136 148 23156 572
rect 22384 120 23156 148
rect 23396 572 24168 600
rect 23396 148 24084 572
rect 24148 148 24168 572
rect 23396 120 24168 148
rect 24408 572 25180 600
rect 24408 148 25096 572
rect 25160 148 25180 572
rect 24408 120 25180 148
rect 25420 572 26192 600
rect 25420 148 26108 572
rect 26172 148 26192 572
rect 25420 120 26192 148
rect 26432 572 27204 600
rect 26432 148 27120 572
rect 27184 148 27204 572
rect 26432 120 27204 148
rect 27444 572 28216 600
rect 27444 148 28132 572
rect 28196 148 28216 572
rect 27444 120 28216 148
rect 28456 572 29228 600
rect 28456 148 29144 572
rect 29208 148 29228 572
rect 28456 120 29228 148
rect 29468 572 30240 600
rect 29468 148 30156 572
rect 30220 148 30240 572
rect 29468 120 30240 148
rect 30480 572 31252 600
rect 30480 148 31168 572
rect 31232 148 31252 572
rect 30480 120 31252 148
rect 31492 572 32264 600
rect 31492 148 32180 572
rect 32244 148 32264 572
rect 31492 120 32264 148
rect -32264 -148 -31492 -120
rect -32264 -572 -31576 -148
rect -31512 -572 -31492 -148
rect -32264 -600 -31492 -572
rect -31252 -148 -30480 -120
rect -31252 -572 -30564 -148
rect -30500 -572 -30480 -148
rect -31252 -600 -30480 -572
rect -30240 -148 -29468 -120
rect -30240 -572 -29552 -148
rect -29488 -572 -29468 -148
rect -30240 -600 -29468 -572
rect -29228 -148 -28456 -120
rect -29228 -572 -28540 -148
rect -28476 -572 -28456 -148
rect -29228 -600 -28456 -572
rect -28216 -148 -27444 -120
rect -28216 -572 -27528 -148
rect -27464 -572 -27444 -148
rect -28216 -600 -27444 -572
rect -27204 -148 -26432 -120
rect -27204 -572 -26516 -148
rect -26452 -572 -26432 -148
rect -27204 -600 -26432 -572
rect -26192 -148 -25420 -120
rect -26192 -572 -25504 -148
rect -25440 -572 -25420 -148
rect -26192 -600 -25420 -572
rect -25180 -148 -24408 -120
rect -25180 -572 -24492 -148
rect -24428 -572 -24408 -148
rect -25180 -600 -24408 -572
rect -24168 -148 -23396 -120
rect -24168 -572 -23480 -148
rect -23416 -572 -23396 -148
rect -24168 -600 -23396 -572
rect -23156 -148 -22384 -120
rect -23156 -572 -22468 -148
rect -22404 -572 -22384 -148
rect -23156 -600 -22384 -572
rect -22144 -148 -21372 -120
rect -22144 -572 -21456 -148
rect -21392 -572 -21372 -148
rect -22144 -600 -21372 -572
rect -21132 -148 -20360 -120
rect -21132 -572 -20444 -148
rect -20380 -572 -20360 -148
rect -21132 -600 -20360 -572
rect -20120 -148 -19348 -120
rect -20120 -572 -19432 -148
rect -19368 -572 -19348 -148
rect -20120 -600 -19348 -572
rect -19108 -148 -18336 -120
rect -19108 -572 -18420 -148
rect -18356 -572 -18336 -148
rect -19108 -600 -18336 -572
rect -18096 -148 -17324 -120
rect -18096 -572 -17408 -148
rect -17344 -572 -17324 -148
rect -18096 -600 -17324 -572
rect -17084 -148 -16312 -120
rect -17084 -572 -16396 -148
rect -16332 -572 -16312 -148
rect -17084 -600 -16312 -572
rect -16072 -148 -15300 -120
rect -16072 -572 -15384 -148
rect -15320 -572 -15300 -148
rect -16072 -600 -15300 -572
rect -15060 -148 -14288 -120
rect -15060 -572 -14372 -148
rect -14308 -572 -14288 -148
rect -15060 -600 -14288 -572
rect -14048 -148 -13276 -120
rect -14048 -572 -13360 -148
rect -13296 -572 -13276 -148
rect -14048 -600 -13276 -572
rect -13036 -148 -12264 -120
rect -13036 -572 -12348 -148
rect -12284 -572 -12264 -148
rect -13036 -600 -12264 -572
rect -12024 -148 -11252 -120
rect -12024 -572 -11336 -148
rect -11272 -572 -11252 -148
rect -12024 -600 -11252 -572
rect -11012 -148 -10240 -120
rect -11012 -572 -10324 -148
rect -10260 -572 -10240 -148
rect -11012 -600 -10240 -572
rect -10000 -148 -9228 -120
rect -10000 -572 -9312 -148
rect -9248 -572 -9228 -148
rect -10000 -600 -9228 -572
rect -8988 -148 -8216 -120
rect -8988 -572 -8300 -148
rect -8236 -572 -8216 -148
rect -8988 -600 -8216 -572
rect -7976 -148 -7204 -120
rect -7976 -572 -7288 -148
rect -7224 -572 -7204 -148
rect -7976 -600 -7204 -572
rect -6964 -148 -6192 -120
rect -6964 -572 -6276 -148
rect -6212 -572 -6192 -148
rect -6964 -600 -6192 -572
rect -5952 -148 -5180 -120
rect -5952 -572 -5264 -148
rect -5200 -572 -5180 -148
rect -5952 -600 -5180 -572
rect -4940 -148 -4168 -120
rect -4940 -572 -4252 -148
rect -4188 -572 -4168 -148
rect -4940 -600 -4168 -572
rect -3928 -148 -3156 -120
rect -3928 -572 -3240 -148
rect -3176 -572 -3156 -148
rect -3928 -600 -3156 -572
rect -2916 -148 -2144 -120
rect -2916 -572 -2228 -148
rect -2164 -572 -2144 -148
rect -2916 -600 -2144 -572
rect -1904 -148 -1132 -120
rect -1904 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -1904 -600 -1132 -572
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect 1132 -148 1904 -120
rect 1132 -572 1820 -148
rect 1884 -572 1904 -148
rect 1132 -600 1904 -572
rect 2144 -148 2916 -120
rect 2144 -572 2832 -148
rect 2896 -572 2916 -148
rect 2144 -600 2916 -572
rect 3156 -148 3928 -120
rect 3156 -572 3844 -148
rect 3908 -572 3928 -148
rect 3156 -600 3928 -572
rect 4168 -148 4940 -120
rect 4168 -572 4856 -148
rect 4920 -572 4940 -148
rect 4168 -600 4940 -572
rect 5180 -148 5952 -120
rect 5180 -572 5868 -148
rect 5932 -572 5952 -148
rect 5180 -600 5952 -572
rect 6192 -148 6964 -120
rect 6192 -572 6880 -148
rect 6944 -572 6964 -148
rect 6192 -600 6964 -572
rect 7204 -148 7976 -120
rect 7204 -572 7892 -148
rect 7956 -572 7976 -148
rect 7204 -600 7976 -572
rect 8216 -148 8988 -120
rect 8216 -572 8904 -148
rect 8968 -572 8988 -148
rect 8216 -600 8988 -572
rect 9228 -148 10000 -120
rect 9228 -572 9916 -148
rect 9980 -572 10000 -148
rect 9228 -600 10000 -572
rect 10240 -148 11012 -120
rect 10240 -572 10928 -148
rect 10992 -572 11012 -148
rect 10240 -600 11012 -572
rect 11252 -148 12024 -120
rect 11252 -572 11940 -148
rect 12004 -572 12024 -148
rect 11252 -600 12024 -572
rect 12264 -148 13036 -120
rect 12264 -572 12952 -148
rect 13016 -572 13036 -148
rect 12264 -600 13036 -572
rect 13276 -148 14048 -120
rect 13276 -572 13964 -148
rect 14028 -572 14048 -148
rect 13276 -600 14048 -572
rect 14288 -148 15060 -120
rect 14288 -572 14976 -148
rect 15040 -572 15060 -148
rect 14288 -600 15060 -572
rect 15300 -148 16072 -120
rect 15300 -572 15988 -148
rect 16052 -572 16072 -148
rect 15300 -600 16072 -572
rect 16312 -148 17084 -120
rect 16312 -572 17000 -148
rect 17064 -572 17084 -148
rect 16312 -600 17084 -572
rect 17324 -148 18096 -120
rect 17324 -572 18012 -148
rect 18076 -572 18096 -148
rect 17324 -600 18096 -572
rect 18336 -148 19108 -120
rect 18336 -572 19024 -148
rect 19088 -572 19108 -148
rect 18336 -600 19108 -572
rect 19348 -148 20120 -120
rect 19348 -572 20036 -148
rect 20100 -572 20120 -148
rect 19348 -600 20120 -572
rect 20360 -148 21132 -120
rect 20360 -572 21048 -148
rect 21112 -572 21132 -148
rect 20360 -600 21132 -572
rect 21372 -148 22144 -120
rect 21372 -572 22060 -148
rect 22124 -572 22144 -148
rect 21372 -600 22144 -572
rect 22384 -148 23156 -120
rect 22384 -572 23072 -148
rect 23136 -572 23156 -148
rect 22384 -600 23156 -572
rect 23396 -148 24168 -120
rect 23396 -572 24084 -148
rect 24148 -572 24168 -148
rect 23396 -600 24168 -572
rect 24408 -148 25180 -120
rect 24408 -572 25096 -148
rect 25160 -572 25180 -148
rect 24408 -600 25180 -572
rect 25420 -148 26192 -120
rect 25420 -572 26108 -148
rect 26172 -572 26192 -148
rect 25420 -600 26192 -572
rect 26432 -148 27204 -120
rect 26432 -572 27120 -148
rect 27184 -572 27204 -148
rect 26432 -600 27204 -572
rect 27444 -148 28216 -120
rect 27444 -572 28132 -148
rect 28196 -572 28216 -148
rect 27444 -600 28216 -572
rect 28456 -148 29228 -120
rect 28456 -572 29144 -148
rect 29208 -572 29228 -148
rect 28456 -600 29228 -572
rect 29468 -148 30240 -120
rect 29468 -572 30156 -148
rect 30220 -572 30240 -148
rect 29468 -600 30240 -572
rect 30480 -148 31252 -120
rect 30480 -572 31168 -148
rect 31232 -572 31252 -148
rect 30480 -600 31252 -572
rect 31492 -148 32264 -120
rect 31492 -572 32180 -148
rect 32244 -572 32264 -148
rect 31492 -600 32264 -572
rect -32264 -868 -31492 -840
rect -32264 -1292 -31576 -868
rect -31512 -1292 -31492 -868
rect -32264 -1320 -31492 -1292
rect -31252 -868 -30480 -840
rect -31252 -1292 -30564 -868
rect -30500 -1292 -30480 -868
rect -31252 -1320 -30480 -1292
rect -30240 -868 -29468 -840
rect -30240 -1292 -29552 -868
rect -29488 -1292 -29468 -868
rect -30240 -1320 -29468 -1292
rect -29228 -868 -28456 -840
rect -29228 -1292 -28540 -868
rect -28476 -1292 -28456 -868
rect -29228 -1320 -28456 -1292
rect -28216 -868 -27444 -840
rect -28216 -1292 -27528 -868
rect -27464 -1292 -27444 -868
rect -28216 -1320 -27444 -1292
rect -27204 -868 -26432 -840
rect -27204 -1292 -26516 -868
rect -26452 -1292 -26432 -868
rect -27204 -1320 -26432 -1292
rect -26192 -868 -25420 -840
rect -26192 -1292 -25504 -868
rect -25440 -1292 -25420 -868
rect -26192 -1320 -25420 -1292
rect -25180 -868 -24408 -840
rect -25180 -1292 -24492 -868
rect -24428 -1292 -24408 -868
rect -25180 -1320 -24408 -1292
rect -24168 -868 -23396 -840
rect -24168 -1292 -23480 -868
rect -23416 -1292 -23396 -868
rect -24168 -1320 -23396 -1292
rect -23156 -868 -22384 -840
rect -23156 -1292 -22468 -868
rect -22404 -1292 -22384 -868
rect -23156 -1320 -22384 -1292
rect -22144 -868 -21372 -840
rect -22144 -1292 -21456 -868
rect -21392 -1292 -21372 -868
rect -22144 -1320 -21372 -1292
rect -21132 -868 -20360 -840
rect -21132 -1292 -20444 -868
rect -20380 -1292 -20360 -868
rect -21132 -1320 -20360 -1292
rect -20120 -868 -19348 -840
rect -20120 -1292 -19432 -868
rect -19368 -1292 -19348 -868
rect -20120 -1320 -19348 -1292
rect -19108 -868 -18336 -840
rect -19108 -1292 -18420 -868
rect -18356 -1292 -18336 -868
rect -19108 -1320 -18336 -1292
rect -18096 -868 -17324 -840
rect -18096 -1292 -17408 -868
rect -17344 -1292 -17324 -868
rect -18096 -1320 -17324 -1292
rect -17084 -868 -16312 -840
rect -17084 -1292 -16396 -868
rect -16332 -1292 -16312 -868
rect -17084 -1320 -16312 -1292
rect -16072 -868 -15300 -840
rect -16072 -1292 -15384 -868
rect -15320 -1292 -15300 -868
rect -16072 -1320 -15300 -1292
rect -15060 -868 -14288 -840
rect -15060 -1292 -14372 -868
rect -14308 -1292 -14288 -868
rect -15060 -1320 -14288 -1292
rect -14048 -868 -13276 -840
rect -14048 -1292 -13360 -868
rect -13296 -1292 -13276 -868
rect -14048 -1320 -13276 -1292
rect -13036 -868 -12264 -840
rect -13036 -1292 -12348 -868
rect -12284 -1292 -12264 -868
rect -13036 -1320 -12264 -1292
rect -12024 -868 -11252 -840
rect -12024 -1292 -11336 -868
rect -11272 -1292 -11252 -868
rect -12024 -1320 -11252 -1292
rect -11012 -868 -10240 -840
rect -11012 -1292 -10324 -868
rect -10260 -1292 -10240 -868
rect -11012 -1320 -10240 -1292
rect -10000 -868 -9228 -840
rect -10000 -1292 -9312 -868
rect -9248 -1292 -9228 -868
rect -10000 -1320 -9228 -1292
rect -8988 -868 -8216 -840
rect -8988 -1292 -8300 -868
rect -8236 -1292 -8216 -868
rect -8988 -1320 -8216 -1292
rect -7976 -868 -7204 -840
rect -7976 -1292 -7288 -868
rect -7224 -1292 -7204 -868
rect -7976 -1320 -7204 -1292
rect -6964 -868 -6192 -840
rect -6964 -1292 -6276 -868
rect -6212 -1292 -6192 -868
rect -6964 -1320 -6192 -1292
rect -5952 -868 -5180 -840
rect -5952 -1292 -5264 -868
rect -5200 -1292 -5180 -868
rect -5952 -1320 -5180 -1292
rect -4940 -868 -4168 -840
rect -4940 -1292 -4252 -868
rect -4188 -1292 -4168 -868
rect -4940 -1320 -4168 -1292
rect -3928 -868 -3156 -840
rect -3928 -1292 -3240 -868
rect -3176 -1292 -3156 -868
rect -3928 -1320 -3156 -1292
rect -2916 -868 -2144 -840
rect -2916 -1292 -2228 -868
rect -2164 -1292 -2144 -868
rect -2916 -1320 -2144 -1292
rect -1904 -868 -1132 -840
rect -1904 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -1904 -1320 -1132 -1292
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect 1132 -868 1904 -840
rect 1132 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 1132 -1320 1904 -1292
rect 2144 -868 2916 -840
rect 2144 -1292 2832 -868
rect 2896 -1292 2916 -868
rect 2144 -1320 2916 -1292
rect 3156 -868 3928 -840
rect 3156 -1292 3844 -868
rect 3908 -1292 3928 -868
rect 3156 -1320 3928 -1292
rect 4168 -868 4940 -840
rect 4168 -1292 4856 -868
rect 4920 -1292 4940 -868
rect 4168 -1320 4940 -1292
rect 5180 -868 5952 -840
rect 5180 -1292 5868 -868
rect 5932 -1292 5952 -868
rect 5180 -1320 5952 -1292
rect 6192 -868 6964 -840
rect 6192 -1292 6880 -868
rect 6944 -1292 6964 -868
rect 6192 -1320 6964 -1292
rect 7204 -868 7976 -840
rect 7204 -1292 7892 -868
rect 7956 -1292 7976 -868
rect 7204 -1320 7976 -1292
rect 8216 -868 8988 -840
rect 8216 -1292 8904 -868
rect 8968 -1292 8988 -868
rect 8216 -1320 8988 -1292
rect 9228 -868 10000 -840
rect 9228 -1292 9916 -868
rect 9980 -1292 10000 -868
rect 9228 -1320 10000 -1292
rect 10240 -868 11012 -840
rect 10240 -1292 10928 -868
rect 10992 -1292 11012 -868
rect 10240 -1320 11012 -1292
rect 11252 -868 12024 -840
rect 11252 -1292 11940 -868
rect 12004 -1292 12024 -868
rect 11252 -1320 12024 -1292
rect 12264 -868 13036 -840
rect 12264 -1292 12952 -868
rect 13016 -1292 13036 -868
rect 12264 -1320 13036 -1292
rect 13276 -868 14048 -840
rect 13276 -1292 13964 -868
rect 14028 -1292 14048 -868
rect 13276 -1320 14048 -1292
rect 14288 -868 15060 -840
rect 14288 -1292 14976 -868
rect 15040 -1292 15060 -868
rect 14288 -1320 15060 -1292
rect 15300 -868 16072 -840
rect 15300 -1292 15988 -868
rect 16052 -1292 16072 -868
rect 15300 -1320 16072 -1292
rect 16312 -868 17084 -840
rect 16312 -1292 17000 -868
rect 17064 -1292 17084 -868
rect 16312 -1320 17084 -1292
rect 17324 -868 18096 -840
rect 17324 -1292 18012 -868
rect 18076 -1292 18096 -868
rect 17324 -1320 18096 -1292
rect 18336 -868 19108 -840
rect 18336 -1292 19024 -868
rect 19088 -1292 19108 -868
rect 18336 -1320 19108 -1292
rect 19348 -868 20120 -840
rect 19348 -1292 20036 -868
rect 20100 -1292 20120 -868
rect 19348 -1320 20120 -1292
rect 20360 -868 21132 -840
rect 20360 -1292 21048 -868
rect 21112 -1292 21132 -868
rect 20360 -1320 21132 -1292
rect 21372 -868 22144 -840
rect 21372 -1292 22060 -868
rect 22124 -1292 22144 -868
rect 21372 -1320 22144 -1292
rect 22384 -868 23156 -840
rect 22384 -1292 23072 -868
rect 23136 -1292 23156 -868
rect 22384 -1320 23156 -1292
rect 23396 -868 24168 -840
rect 23396 -1292 24084 -868
rect 24148 -1292 24168 -868
rect 23396 -1320 24168 -1292
rect 24408 -868 25180 -840
rect 24408 -1292 25096 -868
rect 25160 -1292 25180 -868
rect 24408 -1320 25180 -1292
rect 25420 -868 26192 -840
rect 25420 -1292 26108 -868
rect 26172 -1292 26192 -868
rect 25420 -1320 26192 -1292
rect 26432 -868 27204 -840
rect 26432 -1292 27120 -868
rect 27184 -1292 27204 -868
rect 26432 -1320 27204 -1292
rect 27444 -868 28216 -840
rect 27444 -1292 28132 -868
rect 28196 -1292 28216 -868
rect 27444 -1320 28216 -1292
rect 28456 -868 29228 -840
rect 28456 -1292 29144 -868
rect 29208 -1292 29228 -868
rect 28456 -1320 29228 -1292
rect 29468 -868 30240 -840
rect 29468 -1292 30156 -868
rect 30220 -1292 30240 -868
rect 29468 -1320 30240 -1292
rect 30480 -868 31252 -840
rect 30480 -1292 31168 -868
rect 31232 -1292 31252 -868
rect 30480 -1320 31252 -1292
rect 31492 -868 32264 -840
rect 31492 -1292 32180 -868
rect 32244 -1292 32264 -868
rect 31492 -1320 32264 -1292
rect -32264 -1588 -31492 -1560
rect -32264 -2012 -31576 -1588
rect -31512 -2012 -31492 -1588
rect -32264 -2040 -31492 -2012
rect -31252 -1588 -30480 -1560
rect -31252 -2012 -30564 -1588
rect -30500 -2012 -30480 -1588
rect -31252 -2040 -30480 -2012
rect -30240 -1588 -29468 -1560
rect -30240 -2012 -29552 -1588
rect -29488 -2012 -29468 -1588
rect -30240 -2040 -29468 -2012
rect -29228 -1588 -28456 -1560
rect -29228 -2012 -28540 -1588
rect -28476 -2012 -28456 -1588
rect -29228 -2040 -28456 -2012
rect -28216 -1588 -27444 -1560
rect -28216 -2012 -27528 -1588
rect -27464 -2012 -27444 -1588
rect -28216 -2040 -27444 -2012
rect -27204 -1588 -26432 -1560
rect -27204 -2012 -26516 -1588
rect -26452 -2012 -26432 -1588
rect -27204 -2040 -26432 -2012
rect -26192 -1588 -25420 -1560
rect -26192 -2012 -25504 -1588
rect -25440 -2012 -25420 -1588
rect -26192 -2040 -25420 -2012
rect -25180 -1588 -24408 -1560
rect -25180 -2012 -24492 -1588
rect -24428 -2012 -24408 -1588
rect -25180 -2040 -24408 -2012
rect -24168 -1588 -23396 -1560
rect -24168 -2012 -23480 -1588
rect -23416 -2012 -23396 -1588
rect -24168 -2040 -23396 -2012
rect -23156 -1588 -22384 -1560
rect -23156 -2012 -22468 -1588
rect -22404 -2012 -22384 -1588
rect -23156 -2040 -22384 -2012
rect -22144 -1588 -21372 -1560
rect -22144 -2012 -21456 -1588
rect -21392 -2012 -21372 -1588
rect -22144 -2040 -21372 -2012
rect -21132 -1588 -20360 -1560
rect -21132 -2012 -20444 -1588
rect -20380 -2012 -20360 -1588
rect -21132 -2040 -20360 -2012
rect -20120 -1588 -19348 -1560
rect -20120 -2012 -19432 -1588
rect -19368 -2012 -19348 -1588
rect -20120 -2040 -19348 -2012
rect -19108 -1588 -18336 -1560
rect -19108 -2012 -18420 -1588
rect -18356 -2012 -18336 -1588
rect -19108 -2040 -18336 -2012
rect -18096 -1588 -17324 -1560
rect -18096 -2012 -17408 -1588
rect -17344 -2012 -17324 -1588
rect -18096 -2040 -17324 -2012
rect -17084 -1588 -16312 -1560
rect -17084 -2012 -16396 -1588
rect -16332 -2012 -16312 -1588
rect -17084 -2040 -16312 -2012
rect -16072 -1588 -15300 -1560
rect -16072 -2012 -15384 -1588
rect -15320 -2012 -15300 -1588
rect -16072 -2040 -15300 -2012
rect -15060 -1588 -14288 -1560
rect -15060 -2012 -14372 -1588
rect -14308 -2012 -14288 -1588
rect -15060 -2040 -14288 -2012
rect -14048 -1588 -13276 -1560
rect -14048 -2012 -13360 -1588
rect -13296 -2012 -13276 -1588
rect -14048 -2040 -13276 -2012
rect -13036 -1588 -12264 -1560
rect -13036 -2012 -12348 -1588
rect -12284 -2012 -12264 -1588
rect -13036 -2040 -12264 -2012
rect -12024 -1588 -11252 -1560
rect -12024 -2012 -11336 -1588
rect -11272 -2012 -11252 -1588
rect -12024 -2040 -11252 -2012
rect -11012 -1588 -10240 -1560
rect -11012 -2012 -10324 -1588
rect -10260 -2012 -10240 -1588
rect -11012 -2040 -10240 -2012
rect -10000 -1588 -9228 -1560
rect -10000 -2012 -9312 -1588
rect -9248 -2012 -9228 -1588
rect -10000 -2040 -9228 -2012
rect -8988 -1588 -8216 -1560
rect -8988 -2012 -8300 -1588
rect -8236 -2012 -8216 -1588
rect -8988 -2040 -8216 -2012
rect -7976 -1588 -7204 -1560
rect -7976 -2012 -7288 -1588
rect -7224 -2012 -7204 -1588
rect -7976 -2040 -7204 -2012
rect -6964 -1588 -6192 -1560
rect -6964 -2012 -6276 -1588
rect -6212 -2012 -6192 -1588
rect -6964 -2040 -6192 -2012
rect -5952 -1588 -5180 -1560
rect -5952 -2012 -5264 -1588
rect -5200 -2012 -5180 -1588
rect -5952 -2040 -5180 -2012
rect -4940 -1588 -4168 -1560
rect -4940 -2012 -4252 -1588
rect -4188 -2012 -4168 -1588
rect -4940 -2040 -4168 -2012
rect -3928 -1588 -3156 -1560
rect -3928 -2012 -3240 -1588
rect -3176 -2012 -3156 -1588
rect -3928 -2040 -3156 -2012
rect -2916 -1588 -2144 -1560
rect -2916 -2012 -2228 -1588
rect -2164 -2012 -2144 -1588
rect -2916 -2040 -2144 -2012
rect -1904 -1588 -1132 -1560
rect -1904 -2012 -1216 -1588
rect -1152 -2012 -1132 -1588
rect -1904 -2040 -1132 -2012
rect -892 -1588 -120 -1560
rect -892 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect -892 -2040 -120 -2012
rect 120 -1588 892 -1560
rect 120 -2012 808 -1588
rect 872 -2012 892 -1588
rect 120 -2040 892 -2012
rect 1132 -1588 1904 -1560
rect 1132 -2012 1820 -1588
rect 1884 -2012 1904 -1588
rect 1132 -2040 1904 -2012
rect 2144 -1588 2916 -1560
rect 2144 -2012 2832 -1588
rect 2896 -2012 2916 -1588
rect 2144 -2040 2916 -2012
rect 3156 -1588 3928 -1560
rect 3156 -2012 3844 -1588
rect 3908 -2012 3928 -1588
rect 3156 -2040 3928 -2012
rect 4168 -1588 4940 -1560
rect 4168 -2012 4856 -1588
rect 4920 -2012 4940 -1588
rect 4168 -2040 4940 -2012
rect 5180 -1588 5952 -1560
rect 5180 -2012 5868 -1588
rect 5932 -2012 5952 -1588
rect 5180 -2040 5952 -2012
rect 6192 -1588 6964 -1560
rect 6192 -2012 6880 -1588
rect 6944 -2012 6964 -1588
rect 6192 -2040 6964 -2012
rect 7204 -1588 7976 -1560
rect 7204 -2012 7892 -1588
rect 7956 -2012 7976 -1588
rect 7204 -2040 7976 -2012
rect 8216 -1588 8988 -1560
rect 8216 -2012 8904 -1588
rect 8968 -2012 8988 -1588
rect 8216 -2040 8988 -2012
rect 9228 -1588 10000 -1560
rect 9228 -2012 9916 -1588
rect 9980 -2012 10000 -1588
rect 9228 -2040 10000 -2012
rect 10240 -1588 11012 -1560
rect 10240 -2012 10928 -1588
rect 10992 -2012 11012 -1588
rect 10240 -2040 11012 -2012
rect 11252 -1588 12024 -1560
rect 11252 -2012 11940 -1588
rect 12004 -2012 12024 -1588
rect 11252 -2040 12024 -2012
rect 12264 -1588 13036 -1560
rect 12264 -2012 12952 -1588
rect 13016 -2012 13036 -1588
rect 12264 -2040 13036 -2012
rect 13276 -1588 14048 -1560
rect 13276 -2012 13964 -1588
rect 14028 -2012 14048 -1588
rect 13276 -2040 14048 -2012
rect 14288 -1588 15060 -1560
rect 14288 -2012 14976 -1588
rect 15040 -2012 15060 -1588
rect 14288 -2040 15060 -2012
rect 15300 -1588 16072 -1560
rect 15300 -2012 15988 -1588
rect 16052 -2012 16072 -1588
rect 15300 -2040 16072 -2012
rect 16312 -1588 17084 -1560
rect 16312 -2012 17000 -1588
rect 17064 -2012 17084 -1588
rect 16312 -2040 17084 -2012
rect 17324 -1588 18096 -1560
rect 17324 -2012 18012 -1588
rect 18076 -2012 18096 -1588
rect 17324 -2040 18096 -2012
rect 18336 -1588 19108 -1560
rect 18336 -2012 19024 -1588
rect 19088 -2012 19108 -1588
rect 18336 -2040 19108 -2012
rect 19348 -1588 20120 -1560
rect 19348 -2012 20036 -1588
rect 20100 -2012 20120 -1588
rect 19348 -2040 20120 -2012
rect 20360 -1588 21132 -1560
rect 20360 -2012 21048 -1588
rect 21112 -2012 21132 -1588
rect 20360 -2040 21132 -2012
rect 21372 -1588 22144 -1560
rect 21372 -2012 22060 -1588
rect 22124 -2012 22144 -1588
rect 21372 -2040 22144 -2012
rect 22384 -1588 23156 -1560
rect 22384 -2012 23072 -1588
rect 23136 -2012 23156 -1588
rect 22384 -2040 23156 -2012
rect 23396 -1588 24168 -1560
rect 23396 -2012 24084 -1588
rect 24148 -2012 24168 -1588
rect 23396 -2040 24168 -2012
rect 24408 -1588 25180 -1560
rect 24408 -2012 25096 -1588
rect 25160 -2012 25180 -1588
rect 24408 -2040 25180 -2012
rect 25420 -1588 26192 -1560
rect 25420 -2012 26108 -1588
rect 26172 -2012 26192 -1588
rect 25420 -2040 26192 -2012
rect 26432 -1588 27204 -1560
rect 26432 -2012 27120 -1588
rect 27184 -2012 27204 -1588
rect 26432 -2040 27204 -2012
rect 27444 -1588 28216 -1560
rect 27444 -2012 28132 -1588
rect 28196 -2012 28216 -1588
rect 27444 -2040 28216 -2012
rect 28456 -1588 29228 -1560
rect 28456 -2012 29144 -1588
rect 29208 -2012 29228 -1588
rect 28456 -2040 29228 -2012
rect 29468 -1588 30240 -1560
rect 29468 -2012 30156 -1588
rect 30220 -2012 30240 -1588
rect 29468 -2040 30240 -2012
rect 30480 -1588 31252 -1560
rect 30480 -2012 31168 -1588
rect 31232 -2012 31252 -1588
rect 30480 -2040 31252 -2012
rect 31492 -1588 32264 -1560
rect 31492 -2012 32180 -1588
rect 32244 -2012 32264 -1588
rect 31492 -2040 32264 -2012
rect -32264 -2308 -31492 -2280
rect -32264 -2732 -31576 -2308
rect -31512 -2732 -31492 -2308
rect -32264 -2760 -31492 -2732
rect -31252 -2308 -30480 -2280
rect -31252 -2732 -30564 -2308
rect -30500 -2732 -30480 -2308
rect -31252 -2760 -30480 -2732
rect -30240 -2308 -29468 -2280
rect -30240 -2732 -29552 -2308
rect -29488 -2732 -29468 -2308
rect -30240 -2760 -29468 -2732
rect -29228 -2308 -28456 -2280
rect -29228 -2732 -28540 -2308
rect -28476 -2732 -28456 -2308
rect -29228 -2760 -28456 -2732
rect -28216 -2308 -27444 -2280
rect -28216 -2732 -27528 -2308
rect -27464 -2732 -27444 -2308
rect -28216 -2760 -27444 -2732
rect -27204 -2308 -26432 -2280
rect -27204 -2732 -26516 -2308
rect -26452 -2732 -26432 -2308
rect -27204 -2760 -26432 -2732
rect -26192 -2308 -25420 -2280
rect -26192 -2732 -25504 -2308
rect -25440 -2732 -25420 -2308
rect -26192 -2760 -25420 -2732
rect -25180 -2308 -24408 -2280
rect -25180 -2732 -24492 -2308
rect -24428 -2732 -24408 -2308
rect -25180 -2760 -24408 -2732
rect -24168 -2308 -23396 -2280
rect -24168 -2732 -23480 -2308
rect -23416 -2732 -23396 -2308
rect -24168 -2760 -23396 -2732
rect -23156 -2308 -22384 -2280
rect -23156 -2732 -22468 -2308
rect -22404 -2732 -22384 -2308
rect -23156 -2760 -22384 -2732
rect -22144 -2308 -21372 -2280
rect -22144 -2732 -21456 -2308
rect -21392 -2732 -21372 -2308
rect -22144 -2760 -21372 -2732
rect -21132 -2308 -20360 -2280
rect -21132 -2732 -20444 -2308
rect -20380 -2732 -20360 -2308
rect -21132 -2760 -20360 -2732
rect -20120 -2308 -19348 -2280
rect -20120 -2732 -19432 -2308
rect -19368 -2732 -19348 -2308
rect -20120 -2760 -19348 -2732
rect -19108 -2308 -18336 -2280
rect -19108 -2732 -18420 -2308
rect -18356 -2732 -18336 -2308
rect -19108 -2760 -18336 -2732
rect -18096 -2308 -17324 -2280
rect -18096 -2732 -17408 -2308
rect -17344 -2732 -17324 -2308
rect -18096 -2760 -17324 -2732
rect -17084 -2308 -16312 -2280
rect -17084 -2732 -16396 -2308
rect -16332 -2732 -16312 -2308
rect -17084 -2760 -16312 -2732
rect -16072 -2308 -15300 -2280
rect -16072 -2732 -15384 -2308
rect -15320 -2732 -15300 -2308
rect -16072 -2760 -15300 -2732
rect -15060 -2308 -14288 -2280
rect -15060 -2732 -14372 -2308
rect -14308 -2732 -14288 -2308
rect -15060 -2760 -14288 -2732
rect -14048 -2308 -13276 -2280
rect -14048 -2732 -13360 -2308
rect -13296 -2732 -13276 -2308
rect -14048 -2760 -13276 -2732
rect -13036 -2308 -12264 -2280
rect -13036 -2732 -12348 -2308
rect -12284 -2732 -12264 -2308
rect -13036 -2760 -12264 -2732
rect -12024 -2308 -11252 -2280
rect -12024 -2732 -11336 -2308
rect -11272 -2732 -11252 -2308
rect -12024 -2760 -11252 -2732
rect -11012 -2308 -10240 -2280
rect -11012 -2732 -10324 -2308
rect -10260 -2732 -10240 -2308
rect -11012 -2760 -10240 -2732
rect -10000 -2308 -9228 -2280
rect -10000 -2732 -9312 -2308
rect -9248 -2732 -9228 -2308
rect -10000 -2760 -9228 -2732
rect -8988 -2308 -8216 -2280
rect -8988 -2732 -8300 -2308
rect -8236 -2732 -8216 -2308
rect -8988 -2760 -8216 -2732
rect -7976 -2308 -7204 -2280
rect -7976 -2732 -7288 -2308
rect -7224 -2732 -7204 -2308
rect -7976 -2760 -7204 -2732
rect -6964 -2308 -6192 -2280
rect -6964 -2732 -6276 -2308
rect -6212 -2732 -6192 -2308
rect -6964 -2760 -6192 -2732
rect -5952 -2308 -5180 -2280
rect -5952 -2732 -5264 -2308
rect -5200 -2732 -5180 -2308
rect -5952 -2760 -5180 -2732
rect -4940 -2308 -4168 -2280
rect -4940 -2732 -4252 -2308
rect -4188 -2732 -4168 -2308
rect -4940 -2760 -4168 -2732
rect -3928 -2308 -3156 -2280
rect -3928 -2732 -3240 -2308
rect -3176 -2732 -3156 -2308
rect -3928 -2760 -3156 -2732
rect -2916 -2308 -2144 -2280
rect -2916 -2732 -2228 -2308
rect -2164 -2732 -2144 -2308
rect -2916 -2760 -2144 -2732
rect -1904 -2308 -1132 -2280
rect -1904 -2732 -1216 -2308
rect -1152 -2732 -1132 -2308
rect -1904 -2760 -1132 -2732
rect -892 -2308 -120 -2280
rect -892 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect -892 -2760 -120 -2732
rect 120 -2308 892 -2280
rect 120 -2732 808 -2308
rect 872 -2732 892 -2308
rect 120 -2760 892 -2732
rect 1132 -2308 1904 -2280
rect 1132 -2732 1820 -2308
rect 1884 -2732 1904 -2308
rect 1132 -2760 1904 -2732
rect 2144 -2308 2916 -2280
rect 2144 -2732 2832 -2308
rect 2896 -2732 2916 -2308
rect 2144 -2760 2916 -2732
rect 3156 -2308 3928 -2280
rect 3156 -2732 3844 -2308
rect 3908 -2732 3928 -2308
rect 3156 -2760 3928 -2732
rect 4168 -2308 4940 -2280
rect 4168 -2732 4856 -2308
rect 4920 -2732 4940 -2308
rect 4168 -2760 4940 -2732
rect 5180 -2308 5952 -2280
rect 5180 -2732 5868 -2308
rect 5932 -2732 5952 -2308
rect 5180 -2760 5952 -2732
rect 6192 -2308 6964 -2280
rect 6192 -2732 6880 -2308
rect 6944 -2732 6964 -2308
rect 6192 -2760 6964 -2732
rect 7204 -2308 7976 -2280
rect 7204 -2732 7892 -2308
rect 7956 -2732 7976 -2308
rect 7204 -2760 7976 -2732
rect 8216 -2308 8988 -2280
rect 8216 -2732 8904 -2308
rect 8968 -2732 8988 -2308
rect 8216 -2760 8988 -2732
rect 9228 -2308 10000 -2280
rect 9228 -2732 9916 -2308
rect 9980 -2732 10000 -2308
rect 9228 -2760 10000 -2732
rect 10240 -2308 11012 -2280
rect 10240 -2732 10928 -2308
rect 10992 -2732 11012 -2308
rect 10240 -2760 11012 -2732
rect 11252 -2308 12024 -2280
rect 11252 -2732 11940 -2308
rect 12004 -2732 12024 -2308
rect 11252 -2760 12024 -2732
rect 12264 -2308 13036 -2280
rect 12264 -2732 12952 -2308
rect 13016 -2732 13036 -2308
rect 12264 -2760 13036 -2732
rect 13276 -2308 14048 -2280
rect 13276 -2732 13964 -2308
rect 14028 -2732 14048 -2308
rect 13276 -2760 14048 -2732
rect 14288 -2308 15060 -2280
rect 14288 -2732 14976 -2308
rect 15040 -2732 15060 -2308
rect 14288 -2760 15060 -2732
rect 15300 -2308 16072 -2280
rect 15300 -2732 15988 -2308
rect 16052 -2732 16072 -2308
rect 15300 -2760 16072 -2732
rect 16312 -2308 17084 -2280
rect 16312 -2732 17000 -2308
rect 17064 -2732 17084 -2308
rect 16312 -2760 17084 -2732
rect 17324 -2308 18096 -2280
rect 17324 -2732 18012 -2308
rect 18076 -2732 18096 -2308
rect 17324 -2760 18096 -2732
rect 18336 -2308 19108 -2280
rect 18336 -2732 19024 -2308
rect 19088 -2732 19108 -2308
rect 18336 -2760 19108 -2732
rect 19348 -2308 20120 -2280
rect 19348 -2732 20036 -2308
rect 20100 -2732 20120 -2308
rect 19348 -2760 20120 -2732
rect 20360 -2308 21132 -2280
rect 20360 -2732 21048 -2308
rect 21112 -2732 21132 -2308
rect 20360 -2760 21132 -2732
rect 21372 -2308 22144 -2280
rect 21372 -2732 22060 -2308
rect 22124 -2732 22144 -2308
rect 21372 -2760 22144 -2732
rect 22384 -2308 23156 -2280
rect 22384 -2732 23072 -2308
rect 23136 -2732 23156 -2308
rect 22384 -2760 23156 -2732
rect 23396 -2308 24168 -2280
rect 23396 -2732 24084 -2308
rect 24148 -2732 24168 -2308
rect 23396 -2760 24168 -2732
rect 24408 -2308 25180 -2280
rect 24408 -2732 25096 -2308
rect 25160 -2732 25180 -2308
rect 24408 -2760 25180 -2732
rect 25420 -2308 26192 -2280
rect 25420 -2732 26108 -2308
rect 26172 -2732 26192 -2308
rect 25420 -2760 26192 -2732
rect 26432 -2308 27204 -2280
rect 26432 -2732 27120 -2308
rect 27184 -2732 27204 -2308
rect 26432 -2760 27204 -2732
rect 27444 -2308 28216 -2280
rect 27444 -2732 28132 -2308
rect 28196 -2732 28216 -2308
rect 27444 -2760 28216 -2732
rect 28456 -2308 29228 -2280
rect 28456 -2732 29144 -2308
rect 29208 -2732 29228 -2308
rect 28456 -2760 29228 -2732
rect 29468 -2308 30240 -2280
rect 29468 -2732 30156 -2308
rect 30220 -2732 30240 -2308
rect 29468 -2760 30240 -2732
rect 30480 -2308 31252 -2280
rect 30480 -2732 31168 -2308
rect 31232 -2732 31252 -2308
rect 30480 -2760 31252 -2732
rect 31492 -2308 32264 -2280
rect 31492 -2732 32180 -2308
rect 32244 -2732 32264 -2308
rect 31492 -2760 32264 -2732
rect -32264 -3028 -31492 -3000
rect -32264 -3452 -31576 -3028
rect -31512 -3452 -31492 -3028
rect -32264 -3480 -31492 -3452
rect -31252 -3028 -30480 -3000
rect -31252 -3452 -30564 -3028
rect -30500 -3452 -30480 -3028
rect -31252 -3480 -30480 -3452
rect -30240 -3028 -29468 -3000
rect -30240 -3452 -29552 -3028
rect -29488 -3452 -29468 -3028
rect -30240 -3480 -29468 -3452
rect -29228 -3028 -28456 -3000
rect -29228 -3452 -28540 -3028
rect -28476 -3452 -28456 -3028
rect -29228 -3480 -28456 -3452
rect -28216 -3028 -27444 -3000
rect -28216 -3452 -27528 -3028
rect -27464 -3452 -27444 -3028
rect -28216 -3480 -27444 -3452
rect -27204 -3028 -26432 -3000
rect -27204 -3452 -26516 -3028
rect -26452 -3452 -26432 -3028
rect -27204 -3480 -26432 -3452
rect -26192 -3028 -25420 -3000
rect -26192 -3452 -25504 -3028
rect -25440 -3452 -25420 -3028
rect -26192 -3480 -25420 -3452
rect -25180 -3028 -24408 -3000
rect -25180 -3452 -24492 -3028
rect -24428 -3452 -24408 -3028
rect -25180 -3480 -24408 -3452
rect -24168 -3028 -23396 -3000
rect -24168 -3452 -23480 -3028
rect -23416 -3452 -23396 -3028
rect -24168 -3480 -23396 -3452
rect -23156 -3028 -22384 -3000
rect -23156 -3452 -22468 -3028
rect -22404 -3452 -22384 -3028
rect -23156 -3480 -22384 -3452
rect -22144 -3028 -21372 -3000
rect -22144 -3452 -21456 -3028
rect -21392 -3452 -21372 -3028
rect -22144 -3480 -21372 -3452
rect -21132 -3028 -20360 -3000
rect -21132 -3452 -20444 -3028
rect -20380 -3452 -20360 -3028
rect -21132 -3480 -20360 -3452
rect -20120 -3028 -19348 -3000
rect -20120 -3452 -19432 -3028
rect -19368 -3452 -19348 -3028
rect -20120 -3480 -19348 -3452
rect -19108 -3028 -18336 -3000
rect -19108 -3452 -18420 -3028
rect -18356 -3452 -18336 -3028
rect -19108 -3480 -18336 -3452
rect -18096 -3028 -17324 -3000
rect -18096 -3452 -17408 -3028
rect -17344 -3452 -17324 -3028
rect -18096 -3480 -17324 -3452
rect -17084 -3028 -16312 -3000
rect -17084 -3452 -16396 -3028
rect -16332 -3452 -16312 -3028
rect -17084 -3480 -16312 -3452
rect -16072 -3028 -15300 -3000
rect -16072 -3452 -15384 -3028
rect -15320 -3452 -15300 -3028
rect -16072 -3480 -15300 -3452
rect -15060 -3028 -14288 -3000
rect -15060 -3452 -14372 -3028
rect -14308 -3452 -14288 -3028
rect -15060 -3480 -14288 -3452
rect -14048 -3028 -13276 -3000
rect -14048 -3452 -13360 -3028
rect -13296 -3452 -13276 -3028
rect -14048 -3480 -13276 -3452
rect -13036 -3028 -12264 -3000
rect -13036 -3452 -12348 -3028
rect -12284 -3452 -12264 -3028
rect -13036 -3480 -12264 -3452
rect -12024 -3028 -11252 -3000
rect -12024 -3452 -11336 -3028
rect -11272 -3452 -11252 -3028
rect -12024 -3480 -11252 -3452
rect -11012 -3028 -10240 -3000
rect -11012 -3452 -10324 -3028
rect -10260 -3452 -10240 -3028
rect -11012 -3480 -10240 -3452
rect -10000 -3028 -9228 -3000
rect -10000 -3452 -9312 -3028
rect -9248 -3452 -9228 -3028
rect -10000 -3480 -9228 -3452
rect -8988 -3028 -8216 -3000
rect -8988 -3452 -8300 -3028
rect -8236 -3452 -8216 -3028
rect -8988 -3480 -8216 -3452
rect -7976 -3028 -7204 -3000
rect -7976 -3452 -7288 -3028
rect -7224 -3452 -7204 -3028
rect -7976 -3480 -7204 -3452
rect -6964 -3028 -6192 -3000
rect -6964 -3452 -6276 -3028
rect -6212 -3452 -6192 -3028
rect -6964 -3480 -6192 -3452
rect -5952 -3028 -5180 -3000
rect -5952 -3452 -5264 -3028
rect -5200 -3452 -5180 -3028
rect -5952 -3480 -5180 -3452
rect -4940 -3028 -4168 -3000
rect -4940 -3452 -4252 -3028
rect -4188 -3452 -4168 -3028
rect -4940 -3480 -4168 -3452
rect -3928 -3028 -3156 -3000
rect -3928 -3452 -3240 -3028
rect -3176 -3452 -3156 -3028
rect -3928 -3480 -3156 -3452
rect -2916 -3028 -2144 -3000
rect -2916 -3452 -2228 -3028
rect -2164 -3452 -2144 -3028
rect -2916 -3480 -2144 -3452
rect -1904 -3028 -1132 -3000
rect -1904 -3452 -1216 -3028
rect -1152 -3452 -1132 -3028
rect -1904 -3480 -1132 -3452
rect -892 -3028 -120 -3000
rect -892 -3452 -204 -3028
rect -140 -3452 -120 -3028
rect -892 -3480 -120 -3452
rect 120 -3028 892 -3000
rect 120 -3452 808 -3028
rect 872 -3452 892 -3028
rect 120 -3480 892 -3452
rect 1132 -3028 1904 -3000
rect 1132 -3452 1820 -3028
rect 1884 -3452 1904 -3028
rect 1132 -3480 1904 -3452
rect 2144 -3028 2916 -3000
rect 2144 -3452 2832 -3028
rect 2896 -3452 2916 -3028
rect 2144 -3480 2916 -3452
rect 3156 -3028 3928 -3000
rect 3156 -3452 3844 -3028
rect 3908 -3452 3928 -3028
rect 3156 -3480 3928 -3452
rect 4168 -3028 4940 -3000
rect 4168 -3452 4856 -3028
rect 4920 -3452 4940 -3028
rect 4168 -3480 4940 -3452
rect 5180 -3028 5952 -3000
rect 5180 -3452 5868 -3028
rect 5932 -3452 5952 -3028
rect 5180 -3480 5952 -3452
rect 6192 -3028 6964 -3000
rect 6192 -3452 6880 -3028
rect 6944 -3452 6964 -3028
rect 6192 -3480 6964 -3452
rect 7204 -3028 7976 -3000
rect 7204 -3452 7892 -3028
rect 7956 -3452 7976 -3028
rect 7204 -3480 7976 -3452
rect 8216 -3028 8988 -3000
rect 8216 -3452 8904 -3028
rect 8968 -3452 8988 -3028
rect 8216 -3480 8988 -3452
rect 9228 -3028 10000 -3000
rect 9228 -3452 9916 -3028
rect 9980 -3452 10000 -3028
rect 9228 -3480 10000 -3452
rect 10240 -3028 11012 -3000
rect 10240 -3452 10928 -3028
rect 10992 -3452 11012 -3028
rect 10240 -3480 11012 -3452
rect 11252 -3028 12024 -3000
rect 11252 -3452 11940 -3028
rect 12004 -3452 12024 -3028
rect 11252 -3480 12024 -3452
rect 12264 -3028 13036 -3000
rect 12264 -3452 12952 -3028
rect 13016 -3452 13036 -3028
rect 12264 -3480 13036 -3452
rect 13276 -3028 14048 -3000
rect 13276 -3452 13964 -3028
rect 14028 -3452 14048 -3028
rect 13276 -3480 14048 -3452
rect 14288 -3028 15060 -3000
rect 14288 -3452 14976 -3028
rect 15040 -3452 15060 -3028
rect 14288 -3480 15060 -3452
rect 15300 -3028 16072 -3000
rect 15300 -3452 15988 -3028
rect 16052 -3452 16072 -3028
rect 15300 -3480 16072 -3452
rect 16312 -3028 17084 -3000
rect 16312 -3452 17000 -3028
rect 17064 -3452 17084 -3028
rect 16312 -3480 17084 -3452
rect 17324 -3028 18096 -3000
rect 17324 -3452 18012 -3028
rect 18076 -3452 18096 -3028
rect 17324 -3480 18096 -3452
rect 18336 -3028 19108 -3000
rect 18336 -3452 19024 -3028
rect 19088 -3452 19108 -3028
rect 18336 -3480 19108 -3452
rect 19348 -3028 20120 -3000
rect 19348 -3452 20036 -3028
rect 20100 -3452 20120 -3028
rect 19348 -3480 20120 -3452
rect 20360 -3028 21132 -3000
rect 20360 -3452 21048 -3028
rect 21112 -3452 21132 -3028
rect 20360 -3480 21132 -3452
rect 21372 -3028 22144 -3000
rect 21372 -3452 22060 -3028
rect 22124 -3452 22144 -3028
rect 21372 -3480 22144 -3452
rect 22384 -3028 23156 -3000
rect 22384 -3452 23072 -3028
rect 23136 -3452 23156 -3028
rect 22384 -3480 23156 -3452
rect 23396 -3028 24168 -3000
rect 23396 -3452 24084 -3028
rect 24148 -3452 24168 -3028
rect 23396 -3480 24168 -3452
rect 24408 -3028 25180 -3000
rect 24408 -3452 25096 -3028
rect 25160 -3452 25180 -3028
rect 24408 -3480 25180 -3452
rect 25420 -3028 26192 -3000
rect 25420 -3452 26108 -3028
rect 26172 -3452 26192 -3028
rect 25420 -3480 26192 -3452
rect 26432 -3028 27204 -3000
rect 26432 -3452 27120 -3028
rect 27184 -3452 27204 -3028
rect 26432 -3480 27204 -3452
rect 27444 -3028 28216 -3000
rect 27444 -3452 28132 -3028
rect 28196 -3452 28216 -3028
rect 27444 -3480 28216 -3452
rect 28456 -3028 29228 -3000
rect 28456 -3452 29144 -3028
rect 29208 -3452 29228 -3028
rect 28456 -3480 29228 -3452
rect 29468 -3028 30240 -3000
rect 29468 -3452 30156 -3028
rect 30220 -3452 30240 -3028
rect 29468 -3480 30240 -3452
rect 30480 -3028 31252 -3000
rect 30480 -3452 31168 -3028
rect 31232 -3452 31252 -3028
rect 30480 -3480 31252 -3452
rect 31492 -3028 32264 -3000
rect 31492 -3452 32180 -3028
rect 32244 -3452 32264 -3028
rect 31492 -3480 32264 -3452
rect -32264 -3748 -31492 -3720
rect -32264 -4172 -31576 -3748
rect -31512 -4172 -31492 -3748
rect -32264 -4200 -31492 -4172
rect -31252 -3748 -30480 -3720
rect -31252 -4172 -30564 -3748
rect -30500 -4172 -30480 -3748
rect -31252 -4200 -30480 -4172
rect -30240 -3748 -29468 -3720
rect -30240 -4172 -29552 -3748
rect -29488 -4172 -29468 -3748
rect -30240 -4200 -29468 -4172
rect -29228 -3748 -28456 -3720
rect -29228 -4172 -28540 -3748
rect -28476 -4172 -28456 -3748
rect -29228 -4200 -28456 -4172
rect -28216 -3748 -27444 -3720
rect -28216 -4172 -27528 -3748
rect -27464 -4172 -27444 -3748
rect -28216 -4200 -27444 -4172
rect -27204 -3748 -26432 -3720
rect -27204 -4172 -26516 -3748
rect -26452 -4172 -26432 -3748
rect -27204 -4200 -26432 -4172
rect -26192 -3748 -25420 -3720
rect -26192 -4172 -25504 -3748
rect -25440 -4172 -25420 -3748
rect -26192 -4200 -25420 -4172
rect -25180 -3748 -24408 -3720
rect -25180 -4172 -24492 -3748
rect -24428 -4172 -24408 -3748
rect -25180 -4200 -24408 -4172
rect -24168 -3748 -23396 -3720
rect -24168 -4172 -23480 -3748
rect -23416 -4172 -23396 -3748
rect -24168 -4200 -23396 -4172
rect -23156 -3748 -22384 -3720
rect -23156 -4172 -22468 -3748
rect -22404 -4172 -22384 -3748
rect -23156 -4200 -22384 -4172
rect -22144 -3748 -21372 -3720
rect -22144 -4172 -21456 -3748
rect -21392 -4172 -21372 -3748
rect -22144 -4200 -21372 -4172
rect -21132 -3748 -20360 -3720
rect -21132 -4172 -20444 -3748
rect -20380 -4172 -20360 -3748
rect -21132 -4200 -20360 -4172
rect -20120 -3748 -19348 -3720
rect -20120 -4172 -19432 -3748
rect -19368 -4172 -19348 -3748
rect -20120 -4200 -19348 -4172
rect -19108 -3748 -18336 -3720
rect -19108 -4172 -18420 -3748
rect -18356 -4172 -18336 -3748
rect -19108 -4200 -18336 -4172
rect -18096 -3748 -17324 -3720
rect -18096 -4172 -17408 -3748
rect -17344 -4172 -17324 -3748
rect -18096 -4200 -17324 -4172
rect -17084 -3748 -16312 -3720
rect -17084 -4172 -16396 -3748
rect -16332 -4172 -16312 -3748
rect -17084 -4200 -16312 -4172
rect -16072 -3748 -15300 -3720
rect -16072 -4172 -15384 -3748
rect -15320 -4172 -15300 -3748
rect -16072 -4200 -15300 -4172
rect -15060 -3748 -14288 -3720
rect -15060 -4172 -14372 -3748
rect -14308 -4172 -14288 -3748
rect -15060 -4200 -14288 -4172
rect -14048 -3748 -13276 -3720
rect -14048 -4172 -13360 -3748
rect -13296 -4172 -13276 -3748
rect -14048 -4200 -13276 -4172
rect -13036 -3748 -12264 -3720
rect -13036 -4172 -12348 -3748
rect -12284 -4172 -12264 -3748
rect -13036 -4200 -12264 -4172
rect -12024 -3748 -11252 -3720
rect -12024 -4172 -11336 -3748
rect -11272 -4172 -11252 -3748
rect -12024 -4200 -11252 -4172
rect -11012 -3748 -10240 -3720
rect -11012 -4172 -10324 -3748
rect -10260 -4172 -10240 -3748
rect -11012 -4200 -10240 -4172
rect -10000 -3748 -9228 -3720
rect -10000 -4172 -9312 -3748
rect -9248 -4172 -9228 -3748
rect -10000 -4200 -9228 -4172
rect -8988 -3748 -8216 -3720
rect -8988 -4172 -8300 -3748
rect -8236 -4172 -8216 -3748
rect -8988 -4200 -8216 -4172
rect -7976 -3748 -7204 -3720
rect -7976 -4172 -7288 -3748
rect -7224 -4172 -7204 -3748
rect -7976 -4200 -7204 -4172
rect -6964 -3748 -6192 -3720
rect -6964 -4172 -6276 -3748
rect -6212 -4172 -6192 -3748
rect -6964 -4200 -6192 -4172
rect -5952 -3748 -5180 -3720
rect -5952 -4172 -5264 -3748
rect -5200 -4172 -5180 -3748
rect -5952 -4200 -5180 -4172
rect -4940 -3748 -4168 -3720
rect -4940 -4172 -4252 -3748
rect -4188 -4172 -4168 -3748
rect -4940 -4200 -4168 -4172
rect -3928 -3748 -3156 -3720
rect -3928 -4172 -3240 -3748
rect -3176 -4172 -3156 -3748
rect -3928 -4200 -3156 -4172
rect -2916 -3748 -2144 -3720
rect -2916 -4172 -2228 -3748
rect -2164 -4172 -2144 -3748
rect -2916 -4200 -2144 -4172
rect -1904 -3748 -1132 -3720
rect -1904 -4172 -1216 -3748
rect -1152 -4172 -1132 -3748
rect -1904 -4200 -1132 -4172
rect -892 -3748 -120 -3720
rect -892 -4172 -204 -3748
rect -140 -4172 -120 -3748
rect -892 -4200 -120 -4172
rect 120 -3748 892 -3720
rect 120 -4172 808 -3748
rect 872 -4172 892 -3748
rect 120 -4200 892 -4172
rect 1132 -3748 1904 -3720
rect 1132 -4172 1820 -3748
rect 1884 -4172 1904 -3748
rect 1132 -4200 1904 -4172
rect 2144 -3748 2916 -3720
rect 2144 -4172 2832 -3748
rect 2896 -4172 2916 -3748
rect 2144 -4200 2916 -4172
rect 3156 -3748 3928 -3720
rect 3156 -4172 3844 -3748
rect 3908 -4172 3928 -3748
rect 3156 -4200 3928 -4172
rect 4168 -3748 4940 -3720
rect 4168 -4172 4856 -3748
rect 4920 -4172 4940 -3748
rect 4168 -4200 4940 -4172
rect 5180 -3748 5952 -3720
rect 5180 -4172 5868 -3748
rect 5932 -4172 5952 -3748
rect 5180 -4200 5952 -4172
rect 6192 -3748 6964 -3720
rect 6192 -4172 6880 -3748
rect 6944 -4172 6964 -3748
rect 6192 -4200 6964 -4172
rect 7204 -3748 7976 -3720
rect 7204 -4172 7892 -3748
rect 7956 -4172 7976 -3748
rect 7204 -4200 7976 -4172
rect 8216 -3748 8988 -3720
rect 8216 -4172 8904 -3748
rect 8968 -4172 8988 -3748
rect 8216 -4200 8988 -4172
rect 9228 -3748 10000 -3720
rect 9228 -4172 9916 -3748
rect 9980 -4172 10000 -3748
rect 9228 -4200 10000 -4172
rect 10240 -3748 11012 -3720
rect 10240 -4172 10928 -3748
rect 10992 -4172 11012 -3748
rect 10240 -4200 11012 -4172
rect 11252 -3748 12024 -3720
rect 11252 -4172 11940 -3748
rect 12004 -4172 12024 -3748
rect 11252 -4200 12024 -4172
rect 12264 -3748 13036 -3720
rect 12264 -4172 12952 -3748
rect 13016 -4172 13036 -3748
rect 12264 -4200 13036 -4172
rect 13276 -3748 14048 -3720
rect 13276 -4172 13964 -3748
rect 14028 -4172 14048 -3748
rect 13276 -4200 14048 -4172
rect 14288 -3748 15060 -3720
rect 14288 -4172 14976 -3748
rect 15040 -4172 15060 -3748
rect 14288 -4200 15060 -4172
rect 15300 -3748 16072 -3720
rect 15300 -4172 15988 -3748
rect 16052 -4172 16072 -3748
rect 15300 -4200 16072 -4172
rect 16312 -3748 17084 -3720
rect 16312 -4172 17000 -3748
rect 17064 -4172 17084 -3748
rect 16312 -4200 17084 -4172
rect 17324 -3748 18096 -3720
rect 17324 -4172 18012 -3748
rect 18076 -4172 18096 -3748
rect 17324 -4200 18096 -4172
rect 18336 -3748 19108 -3720
rect 18336 -4172 19024 -3748
rect 19088 -4172 19108 -3748
rect 18336 -4200 19108 -4172
rect 19348 -3748 20120 -3720
rect 19348 -4172 20036 -3748
rect 20100 -4172 20120 -3748
rect 19348 -4200 20120 -4172
rect 20360 -3748 21132 -3720
rect 20360 -4172 21048 -3748
rect 21112 -4172 21132 -3748
rect 20360 -4200 21132 -4172
rect 21372 -3748 22144 -3720
rect 21372 -4172 22060 -3748
rect 22124 -4172 22144 -3748
rect 21372 -4200 22144 -4172
rect 22384 -3748 23156 -3720
rect 22384 -4172 23072 -3748
rect 23136 -4172 23156 -3748
rect 22384 -4200 23156 -4172
rect 23396 -3748 24168 -3720
rect 23396 -4172 24084 -3748
rect 24148 -4172 24168 -3748
rect 23396 -4200 24168 -4172
rect 24408 -3748 25180 -3720
rect 24408 -4172 25096 -3748
rect 25160 -4172 25180 -3748
rect 24408 -4200 25180 -4172
rect 25420 -3748 26192 -3720
rect 25420 -4172 26108 -3748
rect 26172 -4172 26192 -3748
rect 25420 -4200 26192 -4172
rect 26432 -3748 27204 -3720
rect 26432 -4172 27120 -3748
rect 27184 -4172 27204 -3748
rect 26432 -4200 27204 -4172
rect 27444 -3748 28216 -3720
rect 27444 -4172 28132 -3748
rect 28196 -4172 28216 -3748
rect 27444 -4200 28216 -4172
rect 28456 -3748 29228 -3720
rect 28456 -4172 29144 -3748
rect 29208 -4172 29228 -3748
rect 28456 -4200 29228 -4172
rect 29468 -3748 30240 -3720
rect 29468 -4172 30156 -3748
rect 30220 -4172 30240 -3748
rect 29468 -4200 30240 -4172
rect 30480 -3748 31252 -3720
rect 30480 -4172 31168 -3748
rect 31232 -4172 31252 -3748
rect 30480 -4200 31252 -4172
rect 31492 -3748 32264 -3720
rect 31492 -4172 32180 -3748
rect 32244 -4172 32264 -3748
rect 31492 -4200 32264 -4172
rect -32264 -4468 -31492 -4440
rect -32264 -4892 -31576 -4468
rect -31512 -4892 -31492 -4468
rect -32264 -4920 -31492 -4892
rect -31252 -4468 -30480 -4440
rect -31252 -4892 -30564 -4468
rect -30500 -4892 -30480 -4468
rect -31252 -4920 -30480 -4892
rect -30240 -4468 -29468 -4440
rect -30240 -4892 -29552 -4468
rect -29488 -4892 -29468 -4468
rect -30240 -4920 -29468 -4892
rect -29228 -4468 -28456 -4440
rect -29228 -4892 -28540 -4468
rect -28476 -4892 -28456 -4468
rect -29228 -4920 -28456 -4892
rect -28216 -4468 -27444 -4440
rect -28216 -4892 -27528 -4468
rect -27464 -4892 -27444 -4468
rect -28216 -4920 -27444 -4892
rect -27204 -4468 -26432 -4440
rect -27204 -4892 -26516 -4468
rect -26452 -4892 -26432 -4468
rect -27204 -4920 -26432 -4892
rect -26192 -4468 -25420 -4440
rect -26192 -4892 -25504 -4468
rect -25440 -4892 -25420 -4468
rect -26192 -4920 -25420 -4892
rect -25180 -4468 -24408 -4440
rect -25180 -4892 -24492 -4468
rect -24428 -4892 -24408 -4468
rect -25180 -4920 -24408 -4892
rect -24168 -4468 -23396 -4440
rect -24168 -4892 -23480 -4468
rect -23416 -4892 -23396 -4468
rect -24168 -4920 -23396 -4892
rect -23156 -4468 -22384 -4440
rect -23156 -4892 -22468 -4468
rect -22404 -4892 -22384 -4468
rect -23156 -4920 -22384 -4892
rect -22144 -4468 -21372 -4440
rect -22144 -4892 -21456 -4468
rect -21392 -4892 -21372 -4468
rect -22144 -4920 -21372 -4892
rect -21132 -4468 -20360 -4440
rect -21132 -4892 -20444 -4468
rect -20380 -4892 -20360 -4468
rect -21132 -4920 -20360 -4892
rect -20120 -4468 -19348 -4440
rect -20120 -4892 -19432 -4468
rect -19368 -4892 -19348 -4468
rect -20120 -4920 -19348 -4892
rect -19108 -4468 -18336 -4440
rect -19108 -4892 -18420 -4468
rect -18356 -4892 -18336 -4468
rect -19108 -4920 -18336 -4892
rect -18096 -4468 -17324 -4440
rect -18096 -4892 -17408 -4468
rect -17344 -4892 -17324 -4468
rect -18096 -4920 -17324 -4892
rect -17084 -4468 -16312 -4440
rect -17084 -4892 -16396 -4468
rect -16332 -4892 -16312 -4468
rect -17084 -4920 -16312 -4892
rect -16072 -4468 -15300 -4440
rect -16072 -4892 -15384 -4468
rect -15320 -4892 -15300 -4468
rect -16072 -4920 -15300 -4892
rect -15060 -4468 -14288 -4440
rect -15060 -4892 -14372 -4468
rect -14308 -4892 -14288 -4468
rect -15060 -4920 -14288 -4892
rect -14048 -4468 -13276 -4440
rect -14048 -4892 -13360 -4468
rect -13296 -4892 -13276 -4468
rect -14048 -4920 -13276 -4892
rect -13036 -4468 -12264 -4440
rect -13036 -4892 -12348 -4468
rect -12284 -4892 -12264 -4468
rect -13036 -4920 -12264 -4892
rect -12024 -4468 -11252 -4440
rect -12024 -4892 -11336 -4468
rect -11272 -4892 -11252 -4468
rect -12024 -4920 -11252 -4892
rect -11012 -4468 -10240 -4440
rect -11012 -4892 -10324 -4468
rect -10260 -4892 -10240 -4468
rect -11012 -4920 -10240 -4892
rect -10000 -4468 -9228 -4440
rect -10000 -4892 -9312 -4468
rect -9248 -4892 -9228 -4468
rect -10000 -4920 -9228 -4892
rect -8988 -4468 -8216 -4440
rect -8988 -4892 -8300 -4468
rect -8236 -4892 -8216 -4468
rect -8988 -4920 -8216 -4892
rect -7976 -4468 -7204 -4440
rect -7976 -4892 -7288 -4468
rect -7224 -4892 -7204 -4468
rect -7976 -4920 -7204 -4892
rect -6964 -4468 -6192 -4440
rect -6964 -4892 -6276 -4468
rect -6212 -4892 -6192 -4468
rect -6964 -4920 -6192 -4892
rect -5952 -4468 -5180 -4440
rect -5952 -4892 -5264 -4468
rect -5200 -4892 -5180 -4468
rect -5952 -4920 -5180 -4892
rect -4940 -4468 -4168 -4440
rect -4940 -4892 -4252 -4468
rect -4188 -4892 -4168 -4468
rect -4940 -4920 -4168 -4892
rect -3928 -4468 -3156 -4440
rect -3928 -4892 -3240 -4468
rect -3176 -4892 -3156 -4468
rect -3928 -4920 -3156 -4892
rect -2916 -4468 -2144 -4440
rect -2916 -4892 -2228 -4468
rect -2164 -4892 -2144 -4468
rect -2916 -4920 -2144 -4892
rect -1904 -4468 -1132 -4440
rect -1904 -4892 -1216 -4468
rect -1152 -4892 -1132 -4468
rect -1904 -4920 -1132 -4892
rect -892 -4468 -120 -4440
rect -892 -4892 -204 -4468
rect -140 -4892 -120 -4468
rect -892 -4920 -120 -4892
rect 120 -4468 892 -4440
rect 120 -4892 808 -4468
rect 872 -4892 892 -4468
rect 120 -4920 892 -4892
rect 1132 -4468 1904 -4440
rect 1132 -4892 1820 -4468
rect 1884 -4892 1904 -4468
rect 1132 -4920 1904 -4892
rect 2144 -4468 2916 -4440
rect 2144 -4892 2832 -4468
rect 2896 -4892 2916 -4468
rect 2144 -4920 2916 -4892
rect 3156 -4468 3928 -4440
rect 3156 -4892 3844 -4468
rect 3908 -4892 3928 -4468
rect 3156 -4920 3928 -4892
rect 4168 -4468 4940 -4440
rect 4168 -4892 4856 -4468
rect 4920 -4892 4940 -4468
rect 4168 -4920 4940 -4892
rect 5180 -4468 5952 -4440
rect 5180 -4892 5868 -4468
rect 5932 -4892 5952 -4468
rect 5180 -4920 5952 -4892
rect 6192 -4468 6964 -4440
rect 6192 -4892 6880 -4468
rect 6944 -4892 6964 -4468
rect 6192 -4920 6964 -4892
rect 7204 -4468 7976 -4440
rect 7204 -4892 7892 -4468
rect 7956 -4892 7976 -4468
rect 7204 -4920 7976 -4892
rect 8216 -4468 8988 -4440
rect 8216 -4892 8904 -4468
rect 8968 -4892 8988 -4468
rect 8216 -4920 8988 -4892
rect 9228 -4468 10000 -4440
rect 9228 -4892 9916 -4468
rect 9980 -4892 10000 -4468
rect 9228 -4920 10000 -4892
rect 10240 -4468 11012 -4440
rect 10240 -4892 10928 -4468
rect 10992 -4892 11012 -4468
rect 10240 -4920 11012 -4892
rect 11252 -4468 12024 -4440
rect 11252 -4892 11940 -4468
rect 12004 -4892 12024 -4468
rect 11252 -4920 12024 -4892
rect 12264 -4468 13036 -4440
rect 12264 -4892 12952 -4468
rect 13016 -4892 13036 -4468
rect 12264 -4920 13036 -4892
rect 13276 -4468 14048 -4440
rect 13276 -4892 13964 -4468
rect 14028 -4892 14048 -4468
rect 13276 -4920 14048 -4892
rect 14288 -4468 15060 -4440
rect 14288 -4892 14976 -4468
rect 15040 -4892 15060 -4468
rect 14288 -4920 15060 -4892
rect 15300 -4468 16072 -4440
rect 15300 -4892 15988 -4468
rect 16052 -4892 16072 -4468
rect 15300 -4920 16072 -4892
rect 16312 -4468 17084 -4440
rect 16312 -4892 17000 -4468
rect 17064 -4892 17084 -4468
rect 16312 -4920 17084 -4892
rect 17324 -4468 18096 -4440
rect 17324 -4892 18012 -4468
rect 18076 -4892 18096 -4468
rect 17324 -4920 18096 -4892
rect 18336 -4468 19108 -4440
rect 18336 -4892 19024 -4468
rect 19088 -4892 19108 -4468
rect 18336 -4920 19108 -4892
rect 19348 -4468 20120 -4440
rect 19348 -4892 20036 -4468
rect 20100 -4892 20120 -4468
rect 19348 -4920 20120 -4892
rect 20360 -4468 21132 -4440
rect 20360 -4892 21048 -4468
rect 21112 -4892 21132 -4468
rect 20360 -4920 21132 -4892
rect 21372 -4468 22144 -4440
rect 21372 -4892 22060 -4468
rect 22124 -4892 22144 -4468
rect 21372 -4920 22144 -4892
rect 22384 -4468 23156 -4440
rect 22384 -4892 23072 -4468
rect 23136 -4892 23156 -4468
rect 22384 -4920 23156 -4892
rect 23396 -4468 24168 -4440
rect 23396 -4892 24084 -4468
rect 24148 -4892 24168 -4468
rect 23396 -4920 24168 -4892
rect 24408 -4468 25180 -4440
rect 24408 -4892 25096 -4468
rect 25160 -4892 25180 -4468
rect 24408 -4920 25180 -4892
rect 25420 -4468 26192 -4440
rect 25420 -4892 26108 -4468
rect 26172 -4892 26192 -4468
rect 25420 -4920 26192 -4892
rect 26432 -4468 27204 -4440
rect 26432 -4892 27120 -4468
rect 27184 -4892 27204 -4468
rect 26432 -4920 27204 -4892
rect 27444 -4468 28216 -4440
rect 27444 -4892 28132 -4468
rect 28196 -4892 28216 -4468
rect 27444 -4920 28216 -4892
rect 28456 -4468 29228 -4440
rect 28456 -4892 29144 -4468
rect 29208 -4892 29228 -4468
rect 28456 -4920 29228 -4892
rect 29468 -4468 30240 -4440
rect 29468 -4892 30156 -4468
rect 30220 -4892 30240 -4468
rect 29468 -4920 30240 -4892
rect 30480 -4468 31252 -4440
rect 30480 -4892 31168 -4468
rect 31232 -4892 31252 -4468
rect 30480 -4920 31252 -4892
rect 31492 -4468 32264 -4440
rect 31492 -4892 32180 -4468
rect 32244 -4892 32264 -4468
rect 31492 -4920 32264 -4892
rect -32264 -5188 -31492 -5160
rect -32264 -5612 -31576 -5188
rect -31512 -5612 -31492 -5188
rect -32264 -5640 -31492 -5612
rect -31252 -5188 -30480 -5160
rect -31252 -5612 -30564 -5188
rect -30500 -5612 -30480 -5188
rect -31252 -5640 -30480 -5612
rect -30240 -5188 -29468 -5160
rect -30240 -5612 -29552 -5188
rect -29488 -5612 -29468 -5188
rect -30240 -5640 -29468 -5612
rect -29228 -5188 -28456 -5160
rect -29228 -5612 -28540 -5188
rect -28476 -5612 -28456 -5188
rect -29228 -5640 -28456 -5612
rect -28216 -5188 -27444 -5160
rect -28216 -5612 -27528 -5188
rect -27464 -5612 -27444 -5188
rect -28216 -5640 -27444 -5612
rect -27204 -5188 -26432 -5160
rect -27204 -5612 -26516 -5188
rect -26452 -5612 -26432 -5188
rect -27204 -5640 -26432 -5612
rect -26192 -5188 -25420 -5160
rect -26192 -5612 -25504 -5188
rect -25440 -5612 -25420 -5188
rect -26192 -5640 -25420 -5612
rect -25180 -5188 -24408 -5160
rect -25180 -5612 -24492 -5188
rect -24428 -5612 -24408 -5188
rect -25180 -5640 -24408 -5612
rect -24168 -5188 -23396 -5160
rect -24168 -5612 -23480 -5188
rect -23416 -5612 -23396 -5188
rect -24168 -5640 -23396 -5612
rect -23156 -5188 -22384 -5160
rect -23156 -5612 -22468 -5188
rect -22404 -5612 -22384 -5188
rect -23156 -5640 -22384 -5612
rect -22144 -5188 -21372 -5160
rect -22144 -5612 -21456 -5188
rect -21392 -5612 -21372 -5188
rect -22144 -5640 -21372 -5612
rect -21132 -5188 -20360 -5160
rect -21132 -5612 -20444 -5188
rect -20380 -5612 -20360 -5188
rect -21132 -5640 -20360 -5612
rect -20120 -5188 -19348 -5160
rect -20120 -5612 -19432 -5188
rect -19368 -5612 -19348 -5188
rect -20120 -5640 -19348 -5612
rect -19108 -5188 -18336 -5160
rect -19108 -5612 -18420 -5188
rect -18356 -5612 -18336 -5188
rect -19108 -5640 -18336 -5612
rect -18096 -5188 -17324 -5160
rect -18096 -5612 -17408 -5188
rect -17344 -5612 -17324 -5188
rect -18096 -5640 -17324 -5612
rect -17084 -5188 -16312 -5160
rect -17084 -5612 -16396 -5188
rect -16332 -5612 -16312 -5188
rect -17084 -5640 -16312 -5612
rect -16072 -5188 -15300 -5160
rect -16072 -5612 -15384 -5188
rect -15320 -5612 -15300 -5188
rect -16072 -5640 -15300 -5612
rect -15060 -5188 -14288 -5160
rect -15060 -5612 -14372 -5188
rect -14308 -5612 -14288 -5188
rect -15060 -5640 -14288 -5612
rect -14048 -5188 -13276 -5160
rect -14048 -5612 -13360 -5188
rect -13296 -5612 -13276 -5188
rect -14048 -5640 -13276 -5612
rect -13036 -5188 -12264 -5160
rect -13036 -5612 -12348 -5188
rect -12284 -5612 -12264 -5188
rect -13036 -5640 -12264 -5612
rect -12024 -5188 -11252 -5160
rect -12024 -5612 -11336 -5188
rect -11272 -5612 -11252 -5188
rect -12024 -5640 -11252 -5612
rect -11012 -5188 -10240 -5160
rect -11012 -5612 -10324 -5188
rect -10260 -5612 -10240 -5188
rect -11012 -5640 -10240 -5612
rect -10000 -5188 -9228 -5160
rect -10000 -5612 -9312 -5188
rect -9248 -5612 -9228 -5188
rect -10000 -5640 -9228 -5612
rect -8988 -5188 -8216 -5160
rect -8988 -5612 -8300 -5188
rect -8236 -5612 -8216 -5188
rect -8988 -5640 -8216 -5612
rect -7976 -5188 -7204 -5160
rect -7976 -5612 -7288 -5188
rect -7224 -5612 -7204 -5188
rect -7976 -5640 -7204 -5612
rect -6964 -5188 -6192 -5160
rect -6964 -5612 -6276 -5188
rect -6212 -5612 -6192 -5188
rect -6964 -5640 -6192 -5612
rect -5952 -5188 -5180 -5160
rect -5952 -5612 -5264 -5188
rect -5200 -5612 -5180 -5188
rect -5952 -5640 -5180 -5612
rect -4940 -5188 -4168 -5160
rect -4940 -5612 -4252 -5188
rect -4188 -5612 -4168 -5188
rect -4940 -5640 -4168 -5612
rect -3928 -5188 -3156 -5160
rect -3928 -5612 -3240 -5188
rect -3176 -5612 -3156 -5188
rect -3928 -5640 -3156 -5612
rect -2916 -5188 -2144 -5160
rect -2916 -5612 -2228 -5188
rect -2164 -5612 -2144 -5188
rect -2916 -5640 -2144 -5612
rect -1904 -5188 -1132 -5160
rect -1904 -5612 -1216 -5188
rect -1152 -5612 -1132 -5188
rect -1904 -5640 -1132 -5612
rect -892 -5188 -120 -5160
rect -892 -5612 -204 -5188
rect -140 -5612 -120 -5188
rect -892 -5640 -120 -5612
rect 120 -5188 892 -5160
rect 120 -5612 808 -5188
rect 872 -5612 892 -5188
rect 120 -5640 892 -5612
rect 1132 -5188 1904 -5160
rect 1132 -5612 1820 -5188
rect 1884 -5612 1904 -5188
rect 1132 -5640 1904 -5612
rect 2144 -5188 2916 -5160
rect 2144 -5612 2832 -5188
rect 2896 -5612 2916 -5188
rect 2144 -5640 2916 -5612
rect 3156 -5188 3928 -5160
rect 3156 -5612 3844 -5188
rect 3908 -5612 3928 -5188
rect 3156 -5640 3928 -5612
rect 4168 -5188 4940 -5160
rect 4168 -5612 4856 -5188
rect 4920 -5612 4940 -5188
rect 4168 -5640 4940 -5612
rect 5180 -5188 5952 -5160
rect 5180 -5612 5868 -5188
rect 5932 -5612 5952 -5188
rect 5180 -5640 5952 -5612
rect 6192 -5188 6964 -5160
rect 6192 -5612 6880 -5188
rect 6944 -5612 6964 -5188
rect 6192 -5640 6964 -5612
rect 7204 -5188 7976 -5160
rect 7204 -5612 7892 -5188
rect 7956 -5612 7976 -5188
rect 7204 -5640 7976 -5612
rect 8216 -5188 8988 -5160
rect 8216 -5612 8904 -5188
rect 8968 -5612 8988 -5188
rect 8216 -5640 8988 -5612
rect 9228 -5188 10000 -5160
rect 9228 -5612 9916 -5188
rect 9980 -5612 10000 -5188
rect 9228 -5640 10000 -5612
rect 10240 -5188 11012 -5160
rect 10240 -5612 10928 -5188
rect 10992 -5612 11012 -5188
rect 10240 -5640 11012 -5612
rect 11252 -5188 12024 -5160
rect 11252 -5612 11940 -5188
rect 12004 -5612 12024 -5188
rect 11252 -5640 12024 -5612
rect 12264 -5188 13036 -5160
rect 12264 -5612 12952 -5188
rect 13016 -5612 13036 -5188
rect 12264 -5640 13036 -5612
rect 13276 -5188 14048 -5160
rect 13276 -5612 13964 -5188
rect 14028 -5612 14048 -5188
rect 13276 -5640 14048 -5612
rect 14288 -5188 15060 -5160
rect 14288 -5612 14976 -5188
rect 15040 -5612 15060 -5188
rect 14288 -5640 15060 -5612
rect 15300 -5188 16072 -5160
rect 15300 -5612 15988 -5188
rect 16052 -5612 16072 -5188
rect 15300 -5640 16072 -5612
rect 16312 -5188 17084 -5160
rect 16312 -5612 17000 -5188
rect 17064 -5612 17084 -5188
rect 16312 -5640 17084 -5612
rect 17324 -5188 18096 -5160
rect 17324 -5612 18012 -5188
rect 18076 -5612 18096 -5188
rect 17324 -5640 18096 -5612
rect 18336 -5188 19108 -5160
rect 18336 -5612 19024 -5188
rect 19088 -5612 19108 -5188
rect 18336 -5640 19108 -5612
rect 19348 -5188 20120 -5160
rect 19348 -5612 20036 -5188
rect 20100 -5612 20120 -5188
rect 19348 -5640 20120 -5612
rect 20360 -5188 21132 -5160
rect 20360 -5612 21048 -5188
rect 21112 -5612 21132 -5188
rect 20360 -5640 21132 -5612
rect 21372 -5188 22144 -5160
rect 21372 -5612 22060 -5188
rect 22124 -5612 22144 -5188
rect 21372 -5640 22144 -5612
rect 22384 -5188 23156 -5160
rect 22384 -5612 23072 -5188
rect 23136 -5612 23156 -5188
rect 22384 -5640 23156 -5612
rect 23396 -5188 24168 -5160
rect 23396 -5612 24084 -5188
rect 24148 -5612 24168 -5188
rect 23396 -5640 24168 -5612
rect 24408 -5188 25180 -5160
rect 24408 -5612 25096 -5188
rect 25160 -5612 25180 -5188
rect 24408 -5640 25180 -5612
rect 25420 -5188 26192 -5160
rect 25420 -5612 26108 -5188
rect 26172 -5612 26192 -5188
rect 25420 -5640 26192 -5612
rect 26432 -5188 27204 -5160
rect 26432 -5612 27120 -5188
rect 27184 -5612 27204 -5188
rect 26432 -5640 27204 -5612
rect 27444 -5188 28216 -5160
rect 27444 -5612 28132 -5188
rect 28196 -5612 28216 -5188
rect 27444 -5640 28216 -5612
rect 28456 -5188 29228 -5160
rect 28456 -5612 29144 -5188
rect 29208 -5612 29228 -5188
rect 28456 -5640 29228 -5612
rect 29468 -5188 30240 -5160
rect 29468 -5612 30156 -5188
rect 30220 -5612 30240 -5188
rect 29468 -5640 30240 -5612
rect 30480 -5188 31252 -5160
rect 30480 -5612 31168 -5188
rect 31232 -5612 31252 -5188
rect 30480 -5640 31252 -5612
rect 31492 -5188 32264 -5160
rect 31492 -5612 32180 -5188
rect 32244 -5612 32264 -5188
rect 31492 -5640 32264 -5612
<< via3 >>
rect -31576 5188 -31512 5612
rect -30564 5188 -30500 5612
rect -29552 5188 -29488 5612
rect -28540 5188 -28476 5612
rect -27528 5188 -27464 5612
rect -26516 5188 -26452 5612
rect -25504 5188 -25440 5612
rect -24492 5188 -24428 5612
rect -23480 5188 -23416 5612
rect -22468 5188 -22404 5612
rect -21456 5188 -21392 5612
rect -20444 5188 -20380 5612
rect -19432 5188 -19368 5612
rect -18420 5188 -18356 5612
rect -17408 5188 -17344 5612
rect -16396 5188 -16332 5612
rect -15384 5188 -15320 5612
rect -14372 5188 -14308 5612
rect -13360 5188 -13296 5612
rect -12348 5188 -12284 5612
rect -11336 5188 -11272 5612
rect -10324 5188 -10260 5612
rect -9312 5188 -9248 5612
rect -8300 5188 -8236 5612
rect -7288 5188 -7224 5612
rect -6276 5188 -6212 5612
rect -5264 5188 -5200 5612
rect -4252 5188 -4188 5612
rect -3240 5188 -3176 5612
rect -2228 5188 -2164 5612
rect -1216 5188 -1152 5612
rect -204 5188 -140 5612
rect 808 5188 872 5612
rect 1820 5188 1884 5612
rect 2832 5188 2896 5612
rect 3844 5188 3908 5612
rect 4856 5188 4920 5612
rect 5868 5188 5932 5612
rect 6880 5188 6944 5612
rect 7892 5188 7956 5612
rect 8904 5188 8968 5612
rect 9916 5188 9980 5612
rect 10928 5188 10992 5612
rect 11940 5188 12004 5612
rect 12952 5188 13016 5612
rect 13964 5188 14028 5612
rect 14976 5188 15040 5612
rect 15988 5188 16052 5612
rect 17000 5188 17064 5612
rect 18012 5188 18076 5612
rect 19024 5188 19088 5612
rect 20036 5188 20100 5612
rect 21048 5188 21112 5612
rect 22060 5188 22124 5612
rect 23072 5188 23136 5612
rect 24084 5188 24148 5612
rect 25096 5188 25160 5612
rect 26108 5188 26172 5612
rect 27120 5188 27184 5612
rect 28132 5188 28196 5612
rect 29144 5188 29208 5612
rect 30156 5188 30220 5612
rect 31168 5188 31232 5612
rect 32180 5188 32244 5612
rect -31576 4468 -31512 4892
rect -30564 4468 -30500 4892
rect -29552 4468 -29488 4892
rect -28540 4468 -28476 4892
rect -27528 4468 -27464 4892
rect -26516 4468 -26452 4892
rect -25504 4468 -25440 4892
rect -24492 4468 -24428 4892
rect -23480 4468 -23416 4892
rect -22468 4468 -22404 4892
rect -21456 4468 -21392 4892
rect -20444 4468 -20380 4892
rect -19432 4468 -19368 4892
rect -18420 4468 -18356 4892
rect -17408 4468 -17344 4892
rect -16396 4468 -16332 4892
rect -15384 4468 -15320 4892
rect -14372 4468 -14308 4892
rect -13360 4468 -13296 4892
rect -12348 4468 -12284 4892
rect -11336 4468 -11272 4892
rect -10324 4468 -10260 4892
rect -9312 4468 -9248 4892
rect -8300 4468 -8236 4892
rect -7288 4468 -7224 4892
rect -6276 4468 -6212 4892
rect -5264 4468 -5200 4892
rect -4252 4468 -4188 4892
rect -3240 4468 -3176 4892
rect -2228 4468 -2164 4892
rect -1216 4468 -1152 4892
rect -204 4468 -140 4892
rect 808 4468 872 4892
rect 1820 4468 1884 4892
rect 2832 4468 2896 4892
rect 3844 4468 3908 4892
rect 4856 4468 4920 4892
rect 5868 4468 5932 4892
rect 6880 4468 6944 4892
rect 7892 4468 7956 4892
rect 8904 4468 8968 4892
rect 9916 4468 9980 4892
rect 10928 4468 10992 4892
rect 11940 4468 12004 4892
rect 12952 4468 13016 4892
rect 13964 4468 14028 4892
rect 14976 4468 15040 4892
rect 15988 4468 16052 4892
rect 17000 4468 17064 4892
rect 18012 4468 18076 4892
rect 19024 4468 19088 4892
rect 20036 4468 20100 4892
rect 21048 4468 21112 4892
rect 22060 4468 22124 4892
rect 23072 4468 23136 4892
rect 24084 4468 24148 4892
rect 25096 4468 25160 4892
rect 26108 4468 26172 4892
rect 27120 4468 27184 4892
rect 28132 4468 28196 4892
rect 29144 4468 29208 4892
rect 30156 4468 30220 4892
rect 31168 4468 31232 4892
rect 32180 4468 32244 4892
rect -31576 3748 -31512 4172
rect -30564 3748 -30500 4172
rect -29552 3748 -29488 4172
rect -28540 3748 -28476 4172
rect -27528 3748 -27464 4172
rect -26516 3748 -26452 4172
rect -25504 3748 -25440 4172
rect -24492 3748 -24428 4172
rect -23480 3748 -23416 4172
rect -22468 3748 -22404 4172
rect -21456 3748 -21392 4172
rect -20444 3748 -20380 4172
rect -19432 3748 -19368 4172
rect -18420 3748 -18356 4172
rect -17408 3748 -17344 4172
rect -16396 3748 -16332 4172
rect -15384 3748 -15320 4172
rect -14372 3748 -14308 4172
rect -13360 3748 -13296 4172
rect -12348 3748 -12284 4172
rect -11336 3748 -11272 4172
rect -10324 3748 -10260 4172
rect -9312 3748 -9248 4172
rect -8300 3748 -8236 4172
rect -7288 3748 -7224 4172
rect -6276 3748 -6212 4172
rect -5264 3748 -5200 4172
rect -4252 3748 -4188 4172
rect -3240 3748 -3176 4172
rect -2228 3748 -2164 4172
rect -1216 3748 -1152 4172
rect -204 3748 -140 4172
rect 808 3748 872 4172
rect 1820 3748 1884 4172
rect 2832 3748 2896 4172
rect 3844 3748 3908 4172
rect 4856 3748 4920 4172
rect 5868 3748 5932 4172
rect 6880 3748 6944 4172
rect 7892 3748 7956 4172
rect 8904 3748 8968 4172
rect 9916 3748 9980 4172
rect 10928 3748 10992 4172
rect 11940 3748 12004 4172
rect 12952 3748 13016 4172
rect 13964 3748 14028 4172
rect 14976 3748 15040 4172
rect 15988 3748 16052 4172
rect 17000 3748 17064 4172
rect 18012 3748 18076 4172
rect 19024 3748 19088 4172
rect 20036 3748 20100 4172
rect 21048 3748 21112 4172
rect 22060 3748 22124 4172
rect 23072 3748 23136 4172
rect 24084 3748 24148 4172
rect 25096 3748 25160 4172
rect 26108 3748 26172 4172
rect 27120 3748 27184 4172
rect 28132 3748 28196 4172
rect 29144 3748 29208 4172
rect 30156 3748 30220 4172
rect 31168 3748 31232 4172
rect 32180 3748 32244 4172
rect -31576 3028 -31512 3452
rect -30564 3028 -30500 3452
rect -29552 3028 -29488 3452
rect -28540 3028 -28476 3452
rect -27528 3028 -27464 3452
rect -26516 3028 -26452 3452
rect -25504 3028 -25440 3452
rect -24492 3028 -24428 3452
rect -23480 3028 -23416 3452
rect -22468 3028 -22404 3452
rect -21456 3028 -21392 3452
rect -20444 3028 -20380 3452
rect -19432 3028 -19368 3452
rect -18420 3028 -18356 3452
rect -17408 3028 -17344 3452
rect -16396 3028 -16332 3452
rect -15384 3028 -15320 3452
rect -14372 3028 -14308 3452
rect -13360 3028 -13296 3452
rect -12348 3028 -12284 3452
rect -11336 3028 -11272 3452
rect -10324 3028 -10260 3452
rect -9312 3028 -9248 3452
rect -8300 3028 -8236 3452
rect -7288 3028 -7224 3452
rect -6276 3028 -6212 3452
rect -5264 3028 -5200 3452
rect -4252 3028 -4188 3452
rect -3240 3028 -3176 3452
rect -2228 3028 -2164 3452
rect -1216 3028 -1152 3452
rect -204 3028 -140 3452
rect 808 3028 872 3452
rect 1820 3028 1884 3452
rect 2832 3028 2896 3452
rect 3844 3028 3908 3452
rect 4856 3028 4920 3452
rect 5868 3028 5932 3452
rect 6880 3028 6944 3452
rect 7892 3028 7956 3452
rect 8904 3028 8968 3452
rect 9916 3028 9980 3452
rect 10928 3028 10992 3452
rect 11940 3028 12004 3452
rect 12952 3028 13016 3452
rect 13964 3028 14028 3452
rect 14976 3028 15040 3452
rect 15988 3028 16052 3452
rect 17000 3028 17064 3452
rect 18012 3028 18076 3452
rect 19024 3028 19088 3452
rect 20036 3028 20100 3452
rect 21048 3028 21112 3452
rect 22060 3028 22124 3452
rect 23072 3028 23136 3452
rect 24084 3028 24148 3452
rect 25096 3028 25160 3452
rect 26108 3028 26172 3452
rect 27120 3028 27184 3452
rect 28132 3028 28196 3452
rect 29144 3028 29208 3452
rect 30156 3028 30220 3452
rect 31168 3028 31232 3452
rect 32180 3028 32244 3452
rect -31576 2308 -31512 2732
rect -30564 2308 -30500 2732
rect -29552 2308 -29488 2732
rect -28540 2308 -28476 2732
rect -27528 2308 -27464 2732
rect -26516 2308 -26452 2732
rect -25504 2308 -25440 2732
rect -24492 2308 -24428 2732
rect -23480 2308 -23416 2732
rect -22468 2308 -22404 2732
rect -21456 2308 -21392 2732
rect -20444 2308 -20380 2732
rect -19432 2308 -19368 2732
rect -18420 2308 -18356 2732
rect -17408 2308 -17344 2732
rect -16396 2308 -16332 2732
rect -15384 2308 -15320 2732
rect -14372 2308 -14308 2732
rect -13360 2308 -13296 2732
rect -12348 2308 -12284 2732
rect -11336 2308 -11272 2732
rect -10324 2308 -10260 2732
rect -9312 2308 -9248 2732
rect -8300 2308 -8236 2732
rect -7288 2308 -7224 2732
rect -6276 2308 -6212 2732
rect -5264 2308 -5200 2732
rect -4252 2308 -4188 2732
rect -3240 2308 -3176 2732
rect -2228 2308 -2164 2732
rect -1216 2308 -1152 2732
rect -204 2308 -140 2732
rect 808 2308 872 2732
rect 1820 2308 1884 2732
rect 2832 2308 2896 2732
rect 3844 2308 3908 2732
rect 4856 2308 4920 2732
rect 5868 2308 5932 2732
rect 6880 2308 6944 2732
rect 7892 2308 7956 2732
rect 8904 2308 8968 2732
rect 9916 2308 9980 2732
rect 10928 2308 10992 2732
rect 11940 2308 12004 2732
rect 12952 2308 13016 2732
rect 13964 2308 14028 2732
rect 14976 2308 15040 2732
rect 15988 2308 16052 2732
rect 17000 2308 17064 2732
rect 18012 2308 18076 2732
rect 19024 2308 19088 2732
rect 20036 2308 20100 2732
rect 21048 2308 21112 2732
rect 22060 2308 22124 2732
rect 23072 2308 23136 2732
rect 24084 2308 24148 2732
rect 25096 2308 25160 2732
rect 26108 2308 26172 2732
rect 27120 2308 27184 2732
rect 28132 2308 28196 2732
rect 29144 2308 29208 2732
rect 30156 2308 30220 2732
rect 31168 2308 31232 2732
rect 32180 2308 32244 2732
rect -31576 1588 -31512 2012
rect -30564 1588 -30500 2012
rect -29552 1588 -29488 2012
rect -28540 1588 -28476 2012
rect -27528 1588 -27464 2012
rect -26516 1588 -26452 2012
rect -25504 1588 -25440 2012
rect -24492 1588 -24428 2012
rect -23480 1588 -23416 2012
rect -22468 1588 -22404 2012
rect -21456 1588 -21392 2012
rect -20444 1588 -20380 2012
rect -19432 1588 -19368 2012
rect -18420 1588 -18356 2012
rect -17408 1588 -17344 2012
rect -16396 1588 -16332 2012
rect -15384 1588 -15320 2012
rect -14372 1588 -14308 2012
rect -13360 1588 -13296 2012
rect -12348 1588 -12284 2012
rect -11336 1588 -11272 2012
rect -10324 1588 -10260 2012
rect -9312 1588 -9248 2012
rect -8300 1588 -8236 2012
rect -7288 1588 -7224 2012
rect -6276 1588 -6212 2012
rect -5264 1588 -5200 2012
rect -4252 1588 -4188 2012
rect -3240 1588 -3176 2012
rect -2228 1588 -2164 2012
rect -1216 1588 -1152 2012
rect -204 1588 -140 2012
rect 808 1588 872 2012
rect 1820 1588 1884 2012
rect 2832 1588 2896 2012
rect 3844 1588 3908 2012
rect 4856 1588 4920 2012
rect 5868 1588 5932 2012
rect 6880 1588 6944 2012
rect 7892 1588 7956 2012
rect 8904 1588 8968 2012
rect 9916 1588 9980 2012
rect 10928 1588 10992 2012
rect 11940 1588 12004 2012
rect 12952 1588 13016 2012
rect 13964 1588 14028 2012
rect 14976 1588 15040 2012
rect 15988 1588 16052 2012
rect 17000 1588 17064 2012
rect 18012 1588 18076 2012
rect 19024 1588 19088 2012
rect 20036 1588 20100 2012
rect 21048 1588 21112 2012
rect 22060 1588 22124 2012
rect 23072 1588 23136 2012
rect 24084 1588 24148 2012
rect 25096 1588 25160 2012
rect 26108 1588 26172 2012
rect 27120 1588 27184 2012
rect 28132 1588 28196 2012
rect 29144 1588 29208 2012
rect 30156 1588 30220 2012
rect 31168 1588 31232 2012
rect 32180 1588 32244 2012
rect -31576 868 -31512 1292
rect -30564 868 -30500 1292
rect -29552 868 -29488 1292
rect -28540 868 -28476 1292
rect -27528 868 -27464 1292
rect -26516 868 -26452 1292
rect -25504 868 -25440 1292
rect -24492 868 -24428 1292
rect -23480 868 -23416 1292
rect -22468 868 -22404 1292
rect -21456 868 -21392 1292
rect -20444 868 -20380 1292
rect -19432 868 -19368 1292
rect -18420 868 -18356 1292
rect -17408 868 -17344 1292
rect -16396 868 -16332 1292
rect -15384 868 -15320 1292
rect -14372 868 -14308 1292
rect -13360 868 -13296 1292
rect -12348 868 -12284 1292
rect -11336 868 -11272 1292
rect -10324 868 -10260 1292
rect -9312 868 -9248 1292
rect -8300 868 -8236 1292
rect -7288 868 -7224 1292
rect -6276 868 -6212 1292
rect -5264 868 -5200 1292
rect -4252 868 -4188 1292
rect -3240 868 -3176 1292
rect -2228 868 -2164 1292
rect -1216 868 -1152 1292
rect -204 868 -140 1292
rect 808 868 872 1292
rect 1820 868 1884 1292
rect 2832 868 2896 1292
rect 3844 868 3908 1292
rect 4856 868 4920 1292
rect 5868 868 5932 1292
rect 6880 868 6944 1292
rect 7892 868 7956 1292
rect 8904 868 8968 1292
rect 9916 868 9980 1292
rect 10928 868 10992 1292
rect 11940 868 12004 1292
rect 12952 868 13016 1292
rect 13964 868 14028 1292
rect 14976 868 15040 1292
rect 15988 868 16052 1292
rect 17000 868 17064 1292
rect 18012 868 18076 1292
rect 19024 868 19088 1292
rect 20036 868 20100 1292
rect 21048 868 21112 1292
rect 22060 868 22124 1292
rect 23072 868 23136 1292
rect 24084 868 24148 1292
rect 25096 868 25160 1292
rect 26108 868 26172 1292
rect 27120 868 27184 1292
rect 28132 868 28196 1292
rect 29144 868 29208 1292
rect 30156 868 30220 1292
rect 31168 868 31232 1292
rect 32180 868 32244 1292
rect -31576 148 -31512 572
rect -30564 148 -30500 572
rect -29552 148 -29488 572
rect -28540 148 -28476 572
rect -27528 148 -27464 572
rect -26516 148 -26452 572
rect -25504 148 -25440 572
rect -24492 148 -24428 572
rect -23480 148 -23416 572
rect -22468 148 -22404 572
rect -21456 148 -21392 572
rect -20444 148 -20380 572
rect -19432 148 -19368 572
rect -18420 148 -18356 572
rect -17408 148 -17344 572
rect -16396 148 -16332 572
rect -15384 148 -15320 572
rect -14372 148 -14308 572
rect -13360 148 -13296 572
rect -12348 148 -12284 572
rect -11336 148 -11272 572
rect -10324 148 -10260 572
rect -9312 148 -9248 572
rect -8300 148 -8236 572
rect -7288 148 -7224 572
rect -6276 148 -6212 572
rect -5264 148 -5200 572
rect -4252 148 -4188 572
rect -3240 148 -3176 572
rect -2228 148 -2164 572
rect -1216 148 -1152 572
rect -204 148 -140 572
rect 808 148 872 572
rect 1820 148 1884 572
rect 2832 148 2896 572
rect 3844 148 3908 572
rect 4856 148 4920 572
rect 5868 148 5932 572
rect 6880 148 6944 572
rect 7892 148 7956 572
rect 8904 148 8968 572
rect 9916 148 9980 572
rect 10928 148 10992 572
rect 11940 148 12004 572
rect 12952 148 13016 572
rect 13964 148 14028 572
rect 14976 148 15040 572
rect 15988 148 16052 572
rect 17000 148 17064 572
rect 18012 148 18076 572
rect 19024 148 19088 572
rect 20036 148 20100 572
rect 21048 148 21112 572
rect 22060 148 22124 572
rect 23072 148 23136 572
rect 24084 148 24148 572
rect 25096 148 25160 572
rect 26108 148 26172 572
rect 27120 148 27184 572
rect 28132 148 28196 572
rect 29144 148 29208 572
rect 30156 148 30220 572
rect 31168 148 31232 572
rect 32180 148 32244 572
rect -31576 -572 -31512 -148
rect -30564 -572 -30500 -148
rect -29552 -572 -29488 -148
rect -28540 -572 -28476 -148
rect -27528 -572 -27464 -148
rect -26516 -572 -26452 -148
rect -25504 -572 -25440 -148
rect -24492 -572 -24428 -148
rect -23480 -572 -23416 -148
rect -22468 -572 -22404 -148
rect -21456 -572 -21392 -148
rect -20444 -572 -20380 -148
rect -19432 -572 -19368 -148
rect -18420 -572 -18356 -148
rect -17408 -572 -17344 -148
rect -16396 -572 -16332 -148
rect -15384 -572 -15320 -148
rect -14372 -572 -14308 -148
rect -13360 -572 -13296 -148
rect -12348 -572 -12284 -148
rect -11336 -572 -11272 -148
rect -10324 -572 -10260 -148
rect -9312 -572 -9248 -148
rect -8300 -572 -8236 -148
rect -7288 -572 -7224 -148
rect -6276 -572 -6212 -148
rect -5264 -572 -5200 -148
rect -4252 -572 -4188 -148
rect -3240 -572 -3176 -148
rect -2228 -572 -2164 -148
rect -1216 -572 -1152 -148
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect 1820 -572 1884 -148
rect 2832 -572 2896 -148
rect 3844 -572 3908 -148
rect 4856 -572 4920 -148
rect 5868 -572 5932 -148
rect 6880 -572 6944 -148
rect 7892 -572 7956 -148
rect 8904 -572 8968 -148
rect 9916 -572 9980 -148
rect 10928 -572 10992 -148
rect 11940 -572 12004 -148
rect 12952 -572 13016 -148
rect 13964 -572 14028 -148
rect 14976 -572 15040 -148
rect 15988 -572 16052 -148
rect 17000 -572 17064 -148
rect 18012 -572 18076 -148
rect 19024 -572 19088 -148
rect 20036 -572 20100 -148
rect 21048 -572 21112 -148
rect 22060 -572 22124 -148
rect 23072 -572 23136 -148
rect 24084 -572 24148 -148
rect 25096 -572 25160 -148
rect 26108 -572 26172 -148
rect 27120 -572 27184 -148
rect 28132 -572 28196 -148
rect 29144 -572 29208 -148
rect 30156 -572 30220 -148
rect 31168 -572 31232 -148
rect 32180 -572 32244 -148
rect -31576 -1292 -31512 -868
rect -30564 -1292 -30500 -868
rect -29552 -1292 -29488 -868
rect -28540 -1292 -28476 -868
rect -27528 -1292 -27464 -868
rect -26516 -1292 -26452 -868
rect -25504 -1292 -25440 -868
rect -24492 -1292 -24428 -868
rect -23480 -1292 -23416 -868
rect -22468 -1292 -22404 -868
rect -21456 -1292 -21392 -868
rect -20444 -1292 -20380 -868
rect -19432 -1292 -19368 -868
rect -18420 -1292 -18356 -868
rect -17408 -1292 -17344 -868
rect -16396 -1292 -16332 -868
rect -15384 -1292 -15320 -868
rect -14372 -1292 -14308 -868
rect -13360 -1292 -13296 -868
rect -12348 -1292 -12284 -868
rect -11336 -1292 -11272 -868
rect -10324 -1292 -10260 -868
rect -9312 -1292 -9248 -868
rect -8300 -1292 -8236 -868
rect -7288 -1292 -7224 -868
rect -6276 -1292 -6212 -868
rect -5264 -1292 -5200 -868
rect -4252 -1292 -4188 -868
rect -3240 -1292 -3176 -868
rect -2228 -1292 -2164 -868
rect -1216 -1292 -1152 -868
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect 1820 -1292 1884 -868
rect 2832 -1292 2896 -868
rect 3844 -1292 3908 -868
rect 4856 -1292 4920 -868
rect 5868 -1292 5932 -868
rect 6880 -1292 6944 -868
rect 7892 -1292 7956 -868
rect 8904 -1292 8968 -868
rect 9916 -1292 9980 -868
rect 10928 -1292 10992 -868
rect 11940 -1292 12004 -868
rect 12952 -1292 13016 -868
rect 13964 -1292 14028 -868
rect 14976 -1292 15040 -868
rect 15988 -1292 16052 -868
rect 17000 -1292 17064 -868
rect 18012 -1292 18076 -868
rect 19024 -1292 19088 -868
rect 20036 -1292 20100 -868
rect 21048 -1292 21112 -868
rect 22060 -1292 22124 -868
rect 23072 -1292 23136 -868
rect 24084 -1292 24148 -868
rect 25096 -1292 25160 -868
rect 26108 -1292 26172 -868
rect 27120 -1292 27184 -868
rect 28132 -1292 28196 -868
rect 29144 -1292 29208 -868
rect 30156 -1292 30220 -868
rect 31168 -1292 31232 -868
rect 32180 -1292 32244 -868
rect -31576 -2012 -31512 -1588
rect -30564 -2012 -30500 -1588
rect -29552 -2012 -29488 -1588
rect -28540 -2012 -28476 -1588
rect -27528 -2012 -27464 -1588
rect -26516 -2012 -26452 -1588
rect -25504 -2012 -25440 -1588
rect -24492 -2012 -24428 -1588
rect -23480 -2012 -23416 -1588
rect -22468 -2012 -22404 -1588
rect -21456 -2012 -21392 -1588
rect -20444 -2012 -20380 -1588
rect -19432 -2012 -19368 -1588
rect -18420 -2012 -18356 -1588
rect -17408 -2012 -17344 -1588
rect -16396 -2012 -16332 -1588
rect -15384 -2012 -15320 -1588
rect -14372 -2012 -14308 -1588
rect -13360 -2012 -13296 -1588
rect -12348 -2012 -12284 -1588
rect -11336 -2012 -11272 -1588
rect -10324 -2012 -10260 -1588
rect -9312 -2012 -9248 -1588
rect -8300 -2012 -8236 -1588
rect -7288 -2012 -7224 -1588
rect -6276 -2012 -6212 -1588
rect -5264 -2012 -5200 -1588
rect -4252 -2012 -4188 -1588
rect -3240 -2012 -3176 -1588
rect -2228 -2012 -2164 -1588
rect -1216 -2012 -1152 -1588
rect -204 -2012 -140 -1588
rect 808 -2012 872 -1588
rect 1820 -2012 1884 -1588
rect 2832 -2012 2896 -1588
rect 3844 -2012 3908 -1588
rect 4856 -2012 4920 -1588
rect 5868 -2012 5932 -1588
rect 6880 -2012 6944 -1588
rect 7892 -2012 7956 -1588
rect 8904 -2012 8968 -1588
rect 9916 -2012 9980 -1588
rect 10928 -2012 10992 -1588
rect 11940 -2012 12004 -1588
rect 12952 -2012 13016 -1588
rect 13964 -2012 14028 -1588
rect 14976 -2012 15040 -1588
rect 15988 -2012 16052 -1588
rect 17000 -2012 17064 -1588
rect 18012 -2012 18076 -1588
rect 19024 -2012 19088 -1588
rect 20036 -2012 20100 -1588
rect 21048 -2012 21112 -1588
rect 22060 -2012 22124 -1588
rect 23072 -2012 23136 -1588
rect 24084 -2012 24148 -1588
rect 25096 -2012 25160 -1588
rect 26108 -2012 26172 -1588
rect 27120 -2012 27184 -1588
rect 28132 -2012 28196 -1588
rect 29144 -2012 29208 -1588
rect 30156 -2012 30220 -1588
rect 31168 -2012 31232 -1588
rect 32180 -2012 32244 -1588
rect -31576 -2732 -31512 -2308
rect -30564 -2732 -30500 -2308
rect -29552 -2732 -29488 -2308
rect -28540 -2732 -28476 -2308
rect -27528 -2732 -27464 -2308
rect -26516 -2732 -26452 -2308
rect -25504 -2732 -25440 -2308
rect -24492 -2732 -24428 -2308
rect -23480 -2732 -23416 -2308
rect -22468 -2732 -22404 -2308
rect -21456 -2732 -21392 -2308
rect -20444 -2732 -20380 -2308
rect -19432 -2732 -19368 -2308
rect -18420 -2732 -18356 -2308
rect -17408 -2732 -17344 -2308
rect -16396 -2732 -16332 -2308
rect -15384 -2732 -15320 -2308
rect -14372 -2732 -14308 -2308
rect -13360 -2732 -13296 -2308
rect -12348 -2732 -12284 -2308
rect -11336 -2732 -11272 -2308
rect -10324 -2732 -10260 -2308
rect -9312 -2732 -9248 -2308
rect -8300 -2732 -8236 -2308
rect -7288 -2732 -7224 -2308
rect -6276 -2732 -6212 -2308
rect -5264 -2732 -5200 -2308
rect -4252 -2732 -4188 -2308
rect -3240 -2732 -3176 -2308
rect -2228 -2732 -2164 -2308
rect -1216 -2732 -1152 -2308
rect -204 -2732 -140 -2308
rect 808 -2732 872 -2308
rect 1820 -2732 1884 -2308
rect 2832 -2732 2896 -2308
rect 3844 -2732 3908 -2308
rect 4856 -2732 4920 -2308
rect 5868 -2732 5932 -2308
rect 6880 -2732 6944 -2308
rect 7892 -2732 7956 -2308
rect 8904 -2732 8968 -2308
rect 9916 -2732 9980 -2308
rect 10928 -2732 10992 -2308
rect 11940 -2732 12004 -2308
rect 12952 -2732 13016 -2308
rect 13964 -2732 14028 -2308
rect 14976 -2732 15040 -2308
rect 15988 -2732 16052 -2308
rect 17000 -2732 17064 -2308
rect 18012 -2732 18076 -2308
rect 19024 -2732 19088 -2308
rect 20036 -2732 20100 -2308
rect 21048 -2732 21112 -2308
rect 22060 -2732 22124 -2308
rect 23072 -2732 23136 -2308
rect 24084 -2732 24148 -2308
rect 25096 -2732 25160 -2308
rect 26108 -2732 26172 -2308
rect 27120 -2732 27184 -2308
rect 28132 -2732 28196 -2308
rect 29144 -2732 29208 -2308
rect 30156 -2732 30220 -2308
rect 31168 -2732 31232 -2308
rect 32180 -2732 32244 -2308
rect -31576 -3452 -31512 -3028
rect -30564 -3452 -30500 -3028
rect -29552 -3452 -29488 -3028
rect -28540 -3452 -28476 -3028
rect -27528 -3452 -27464 -3028
rect -26516 -3452 -26452 -3028
rect -25504 -3452 -25440 -3028
rect -24492 -3452 -24428 -3028
rect -23480 -3452 -23416 -3028
rect -22468 -3452 -22404 -3028
rect -21456 -3452 -21392 -3028
rect -20444 -3452 -20380 -3028
rect -19432 -3452 -19368 -3028
rect -18420 -3452 -18356 -3028
rect -17408 -3452 -17344 -3028
rect -16396 -3452 -16332 -3028
rect -15384 -3452 -15320 -3028
rect -14372 -3452 -14308 -3028
rect -13360 -3452 -13296 -3028
rect -12348 -3452 -12284 -3028
rect -11336 -3452 -11272 -3028
rect -10324 -3452 -10260 -3028
rect -9312 -3452 -9248 -3028
rect -8300 -3452 -8236 -3028
rect -7288 -3452 -7224 -3028
rect -6276 -3452 -6212 -3028
rect -5264 -3452 -5200 -3028
rect -4252 -3452 -4188 -3028
rect -3240 -3452 -3176 -3028
rect -2228 -3452 -2164 -3028
rect -1216 -3452 -1152 -3028
rect -204 -3452 -140 -3028
rect 808 -3452 872 -3028
rect 1820 -3452 1884 -3028
rect 2832 -3452 2896 -3028
rect 3844 -3452 3908 -3028
rect 4856 -3452 4920 -3028
rect 5868 -3452 5932 -3028
rect 6880 -3452 6944 -3028
rect 7892 -3452 7956 -3028
rect 8904 -3452 8968 -3028
rect 9916 -3452 9980 -3028
rect 10928 -3452 10992 -3028
rect 11940 -3452 12004 -3028
rect 12952 -3452 13016 -3028
rect 13964 -3452 14028 -3028
rect 14976 -3452 15040 -3028
rect 15988 -3452 16052 -3028
rect 17000 -3452 17064 -3028
rect 18012 -3452 18076 -3028
rect 19024 -3452 19088 -3028
rect 20036 -3452 20100 -3028
rect 21048 -3452 21112 -3028
rect 22060 -3452 22124 -3028
rect 23072 -3452 23136 -3028
rect 24084 -3452 24148 -3028
rect 25096 -3452 25160 -3028
rect 26108 -3452 26172 -3028
rect 27120 -3452 27184 -3028
rect 28132 -3452 28196 -3028
rect 29144 -3452 29208 -3028
rect 30156 -3452 30220 -3028
rect 31168 -3452 31232 -3028
rect 32180 -3452 32244 -3028
rect -31576 -4172 -31512 -3748
rect -30564 -4172 -30500 -3748
rect -29552 -4172 -29488 -3748
rect -28540 -4172 -28476 -3748
rect -27528 -4172 -27464 -3748
rect -26516 -4172 -26452 -3748
rect -25504 -4172 -25440 -3748
rect -24492 -4172 -24428 -3748
rect -23480 -4172 -23416 -3748
rect -22468 -4172 -22404 -3748
rect -21456 -4172 -21392 -3748
rect -20444 -4172 -20380 -3748
rect -19432 -4172 -19368 -3748
rect -18420 -4172 -18356 -3748
rect -17408 -4172 -17344 -3748
rect -16396 -4172 -16332 -3748
rect -15384 -4172 -15320 -3748
rect -14372 -4172 -14308 -3748
rect -13360 -4172 -13296 -3748
rect -12348 -4172 -12284 -3748
rect -11336 -4172 -11272 -3748
rect -10324 -4172 -10260 -3748
rect -9312 -4172 -9248 -3748
rect -8300 -4172 -8236 -3748
rect -7288 -4172 -7224 -3748
rect -6276 -4172 -6212 -3748
rect -5264 -4172 -5200 -3748
rect -4252 -4172 -4188 -3748
rect -3240 -4172 -3176 -3748
rect -2228 -4172 -2164 -3748
rect -1216 -4172 -1152 -3748
rect -204 -4172 -140 -3748
rect 808 -4172 872 -3748
rect 1820 -4172 1884 -3748
rect 2832 -4172 2896 -3748
rect 3844 -4172 3908 -3748
rect 4856 -4172 4920 -3748
rect 5868 -4172 5932 -3748
rect 6880 -4172 6944 -3748
rect 7892 -4172 7956 -3748
rect 8904 -4172 8968 -3748
rect 9916 -4172 9980 -3748
rect 10928 -4172 10992 -3748
rect 11940 -4172 12004 -3748
rect 12952 -4172 13016 -3748
rect 13964 -4172 14028 -3748
rect 14976 -4172 15040 -3748
rect 15988 -4172 16052 -3748
rect 17000 -4172 17064 -3748
rect 18012 -4172 18076 -3748
rect 19024 -4172 19088 -3748
rect 20036 -4172 20100 -3748
rect 21048 -4172 21112 -3748
rect 22060 -4172 22124 -3748
rect 23072 -4172 23136 -3748
rect 24084 -4172 24148 -3748
rect 25096 -4172 25160 -3748
rect 26108 -4172 26172 -3748
rect 27120 -4172 27184 -3748
rect 28132 -4172 28196 -3748
rect 29144 -4172 29208 -3748
rect 30156 -4172 30220 -3748
rect 31168 -4172 31232 -3748
rect 32180 -4172 32244 -3748
rect -31576 -4892 -31512 -4468
rect -30564 -4892 -30500 -4468
rect -29552 -4892 -29488 -4468
rect -28540 -4892 -28476 -4468
rect -27528 -4892 -27464 -4468
rect -26516 -4892 -26452 -4468
rect -25504 -4892 -25440 -4468
rect -24492 -4892 -24428 -4468
rect -23480 -4892 -23416 -4468
rect -22468 -4892 -22404 -4468
rect -21456 -4892 -21392 -4468
rect -20444 -4892 -20380 -4468
rect -19432 -4892 -19368 -4468
rect -18420 -4892 -18356 -4468
rect -17408 -4892 -17344 -4468
rect -16396 -4892 -16332 -4468
rect -15384 -4892 -15320 -4468
rect -14372 -4892 -14308 -4468
rect -13360 -4892 -13296 -4468
rect -12348 -4892 -12284 -4468
rect -11336 -4892 -11272 -4468
rect -10324 -4892 -10260 -4468
rect -9312 -4892 -9248 -4468
rect -8300 -4892 -8236 -4468
rect -7288 -4892 -7224 -4468
rect -6276 -4892 -6212 -4468
rect -5264 -4892 -5200 -4468
rect -4252 -4892 -4188 -4468
rect -3240 -4892 -3176 -4468
rect -2228 -4892 -2164 -4468
rect -1216 -4892 -1152 -4468
rect -204 -4892 -140 -4468
rect 808 -4892 872 -4468
rect 1820 -4892 1884 -4468
rect 2832 -4892 2896 -4468
rect 3844 -4892 3908 -4468
rect 4856 -4892 4920 -4468
rect 5868 -4892 5932 -4468
rect 6880 -4892 6944 -4468
rect 7892 -4892 7956 -4468
rect 8904 -4892 8968 -4468
rect 9916 -4892 9980 -4468
rect 10928 -4892 10992 -4468
rect 11940 -4892 12004 -4468
rect 12952 -4892 13016 -4468
rect 13964 -4892 14028 -4468
rect 14976 -4892 15040 -4468
rect 15988 -4892 16052 -4468
rect 17000 -4892 17064 -4468
rect 18012 -4892 18076 -4468
rect 19024 -4892 19088 -4468
rect 20036 -4892 20100 -4468
rect 21048 -4892 21112 -4468
rect 22060 -4892 22124 -4468
rect 23072 -4892 23136 -4468
rect 24084 -4892 24148 -4468
rect 25096 -4892 25160 -4468
rect 26108 -4892 26172 -4468
rect 27120 -4892 27184 -4468
rect 28132 -4892 28196 -4468
rect 29144 -4892 29208 -4468
rect 30156 -4892 30220 -4468
rect 31168 -4892 31232 -4468
rect 32180 -4892 32244 -4468
rect -31576 -5612 -31512 -5188
rect -30564 -5612 -30500 -5188
rect -29552 -5612 -29488 -5188
rect -28540 -5612 -28476 -5188
rect -27528 -5612 -27464 -5188
rect -26516 -5612 -26452 -5188
rect -25504 -5612 -25440 -5188
rect -24492 -5612 -24428 -5188
rect -23480 -5612 -23416 -5188
rect -22468 -5612 -22404 -5188
rect -21456 -5612 -21392 -5188
rect -20444 -5612 -20380 -5188
rect -19432 -5612 -19368 -5188
rect -18420 -5612 -18356 -5188
rect -17408 -5612 -17344 -5188
rect -16396 -5612 -16332 -5188
rect -15384 -5612 -15320 -5188
rect -14372 -5612 -14308 -5188
rect -13360 -5612 -13296 -5188
rect -12348 -5612 -12284 -5188
rect -11336 -5612 -11272 -5188
rect -10324 -5612 -10260 -5188
rect -9312 -5612 -9248 -5188
rect -8300 -5612 -8236 -5188
rect -7288 -5612 -7224 -5188
rect -6276 -5612 -6212 -5188
rect -5264 -5612 -5200 -5188
rect -4252 -5612 -4188 -5188
rect -3240 -5612 -3176 -5188
rect -2228 -5612 -2164 -5188
rect -1216 -5612 -1152 -5188
rect -204 -5612 -140 -5188
rect 808 -5612 872 -5188
rect 1820 -5612 1884 -5188
rect 2832 -5612 2896 -5188
rect 3844 -5612 3908 -5188
rect 4856 -5612 4920 -5188
rect 5868 -5612 5932 -5188
rect 6880 -5612 6944 -5188
rect 7892 -5612 7956 -5188
rect 8904 -5612 8968 -5188
rect 9916 -5612 9980 -5188
rect 10928 -5612 10992 -5188
rect 11940 -5612 12004 -5188
rect 12952 -5612 13016 -5188
rect 13964 -5612 14028 -5188
rect 14976 -5612 15040 -5188
rect 15988 -5612 16052 -5188
rect 17000 -5612 17064 -5188
rect 18012 -5612 18076 -5188
rect 19024 -5612 19088 -5188
rect 20036 -5612 20100 -5188
rect 21048 -5612 21112 -5188
rect 22060 -5612 22124 -5188
rect 23072 -5612 23136 -5188
rect 24084 -5612 24148 -5188
rect 25096 -5612 25160 -5188
rect 26108 -5612 26172 -5188
rect 27120 -5612 27184 -5188
rect 28132 -5612 28196 -5188
rect 29144 -5612 29208 -5188
rect 30156 -5612 30220 -5188
rect 31168 -5612 31232 -5188
rect 32180 -5612 32244 -5188
<< mimcap >>
rect -32224 5560 -31824 5600
rect -32224 5240 -32184 5560
rect -31864 5240 -31824 5560
rect -32224 5200 -31824 5240
rect -31212 5560 -30812 5600
rect -31212 5240 -31172 5560
rect -30852 5240 -30812 5560
rect -31212 5200 -30812 5240
rect -30200 5560 -29800 5600
rect -30200 5240 -30160 5560
rect -29840 5240 -29800 5560
rect -30200 5200 -29800 5240
rect -29188 5560 -28788 5600
rect -29188 5240 -29148 5560
rect -28828 5240 -28788 5560
rect -29188 5200 -28788 5240
rect -28176 5560 -27776 5600
rect -28176 5240 -28136 5560
rect -27816 5240 -27776 5560
rect -28176 5200 -27776 5240
rect -27164 5560 -26764 5600
rect -27164 5240 -27124 5560
rect -26804 5240 -26764 5560
rect -27164 5200 -26764 5240
rect -26152 5560 -25752 5600
rect -26152 5240 -26112 5560
rect -25792 5240 -25752 5560
rect -26152 5200 -25752 5240
rect -25140 5560 -24740 5600
rect -25140 5240 -25100 5560
rect -24780 5240 -24740 5560
rect -25140 5200 -24740 5240
rect -24128 5560 -23728 5600
rect -24128 5240 -24088 5560
rect -23768 5240 -23728 5560
rect -24128 5200 -23728 5240
rect -23116 5560 -22716 5600
rect -23116 5240 -23076 5560
rect -22756 5240 -22716 5560
rect -23116 5200 -22716 5240
rect -22104 5560 -21704 5600
rect -22104 5240 -22064 5560
rect -21744 5240 -21704 5560
rect -22104 5200 -21704 5240
rect -21092 5560 -20692 5600
rect -21092 5240 -21052 5560
rect -20732 5240 -20692 5560
rect -21092 5200 -20692 5240
rect -20080 5560 -19680 5600
rect -20080 5240 -20040 5560
rect -19720 5240 -19680 5560
rect -20080 5200 -19680 5240
rect -19068 5560 -18668 5600
rect -19068 5240 -19028 5560
rect -18708 5240 -18668 5560
rect -19068 5200 -18668 5240
rect -18056 5560 -17656 5600
rect -18056 5240 -18016 5560
rect -17696 5240 -17656 5560
rect -18056 5200 -17656 5240
rect -17044 5560 -16644 5600
rect -17044 5240 -17004 5560
rect -16684 5240 -16644 5560
rect -17044 5200 -16644 5240
rect -16032 5560 -15632 5600
rect -16032 5240 -15992 5560
rect -15672 5240 -15632 5560
rect -16032 5200 -15632 5240
rect -15020 5560 -14620 5600
rect -15020 5240 -14980 5560
rect -14660 5240 -14620 5560
rect -15020 5200 -14620 5240
rect -14008 5560 -13608 5600
rect -14008 5240 -13968 5560
rect -13648 5240 -13608 5560
rect -14008 5200 -13608 5240
rect -12996 5560 -12596 5600
rect -12996 5240 -12956 5560
rect -12636 5240 -12596 5560
rect -12996 5200 -12596 5240
rect -11984 5560 -11584 5600
rect -11984 5240 -11944 5560
rect -11624 5240 -11584 5560
rect -11984 5200 -11584 5240
rect -10972 5560 -10572 5600
rect -10972 5240 -10932 5560
rect -10612 5240 -10572 5560
rect -10972 5200 -10572 5240
rect -9960 5560 -9560 5600
rect -9960 5240 -9920 5560
rect -9600 5240 -9560 5560
rect -9960 5200 -9560 5240
rect -8948 5560 -8548 5600
rect -8948 5240 -8908 5560
rect -8588 5240 -8548 5560
rect -8948 5200 -8548 5240
rect -7936 5560 -7536 5600
rect -7936 5240 -7896 5560
rect -7576 5240 -7536 5560
rect -7936 5200 -7536 5240
rect -6924 5560 -6524 5600
rect -6924 5240 -6884 5560
rect -6564 5240 -6524 5560
rect -6924 5200 -6524 5240
rect -5912 5560 -5512 5600
rect -5912 5240 -5872 5560
rect -5552 5240 -5512 5560
rect -5912 5200 -5512 5240
rect -4900 5560 -4500 5600
rect -4900 5240 -4860 5560
rect -4540 5240 -4500 5560
rect -4900 5200 -4500 5240
rect -3888 5560 -3488 5600
rect -3888 5240 -3848 5560
rect -3528 5240 -3488 5560
rect -3888 5200 -3488 5240
rect -2876 5560 -2476 5600
rect -2876 5240 -2836 5560
rect -2516 5240 -2476 5560
rect -2876 5200 -2476 5240
rect -1864 5560 -1464 5600
rect -1864 5240 -1824 5560
rect -1504 5240 -1464 5560
rect -1864 5200 -1464 5240
rect -852 5560 -452 5600
rect -852 5240 -812 5560
rect -492 5240 -452 5560
rect -852 5200 -452 5240
rect 160 5560 560 5600
rect 160 5240 200 5560
rect 520 5240 560 5560
rect 160 5200 560 5240
rect 1172 5560 1572 5600
rect 1172 5240 1212 5560
rect 1532 5240 1572 5560
rect 1172 5200 1572 5240
rect 2184 5560 2584 5600
rect 2184 5240 2224 5560
rect 2544 5240 2584 5560
rect 2184 5200 2584 5240
rect 3196 5560 3596 5600
rect 3196 5240 3236 5560
rect 3556 5240 3596 5560
rect 3196 5200 3596 5240
rect 4208 5560 4608 5600
rect 4208 5240 4248 5560
rect 4568 5240 4608 5560
rect 4208 5200 4608 5240
rect 5220 5560 5620 5600
rect 5220 5240 5260 5560
rect 5580 5240 5620 5560
rect 5220 5200 5620 5240
rect 6232 5560 6632 5600
rect 6232 5240 6272 5560
rect 6592 5240 6632 5560
rect 6232 5200 6632 5240
rect 7244 5560 7644 5600
rect 7244 5240 7284 5560
rect 7604 5240 7644 5560
rect 7244 5200 7644 5240
rect 8256 5560 8656 5600
rect 8256 5240 8296 5560
rect 8616 5240 8656 5560
rect 8256 5200 8656 5240
rect 9268 5560 9668 5600
rect 9268 5240 9308 5560
rect 9628 5240 9668 5560
rect 9268 5200 9668 5240
rect 10280 5560 10680 5600
rect 10280 5240 10320 5560
rect 10640 5240 10680 5560
rect 10280 5200 10680 5240
rect 11292 5560 11692 5600
rect 11292 5240 11332 5560
rect 11652 5240 11692 5560
rect 11292 5200 11692 5240
rect 12304 5560 12704 5600
rect 12304 5240 12344 5560
rect 12664 5240 12704 5560
rect 12304 5200 12704 5240
rect 13316 5560 13716 5600
rect 13316 5240 13356 5560
rect 13676 5240 13716 5560
rect 13316 5200 13716 5240
rect 14328 5560 14728 5600
rect 14328 5240 14368 5560
rect 14688 5240 14728 5560
rect 14328 5200 14728 5240
rect 15340 5560 15740 5600
rect 15340 5240 15380 5560
rect 15700 5240 15740 5560
rect 15340 5200 15740 5240
rect 16352 5560 16752 5600
rect 16352 5240 16392 5560
rect 16712 5240 16752 5560
rect 16352 5200 16752 5240
rect 17364 5560 17764 5600
rect 17364 5240 17404 5560
rect 17724 5240 17764 5560
rect 17364 5200 17764 5240
rect 18376 5560 18776 5600
rect 18376 5240 18416 5560
rect 18736 5240 18776 5560
rect 18376 5200 18776 5240
rect 19388 5560 19788 5600
rect 19388 5240 19428 5560
rect 19748 5240 19788 5560
rect 19388 5200 19788 5240
rect 20400 5560 20800 5600
rect 20400 5240 20440 5560
rect 20760 5240 20800 5560
rect 20400 5200 20800 5240
rect 21412 5560 21812 5600
rect 21412 5240 21452 5560
rect 21772 5240 21812 5560
rect 21412 5200 21812 5240
rect 22424 5560 22824 5600
rect 22424 5240 22464 5560
rect 22784 5240 22824 5560
rect 22424 5200 22824 5240
rect 23436 5560 23836 5600
rect 23436 5240 23476 5560
rect 23796 5240 23836 5560
rect 23436 5200 23836 5240
rect 24448 5560 24848 5600
rect 24448 5240 24488 5560
rect 24808 5240 24848 5560
rect 24448 5200 24848 5240
rect 25460 5560 25860 5600
rect 25460 5240 25500 5560
rect 25820 5240 25860 5560
rect 25460 5200 25860 5240
rect 26472 5560 26872 5600
rect 26472 5240 26512 5560
rect 26832 5240 26872 5560
rect 26472 5200 26872 5240
rect 27484 5560 27884 5600
rect 27484 5240 27524 5560
rect 27844 5240 27884 5560
rect 27484 5200 27884 5240
rect 28496 5560 28896 5600
rect 28496 5240 28536 5560
rect 28856 5240 28896 5560
rect 28496 5200 28896 5240
rect 29508 5560 29908 5600
rect 29508 5240 29548 5560
rect 29868 5240 29908 5560
rect 29508 5200 29908 5240
rect 30520 5560 30920 5600
rect 30520 5240 30560 5560
rect 30880 5240 30920 5560
rect 30520 5200 30920 5240
rect 31532 5560 31932 5600
rect 31532 5240 31572 5560
rect 31892 5240 31932 5560
rect 31532 5200 31932 5240
rect -32224 4840 -31824 4880
rect -32224 4520 -32184 4840
rect -31864 4520 -31824 4840
rect -32224 4480 -31824 4520
rect -31212 4840 -30812 4880
rect -31212 4520 -31172 4840
rect -30852 4520 -30812 4840
rect -31212 4480 -30812 4520
rect -30200 4840 -29800 4880
rect -30200 4520 -30160 4840
rect -29840 4520 -29800 4840
rect -30200 4480 -29800 4520
rect -29188 4840 -28788 4880
rect -29188 4520 -29148 4840
rect -28828 4520 -28788 4840
rect -29188 4480 -28788 4520
rect -28176 4840 -27776 4880
rect -28176 4520 -28136 4840
rect -27816 4520 -27776 4840
rect -28176 4480 -27776 4520
rect -27164 4840 -26764 4880
rect -27164 4520 -27124 4840
rect -26804 4520 -26764 4840
rect -27164 4480 -26764 4520
rect -26152 4840 -25752 4880
rect -26152 4520 -26112 4840
rect -25792 4520 -25752 4840
rect -26152 4480 -25752 4520
rect -25140 4840 -24740 4880
rect -25140 4520 -25100 4840
rect -24780 4520 -24740 4840
rect -25140 4480 -24740 4520
rect -24128 4840 -23728 4880
rect -24128 4520 -24088 4840
rect -23768 4520 -23728 4840
rect -24128 4480 -23728 4520
rect -23116 4840 -22716 4880
rect -23116 4520 -23076 4840
rect -22756 4520 -22716 4840
rect -23116 4480 -22716 4520
rect -22104 4840 -21704 4880
rect -22104 4520 -22064 4840
rect -21744 4520 -21704 4840
rect -22104 4480 -21704 4520
rect -21092 4840 -20692 4880
rect -21092 4520 -21052 4840
rect -20732 4520 -20692 4840
rect -21092 4480 -20692 4520
rect -20080 4840 -19680 4880
rect -20080 4520 -20040 4840
rect -19720 4520 -19680 4840
rect -20080 4480 -19680 4520
rect -19068 4840 -18668 4880
rect -19068 4520 -19028 4840
rect -18708 4520 -18668 4840
rect -19068 4480 -18668 4520
rect -18056 4840 -17656 4880
rect -18056 4520 -18016 4840
rect -17696 4520 -17656 4840
rect -18056 4480 -17656 4520
rect -17044 4840 -16644 4880
rect -17044 4520 -17004 4840
rect -16684 4520 -16644 4840
rect -17044 4480 -16644 4520
rect -16032 4840 -15632 4880
rect -16032 4520 -15992 4840
rect -15672 4520 -15632 4840
rect -16032 4480 -15632 4520
rect -15020 4840 -14620 4880
rect -15020 4520 -14980 4840
rect -14660 4520 -14620 4840
rect -15020 4480 -14620 4520
rect -14008 4840 -13608 4880
rect -14008 4520 -13968 4840
rect -13648 4520 -13608 4840
rect -14008 4480 -13608 4520
rect -12996 4840 -12596 4880
rect -12996 4520 -12956 4840
rect -12636 4520 -12596 4840
rect -12996 4480 -12596 4520
rect -11984 4840 -11584 4880
rect -11984 4520 -11944 4840
rect -11624 4520 -11584 4840
rect -11984 4480 -11584 4520
rect -10972 4840 -10572 4880
rect -10972 4520 -10932 4840
rect -10612 4520 -10572 4840
rect -10972 4480 -10572 4520
rect -9960 4840 -9560 4880
rect -9960 4520 -9920 4840
rect -9600 4520 -9560 4840
rect -9960 4480 -9560 4520
rect -8948 4840 -8548 4880
rect -8948 4520 -8908 4840
rect -8588 4520 -8548 4840
rect -8948 4480 -8548 4520
rect -7936 4840 -7536 4880
rect -7936 4520 -7896 4840
rect -7576 4520 -7536 4840
rect -7936 4480 -7536 4520
rect -6924 4840 -6524 4880
rect -6924 4520 -6884 4840
rect -6564 4520 -6524 4840
rect -6924 4480 -6524 4520
rect -5912 4840 -5512 4880
rect -5912 4520 -5872 4840
rect -5552 4520 -5512 4840
rect -5912 4480 -5512 4520
rect -4900 4840 -4500 4880
rect -4900 4520 -4860 4840
rect -4540 4520 -4500 4840
rect -4900 4480 -4500 4520
rect -3888 4840 -3488 4880
rect -3888 4520 -3848 4840
rect -3528 4520 -3488 4840
rect -3888 4480 -3488 4520
rect -2876 4840 -2476 4880
rect -2876 4520 -2836 4840
rect -2516 4520 -2476 4840
rect -2876 4480 -2476 4520
rect -1864 4840 -1464 4880
rect -1864 4520 -1824 4840
rect -1504 4520 -1464 4840
rect -1864 4480 -1464 4520
rect -852 4840 -452 4880
rect -852 4520 -812 4840
rect -492 4520 -452 4840
rect -852 4480 -452 4520
rect 160 4840 560 4880
rect 160 4520 200 4840
rect 520 4520 560 4840
rect 160 4480 560 4520
rect 1172 4840 1572 4880
rect 1172 4520 1212 4840
rect 1532 4520 1572 4840
rect 1172 4480 1572 4520
rect 2184 4840 2584 4880
rect 2184 4520 2224 4840
rect 2544 4520 2584 4840
rect 2184 4480 2584 4520
rect 3196 4840 3596 4880
rect 3196 4520 3236 4840
rect 3556 4520 3596 4840
rect 3196 4480 3596 4520
rect 4208 4840 4608 4880
rect 4208 4520 4248 4840
rect 4568 4520 4608 4840
rect 4208 4480 4608 4520
rect 5220 4840 5620 4880
rect 5220 4520 5260 4840
rect 5580 4520 5620 4840
rect 5220 4480 5620 4520
rect 6232 4840 6632 4880
rect 6232 4520 6272 4840
rect 6592 4520 6632 4840
rect 6232 4480 6632 4520
rect 7244 4840 7644 4880
rect 7244 4520 7284 4840
rect 7604 4520 7644 4840
rect 7244 4480 7644 4520
rect 8256 4840 8656 4880
rect 8256 4520 8296 4840
rect 8616 4520 8656 4840
rect 8256 4480 8656 4520
rect 9268 4840 9668 4880
rect 9268 4520 9308 4840
rect 9628 4520 9668 4840
rect 9268 4480 9668 4520
rect 10280 4840 10680 4880
rect 10280 4520 10320 4840
rect 10640 4520 10680 4840
rect 10280 4480 10680 4520
rect 11292 4840 11692 4880
rect 11292 4520 11332 4840
rect 11652 4520 11692 4840
rect 11292 4480 11692 4520
rect 12304 4840 12704 4880
rect 12304 4520 12344 4840
rect 12664 4520 12704 4840
rect 12304 4480 12704 4520
rect 13316 4840 13716 4880
rect 13316 4520 13356 4840
rect 13676 4520 13716 4840
rect 13316 4480 13716 4520
rect 14328 4840 14728 4880
rect 14328 4520 14368 4840
rect 14688 4520 14728 4840
rect 14328 4480 14728 4520
rect 15340 4840 15740 4880
rect 15340 4520 15380 4840
rect 15700 4520 15740 4840
rect 15340 4480 15740 4520
rect 16352 4840 16752 4880
rect 16352 4520 16392 4840
rect 16712 4520 16752 4840
rect 16352 4480 16752 4520
rect 17364 4840 17764 4880
rect 17364 4520 17404 4840
rect 17724 4520 17764 4840
rect 17364 4480 17764 4520
rect 18376 4840 18776 4880
rect 18376 4520 18416 4840
rect 18736 4520 18776 4840
rect 18376 4480 18776 4520
rect 19388 4840 19788 4880
rect 19388 4520 19428 4840
rect 19748 4520 19788 4840
rect 19388 4480 19788 4520
rect 20400 4840 20800 4880
rect 20400 4520 20440 4840
rect 20760 4520 20800 4840
rect 20400 4480 20800 4520
rect 21412 4840 21812 4880
rect 21412 4520 21452 4840
rect 21772 4520 21812 4840
rect 21412 4480 21812 4520
rect 22424 4840 22824 4880
rect 22424 4520 22464 4840
rect 22784 4520 22824 4840
rect 22424 4480 22824 4520
rect 23436 4840 23836 4880
rect 23436 4520 23476 4840
rect 23796 4520 23836 4840
rect 23436 4480 23836 4520
rect 24448 4840 24848 4880
rect 24448 4520 24488 4840
rect 24808 4520 24848 4840
rect 24448 4480 24848 4520
rect 25460 4840 25860 4880
rect 25460 4520 25500 4840
rect 25820 4520 25860 4840
rect 25460 4480 25860 4520
rect 26472 4840 26872 4880
rect 26472 4520 26512 4840
rect 26832 4520 26872 4840
rect 26472 4480 26872 4520
rect 27484 4840 27884 4880
rect 27484 4520 27524 4840
rect 27844 4520 27884 4840
rect 27484 4480 27884 4520
rect 28496 4840 28896 4880
rect 28496 4520 28536 4840
rect 28856 4520 28896 4840
rect 28496 4480 28896 4520
rect 29508 4840 29908 4880
rect 29508 4520 29548 4840
rect 29868 4520 29908 4840
rect 29508 4480 29908 4520
rect 30520 4840 30920 4880
rect 30520 4520 30560 4840
rect 30880 4520 30920 4840
rect 30520 4480 30920 4520
rect 31532 4840 31932 4880
rect 31532 4520 31572 4840
rect 31892 4520 31932 4840
rect 31532 4480 31932 4520
rect -32224 4120 -31824 4160
rect -32224 3800 -32184 4120
rect -31864 3800 -31824 4120
rect -32224 3760 -31824 3800
rect -31212 4120 -30812 4160
rect -31212 3800 -31172 4120
rect -30852 3800 -30812 4120
rect -31212 3760 -30812 3800
rect -30200 4120 -29800 4160
rect -30200 3800 -30160 4120
rect -29840 3800 -29800 4120
rect -30200 3760 -29800 3800
rect -29188 4120 -28788 4160
rect -29188 3800 -29148 4120
rect -28828 3800 -28788 4120
rect -29188 3760 -28788 3800
rect -28176 4120 -27776 4160
rect -28176 3800 -28136 4120
rect -27816 3800 -27776 4120
rect -28176 3760 -27776 3800
rect -27164 4120 -26764 4160
rect -27164 3800 -27124 4120
rect -26804 3800 -26764 4120
rect -27164 3760 -26764 3800
rect -26152 4120 -25752 4160
rect -26152 3800 -26112 4120
rect -25792 3800 -25752 4120
rect -26152 3760 -25752 3800
rect -25140 4120 -24740 4160
rect -25140 3800 -25100 4120
rect -24780 3800 -24740 4120
rect -25140 3760 -24740 3800
rect -24128 4120 -23728 4160
rect -24128 3800 -24088 4120
rect -23768 3800 -23728 4120
rect -24128 3760 -23728 3800
rect -23116 4120 -22716 4160
rect -23116 3800 -23076 4120
rect -22756 3800 -22716 4120
rect -23116 3760 -22716 3800
rect -22104 4120 -21704 4160
rect -22104 3800 -22064 4120
rect -21744 3800 -21704 4120
rect -22104 3760 -21704 3800
rect -21092 4120 -20692 4160
rect -21092 3800 -21052 4120
rect -20732 3800 -20692 4120
rect -21092 3760 -20692 3800
rect -20080 4120 -19680 4160
rect -20080 3800 -20040 4120
rect -19720 3800 -19680 4120
rect -20080 3760 -19680 3800
rect -19068 4120 -18668 4160
rect -19068 3800 -19028 4120
rect -18708 3800 -18668 4120
rect -19068 3760 -18668 3800
rect -18056 4120 -17656 4160
rect -18056 3800 -18016 4120
rect -17696 3800 -17656 4120
rect -18056 3760 -17656 3800
rect -17044 4120 -16644 4160
rect -17044 3800 -17004 4120
rect -16684 3800 -16644 4120
rect -17044 3760 -16644 3800
rect -16032 4120 -15632 4160
rect -16032 3800 -15992 4120
rect -15672 3800 -15632 4120
rect -16032 3760 -15632 3800
rect -15020 4120 -14620 4160
rect -15020 3800 -14980 4120
rect -14660 3800 -14620 4120
rect -15020 3760 -14620 3800
rect -14008 4120 -13608 4160
rect -14008 3800 -13968 4120
rect -13648 3800 -13608 4120
rect -14008 3760 -13608 3800
rect -12996 4120 -12596 4160
rect -12996 3800 -12956 4120
rect -12636 3800 -12596 4120
rect -12996 3760 -12596 3800
rect -11984 4120 -11584 4160
rect -11984 3800 -11944 4120
rect -11624 3800 -11584 4120
rect -11984 3760 -11584 3800
rect -10972 4120 -10572 4160
rect -10972 3800 -10932 4120
rect -10612 3800 -10572 4120
rect -10972 3760 -10572 3800
rect -9960 4120 -9560 4160
rect -9960 3800 -9920 4120
rect -9600 3800 -9560 4120
rect -9960 3760 -9560 3800
rect -8948 4120 -8548 4160
rect -8948 3800 -8908 4120
rect -8588 3800 -8548 4120
rect -8948 3760 -8548 3800
rect -7936 4120 -7536 4160
rect -7936 3800 -7896 4120
rect -7576 3800 -7536 4120
rect -7936 3760 -7536 3800
rect -6924 4120 -6524 4160
rect -6924 3800 -6884 4120
rect -6564 3800 -6524 4120
rect -6924 3760 -6524 3800
rect -5912 4120 -5512 4160
rect -5912 3800 -5872 4120
rect -5552 3800 -5512 4120
rect -5912 3760 -5512 3800
rect -4900 4120 -4500 4160
rect -4900 3800 -4860 4120
rect -4540 3800 -4500 4120
rect -4900 3760 -4500 3800
rect -3888 4120 -3488 4160
rect -3888 3800 -3848 4120
rect -3528 3800 -3488 4120
rect -3888 3760 -3488 3800
rect -2876 4120 -2476 4160
rect -2876 3800 -2836 4120
rect -2516 3800 -2476 4120
rect -2876 3760 -2476 3800
rect -1864 4120 -1464 4160
rect -1864 3800 -1824 4120
rect -1504 3800 -1464 4120
rect -1864 3760 -1464 3800
rect -852 4120 -452 4160
rect -852 3800 -812 4120
rect -492 3800 -452 4120
rect -852 3760 -452 3800
rect 160 4120 560 4160
rect 160 3800 200 4120
rect 520 3800 560 4120
rect 160 3760 560 3800
rect 1172 4120 1572 4160
rect 1172 3800 1212 4120
rect 1532 3800 1572 4120
rect 1172 3760 1572 3800
rect 2184 4120 2584 4160
rect 2184 3800 2224 4120
rect 2544 3800 2584 4120
rect 2184 3760 2584 3800
rect 3196 4120 3596 4160
rect 3196 3800 3236 4120
rect 3556 3800 3596 4120
rect 3196 3760 3596 3800
rect 4208 4120 4608 4160
rect 4208 3800 4248 4120
rect 4568 3800 4608 4120
rect 4208 3760 4608 3800
rect 5220 4120 5620 4160
rect 5220 3800 5260 4120
rect 5580 3800 5620 4120
rect 5220 3760 5620 3800
rect 6232 4120 6632 4160
rect 6232 3800 6272 4120
rect 6592 3800 6632 4120
rect 6232 3760 6632 3800
rect 7244 4120 7644 4160
rect 7244 3800 7284 4120
rect 7604 3800 7644 4120
rect 7244 3760 7644 3800
rect 8256 4120 8656 4160
rect 8256 3800 8296 4120
rect 8616 3800 8656 4120
rect 8256 3760 8656 3800
rect 9268 4120 9668 4160
rect 9268 3800 9308 4120
rect 9628 3800 9668 4120
rect 9268 3760 9668 3800
rect 10280 4120 10680 4160
rect 10280 3800 10320 4120
rect 10640 3800 10680 4120
rect 10280 3760 10680 3800
rect 11292 4120 11692 4160
rect 11292 3800 11332 4120
rect 11652 3800 11692 4120
rect 11292 3760 11692 3800
rect 12304 4120 12704 4160
rect 12304 3800 12344 4120
rect 12664 3800 12704 4120
rect 12304 3760 12704 3800
rect 13316 4120 13716 4160
rect 13316 3800 13356 4120
rect 13676 3800 13716 4120
rect 13316 3760 13716 3800
rect 14328 4120 14728 4160
rect 14328 3800 14368 4120
rect 14688 3800 14728 4120
rect 14328 3760 14728 3800
rect 15340 4120 15740 4160
rect 15340 3800 15380 4120
rect 15700 3800 15740 4120
rect 15340 3760 15740 3800
rect 16352 4120 16752 4160
rect 16352 3800 16392 4120
rect 16712 3800 16752 4120
rect 16352 3760 16752 3800
rect 17364 4120 17764 4160
rect 17364 3800 17404 4120
rect 17724 3800 17764 4120
rect 17364 3760 17764 3800
rect 18376 4120 18776 4160
rect 18376 3800 18416 4120
rect 18736 3800 18776 4120
rect 18376 3760 18776 3800
rect 19388 4120 19788 4160
rect 19388 3800 19428 4120
rect 19748 3800 19788 4120
rect 19388 3760 19788 3800
rect 20400 4120 20800 4160
rect 20400 3800 20440 4120
rect 20760 3800 20800 4120
rect 20400 3760 20800 3800
rect 21412 4120 21812 4160
rect 21412 3800 21452 4120
rect 21772 3800 21812 4120
rect 21412 3760 21812 3800
rect 22424 4120 22824 4160
rect 22424 3800 22464 4120
rect 22784 3800 22824 4120
rect 22424 3760 22824 3800
rect 23436 4120 23836 4160
rect 23436 3800 23476 4120
rect 23796 3800 23836 4120
rect 23436 3760 23836 3800
rect 24448 4120 24848 4160
rect 24448 3800 24488 4120
rect 24808 3800 24848 4120
rect 24448 3760 24848 3800
rect 25460 4120 25860 4160
rect 25460 3800 25500 4120
rect 25820 3800 25860 4120
rect 25460 3760 25860 3800
rect 26472 4120 26872 4160
rect 26472 3800 26512 4120
rect 26832 3800 26872 4120
rect 26472 3760 26872 3800
rect 27484 4120 27884 4160
rect 27484 3800 27524 4120
rect 27844 3800 27884 4120
rect 27484 3760 27884 3800
rect 28496 4120 28896 4160
rect 28496 3800 28536 4120
rect 28856 3800 28896 4120
rect 28496 3760 28896 3800
rect 29508 4120 29908 4160
rect 29508 3800 29548 4120
rect 29868 3800 29908 4120
rect 29508 3760 29908 3800
rect 30520 4120 30920 4160
rect 30520 3800 30560 4120
rect 30880 3800 30920 4120
rect 30520 3760 30920 3800
rect 31532 4120 31932 4160
rect 31532 3800 31572 4120
rect 31892 3800 31932 4120
rect 31532 3760 31932 3800
rect -32224 3400 -31824 3440
rect -32224 3080 -32184 3400
rect -31864 3080 -31824 3400
rect -32224 3040 -31824 3080
rect -31212 3400 -30812 3440
rect -31212 3080 -31172 3400
rect -30852 3080 -30812 3400
rect -31212 3040 -30812 3080
rect -30200 3400 -29800 3440
rect -30200 3080 -30160 3400
rect -29840 3080 -29800 3400
rect -30200 3040 -29800 3080
rect -29188 3400 -28788 3440
rect -29188 3080 -29148 3400
rect -28828 3080 -28788 3400
rect -29188 3040 -28788 3080
rect -28176 3400 -27776 3440
rect -28176 3080 -28136 3400
rect -27816 3080 -27776 3400
rect -28176 3040 -27776 3080
rect -27164 3400 -26764 3440
rect -27164 3080 -27124 3400
rect -26804 3080 -26764 3400
rect -27164 3040 -26764 3080
rect -26152 3400 -25752 3440
rect -26152 3080 -26112 3400
rect -25792 3080 -25752 3400
rect -26152 3040 -25752 3080
rect -25140 3400 -24740 3440
rect -25140 3080 -25100 3400
rect -24780 3080 -24740 3400
rect -25140 3040 -24740 3080
rect -24128 3400 -23728 3440
rect -24128 3080 -24088 3400
rect -23768 3080 -23728 3400
rect -24128 3040 -23728 3080
rect -23116 3400 -22716 3440
rect -23116 3080 -23076 3400
rect -22756 3080 -22716 3400
rect -23116 3040 -22716 3080
rect -22104 3400 -21704 3440
rect -22104 3080 -22064 3400
rect -21744 3080 -21704 3400
rect -22104 3040 -21704 3080
rect -21092 3400 -20692 3440
rect -21092 3080 -21052 3400
rect -20732 3080 -20692 3400
rect -21092 3040 -20692 3080
rect -20080 3400 -19680 3440
rect -20080 3080 -20040 3400
rect -19720 3080 -19680 3400
rect -20080 3040 -19680 3080
rect -19068 3400 -18668 3440
rect -19068 3080 -19028 3400
rect -18708 3080 -18668 3400
rect -19068 3040 -18668 3080
rect -18056 3400 -17656 3440
rect -18056 3080 -18016 3400
rect -17696 3080 -17656 3400
rect -18056 3040 -17656 3080
rect -17044 3400 -16644 3440
rect -17044 3080 -17004 3400
rect -16684 3080 -16644 3400
rect -17044 3040 -16644 3080
rect -16032 3400 -15632 3440
rect -16032 3080 -15992 3400
rect -15672 3080 -15632 3400
rect -16032 3040 -15632 3080
rect -15020 3400 -14620 3440
rect -15020 3080 -14980 3400
rect -14660 3080 -14620 3400
rect -15020 3040 -14620 3080
rect -14008 3400 -13608 3440
rect -14008 3080 -13968 3400
rect -13648 3080 -13608 3400
rect -14008 3040 -13608 3080
rect -12996 3400 -12596 3440
rect -12996 3080 -12956 3400
rect -12636 3080 -12596 3400
rect -12996 3040 -12596 3080
rect -11984 3400 -11584 3440
rect -11984 3080 -11944 3400
rect -11624 3080 -11584 3400
rect -11984 3040 -11584 3080
rect -10972 3400 -10572 3440
rect -10972 3080 -10932 3400
rect -10612 3080 -10572 3400
rect -10972 3040 -10572 3080
rect -9960 3400 -9560 3440
rect -9960 3080 -9920 3400
rect -9600 3080 -9560 3400
rect -9960 3040 -9560 3080
rect -8948 3400 -8548 3440
rect -8948 3080 -8908 3400
rect -8588 3080 -8548 3400
rect -8948 3040 -8548 3080
rect -7936 3400 -7536 3440
rect -7936 3080 -7896 3400
rect -7576 3080 -7536 3400
rect -7936 3040 -7536 3080
rect -6924 3400 -6524 3440
rect -6924 3080 -6884 3400
rect -6564 3080 -6524 3400
rect -6924 3040 -6524 3080
rect -5912 3400 -5512 3440
rect -5912 3080 -5872 3400
rect -5552 3080 -5512 3400
rect -5912 3040 -5512 3080
rect -4900 3400 -4500 3440
rect -4900 3080 -4860 3400
rect -4540 3080 -4500 3400
rect -4900 3040 -4500 3080
rect -3888 3400 -3488 3440
rect -3888 3080 -3848 3400
rect -3528 3080 -3488 3400
rect -3888 3040 -3488 3080
rect -2876 3400 -2476 3440
rect -2876 3080 -2836 3400
rect -2516 3080 -2476 3400
rect -2876 3040 -2476 3080
rect -1864 3400 -1464 3440
rect -1864 3080 -1824 3400
rect -1504 3080 -1464 3400
rect -1864 3040 -1464 3080
rect -852 3400 -452 3440
rect -852 3080 -812 3400
rect -492 3080 -452 3400
rect -852 3040 -452 3080
rect 160 3400 560 3440
rect 160 3080 200 3400
rect 520 3080 560 3400
rect 160 3040 560 3080
rect 1172 3400 1572 3440
rect 1172 3080 1212 3400
rect 1532 3080 1572 3400
rect 1172 3040 1572 3080
rect 2184 3400 2584 3440
rect 2184 3080 2224 3400
rect 2544 3080 2584 3400
rect 2184 3040 2584 3080
rect 3196 3400 3596 3440
rect 3196 3080 3236 3400
rect 3556 3080 3596 3400
rect 3196 3040 3596 3080
rect 4208 3400 4608 3440
rect 4208 3080 4248 3400
rect 4568 3080 4608 3400
rect 4208 3040 4608 3080
rect 5220 3400 5620 3440
rect 5220 3080 5260 3400
rect 5580 3080 5620 3400
rect 5220 3040 5620 3080
rect 6232 3400 6632 3440
rect 6232 3080 6272 3400
rect 6592 3080 6632 3400
rect 6232 3040 6632 3080
rect 7244 3400 7644 3440
rect 7244 3080 7284 3400
rect 7604 3080 7644 3400
rect 7244 3040 7644 3080
rect 8256 3400 8656 3440
rect 8256 3080 8296 3400
rect 8616 3080 8656 3400
rect 8256 3040 8656 3080
rect 9268 3400 9668 3440
rect 9268 3080 9308 3400
rect 9628 3080 9668 3400
rect 9268 3040 9668 3080
rect 10280 3400 10680 3440
rect 10280 3080 10320 3400
rect 10640 3080 10680 3400
rect 10280 3040 10680 3080
rect 11292 3400 11692 3440
rect 11292 3080 11332 3400
rect 11652 3080 11692 3400
rect 11292 3040 11692 3080
rect 12304 3400 12704 3440
rect 12304 3080 12344 3400
rect 12664 3080 12704 3400
rect 12304 3040 12704 3080
rect 13316 3400 13716 3440
rect 13316 3080 13356 3400
rect 13676 3080 13716 3400
rect 13316 3040 13716 3080
rect 14328 3400 14728 3440
rect 14328 3080 14368 3400
rect 14688 3080 14728 3400
rect 14328 3040 14728 3080
rect 15340 3400 15740 3440
rect 15340 3080 15380 3400
rect 15700 3080 15740 3400
rect 15340 3040 15740 3080
rect 16352 3400 16752 3440
rect 16352 3080 16392 3400
rect 16712 3080 16752 3400
rect 16352 3040 16752 3080
rect 17364 3400 17764 3440
rect 17364 3080 17404 3400
rect 17724 3080 17764 3400
rect 17364 3040 17764 3080
rect 18376 3400 18776 3440
rect 18376 3080 18416 3400
rect 18736 3080 18776 3400
rect 18376 3040 18776 3080
rect 19388 3400 19788 3440
rect 19388 3080 19428 3400
rect 19748 3080 19788 3400
rect 19388 3040 19788 3080
rect 20400 3400 20800 3440
rect 20400 3080 20440 3400
rect 20760 3080 20800 3400
rect 20400 3040 20800 3080
rect 21412 3400 21812 3440
rect 21412 3080 21452 3400
rect 21772 3080 21812 3400
rect 21412 3040 21812 3080
rect 22424 3400 22824 3440
rect 22424 3080 22464 3400
rect 22784 3080 22824 3400
rect 22424 3040 22824 3080
rect 23436 3400 23836 3440
rect 23436 3080 23476 3400
rect 23796 3080 23836 3400
rect 23436 3040 23836 3080
rect 24448 3400 24848 3440
rect 24448 3080 24488 3400
rect 24808 3080 24848 3400
rect 24448 3040 24848 3080
rect 25460 3400 25860 3440
rect 25460 3080 25500 3400
rect 25820 3080 25860 3400
rect 25460 3040 25860 3080
rect 26472 3400 26872 3440
rect 26472 3080 26512 3400
rect 26832 3080 26872 3400
rect 26472 3040 26872 3080
rect 27484 3400 27884 3440
rect 27484 3080 27524 3400
rect 27844 3080 27884 3400
rect 27484 3040 27884 3080
rect 28496 3400 28896 3440
rect 28496 3080 28536 3400
rect 28856 3080 28896 3400
rect 28496 3040 28896 3080
rect 29508 3400 29908 3440
rect 29508 3080 29548 3400
rect 29868 3080 29908 3400
rect 29508 3040 29908 3080
rect 30520 3400 30920 3440
rect 30520 3080 30560 3400
rect 30880 3080 30920 3400
rect 30520 3040 30920 3080
rect 31532 3400 31932 3440
rect 31532 3080 31572 3400
rect 31892 3080 31932 3400
rect 31532 3040 31932 3080
rect -32224 2680 -31824 2720
rect -32224 2360 -32184 2680
rect -31864 2360 -31824 2680
rect -32224 2320 -31824 2360
rect -31212 2680 -30812 2720
rect -31212 2360 -31172 2680
rect -30852 2360 -30812 2680
rect -31212 2320 -30812 2360
rect -30200 2680 -29800 2720
rect -30200 2360 -30160 2680
rect -29840 2360 -29800 2680
rect -30200 2320 -29800 2360
rect -29188 2680 -28788 2720
rect -29188 2360 -29148 2680
rect -28828 2360 -28788 2680
rect -29188 2320 -28788 2360
rect -28176 2680 -27776 2720
rect -28176 2360 -28136 2680
rect -27816 2360 -27776 2680
rect -28176 2320 -27776 2360
rect -27164 2680 -26764 2720
rect -27164 2360 -27124 2680
rect -26804 2360 -26764 2680
rect -27164 2320 -26764 2360
rect -26152 2680 -25752 2720
rect -26152 2360 -26112 2680
rect -25792 2360 -25752 2680
rect -26152 2320 -25752 2360
rect -25140 2680 -24740 2720
rect -25140 2360 -25100 2680
rect -24780 2360 -24740 2680
rect -25140 2320 -24740 2360
rect -24128 2680 -23728 2720
rect -24128 2360 -24088 2680
rect -23768 2360 -23728 2680
rect -24128 2320 -23728 2360
rect -23116 2680 -22716 2720
rect -23116 2360 -23076 2680
rect -22756 2360 -22716 2680
rect -23116 2320 -22716 2360
rect -22104 2680 -21704 2720
rect -22104 2360 -22064 2680
rect -21744 2360 -21704 2680
rect -22104 2320 -21704 2360
rect -21092 2680 -20692 2720
rect -21092 2360 -21052 2680
rect -20732 2360 -20692 2680
rect -21092 2320 -20692 2360
rect -20080 2680 -19680 2720
rect -20080 2360 -20040 2680
rect -19720 2360 -19680 2680
rect -20080 2320 -19680 2360
rect -19068 2680 -18668 2720
rect -19068 2360 -19028 2680
rect -18708 2360 -18668 2680
rect -19068 2320 -18668 2360
rect -18056 2680 -17656 2720
rect -18056 2360 -18016 2680
rect -17696 2360 -17656 2680
rect -18056 2320 -17656 2360
rect -17044 2680 -16644 2720
rect -17044 2360 -17004 2680
rect -16684 2360 -16644 2680
rect -17044 2320 -16644 2360
rect -16032 2680 -15632 2720
rect -16032 2360 -15992 2680
rect -15672 2360 -15632 2680
rect -16032 2320 -15632 2360
rect -15020 2680 -14620 2720
rect -15020 2360 -14980 2680
rect -14660 2360 -14620 2680
rect -15020 2320 -14620 2360
rect -14008 2680 -13608 2720
rect -14008 2360 -13968 2680
rect -13648 2360 -13608 2680
rect -14008 2320 -13608 2360
rect -12996 2680 -12596 2720
rect -12996 2360 -12956 2680
rect -12636 2360 -12596 2680
rect -12996 2320 -12596 2360
rect -11984 2680 -11584 2720
rect -11984 2360 -11944 2680
rect -11624 2360 -11584 2680
rect -11984 2320 -11584 2360
rect -10972 2680 -10572 2720
rect -10972 2360 -10932 2680
rect -10612 2360 -10572 2680
rect -10972 2320 -10572 2360
rect -9960 2680 -9560 2720
rect -9960 2360 -9920 2680
rect -9600 2360 -9560 2680
rect -9960 2320 -9560 2360
rect -8948 2680 -8548 2720
rect -8948 2360 -8908 2680
rect -8588 2360 -8548 2680
rect -8948 2320 -8548 2360
rect -7936 2680 -7536 2720
rect -7936 2360 -7896 2680
rect -7576 2360 -7536 2680
rect -7936 2320 -7536 2360
rect -6924 2680 -6524 2720
rect -6924 2360 -6884 2680
rect -6564 2360 -6524 2680
rect -6924 2320 -6524 2360
rect -5912 2680 -5512 2720
rect -5912 2360 -5872 2680
rect -5552 2360 -5512 2680
rect -5912 2320 -5512 2360
rect -4900 2680 -4500 2720
rect -4900 2360 -4860 2680
rect -4540 2360 -4500 2680
rect -4900 2320 -4500 2360
rect -3888 2680 -3488 2720
rect -3888 2360 -3848 2680
rect -3528 2360 -3488 2680
rect -3888 2320 -3488 2360
rect -2876 2680 -2476 2720
rect -2876 2360 -2836 2680
rect -2516 2360 -2476 2680
rect -2876 2320 -2476 2360
rect -1864 2680 -1464 2720
rect -1864 2360 -1824 2680
rect -1504 2360 -1464 2680
rect -1864 2320 -1464 2360
rect -852 2680 -452 2720
rect -852 2360 -812 2680
rect -492 2360 -452 2680
rect -852 2320 -452 2360
rect 160 2680 560 2720
rect 160 2360 200 2680
rect 520 2360 560 2680
rect 160 2320 560 2360
rect 1172 2680 1572 2720
rect 1172 2360 1212 2680
rect 1532 2360 1572 2680
rect 1172 2320 1572 2360
rect 2184 2680 2584 2720
rect 2184 2360 2224 2680
rect 2544 2360 2584 2680
rect 2184 2320 2584 2360
rect 3196 2680 3596 2720
rect 3196 2360 3236 2680
rect 3556 2360 3596 2680
rect 3196 2320 3596 2360
rect 4208 2680 4608 2720
rect 4208 2360 4248 2680
rect 4568 2360 4608 2680
rect 4208 2320 4608 2360
rect 5220 2680 5620 2720
rect 5220 2360 5260 2680
rect 5580 2360 5620 2680
rect 5220 2320 5620 2360
rect 6232 2680 6632 2720
rect 6232 2360 6272 2680
rect 6592 2360 6632 2680
rect 6232 2320 6632 2360
rect 7244 2680 7644 2720
rect 7244 2360 7284 2680
rect 7604 2360 7644 2680
rect 7244 2320 7644 2360
rect 8256 2680 8656 2720
rect 8256 2360 8296 2680
rect 8616 2360 8656 2680
rect 8256 2320 8656 2360
rect 9268 2680 9668 2720
rect 9268 2360 9308 2680
rect 9628 2360 9668 2680
rect 9268 2320 9668 2360
rect 10280 2680 10680 2720
rect 10280 2360 10320 2680
rect 10640 2360 10680 2680
rect 10280 2320 10680 2360
rect 11292 2680 11692 2720
rect 11292 2360 11332 2680
rect 11652 2360 11692 2680
rect 11292 2320 11692 2360
rect 12304 2680 12704 2720
rect 12304 2360 12344 2680
rect 12664 2360 12704 2680
rect 12304 2320 12704 2360
rect 13316 2680 13716 2720
rect 13316 2360 13356 2680
rect 13676 2360 13716 2680
rect 13316 2320 13716 2360
rect 14328 2680 14728 2720
rect 14328 2360 14368 2680
rect 14688 2360 14728 2680
rect 14328 2320 14728 2360
rect 15340 2680 15740 2720
rect 15340 2360 15380 2680
rect 15700 2360 15740 2680
rect 15340 2320 15740 2360
rect 16352 2680 16752 2720
rect 16352 2360 16392 2680
rect 16712 2360 16752 2680
rect 16352 2320 16752 2360
rect 17364 2680 17764 2720
rect 17364 2360 17404 2680
rect 17724 2360 17764 2680
rect 17364 2320 17764 2360
rect 18376 2680 18776 2720
rect 18376 2360 18416 2680
rect 18736 2360 18776 2680
rect 18376 2320 18776 2360
rect 19388 2680 19788 2720
rect 19388 2360 19428 2680
rect 19748 2360 19788 2680
rect 19388 2320 19788 2360
rect 20400 2680 20800 2720
rect 20400 2360 20440 2680
rect 20760 2360 20800 2680
rect 20400 2320 20800 2360
rect 21412 2680 21812 2720
rect 21412 2360 21452 2680
rect 21772 2360 21812 2680
rect 21412 2320 21812 2360
rect 22424 2680 22824 2720
rect 22424 2360 22464 2680
rect 22784 2360 22824 2680
rect 22424 2320 22824 2360
rect 23436 2680 23836 2720
rect 23436 2360 23476 2680
rect 23796 2360 23836 2680
rect 23436 2320 23836 2360
rect 24448 2680 24848 2720
rect 24448 2360 24488 2680
rect 24808 2360 24848 2680
rect 24448 2320 24848 2360
rect 25460 2680 25860 2720
rect 25460 2360 25500 2680
rect 25820 2360 25860 2680
rect 25460 2320 25860 2360
rect 26472 2680 26872 2720
rect 26472 2360 26512 2680
rect 26832 2360 26872 2680
rect 26472 2320 26872 2360
rect 27484 2680 27884 2720
rect 27484 2360 27524 2680
rect 27844 2360 27884 2680
rect 27484 2320 27884 2360
rect 28496 2680 28896 2720
rect 28496 2360 28536 2680
rect 28856 2360 28896 2680
rect 28496 2320 28896 2360
rect 29508 2680 29908 2720
rect 29508 2360 29548 2680
rect 29868 2360 29908 2680
rect 29508 2320 29908 2360
rect 30520 2680 30920 2720
rect 30520 2360 30560 2680
rect 30880 2360 30920 2680
rect 30520 2320 30920 2360
rect 31532 2680 31932 2720
rect 31532 2360 31572 2680
rect 31892 2360 31932 2680
rect 31532 2320 31932 2360
rect -32224 1960 -31824 2000
rect -32224 1640 -32184 1960
rect -31864 1640 -31824 1960
rect -32224 1600 -31824 1640
rect -31212 1960 -30812 2000
rect -31212 1640 -31172 1960
rect -30852 1640 -30812 1960
rect -31212 1600 -30812 1640
rect -30200 1960 -29800 2000
rect -30200 1640 -30160 1960
rect -29840 1640 -29800 1960
rect -30200 1600 -29800 1640
rect -29188 1960 -28788 2000
rect -29188 1640 -29148 1960
rect -28828 1640 -28788 1960
rect -29188 1600 -28788 1640
rect -28176 1960 -27776 2000
rect -28176 1640 -28136 1960
rect -27816 1640 -27776 1960
rect -28176 1600 -27776 1640
rect -27164 1960 -26764 2000
rect -27164 1640 -27124 1960
rect -26804 1640 -26764 1960
rect -27164 1600 -26764 1640
rect -26152 1960 -25752 2000
rect -26152 1640 -26112 1960
rect -25792 1640 -25752 1960
rect -26152 1600 -25752 1640
rect -25140 1960 -24740 2000
rect -25140 1640 -25100 1960
rect -24780 1640 -24740 1960
rect -25140 1600 -24740 1640
rect -24128 1960 -23728 2000
rect -24128 1640 -24088 1960
rect -23768 1640 -23728 1960
rect -24128 1600 -23728 1640
rect -23116 1960 -22716 2000
rect -23116 1640 -23076 1960
rect -22756 1640 -22716 1960
rect -23116 1600 -22716 1640
rect -22104 1960 -21704 2000
rect -22104 1640 -22064 1960
rect -21744 1640 -21704 1960
rect -22104 1600 -21704 1640
rect -21092 1960 -20692 2000
rect -21092 1640 -21052 1960
rect -20732 1640 -20692 1960
rect -21092 1600 -20692 1640
rect -20080 1960 -19680 2000
rect -20080 1640 -20040 1960
rect -19720 1640 -19680 1960
rect -20080 1600 -19680 1640
rect -19068 1960 -18668 2000
rect -19068 1640 -19028 1960
rect -18708 1640 -18668 1960
rect -19068 1600 -18668 1640
rect -18056 1960 -17656 2000
rect -18056 1640 -18016 1960
rect -17696 1640 -17656 1960
rect -18056 1600 -17656 1640
rect -17044 1960 -16644 2000
rect -17044 1640 -17004 1960
rect -16684 1640 -16644 1960
rect -17044 1600 -16644 1640
rect -16032 1960 -15632 2000
rect -16032 1640 -15992 1960
rect -15672 1640 -15632 1960
rect -16032 1600 -15632 1640
rect -15020 1960 -14620 2000
rect -15020 1640 -14980 1960
rect -14660 1640 -14620 1960
rect -15020 1600 -14620 1640
rect -14008 1960 -13608 2000
rect -14008 1640 -13968 1960
rect -13648 1640 -13608 1960
rect -14008 1600 -13608 1640
rect -12996 1960 -12596 2000
rect -12996 1640 -12956 1960
rect -12636 1640 -12596 1960
rect -12996 1600 -12596 1640
rect -11984 1960 -11584 2000
rect -11984 1640 -11944 1960
rect -11624 1640 -11584 1960
rect -11984 1600 -11584 1640
rect -10972 1960 -10572 2000
rect -10972 1640 -10932 1960
rect -10612 1640 -10572 1960
rect -10972 1600 -10572 1640
rect -9960 1960 -9560 2000
rect -9960 1640 -9920 1960
rect -9600 1640 -9560 1960
rect -9960 1600 -9560 1640
rect -8948 1960 -8548 2000
rect -8948 1640 -8908 1960
rect -8588 1640 -8548 1960
rect -8948 1600 -8548 1640
rect -7936 1960 -7536 2000
rect -7936 1640 -7896 1960
rect -7576 1640 -7536 1960
rect -7936 1600 -7536 1640
rect -6924 1960 -6524 2000
rect -6924 1640 -6884 1960
rect -6564 1640 -6524 1960
rect -6924 1600 -6524 1640
rect -5912 1960 -5512 2000
rect -5912 1640 -5872 1960
rect -5552 1640 -5512 1960
rect -5912 1600 -5512 1640
rect -4900 1960 -4500 2000
rect -4900 1640 -4860 1960
rect -4540 1640 -4500 1960
rect -4900 1600 -4500 1640
rect -3888 1960 -3488 2000
rect -3888 1640 -3848 1960
rect -3528 1640 -3488 1960
rect -3888 1600 -3488 1640
rect -2876 1960 -2476 2000
rect -2876 1640 -2836 1960
rect -2516 1640 -2476 1960
rect -2876 1600 -2476 1640
rect -1864 1960 -1464 2000
rect -1864 1640 -1824 1960
rect -1504 1640 -1464 1960
rect -1864 1600 -1464 1640
rect -852 1960 -452 2000
rect -852 1640 -812 1960
rect -492 1640 -452 1960
rect -852 1600 -452 1640
rect 160 1960 560 2000
rect 160 1640 200 1960
rect 520 1640 560 1960
rect 160 1600 560 1640
rect 1172 1960 1572 2000
rect 1172 1640 1212 1960
rect 1532 1640 1572 1960
rect 1172 1600 1572 1640
rect 2184 1960 2584 2000
rect 2184 1640 2224 1960
rect 2544 1640 2584 1960
rect 2184 1600 2584 1640
rect 3196 1960 3596 2000
rect 3196 1640 3236 1960
rect 3556 1640 3596 1960
rect 3196 1600 3596 1640
rect 4208 1960 4608 2000
rect 4208 1640 4248 1960
rect 4568 1640 4608 1960
rect 4208 1600 4608 1640
rect 5220 1960 5620 2000
rect 5220 1640 5260 1960
rect 5580 1640 5620 1960
rect 5220 1600 5620 1640
rect 6232 1960 6632 2000
rect 6232 1640 6272 1960
rect 6592 1640 6632 1960
rect 6232 1600 6632 1640
rect 7244 1960 7644 2000
rect 7244 1640 7284 1960
rect 7604 1640 7644 1960
rect 7244 1600 7644 1640
rect 8256 1960 8656 2000
rect 8256 1640 8296 1960
rect 8616 1640 8656 1960
rect 8256 1600 8656 1640
rect 9268 1960 9668 2000
rect 9268 1640 9308 1960
rect 9628 1640 9668 1960
rect 9268 1600 9668 1640
rect 10280 1960 10680 2000
rect 10280 1640 10320 1960
rect 10640 1640 10680 1960
rect 10280 1600 10680 1640
rect 11292 1960 11692 2000
rect 11292 1640 11332 1960
rect 11652 1640 11692 1960
rect 11292 1600 11692 1640
rect 12304 1960 12704 2000
rect 12304 1640 12344 1960
rect 12664 1640 12704 1960
rect 12304 1600 12704 1640
rect 13316 1960 13716 2000
rect 13316 1640 13356 1960
rect 13676 1640 13716 1960
rect 13316 1600 13716 1640
rect 14328 1960 14728 2000
rect 14328 1640 14368 1960
rect 14688 1640 14728 1960
rect 14328 1600 14728 1640
rect 15340 1960 15740 2000
rect 15340 1640 15380 1960
rect 15700 1640 15740 1960
rect 15340 1600 15740 1640
rect 16352 1960 16752 2000
rect 16352 1640 16392 1960
rect 16712 1640 16752 1960
rect 16352 1600 16752 1640
rect 17364 1960 17764 2000
rect 17364 1640 17404 1960
rect 17724 1640 17764 1960
rect 17364 1600 17764 1640
rect 18376 1960 18776 2000
rect 18376 1640 18416 1960
rect 18736 1640 18776 1960
rect 18376 1600 18776 1640
rect 19388 1960 19788 2000
rect 19388 1640 19428 1960
rect 19748 1640 19788 1960
rect 19388 1600 19788 1640
rect 20400 1960 20800 2000
rect 20400 1640 20440 1960
rect 20760 1640 20800 1960
rect 20400 1600 20800 1640
rect 21412 1960 21812 2000
rect 21412 1640 21452 1960
rect 21772 1640 21812 1960
rect 21412 1600 21812 1640
rect 22424 1960 22824 2000
rect 22424 1640 22464 1960
rect 22784 1640 22824 1960
rect 22424 1600 22824 1640
rect 23436 1960 23836 2000
rect 23436 1640 23476 1960
rect 23796 1640 23836 1960
rect 23436 1600 23836 1640
rect 24448 1960 24848 2000
rect 24448 1640 24488 1960
rect 24808 1640 24848 1960
rect 24448 1600 24848 1640
rect 25460 1960 25860 2000
rect 25460 1640 25500 1960
rect 25820 1640 25860 1960
rect 25460 1600 25860 1640
rect 26472 1960 26872 2000
rect 26472 1640 26512 1960
rect 26832 1640 26872 1960
rect 26472 1600 26872 1640
rect 27484 1960 27884 2000
rect 27484 1640 27524 1960
rect 27844 1640 27884 1960
rect 27484 1600 27884 1640
rect 28496 1960 28896 2000
rect 28496 1640 28536 1960
rect 28856 1640 28896 1960
rect 28496 1600 28896 1640
rect 29508 1960 29908 2000
rect 29508 1640 29548 1960
rect 29868 1640 29908 1960
rect 29508 1600 29908 1640
rect 30520 1960 30920 2000
rect 30520 1640 30560 1960
rect 30880 1640 30920 1960
rect 30520 1600 30920 1640
rect 31532 1960 31932 2000
rect 31532 1640 31572 1960
rect 31892 1640 31932 1960
rect 31532 1600 31932 1640
rect -32224 1240 -31824 1280
rect -32224 920 -32184 1240
rect -31864 920 -31824 1240
rect -32224 880 -31824 920
rect -31212 1240 -30812 1280
rect -31212 920 -31172 1240
rect -30852 920 -30812 1240
rect -31212 880 -30812 920
rect -30200 1240 -29800 1280
rect -30200 920 -30160 1240
rect -29840 920 -29800 1240
rect -30200 880 -29800 920
rect -29188 1240 -28788 1280
rect -29188 920 -29148 1240
rect -28828 920 -28788 1240
rect -29188 880 -28788 920
rect -28176 1240 -27776 1280
rect -28176 920 -28136 1240
rect -27816 920 -27776 1240
rect -28176 880 -27776 920
rect -27164 1240 -26764 1280
rect -27164 920 -27124 1240
rect -26804 920 -26764 1240
rect -27164 880 -26764 920
rect -26152 1240 -25752 1280
rect -26152 920 -26112 1240
rect -25792 920 -25752 1240
rect -26152 880 -25752 920
rect -25140 1240 -24740 1280
rect -25140 920 -25100 1240
rect -24780 920 -24740 1240
rect -25140 880 -24740 920
rect -24128 1240 -23728 1280
rect -24128 920 -24088 1240
rect -23768 920 -23728 1240
rect -24128 880 -23728 920
rect -23116 1240 -22716 1280
rect -23116 920 -23076 1240
rect -22756 920 -22716 1240
rect -23116 880 -22716 920
rect -22104 1240 -21704 1280
rect -22104 920 -22064 1240
rect -21744 920 -21704 1240
rect -22104 880 -21704 920
rect -21092 1240 -20692 1280
rect -21092 920 -21052 1240
rect -20732 920 -20692 1240
rect -21092 880 -20692 920
rect -20080 1240 -19680 1280
rect -20080 920 -20040 1240
rect -19720 920 -19680 1240
rect -20080 880 -19680 920
rect -19068 1240 -18668 1280
rect -19068 920 -19028 1240
rect -18708 920 -18668 1240
rect -19068 880 -18668 920
rect -18056 1240 -17656 1280
rect -18056 920 -18016 1240
rect -17696 920 -17656 1240
rect -18056 880 -17656 920
rect -17044 1240 -16644 1280
rect -17044 920 -17004 1240
rect -16684 920 -16644 1240
rect -17044 880 -16644 920
rect -16032 1240 -15632 1280
rect -16032 920 -15992 1240
rect -15672 920 -15632 1240
rect -16032 880 -15632 920
rect -15020 1240 -14620 1280
rect -15020 920 -14980 1240
rect -14660 920 -14620 1240
rect -15020 880 -14620 920
rect -14008 1240 -13608 1280
rect -14008 920 -13968 1240
rect -13648 920 -13608 1240
rect -14008 880 -13608 920
rect -12996 1240 -12596 1280
rect -12996 920 -12956 1240
rect -12636 920 -12596 1240
rect -12996 880 -12596 920
rect -11984 1240 -11584 1280
rect -11984 920 -11944 1240
rect -11624 920 -11584 1240
rect -11984 880 -11584 920
rect -10972 1240 -10572 1280
rect -10972 920 -10932 1240
rect -10612 920 -10572 1240
rect -10972 880 -10572 920
rect -9960 1240 -9560 1280
rect -9960 920 -9920 1240
rect -9600 920 -9560 1240
rect -9960 880 -9560 920
rect -8948 1240 -8548 1280
rect -8948 920 -8908 1240
rect -8588 920 -8548 1240
rect -8948 880 -8548 920
rect -7936 1240 -7536 1280
rect -7936 920 -7896 1240
rect -7576 920 -7536 1240
rect -7936 880 -7536 920
rect -6924 1240 -6524 1280
rect -6924 920 -6884 1240
rect -6564 920 -6524 1240
rect -6924 880 -6524 920
rect -5912 1240 -5512 1280
rect -5912 920 -5872 1240
rect -5552 920 -5512 1240
rect -5912 880 -5512 920
rect -4900 1240 -4500 1280
rect -4900 920 -4860 1240
rect -4540 920 -4500 1240
rect -4900 880 -4500 920
rect -3888 1240 -3488 1280
rect -3888 920 -3848 1240
rect -3528 920 -3488 1240
rect -3888 880 -3488 920
rect -2876 1240 -2476 1280
rect -2876 920 -2836 1240
rect -2516 920 -2476 1240
rect -2876 880 -2476 920
rect -1864 1240 -1464 1280
rect -1864 920 -1824 1240
rect -1504 920 -1464 1240
rect -1864 880 -1464 920
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect 1172 1240 1572 1280
rect 1172 920 1212 1240
rect 1532 920 1572 1240
rect 1172 880 1572 920
rect 2184 1240 2584 1280
rect 2184 920 2224 1240
rect 2544 920 2584 1240
rect 2184 880 2584 920
rect 3196 1240 3596 1280
rect 3196 920 3236 1240
rect 3556 920 3596 1240
rect 3196 880 3596 920
rect 4208 1240 4608 1280
rect 4208 920 4248 1240
rect 4568 920 4608 1240
rect 4208 880 4608 920
rect 5220 1240 5620 1280
rect 5220 920 5260 1240
rect 5580 920 5620 1240
rect 5220 880 5620 920
rect 6232 1240 6632 1280
rect 6232 920 6272 1240
rect 6592 920 6632 1240
rect 6232 880 6632 920
rect 7244 1240 7644 1280
rect 7244 920 7284 1240
rect 7604 920 7644 1240
rect 7244 880 7644 920
rect 8256 1240 8656 1280
rect 8256 920 8296 1240
rect 8616 920 8656 1240
rect 8256 880 8656 920
rect 9268 1240 9668 1280
rect 9268 920 9308 1240
rect 9628 920 9668 1240
rect 9268 880 9668 920
rect 10280 1240 10680 1280
rect 10280 920 10320 1240
rect 10640 920 10680 1240
rect 10280 880 10680 920
rect 11292 1240 11692 1280
rect 11292 920 11332 1240
rect 11652 920 11692 1240
rect 11292 880 11692 920
rect 12304 1240 12704 1280
rect 12304 920 12344 1240
rect 12664 920 12704 1240
rect 12304 880 12704 920
rect 13316 1240 13716 1280
rect 13316 920 13356 1240
rect 13676 920 13716 1240
rect 13316 880 13716 920
rect 14328 1240 14728 1280
rect 14328 920 14368 1240
rect 14688 920 14728 1240
rect 14328 880 14728 920
rect 15340 1240 15740 1280
rect 15340 920 15380 1240
rect 15700 920 15740 1240
rect 15340 880 15740 920
rect 16352 1240 16752 1280
rect 16352 920 16392 1240
rect 16712 920 16752 1240
rect 16352 880 16752 920
rect 17364 1240 17764 1280
rect 17364 920 17404 1240
rect 17724 920 17764 1240
rect 17364 880 17764 920
rect 18376 1240 18776 1280
rect 18376 920 18416 1240
rect 18736 920 18776 1240
rect 18376 880 18776 920
rect 19388 1240 19788 1280
rect 19388 920 19428 1240
rect 19748 920 19788 1240
rect 19388 880 19788 920
rect 20400 1240 20800 1280
rect 20400 920 20440 1240
rect 20760 920 20800 1240
rect 20400 880 20800 920
rect 21412 1240 21812 1280
rect 21412 920 21452 1240
rect 21772 920 21812 1240
rect 21412 880 21812 920
rect 22424 1240 22824 1280
rect 22424 920 22464 1240
rect 22784 920 22824 1240
rect 22424 880 22824 920
rect 23436 1240 23836 1280
rect 23436 920 23476 1240
rect 23796 920 23836 1240
rect 23436 880 23836 920
rect 24448 1240 24848 1280
rect 24448 920 24488 1240
rect 24808 920 24848 1240
rect 24448 880 24848 920
rect 25460 1240 25860 1280
rect 25460 920 25500 1240
rect 25820 920 25860 1240
rect 25460 880 25860 920
rect 26472 1240 26872 1280
rect 26472 920 26512 1240
rect 26832 920 26872 1240
rect 26472 880 26872 920
rect 27484 1240 27884 1280
rect 27484 920 27524 1240
rect 27844 920 27884 1240
rect 27484 880 27884 920
rect 28496 1240 28896 1280
rect 28496 920 28536 1240
rect 28856 920 28896 1240
rect 28496 880 28896 920
rect 29508 1240 29908 1280
rect 29508 920 29548 1240
rect 29868 920 29908 1240
rect 29508 880 29908 920
rect 30520 1240 30920 1280
rect 30520 920 30560 1240
rect 30880 920 30920 1240
rect 30520 880 30920 920
rect 31532 1240 31932 1280
rect 31532 920 31572 1240
rect 31892 920 31932 1240
rect 31532 880 31932 920
rect -32224 520 -31824 560
rect -32224 200 -32184 520
rect -31864 200 -31824 520
rect -32224 160 -31824 200
rect -31212 520 -30812 560
rect -31212 200 -31172 520
rect -30852 200 -30812 520
rect -31212 160 -30812 200
rect -30200 520 -29800 560
rect -30200 200 -30160 520
rect -29840 200 -29800 520
rect -30200 160 -29800 200
rect -29188 520 -28788 560
rect -29188 200 -29148 520
rect -28828 200 -28788 520
rect -29188 160 -28788 200
rect -28176 520 -27776 560
rect -28176 200 -28136 520
rect -27816 200 -27776 520
rect -28176 160 -27776 200
rect -27164 520 -26764 560
rect -27164 200 -27124 520
rect -26804 200 -26764 520
rect -27164 160 -26764 200
rect -26152 520 -25752 560
rect -26152 200 -26112 520
rect -25792 200 -25752 520
rect -26152 160 -25752 200
rect -25140 520 -24740 560
rect -25140 200 -25100 520
rect -24780 200 -24740 520
rect -25140 160 -24740 200
rect -24128 520 -23728 560
rect -24128 200 -24088 520
rect -23768 200 -23728 520
rect -24128 160 -23728 200
rect -23116 520 -22716 560
rect -23116 200 -23076 520
rect -22756 200 -22716 520
rect -23116 160 -22716 200
rect -22104 520 -21704 560
rect -22104 200 -22064 520
rect -21744 200 -21704 520
rect -22104 160 -21704 200
rect -21092 520 -20692 560
rect -21092 200 -21052 520
rect -20732 200 -20692 520
rect -21092 160 -20692 200
rect -20080 520 -19680 560
rect -20080 200 -20040 520
rect -19720 200 -19680 520
rect -20080 160 -19680 200
rect -19068 520 -18668 560
rect -19068 200 -19028 520
rect -18708 200 -18668 520
rect -19068 160 -18668 200
rect -18056 520 -17656 560
rect -18056 200 -18016 520
rect -17696 200 -17656 520
rect -18056 160 -17656 200
rect -17044 520 -16644 560
rect -17044 200 -17004 520
rect -16684 200 -16644 520
rect -17044 160 -16644 200
rect -16032 520 -15632 560
rect -16032 200 -15992 520
rect -15672 200 -15632 520
rect -16032 160 -15632 200
rect -15020 520 -14620 560
rect -15020 200 -14980 520
rect -14660 200 -14620 520
rect -15020 160 -14620 200
rect -14008 520 -13608 560
rect -14008 200 -13968 520
rect -13648 200 -13608 520
rect -14008 160 -13608 200
rect -12996 520 -12596 560
rect -12996 200 -12956 520
rect -12636 200 -12596 520
rect -12996 160 -12596 200
rect -11984 520 -11584 560
rect -11984 200 -11944 520
rect -11624 200 -11584 520
rect -11984 160 -11584 200
rect -10972 520 -10572 560
rect -10972 200 -10932 520
rect -10612 200 -10572 520
rect -10972 160 -10572 200
rect -9960 520 -9560 560
rect -9960 200 -9920 520
rect -9600 200 -9560 520
rect -9960 160 -9560 200
rect -8948 520 -8548 560
rect -8948 200 -8908 520
rect -8588 200 -8548 520
rect -8948 160 -8548 200
rect -7936 520 -7536 560
rect -7936 200 -7896 520
rect -7576 200 -7536 520
rect -7936 160 -7536 200
rect -6924 520 -6524 560
rect -6924 200 -6884 520
rect -6564 200 -6524 520
rect -6924 160 -6524 200
rect -5912 520 -5512 560
rect -5912 200 -5872 520
rect -5552 200 -5512 520
rect -5912 160 -5512 200
rect -4900 520 -4500 560
rect -4900 200 -4860 520
rect -4540 200 -4500 520
rect -4900 160 -4500 200
rect -3888 520 -3488 560
rect -3888 200 -3848 520
rect -3528 200 -3488 520
rect -3888 160 -3488 200
rect -2876 520 -2476 560
rect -2876 200 -2836 520
rect -2516 200 -2476 520
rect -2876 160 -2476 200
rect -1864 520 -1464 560
rect -1864 200 -1824 520
rect -1504 200 -1464 520
rect -1864 160 -1464 200
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect 1172 520 1572 560
rect 1172 200 1212 520
rect 1532 200 1572 520
rect 1172 160 1572 200
rect 2184 520 2584 560
rect 2184 200 2224 520
rect 2544 200 2584 520
rect 2184 160 2584 200
rect 3196 520 3596 560
rect 3196 200 3236 520
rect 3556 200 3596 520
rect 3196 160 3596 200
rect 4208 520 4608 560
rect 4208 200 4248 520
rect 4568 200 4608 520
rect 4208 160 4608 200
rect 5220 520 5620 560
rect 5220 200 5260 520
rect 5580 200 5620 520
rect 5220 160 5620 200
rect 6232 520 6632 560
rect 6232 200 6272 520
rect 6592 200 6632 520
rect 6232 160 6632 200
rect 7244 520 7644 560
rect 7244 200 7284 520
rect 7604 200 7644 520
rect 7244 160 7644 200
rect 8256 520 8656 560
rect 8256 200 8296 520
rect 8616 200 8656 520
rect 8256 160 8656 200
rect 9268 520 9668 560
rect 9268 200 9308 520
rect 9628 200 9668 520
rect 9268 160 9668 200
rect 10280 520 10680 560
rect 10280 200 10320 520
rect 10640 200 10680 520
rect 10280 160 10680 200
rect 11292 520 11692 560
rect 11292 200 11332 520
rect 11652 200 11692 520
rect 11292 160 11692 200
rect 12304 520 12704 560
rect 12304 200 12344 520
rect 12664 200 12704 520
rect 12304 160 12704 200
rect 13316 520 13716 560
rect 13316 200 13356 520
rect 13676 200 13716 520
rect 13316 160 13716 200
rect 14328 520 14728 560
rect 14328 200 14368 520
rect 14688 200 14728 520
rect 14328 160 14728 200
rect 15340 520 15740 560
rect 15340 200 15380 520
rect 15700 200 15740 520
rect 15340 160 15740 200
rect 16352 520 16752 560
rect 16352 200 16392 520
rect 16712 200 16752 520
rect 16352 160 16752 200
rect 17364 520 17764 560
rect 17364 200 17404 520
rect 17724 200 17764 520
rect 17364 160 17764 200
rect 18376 520 18776 560
rect 18376 200 18416 520
rect 18736 200 18776 520
rect 18376 160 18776 200
rect 19388 520 19788 560
rect 19388 200 19428 520
rect 19748 200 19788 520
rect 19388 160 19788 200
rect 20400 520 20800 560
rect 20400 200 20440 520
rect 20760 200 20800 520
rect 20400 160 20800 200
rect 21412 520 21812 560
rect 21412 200 21452 520
rect 21772 200 21812 520
rect 21412 160 21812 200
rect 22424 520 22824 560
rect 22424 200 22464 520
rect 22784 200 22824 520
rect 22424 160 22824 200
rect 23436 520 23836 560
rect 23436 200 23476 520
rect 23796 200 23836 520
rect 23436 160 23836 200
rect 24448 520 24848 560
rect 24448 200 24488 520
rect 24808 200 24848 520
rect 24448 160 24848 200
rect 25460 520 25860 560
rect 25460 200 25500 520
rect 25820 200 25860 520
rect 25460 160 25860 200
rect 26472 520 26872 560
rect 26472 200 26512 520
rect 26832 200 26872 520
rect 26472 160 26872 200
rect 27484 520 27884 560
rect 27484 200 27524 520
rect 27844 200 27884 520
rect 27484 160 27884 200
rect 28496 520 28896 560
rect 28496 200 28536 520
rect 28856 200 28896 520
rect 28496 160 28896 200
rect 29508 520 29908 560
rect 29508 200 29548 520
rect 29868 200 29908 520
rect 29508 160 29908 200
rect 30520 520 30920 560
rect 30520 200 30560 520
rect 30880 200 30920 520
rect 30520 160 30920 200
rect 31532 520 31932 560
rect 31532 200 31572 520
rect 31892 200 31932 520
rect 31532 160 31932 200
rect -32224 -200 -31824 -160
rect -32224 -520 -32184 -200
rect -31864 -520 -31824 -200
rect -32224 -560 -31824 -520
rect -31212 -200 -30812 -160
rect -31212 -520 -31172 -200
rect -30852 -520 -30812 -200
rect -31212 -560 -30812 -520
rect -30200 -200 -29800 -160
rect -30200 -520 -30160 -200
rect -29840 -520 -29800 -200
rect -30200 -560 -29800 -520
rect -29188 -200 -28788 -160
rect -29188 -520 -29148 -200
rect -28828 -520 -28788 -200
rect -29188 -560 -28788 -520
rect -28176 -200 -27776 -160
rect -28176 -520 -28136 -200
rect -27816 -520 -27776 -200
rect -28176 -560 -27776 -520
rect -27164 -200 -26764 -160
rect -27164 -520 -27124 -200
rect -26804 -520 -26764 -200
rect -27164 -560 -26764 -520
rect -26152 -200 -25752 -160
rect -26152 -520 -26112 -200
rect -25792 -520 -25752 -200
rect -26152 -560 -25752 -520
rect -25140 -200 -24740 -160
rect -25140 -520 -25100 -200
rect -24780 -520 -24740 -200
rect -25140 -560 -24740 -520
rect -24128 -200 -23728 -160
rect -24128 -520 -24088 -200
rect -23768 -520 -23728 -200
rect -24128 -560 -23728 -520
rect -23116 -200 -22716 -160
rect -23116 -520 -23076 -200
rect -22756 -520 -22716 -200
rect -23116 -560 -22716 -520
rect -22104 -200 -21704 -160
rect -22104 -520 -22064 -200
rect -21744 -520 -21704 -200
rect -22104 -560 -21704 -520
rect -21092 -200 -20692 -160
rect -21092 -520 -21052 -200
rect -20732 -520 -20692 -200
rect -21092 -560 -20692 -520
rect -20080 -200 -19680 -160
rect -20080 -520 -20040 -200
rect -19720 -520 -19680 -200
rect -20080 -560 -19680 -520
rect -19068 -200 -18668 -160
rect -19068 -520 -19028 -200
rect -18708 -520 -18668 -200
rect -19068 -560 -18668 -520
rect -18056 -200 -17656 -160
rect -18056 -520 -18016 -200
rect -17696 -520 -17656 -200
rect -18056 -560 -17656 -520
rect -17044 -200 -16644 -160
rect -17044 -520 -17004 -200
rect -16684 -520 -16644 -200
rect -17044 -560 -16644 -520
rect -16032 -200 -15632 -160
rect -16032 -520 -15992 -200
rect -15672 -520 -15632 -200
rect -16032 -560 -15632 -520
rect -15020 -200 -14620 -160
rect -15020 -520 -14980 -200
rect -14660 -520 -14620 -200
rect -15020 -560 -14620 -520
rect -14008 -200 -13608 -160
rect -14008 -520 -13968 -200
rect -13648 -520 -13608 -200
rect -14008 -560 -13608 -520
rect -12996 -200 -12596 -160
rect -12996 -520 -12956 -200
rect -12636 -520 -12596 -200
rect -12996 -560 -12596 -520
rect -11984 -200 -11584 -160
rect -11984 -520 -11944 -200
rect -11624 -520 -11584 -200
rect -11984 -560 -11584 -520
rect -10972 -200 -10572 -160
rect -10972 -520 -10932 -200
rect -10612 -520 -10572 -200
rect -10972 -560 -10572 -520
rect -9960 -200 -9560 -160
rect -9960 -520 -9920 -200
rect -9600 -520 -9560 -200
rect -9960 -560 -9560 -520
rect -8948 -200 -8548 -160
rect -8948 -520 -8908 -200
rect -8588 -520 -8548 -200
rect -8948 -560 -8548 -520
rect -7936 -200 -7536 -160
rect -7936 -520 -7896 -200
rect -7576 -520 -7536 -200
rect -7936 -560 -7536 -520
rect -6924 -200 -6524 -160
rect -6924 -520 -6884 -200
rect -6564 -520 -6524 -200
rect -6924 -560 -6524 -520
rect -5912 -200 -5512 -160
rect -5912 -520 -5872 -200
rect -5552 -520 -5512 -200
rect -5912 -560 -5512 -520
rect -4900 -200 -4500 -160
rect -4900 -520 -4860 -200
rect -4540 -520 -4500 -200
rect -4900 -560 -4500 -520
rect -3888 -200 -3488 -160
rect -3888 -520 -3848 -200
rect -3528 -520 -3488 -200
rect -3888 -560 -3488 -520
rect -2876 -200 -2476 -160
rect -2876 -520 -2836 -200
rect -2516 -520 -2476 -200
rect -2876 -560 -2476 -520
rect -1864 -200 -1464 -160
rect -1864 -520 -1824 -200
rect -1504 -520 -1464 -200
rect -1864 -560 -1464 -520
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect 1172 -200 1572 -160
rect 1172 -520 1212 -200
rect 1532 -520 1572 -200
rect 1172 -560 1572 -520
rect 2184 -200 2584 -160
rect 2184 -520 2224 -200
rect 2544 -520 2584 -200
rect 2184 -560 2584 -520
rect 3196 -200 3596 -160
rect 3196 -520 3236 -200
rect 3556 -520 3596 -200
rect 3196 -560 3596 -520
rect 4208 -200 4608 -160
rect 4208 -520 4248 -200
rect 4568 -520 4608 -200
rect 4208 -560 4608 -520
rect 5220 -200 5620 -160
rect 5220 -520 5260 -200
rect 5580 -520 5620 -200
rect 5220 -560 5620 -520
rect 6232 -200 6632 -160
rect 6232 -520 6272 -200
rect 6592 -520 6632 -200
rect 6232 -560 6632 -520
rect 7244 -200 7644 -160
rect 7244 -520 7284 -200
rect 7604 -520 7644 -200
rect 7244 -560 7644 -520
rect 8256 -200 8656 -160
rect 8256 -520 8296 -200
rect 8616 -520 8656 -200
rect 8256 -560 8656 -520
rect 9268 -200 9668 -160
rect 9268 -520 9308 -200
rect 9628 -520 9668 -200
rect 9268 -560 9668 -520
rect 10280 -200 10680 -160
rect 10280 -520 10320 -200
rect 10640 -520 10680 -200
rect 10280 -560 10680 -520
rect 11292 -200 11692 -160
rect 11292 -520 11332 -200
rect 11652 -520 11692 -200
rect 11292 -560 11692 -520
rect 12304 -200 12704 -160
rect 12304 -520 12344 -200
rect 12664 -520 12704 -200
rect 12304 -560 12704 -520
rect 13316 -200 13716 -160
rect 13316 -520 13356 -200
rect 13676 -520 13716 -200
rect 13316 -560 13716 -520
rect 14328 -200 14728 -160
rect 14328 -520 14368 -200
rect 14688 -520 14728 -200
rect 14328 -560 14728 -520
rect 15340 -200 15740 -160
rect 15340 -520 15380 -200
rect 15700 -520 15740 -200
rect 15340 -560 15740 -520
rect 16352 -200 16752 -160
rect 16352 -520 16392 -200
rect 16712 -520 16752 -200
rect 16352 -560 16752 -520
rect 17364 -200 17764 -160
rect 17364 -520 17404 -200
rect 17724 -520 17764 -200
rect 17364 -560 17764 -520
rect 18376 -200 18776 -160
rect 18376 -520 18416 -200
rect 18736 -520 18776 -200
rect 18376 -560 18776 -520
rect 19388 -200 19788 -160
rect 19388 -520 19428 -200
rect 19748 -520 19788 -200
rect 19388 -560 19788 -520
rect 20400 -200 20800 -160
rect 20400 -520 20440 -200
rect 20760 -520 20800 -200
rect 20400 -560 20800 -520
rect 21412 -200 21812 -160
rect 21412 -520 21452 -200
rect 21772 -520 21812 -200
rect 21412 -560 21812 -520
rect 22424 -200 22824 -160
rect 22424 -520 22464 -200
rect 22784 -520 22824 -200
rect 22424 -560 22824 -520
rect 23436 -200 23836 -160
rect 23436 -520 23476 -200
rect 23796 -520 23836 -200
rect 23436 -560 23836 -520
rect 24448 -200 24848 -160
rect 24448 -520 24488 -200
rect 24808 -520 24848 -200
rect 24448 -560 24848 -520
rect 25460 -200 25860 -160
rect 25460 -520 25500 -200
rect 25820 -520 25860 -200
rect 25460 -560 25860 -520
rect 26472 -200 26872 -160
rect 26472 -520 26512 -200
rect 26832 -520 26872 -200
rect 26472 -560 26872 -520
rect 27484 -200 27884 -160
rect 27484 -520 27524 -200
rect 27844 -520 27884 -200
rect 27484 -560 27884 -520
rect 28496 -200 28896 -160
rect 28496 -520 28536 -200
rect 28856 -520 28896 -200
rect 28496 -560 28896 -520
rect 29508 -200 29908 -160
rect 29508 -520 29548 -200
rect 29868 -520 29908 -200
rect 29508 -560 29908 -520
rect 30520 -200 30920 -160
rect 30520 -520 30560 -200
rect 30880 -520 30920 -200
rect 30520 -560 30920 -520
rect 31532 -200 31932 -160
rect 31532 -520 31572 -200
rect 31892 -520 31932 -200
rect 31532 -560 31932 -520
rect -32224 -920 -31824 -880
rect -32224 -1240 -32184 -920
rect -31864 -1240 -31824 -920
rect -32224 -1280 -31824 -1240
rect -31212 -920 -30812 -880
rect -31212 -1240 -31172 -920
rect -30852 -1240 -30812 -920
rect -31212 -1280 -30812 -1240
rect -30200 -920 -29800 -880
rect -30200 -1240 -30160 -920
rect -29840 -1240 -29800 -920
rect -30200 -1280 -29800 -1240
rect -29188 -920 -28788 -880
rect -29188 -1240 -29148 -920
rect -28828 -1240 -28788 -920
rect -29188 -1280 -28788 -1240
rect -28176 -920 -27776 -880
rect -28176 -1240 -28136 -920
rect -27816 -1240 -27776 -920
rect -28176 -1280 -27776 -1240
rect -27164 -920 -26764 -880
rect -27164 -1240 -27124 -920
rect -26804 -1240 -26764 -920
rect -27164 -1280 -26764 -1240
rect -26152 -920 -25752 -880
rect -26152 -1240 -26112 -920
rect -25792 -1240 -25752 -920
rect -26152 -1280 -25752 -1240
rect -25140 -920 -24740 -880
rect -25140 -1240 -25100 -920
rect -24780 -1240 -24740 -920
rect -25140 -1280 -24740 -1240
rect -24128 -920 -23728 -880
rect -24128 -1240 -24088 -920
rect -23768 -1240 -23728 -920
rect -24128 -1280 -23728 -1240
rect -23116 -920 -22716 -880
rect -23116 -1240 -23076 -920
rect -22756 -1240 -22716 -920
rect -23116 -1280 -22716 -1240
rect -22104 -920 -21704 -880
rect -22104 -1240 -22064 -920
rect -21744 -1240 -21704 -920
rect -22104 -1280 -21704 -1240
rect -21092 -920 -20692 -880
rect -21092 -1240 -21052 -920
rect -20732 -1240 -20692 -920
rect -21092 -1280 -20692 -1240
rect -20080 -920 -19680 -880
rect -20080 -1240 -20040 -920
rect -19720 -1240 -19680 -920
rect -20080 -1280 -19680 -1240
rect -19068 -920 -18668 -880
rect -19068 -1240 -19028 -920
rect -18708 -1240 -18668 -920
rect -19068 -1280 -18668 -1240
rect -18056 -920 -17656 -880
rect -18056 -1240 -18016 -920
rect -17696 -1240 -17656 -920
rect -18056 -1280 -17656 -1240
rect -17044 -920 -16644 -880
rect -17044 -1240 -17004 -920
rect -16684 -1240 -16644 -920
rect -17044 -1280 -16644 -1240
rect -16032 -920 -15632 -880
rect -16032 -1240 -15992 -920
rect -15672 -1240 -15632 -920
rect -16032 -1280 -15632 -1240
rect -15020 -920 -14620 -880
rect -15020 -1240 -14980 -920
rect -14660 -1240 -14620 -920
rect -15020 -1280 -14620 -1240
rect -14008 -920 -13608 -880
rect -14008 -1240 -13968 -920
rect -13648 -1240 -13608 -920
rect -14008 -1280 -13608 -1240
rect -12996 -920 -12596 -880
rect -12996 -1240 -12956 -920
rect -12636 -1240 -12596 -920
rect -12996 -1280 -12596 -1240
rect -11984 -920 -11584 -880
rect -11984 -1240 -11944 -920
rect -11624 -1240 -11584 -920
rect -11984 -1280 -11584 -1240
rect -10972 -920 -10572 -880
rect -10972 -1240 -10932 -920
rect -10612 -1240 -10572 -920
rect -10972 -1280 -10572 -1240
rect -9960 -920 -9560 -880
rect -9960 -1240 -9920 -920
rect -9600 -1240 -9560 -920
rect -9960 -1280 -9560 -1240
rect -8948 -920 -8548 -880
rect -8948 -1240 -8908 -920
rect -8588 -1240 -8548 -920
rect -8948 -1280 -8548 -1240
rect -7936 -920 -7536 -880
rect -7936 -1240 -7896 -920
rect -7576 -1240 -7536 -920
rect -7936 -1280 -7536 -1240
rect -6924 -920 -6524 -880
rect -6924 -1240 -6884 -920
rect -6564 -1240 -6524 -920
rect -6924 -1280 -6524 -1240
rect -5912 -920 -5512 -880
rect -5912 -1240 -5872 -920
rect -5552 -1240 -5512 -920
rect -5912 -1280 -5512 -1240
rect -4900 -920 -4500 -880
rect -4900 -1240 -4860 -920
rect -4540 -1240 -4500 -920
rect -4900 -1280 -4500 -1240
rect -3888 -920 -3488 -880
rect -3888 -1240 -3848 -920
rect -3528 -1240 -3488 -920
rect -3888 -1280 -3488 -1240
rect -2876 -920 -2476 -880
rect -2876 -1240 -2836 -920
rect -2516 -1240 -2476 -920
rect -2876 -1280 -2476 -1240
rect -1864 -920 -1464 -880
rect -1864 -1240 -1824 -920
rect -1504 -1240 -1464 -920
rect -1864 -1280 -1464 -1240
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect 1172 -920 1572 -880
rect 1172 -1240 1212 -920
rect 1532 -1240 1572 -920
rect 1172 -1280 1572 -1240
rect 2184 -920 2584 -880
rect 2184 -1240 2224 -920
rect 2544 -1240 2584 -920
rect 2184 -1280 2584 -1240
rect 3196 -920 3596 -880
rect 3196 -1240 3236 -920
rect 3556 -1240 3596 -920
rect 3196 -1280 3596 -1240
rect 4208 -920 4608 -880
rect 4208 -1240 4248 -920
rect 4568 -1240 4608 -920
rect 4208 -1280 4608 -1240
rect 5220 -920 5620 -880
rect 5220 -1240 5260 -920
rect 5580 -1240 5620 -920
rect 5220 -1280 5620 -1240
rect 6232 -920 6632 -880
rect 6232 -1240 6272 -920
rect 6592 -1240 6632 -920
rect 6232 -1280 6632 -1240
rect 7244 -920 7644 -880
rect 7244 -1240 7284 -920
rect 7604 -1240 7644 -920
rect 7244 -1280 7644 -1240
rect 8256 -920 8656 -880
rect 8256 -1240 8296 -920
rect 8616 -1240 8656 -920
rect 8256 -1280 8656 -1240
rect 9268 -920 9668 -880
rect 9268 -1240 9308 -920
rect 9628 -1240 9668 -920
rect 9268 -1280 9668 -1240
rect 10280 -920 10680 -880
rect 10280 -1240 10320 -920
rect 10640 -1240 10680 -920
rect 10280 -1280 10680 -1240
rect 11292 -920 11692 -880
rect 11292 -1240 11332 -920
rect 11652 -1240 11692 -920
rect 11292 -1280 11692 -1240
rect 12304 -920 12704 -880
rect 12304 -1240 12344 -920
rect 12664 -1240 12704 -920
rect 12304 -1280 12704 -1240
rect 13316 -920 13716 -880
rect 13316 -1240 13356 -920
rect 13676 -1240 13716 -920
rect 13316 -1280 13716 -1240
rect 14328 -920 14728 -880
rect 14328 -1240 14368 -920
rect 14688 -1240 14728 -920
rect 14328 -1280 14728 -1240
rect 15340 -920 15740 -880
rect 15340 -1240 15380 -920
rect 15700 -1240 15740 -920
rect 15340 -1280 15740 -1240
rect 16352 -920 16752 -880
rect 16352 -1240 16392 -920
rect 16712 -1240 16752 -920
rect 16352 -1280 16752 -1240
rect 17364 -920 17764 -880
rect 17364 -1240 17404 -920
rect 17724 -1240 17764 -920
rect 17364 -1280 17764 -1240
rect 18376 -920 18776 -880
rect 18376 -1240 18416 -920
rect 18736 -1240 18776 -920
rect 18376 -1280 18776 -1240
rect 19388 -920 19788 -880
rect 19388 -1240 19428 -920
rect 19748 -1240 19788 -920
rect 19388 -1280 19788 -1240
rect 20400 -920 20800 -880
rect 20400 -1240 20440 -920
rect 20760 -1240 20800 -920
rect 20400 -1280 20800 -1240
rect 21412 -920 21812 -880
rect 21412 -1240 21452 -920
rect 21772 -1240 21812 -920
rect 21412 -1280 21812 -1240
rect 22424 -920 22824 -880
rect 22424 -1240 22464 -920
rect 22784 -1240 22824 -920
rect 22424 -1280 22824 -1240
rect 23436 -920 23836 -880
rect 23436 -1240 23476 -920
rect 23796 -1240 23836 -920
rect 23436 -1280 23836 -1240
rect 24448 -920 24848 -880
rect 24448 -1240 24488 -920
rect 24808 -1240 24848 -920
rect 24448 -1280 24848 -1240
rect 25460 -920 25860 -880
rect 25460 -1240 25500 -920
rect 25820 -1240 25860 -920
rect 25460 -1280 25860 -1240
rect 26472 -920 26872 -880
rect 26472 -1240 26512 -920
rect 26832 -1240 26872 -920
rect 26472 -1280 26872 -1240
rect 27484 -920 27884 -880
rect 27484 -1240 27524 -920
rect 27844 -1240 27884 -920
rect 27484 -1280 27884 -1240
rect 28496 -920 28896 -880
rect 28496 -1240 28536 -920
rect 28856 -1240 28896 -920
rect 28496 -1280 28896 -1240
rect 29508 -920 29908 -880
rect 29508 -1240 29548 -920
rect 29868 -1240 29908 -920
rect 29508 -1280 29908 -1240
rect 30520 -920 30920 -880
rect 30520 -1240 30560 -920
rect 30880 -1240 30920 -920
rect 30520 -1280 30920 -1240
rect 31532 -920 31932 -880
rect 31532 -1240 31572 -920
rect 31892 -1240 31932 -920
rect 31532 -1280 31932 -1240
rect -32224 -1640 -31824 -1600
rect -32224 -1960 -32184 -1640
rect -31864 -1960 -31824 -1640
rect -32224 -2000 -31824 -1960
rect -31212 -1640 -30812 -1600
rect -31212 -1960 -31172 -1640
rect -30852 -1960 -30812 -1640
rect -31212 -2000 -30812 -1960
rect -30200 -1640 -29800 -1600
rect -30200 -1960 -30160 -1640
rect -29840 -1960 -29800 -1640
rect -30200 -2000 -29800 -1960
rect -29188 -1640 -28788 -1600
rect -29188 -1960 -29148 -1640
rect -28828 -1960 -28788 -1640
rect -29188 -2000 -28788 -1960
rect -28176 -1640 -27776 -1600
rect -28176 -1960 -28136 -1640
rect -27816 -1960 -27776 -1640
rect -28176 -2000 -27776 -1960
rect -27164 -1640 -26764 -1600
rect -27164 -1960 -27124 -1640
rect -26804 -1960 -26764 -1640
rect -27164 -2000 -26764 -1960
rect -26152 -1640 -25752 -1600
rect -26152 -1960 -26112 -1640
rect -25792 -1960 -25752 -1640
rect -26152 -2000 -25752 -1960
rect -25140 -1640 -24740 -1600
rect -25140 -1960 -25100 -1640
rect -24780 -1960 -24740 -1640
rect -25140 -2000 -24740 -1960
rect -24128 -1640 -23728 -1600
rect -24128 -1960 -24088 -1640
rect -23768 -1960 -23728 -1640
rect -24128 -2000 -23728 -1960
rect -23116 -1640 -22716 -1600
rect -23116 -1960 -23076 -1640
rect -22756 -1960 -22716 -1640
rect -23116 -2000 -22716 -1960
rect -22104 -1640 -21704 -1600
rect -22104 -1960 -22064 -1640
rect -21744 -1960 -21704 -1640
rect -22104 -2000 -21704 -1960
rect -21092 -1640 -20692 -1600
rect -21092 -1960 -21052 -1640
rect -20732 -1960 -20692 -1640
rect -21092 -2000 -20692 -1960
rect -20080 -1640 -19680 -1600
rect -20080 -1960 -20040 -1640
rect -19720 -1960 -19680 -1640
rect -20080 -2000 -19680 -1960
rect -19068 -1640 -18668 -1600
rect -19068 -1960 -19028 -1640
rect -18708 -1960 -18668 -1640
rect -19068 -2000 -18668 -1960
rect -18056 -1640 -17656 -1600
rect -18056 -1960 -18016 -1640
rect -17696 -1960 -17656 -1640
rect -18056 -2000 -17656 -1960
rect -17044 -1640 -16644 -1600
rect -17044 -1960 -17004 -1640
rect -16684 -1960 -16644 -1640
rect -17044 -2000 -16644 -1960
rect -16032 -1640 -15632 -1600
rect -16032 -1960 -15992 -1640
rect -15672 -1960 -15632 -1640
rect -16032 -2000 -15632 -1960
rect -15020 -1640 -14620 -1600
rect -15020 -1960 -14980 -1640
rect -14660 -1960 -14620 -1640
rect -15020 -2000 -14620 -1960
rect -14008 -1640 -13608 -1600
rect -14008 -1960 -13968 -1640
rect -13648 -1960 -13608 -1640
rect -14008 -2000 -13608 -1960
rect -12996 -1640 -12596 -1600
rect -12996 -1960 -12956 -1640
rect -12636 -1960 -12596 -1640
rect -12996 -2000 -12596 -1960
rect -11984 -1640 -11584 -1600
rect -11984 -1960 -11944 -1640
rect -11624 -1960 -11584 -1640
rect -11984 -2000 -11584 -1960
rect -10972 -1640 -10572 -1600
rect -10972 -1960 -10932 -1640
rect -10612 -1960 -10572 -1640
rect -10972 -2000 -10572 -1960
rect -9960 -1640 -9560 -1600
rect -9960 -1960 -9920 -1640
rect -9600 -1960 -9560 -1640
rect -9960 -2000 -9560 -1960
rect -8948 -1640 -8548 -1600
rect -8948 -1960 -8908 -1640
rect -8588 -1960 -8548 -1640
rect -8948 -2000 -8548 -1960
rect -7936 -1640 -7536 -1600
rect -7936 -1960 -7896 -1640
rect -7576 -1960 -7536 -1640
rect -7936 -2000 -7536 -1960
rect -6924 -1640 -6524 -1600
rect -6924 -1960 -6884 -1640
rect -6564 -1960 -6524 -1640
rect -6924 -2000 -6524 -1960
rect -5912 -1640 -5512 -1600
rect -5912 -1960 -5872 -1640
rect -5552 -1960 -5512 -1640
rect -5912 -2000 -5512 -1960
rect -4900 -1640 -4500 -1600
rect -4900 -1960 -4860 -1640
rect -4540 -1960 -4500 -1640
rect -4900 -2000 -4500 -1960
rect -3888 -1640 -3488 -1600
rect -3888 -1960 -3848 -1640
rect -3528 -1960 -3488 -1640
rect -3888 -2000 -3488 -1960
rect -2876 -1640 -2476 -1600
rect -2876 -1960 -2836 -1640
rect -2516 -1960 -2476 -1640
rect -2876 -2000 -2476 -1960
rect -1864 -1640 -1464 -1600
rect -1864 -1960 -1824 -1640
rect -1504 -1960 -1464 -1640
rect -1864 -2000 -1464 -1960
rect -852 -1640 -452 -1600
rect -852 -1960 -812 -1640
rect -492 -1960 -452 -1640
rect -852 -2000 -452 -1960
rect 160 -1640 560 -1600
rect 160 -1960 200 -1640
rect 520 -1960 560 -1640
rect 160 -2000 560 -1960
rect 1172 -1640 1572 -1600
rect 1172 -1960 1212 -1640
rect 1532 -1960 1572 -1640
rect 1172 -2000 1572 -1960
rect 2184 -1640 2584 -1600
rect 2184 -1960 2224 -1640
rect 2544 -1960 2584 -1640
rect 2184 -2000 2584 -1960
rect 3196 -1640 3596 -1600
rect 3196 -1960 3236 -1640
rect 3556 -1960 3596 -1640
rect 3196 -2000 3596 -1960
rect 4208 -1640 4608 -1600
rect 4208 -1960 4248 -1640
rect 4568 -1960 4608 -1640
rect 4208 -2000 4608 -1960
rect 5220 -1640 5620 -1600
rect 5220 -1960 5260 -1640
rect 5580 -1960 5620 -1640
rect 5220 -2000 5620 -1960
rect 6232 -1640 6632 -1600
rect 6232 -1960 6272 -1640
rect 6592 -1960 6632 -1640
rect 6232 -2000 6632 -1960
rect 7244 -1640 7644 -1600
rect 7244 -1960 7284 -1640
rect 7604 -1960 7644 -1640
rect 7244 -2000 7644 -1960
rect 8256 -1640 8656 -1600
rect 8256 -1960 8296 -1640
rect 8616 -1960 8656 -1640
rect 8256 -2000 8656 -1960
rect 9268 -1640 9668 -1600
rect 9268 -1960 9308 -1640
rect 9628 -1960 9668 -1640
rect 9268 -2000 9668 -1960
rect 10280 -1640 10680 -1600
rect 10280 -1960 10320 -1640
rect 10640 -1960 10680 -1640
rect 10280 -2000 10680 -1960
rect 11292 -1640 11692 -1600
rect 11292 -1960 11332 -1640
rect 11652 -1960 11692 -1640
rect 11292 -2000 11692 -1960
rect 12304 -1640 12704 -1600
rect 12304 -1960 12344 -1640
rect 12664 -1960 12704 -1640
rect 12304 -2000 12704 -1960
rect 13316 -1640 13716 -1600
rect 13316 -1960 13356 -1640
rect 13676 -1960 13716 -1640
rect 13316 -2000 13716 -1960
rect 14328 -1640 14728 -1600
rect 14328 -1960 14368 -1640
rect 14688 -1960 14728 -1640
rect 14328 -2000 14728 -1960
rect 15340 -1640 15740 -1600
rect 15340 -1960 15380 -1640
rect 15700 -1960 15740 -1640
rect 15340 -2000 15740 -1960
rect 16352 -1640 16752 -1600
rect 16352 -1960 16392 -1640
rect 16712 -1960 16752 -1640
rect 16352 -2000 16752 -1960
rect 17364 -1640 17764 -1600
rect 17364 -1960 17404 -1640
rect 17724 -1960 17764 -1640
rect 17364 -2000 17764 -1960
rect 18376 -1640 18776 -1600
rect 18376 -1960 18416 -1640
rect 18736 -1960 18776 -1640
rect 18376 -2000 18776 -1960
rect 19388 -1640 19788 -1600
rect 19388 -1960 19428 -1640
rect 19748 -1960 19788 -1640
rect 19388 -2000 19788 -1960
rect 20400 -1640 20800 -1600
rect 20400 -1960 20440 -1640
rect 20760 -1960 20800 -1640
rect 20400 -2000 20800 -1960
rect 21412 -1640 21812 -1600
rect 21412 -1960 21452 -1640
rect 21772 -1960 21812 -1640
rect 21412 -2000 21812 -1960
rect 22424 -1640 22824 -1600
rect 22424 -1960 22464 -1640
rect 22784 -1960 22824 -1640
rect 22424 -2000 22824 -1960
rect 23436 -1640 23836 -1600
rect 23436 -1960 23476 -1640
rect 23796 -1960 23836 -1640
rect 23436 -2000 23836 -1960
rect 24448 -1640 24848 -1600
rect 24448 -1960 24488 -1640
rect 24808 -1960 24848 -1640
rect 24448 -2000 24848 -1960
rect 25460 -1640 25860 -1600
rect 25460 -1960 25500 -1640
rect 25820 -1960 25860 -1640
rect 25460 -2000 25860 -1960
rect 26472 -1640 26872 -1600
rect 26472 -1960 26512 -1640
rect 26832 -1960 26872 -1640
rect 26472 -2000 26872 -1960
rect 27484 -1640 27884 -1600
rect 27484 -1960 27524 -1640
rect 27844 -1960 27884 -1640
rect 27484 -2000 27884 -1960
rect 28496 -1640 28896 -1600
rect 28496 -1960 28536 -1640
rect 28856 -1960 28896 -1640
rect 28496 -2000 28896 -1960
rect 29508 -1640 29908 -1600
rect 29508 -1960 29548 -1640
rect 29868 -1960 29908 -1640
rect 29508 -2000 29908 -1960
rect 30520 -1640 30920 -1600
rect 30520 -1960 30560 -1640
rect 30880 -1960 30920 -1640
rect 30520 -2000 30920 -1960
rect 31532 -1640 31932 -1600
rect 31532 -1960 31572 -1640
rect 31892 -1960 31932 -1640
rect 31532 -2000 31932 -1960
rect -32224 -2360 -31824 -2320
rect -32224 -2680 -32184 -2360
rect -31864 -2680 -31824 -2360
rect -32224 -2720 -31824 -2680
rect -31212 -2360 -30812 -2320
rect -31212 -2680 -31172 -2360
rect -30852 -2680 -30812 -2360
rect -31212 -2720 -30812 -2680
rect -30200 -2360 -29800 -2320
rect -30200 -2680 -30160 -2360
rect -29840 -2680 -29800 -2360
rect -30200 -2720 -29800 -2680
rect -29188 -2360 -28788 -2320
rect -29188 -2680 -29148 -2360
rect -28828 -2680 -28788 -2360
rect -29188 -2720 -28788 -2680
rect -28176 -2360 -27776 -2320
rect -28176 -2680 -28136 -2360
rect -27816 -2680 -27776 -2360
rect -28176 -2720 -27776 -2680
rect -27164 -2360 -26764 -2320
rect -27164 -2680 -27124 -2360
rect -26804 -2680 -26764 -2360
rect -27164 -2720 -26764 -2680
rect -26152 -2360 -25752 -2320
rect -26152 -2680 -26112 -2360
rect -25792 -2680 -25752 -2360
rect -26152 -2720 -25752 -2680
rect -25140 -2360 -24740 -2320
rect -25140 -2680 -25100 -2360
rect -24780 -2680 -24740 -2360
rect -25140 -2720 -24740 -2680
rect -24128 -2360 -23728 -2320
rect -24128 -2680 -24088 -2360
rect -23768 -2680 -23728 -2360
rect -24128 -2720 -23728 -2680
rect -23116 -2360 -22716 -2320
rect -23116 -2680 -23076 -2360
rect -22756 -2680 -22716 -2360
rect -23116 -2720 -22716 -2680
rect -22104 -2360 -21704 -2320
rect -22104 -2680 -22064 -2360
rect -21744 -2680 -21704 -2360
rect -22104 -2720 -21704 -2680
rect -21092 -2360 -20692 -2320
rect -21092 -2680 -21052 -2360
rect -20732 -2680 -20692 -2360
rect -21092 -2720 -20692 -2680
rect -20080 -2360 -19680 -2320
rect -20080 -2680 -20040 -2360
rect -19720 -2680 -19680 -2360
rect -20080 -2720 -19680 -2680
rect -19068 -2360 -18668 -2320
rect -19068 -2680 -19028 -2360
rect -18708 -2680 -18668 -2360
rect -19068 -2720 -18668 -2680
rect -18056 -2360 -17656 -2320
rect -18056 -2680 -18016 -2360
rect -17696 -2680 -17656 -2360
rect -18056 -2720 -17656 -2680
rect -17044 -2360 -16644 -2320
rect -17044 -2680 -17004 -2360
rect -16684 -2680 -16644 -2360
rect -17044 -2720 -16644 -2680
rect -16032 -2360 -15632 -2320
rect -16032 -2680 -15992 -2360
rect -15672 -2680 -15632 -2360
rect -16032 -2720 -15632 -2680
rect -15020 -2360 -14620 -2320
rect -15020 -2680 -14980 -2360
rect -14660 -2680 -14620 -2360
rect -15020 -2720 -14620 -2680
rect -14008 -2360 -13608 -2320
rect -14008 -2680 -13968 -2360
rect -13648 -2680 -13608 -2360
rect -14008 -2720 -13608 -2680
rect -12996 -2360 -12596 -2320
rect -12996 -2680 -12956 -2360
rect -12636 -2680 -12596 -2360
rect -12996 -2720 -12596 -2680
rect -11984 -2360 -11584 -2320
rect -11984 -2680 -11944 -2360
rect -11624 -2680 -11584 -2360
rect -11984 -2720 -11584 -2680
rect -10972 -2360 -10572 -2320
rect -10972 -2680 -10932 -2360
rect -10612 -2680 -10572 -2360
rect -10972 -2720 -10572 -2680
rect -9960 -2360 -9560 -2320
rect -9960 -2680 -9920 -2360
rect -9600 -2680 -9560 -2360
rect -9960 -2720 -9560 -2680
rect -8948 -2360 -8548 -2320
rect -8948 -2680 -8908 -2360
rect -8588 -2680 -8548 -2360
rect -8948 -2720 -8548 -2680
rect -7936 -2360 -7536 -2320
rect -7936 -2680 -7896 -2360
rect -7576 -2680 -7536 -2360
rect -7936 -2720 -7536 -2680
rect -6924 -2360 -6524 -2320
rect -6924 -2680 -6884 -2360
rect -6564 -2680 -6524 -2360
rect -6924 -2720 -6524 -2680
rect -5912 -2360 -5512 -2320
rect -5912 -2680 -5872 -2360
rect -5552 -2680 -5512 -2360
rect -5912 -2720 -5512 -2680
rect -4900 -2360 -4500 -2320
rect -4900 -2680 -4860 -2360
rect -4540 -2680 -4500 -2360
rect -4900 -2720 -4500 -2680
rect -3888 -2360 -3488 -2320
rect -3888 -2680 -3848 -2360
rect -3528 -2680 -3488 -2360
rect -3888 -2720 -3488 -2680
rect -2876 -2360 -2476 -2320
rect -2876 -2680 -2836 -2360
rect -2516 -2680 -2476 -2360
rect -2876 -2720 -2476 -2680
rect -1864 -2360 -1464 -2320
rect -1864 -2680 -1824 -2360
rect -1504 -2680 -1464 -2360
rect -1864 -2720 -1464 -2680
rect -852 -2360 -452 -2320
rect -852 -2680 -812 -2360
rect -492 -2680 -452 -2360
rect -852 -2720 -452 -2680
rect 160 -2360 560 -2320
rect 160 -2680 200 -2360
rect 520 -2680 560 -2360
rect 160 -2720 560 -2680
rect 1172 -2360 1572 -2320
rect 1172 -2680 1212 -2360
rect 1532 -2680 1572 -2360
rect 1172 -2720 1572 -2680
rect 2184 -2360 2584 -2320
rect 2184 -2680 2224 -2360
rect 2544 -2680 2584 -2360
rect 2184 -2720 2584 -2680
rect 3196 -2360 3596 -2320
rect 3196 -2680 3236 -2360
rect 3556 -2680 3596 -2360
rect 3196 -2720 3596 -2680
rect 4208 -2360 4608 -2320
rect 4208 -2680 4248 -2360
rect 4568 -2680 4608 -2360
rect 4208 -2720 4608 -2680
rect 5220 -2360 5620 -2320
rect 5220 -2680 5260 -2360
rect 5580 -2680 5620 -2360
rect 5220 -2720 5620 -2680
rect 6232 -2360 6632 -2320
rect 6232 -2680 6272 -2360
rect 6592 -2680 6632 -2360
rect 6232 -2720 6632 -2680
rect 7244 -2360 7644 -2320
rect 7244 -2680 7284 -2360
rect 7604 -2680 7644 -2360
rect 7244 -2720 7644 -2680
rect 8256 -2360 8656 -2320
rect 8256 -2680 8296 -2360
rect 8616 -2680 8656 -2360
rect 8256 -2720 8656 -2680
rect 9268 -2360 9668 -2320
rect 9268 -2680 9308 -2360
rect 9628 -2680 9668 -2360
rect 9268 -2720 9668 -2680
rect 10280 -2360 10680 -2320
rect 10280 -2680 10320 -2360
rect 10640 -2680 10680 -2360
rect 10280 -2720 10680 -2680
rect 11292 -2360 11692 -2320
rect 11292 -2680 11332 -2360
rect 11652 -2680 11692 -2360
rect 11292 -2720 11692 -2680
rect 12304 -2360 12704 -2320
rect 12304 -2680 12344 -2360
rect 12664 -2680 12704 -2360
rect 12304 -2720 12704 -2680
rect 13316 -2360 13716 -2320
rect 13316 -2680 13356 -2360
rect 13676 -2680 13716 -2360
rect 13316 -2720 13716 -2680
rect 14328 -2360 14728 -2320
rect 14328 -2680 14368 -2360
rect 14688 -2680 14728 -2360
rect 14328 -2720 14728 -2680
rect 15340 -2360 15740 -2320
rect 15340 -2680 15380 -2360
rect 15700 -2680 15740 -2360
rect 15340 -2720 15740 -2680
rect 16352 -2360 16752 -2320
rect 16352 -2680 16392 -2360
rect 16712 -2680 16752 -2360
rect 16352 -2720 16752 -2680
rect 17364 -2360 17764 -2320
rect 17364 -2680 17404 -2360
rect 17724 -2680 17764 -2360
rect 17364 -2720 17764 -2680
rect 18376 -2360 18776 -2320
rect 18376 -2680 18416 -2360
rect 18736 -2680 18776 -2360
rect 18376 -2720 18776 -2680
rect 19388 -2360 19788 -2320
rect 19388 -2680 19428 -2360
rect 19748 -2680 19788 -2360
rect 19388 -2720 19788 -2680
rect 20400 -2360 20800 -2320
rect 20400 -2680 20440 -2360
rect 20760 -2680 20800 -2360
rect 20400 -2720 20800 -2680
rect 21412 -2360 21812 -2320
rect 21412 -2680 21452 -2360
rect 21772 -2680 21812 -2360
rect 21412 -2720 21812 -2680
rect 22424 -2360 22824 -2320
rect 22424 -2680 22464 -2360
rect 22784 -2680 22824 -2360
rect 22424 -2720 22824 -2680
rect 23436 -2360 23836 -2320
rect 23436 -2680 23476 -2360
rect 23796 -2680 23836 -2360
rect 23436 -2720 23836 -2680
rect 24448 -2360 24848 -2320
rect 24448 -2680 24488 -2360
rect 24808 -2680 24848 -2360
rect 24448 -2720 24848 -2680
rect 25460 -2360 25860 -2320
rect 25460 -2680 25500 -2360
rect 25820 -2680 25860 -2360
rect 25460 -2720 25860 -2680
rect 26472 -2360 26872 -2320
rect 26472 -2680 26512 -2360
rect 26832 -2680 26872 -2360
rect 26472 -2720 26872 -2680
rect 27484 -2360 27884 -2320
rect 27484 -2680 27524 -2360
rect 27844 -2680 27884 -2360
rect 27484 -2720 27884 -2680
rect 28496 -2360 28896 -2320
rect 28496 -2680 28536 -2360
rect 28856 -2680 28896 -2360
rect 28496 -2720 28896 -2680
rect 29508 -2360 29908 -2320
rect 29508 -2680 29548 -2360
rect 29868 -2680 29908 -2360
rect 29508 -2720 29908 -2680
rect 30520 -2360 30920 -2320
rect 30520 -2680 30560 -2360
rect 30880 -2680 30920 -2360
rect 30520 -2720 30920 -2680
rect 31532 -2360 31932 -2320
rect 31532 -2680 31572 -2360
rect 31892 -2680 31932 -2360
rect 31532 -2720 31932 -2680
rect -32224 -3080 -31824 -3040
rect -32224 -3400 -32184 -3080
rect -31864 -3400 -31824 -3080
rect -32224 -3440 -31824 -3400
rect -31212 -3080 -30812 -3040
rect -31212 -3400 -31172 -3080
rect -30852 -3400 -30812 -3080
rect -31212 -3440 -30812 -3400
rect -30200 -3080 -29800 -3040
rect -30200 -3400 -30160 -3080
rect -29840 -3400 -29800 -3080
rect -30200 -3440 -29800 -3400
rect -29188 -3080 -28788 -3040
rect -29188 -3400 -29148 -3080
rect -28828 -3400 -28788 -3080
rect -29188 -3440 -28788 -3400
rect -28176 -3080 -27776 -3040
rect -28176 -3400 -28136 -3080
rect -27816 -3400 -27776 -3080
rect -28176 -3440 -27776 -3400
rect -27164 -3080 -26764 -3040
rect -27164 -3400 -27124 -3080
rect -26804 -3400 -26764 -3080
rect -27164 -3440 -26764 -3400
rect -26152 -3080 -25752 -3040
rect -26152 -3400 -26112 -3080
rect -25792 -3400 -25752 -3080
rect -26152 -3440 -25752 -3400
rect -25140 -3080 -24740 -3040
rect -25140 -3400 -25100 -3080
rect -24780 -3400 -24740 -3080
rect -25140 -3440 -24740 -3400
rect -24128 -3080 -23728 -3040
rect -24128 -3400 -24088 -3080
rect -23768 -3400 -23728 -3080
rect -24128 -3440 -23728 -3400
rect -23116 -3080 -22716 -3040
rect -23116 -3400 -23076 -3080
rect -22756 -3400 -22716 -3080
rect -23116 -3440 -22716 -3400
rect -22104 -3080 -21704 -3040
rect -22104 -3400 -22064 -3080
rect -21744 -3400 -21704 -3080
rect -22104 -3440 -21704 -3400
rect -21092 -3080 -20692 -3040
rect -21092 -3400 -21052 -3080
rect -20732 -3400 -20692 -3080
rect -21092 -3440 -20692 -3400
rect -20080 -3080 -19680 -3040
rect -20080 -3400 -20040 -3080
rect -19720 -3400 -19680 -3080
rect -20080 -3440 -19680 -3400
rect -19068 -3080 -18668 -3040
rect -19068 -3400 -19028 -3080
rect -18708 -3400 -18668 -3080
rect -19068 -3440 -18668 -3400
rect -18056 -3080 -17656 -3040
rect -18056 -3400 -18016 -3080
rect -17696 -3400 -17656 -3080
rect -18056 -3440 -17656 -3400
rect -17044 -3080 -16644 -3040
rect -17044 -3400 -17004 -3080
rect -16684 -3400 -16644 -3080
rect -17044 -3440 -16644 -3400
rect -16032 -3080 -15632 -3040
rect -16032 -3400 -15992 -3080
rect -15672 -3400 -15632 -3080
rect -16032 -3440 -15632 -3400
rect -15020 -3080 -14620 -3040
rect -15020 -3400 -14980 -3080
rect -14660 -3400 -14620 -3080
rect -15020 -3440 -14620 -3400
rect -14008 -3080 -13608 -3040
rect -14008 -3400 -13968 -3080
rect -13648 -3400 -13608 -3080
rect -14008 -3440 -13608 -3400
rect -12996 -3080 -12596 -3040
rect -12996 -3400 -12956 -3080
rect -12636 -3400 -12596 -3080
rect -12996 -3440 -12596 -3400
rect -11984 -3080 -11584 -3040
rect -11984 -3400 -11944 -3080
rect -11624 -3400 -11584 -3080
rect -11984 -3440 -11584 -3400
rect -10972 -3080 -10572 -3040
rect -10972 -3400 -10932 -3080
rect -10612 -3400 -10572 -3080
rect -10972 -3440 -10572 -3400
rect -9960 -3080 -9560 -3040
rect -9960 -3400 -9920 -3080
rect -9600 -3400 -9560 -3080
rect -9960 -3440 -9560 -3400
rect -8948 -3080 -8548 -3040
rect -8948 -3400 -8908 -3080
rect -8588 -3400 -8548 -3080
rect -8948 -3440 -8548 -3400
rect -7936 -3080 -7536 -3040
rect -7936 -3400 -7896 -3080
rect -7576 -3400 -7536 -3080
rect -7936 -3440 -7536 -3400
rect -6924 -3080 -6524 -3040
rect -6924 -3400 -6884 -3080
rect -6564 -3400 -6524 -3080
rect -6924 -3440 -6524 -3400
rect -5912 -3080 -5512 -3040
rect -5912 -3400 -5872 -3080
rect -5552 -3400 -5512 -3080
rect -5912 -3440 -5512 -3400
rect -4900 -3080 -4500 -3040
rect -4900 -3400 -4860 -3080
rect -4540 -3400 -4500 -3080
rect -4900 -3440 -4500 -3400
rect -3888 -3080 -3488 -3040
rect -3888 -3400 -3848 -3080
rect -3528 -3400 -3488 -3080
rect -3888 -3440 -3488 -3400
rect -2876 -3080 -2476 -3040
rect -2876 -3400 -2836 -3080
rect -2516 -3400 -2476 -3080
rect -2876 -3440 -2476 -3400
rect -1864 -3080 -1464 -3040
rect -1864 -3400 -1824 -3080
rect -1504 -3400 -1464 -3080
rect -1864 -3440 -1464 -3400
rect -852 -3080 -452 -3040
rect -852 -3400 -812 -3080
rect -492 -3400 -452 -3080
rect -852 -3440 -452 -3400
rect 160 -3080 560 -3040
rect 160 -3400 200 -3080
rect 520 -3400 560 -3080
rect 160 -3440 560 -3400
rect 1172 -3080 1572 -3040
rect 1172 -3400 1212 -3080
rect 1532 -3400 1572 -3080
rect 1172 -3440 1572 -3400
rect 2184 -3080 2584 -3040
rect 2184 -3400 2224 -3080
rect 2544 -3400 2584 -3080
rect 2184 -3440 2584 -3400
rect 3196 -3080 3596 -3040
rect 3196 -3400 3236 -3080
rect 3556 -3400 3596 -3080
rect 3196 -3440 3596 -3400
rect 4208 -3080 4608 -3040
rect 4208 -3400 4248 -3080
rect 4568 -3400 4608 -3080
rect 4208 -3440 4608 -3400
rect 5220 -3080 5620 -3040
rect 5220 -3400 5260 -3080
rect 5580 -3400 5620 -3080
rect 5220 -3440 5620 -3400
rect 6232 -3080 6632 -3040
rect 6232 -3400 6272 -3080
rect 6592 -3400 6632 -3080
rect 6232 -3440 6632 -3400
rect 7244 -3080 7644 -3040
rect 7244 -3400 7284 -3080
rect 7604 -3400 7644 -3080
rect 7244 -3440 7644 -3400
rect 8256 -3080 8656 -3040
rect 8256 -3400 8296 -3080
rect 8616 -3400 8656 -3080
rect 8256 -3440 8656 -3400
rect 9268 -3080 9668 -3040
rect 9268 -3400 9308 -3080
rect 9628 -3400 9668 -3080
rect 9268 -3440 9668 -3400
rect 10280 -3080 10680 -3040
rect 10280 -3400 10320 -3080
rect 10640 -3400 10680 -3080
rect 10280 -3440 10680 -3400
rect 11292 -3080 11692 -3040
rect 11292 -3400 11332 -3080
rect 11652 -3400 11692 -3080
rect 11292 -3440 11692 -3400
rect 12304 -3080 12704 -3040
rect 12304 -3400 12344 -3080
rect 12664 -3400 12704 -3080
rect 12304 -3440 12704 -3400
rect 13316 -3080 13716 -3040
rect 13316 -3400 13356 -3080
rect 13676 -3400 13716 -3080
rect 13316 -3440 13716 -3400
rect 14328 -3080 14728 -3040
rect 14328 -3400 14368 -3080
rect 14688 -3400 14728 -3080
rect 14328 -3440 14728 -3400
rect 15340 -3080 15740 -3040
rect 15340 -3400 15380 -3080
rect 15700 -3400 15740 -3080
rect 15340 -3440 15740 -3400
rect 16352 -3080 16752 -3040
rect 16352 -3400 16392 -3080
rect 16712 -3400 16752 -3080
rect 16352 -3440 16752 -3400
rect 17364 -3080 17764 -3040
rect 17364 -3400 17404 -3080
rect 17724 -3400 17764 -3080
rect 17364 -3440 17764 -3400
rect 18376 -3080 18776 -3040
rect 18376 -3400 18416 -3080
rect 18736 -3400 18776 -3080
rect 18376 -3440 18776 -3400
rect 19388 -3080 19788 -3040
rect 19388 -3400 19428 -3080
rect 19748 -3400 19788 -3080
rect 19388 -3440 19788 -3400
rect 20400 -3080 20800 -3040
rect 20400 -3400 20440 -3080
rect 20760 -3400 20800 -3080
rect 20400 -3440 20800 -3400
rect 21412 -3080 21812 -3040
rect 21412 -3400 21452 -3080
rect 21772 -3400 21812 -3080
rect 21412 -3440 21812 -3400
rect 22424 -3080 22824 -3040
rect 22424 -3400 22464 -3080
rect 22784 -3400 22824 -3080
rect 22424 -3440 22824 -3400
rect 23436 -3080 23836 -3040
rect 23436 -3400 23476 -3080
rect 23796 -3400 23836 -3080
rect 23436 -3440 23836 -3400
rect 24448 -3080 24848 -3040
rect 24448 -3400 24488 -3080
rect 24808 -3400 24848 -3080
rect 24448 -3440 24848 -3400
rect 25460 -3080 25860 -3040
rect 25460 -3400 25500 -3080
rect 25820 -3400 25860 -3080
rect 25460 -3440 25860 -3400
rect 26472 -3080 26872 -3040
rect 26472 -3400 26512 -3080
rect 26832 -3400 26872 -3080
rect 26472 -3440 26872 -3400
rect 27484 -3080 27884 -3040
rect 27484 -3400 27524 -3080
rect 27844 -3400 27884 -3080
rect 27484 -3440 27884 -3400
rect 28496 -3080 28896 -3040
rect 28496 -3400 28536 -3080
rect 28856 -3400 28896 -3080
rect 28496 -3440 28896 -3400
rect 29508 -3080 29908 -3040
rect 29508 -3400 29548 -3080
rect 29868 -3400 29908 -3080
rect 29508 -3440 29908 -3400
rect 30520 -3080 30920 -3040
rect 30520 -3400 30560 -3080
rect 30880 -3400 30920 -3080
rect 30520 -3440 30920 -3400
rect 31532 -3080 31932 -3040
rect 31532 -3400 31572 -3080
rect 31892 -3400 31932 -3080
rect 31532 -3440 31932 -3400
rect -32224 -3800 -31824 -3760
rect -32224 -4120 -32184 -3800
rect -31864 -4120 -31824 -3800
rect -32224 -4160 -31824 -4120
rect -31212 -3800 -30812 -3760
rect -31212 -4120 -31172 -3800
rect -30852 -4120 -30812 -3800
rect -31212 -4160 -30812 -4120
rect -30200 -3800 -29800 -3760
rect -30200 -4120 -30160 -3800
rect -29840 -4120 -29800 -3800
rect -30200 -4160 -29800 -4120
rect -29188 -3800 -28788 -3760
rect -29188 -4120 -29148 -3800
rect -28828 -4120 -28788 -3800
rect -29188 -4160 -28788 -4120
rect -28176 -3800 -27776 -3760
rect -28176 -4120 -28136 -3800
rect -27816 -4120 -27776 -3800
rect -28176 -4160 -27776 -4120
rect -27164 -3800 -26764 -3760
rect -27164 -4120 -27124 -3800
rect -26804 -4120 -26764 -3800
rect -27164 -4160 -26764 -4120
rect -26152 -3800 -25752 -3760
rect -26152 -4120 -26112 -3800
rect -25792 -4120 -25752 -3800
rect -26152 -4160 -25752 -4120
rect -25140 -3800 -24740 -3760
rect -25140 -4120 -25100 -3800
rect -24780 -4120 -24740 -3800
rect -25140 -4160 -24740 -4120
rect -24128 -3800 -23728 -3760
rect -24128 -4120 -24088 -3800
rect -23768 -4120 -23728 -3800
rect -24128 -4160 -23728 -4120
rect -23116 -3800 -22716 -3760
rect -23116 -4120 -23076 -3800
rect -22756 -4120 -22716 -3800
rect -23116 -4160 -22716 -4120
rect -22104 -3800 -21704 -3760
rect -22104 -4120 -22064 -3800
rect -21744 -4120 -21704 -3800
rect -22104 -4160 -21704 -4120
rect -21092 -3800 -20692 -3760
rect -21092 -4120 -21052 -3800
rect -20732 -4120 -20692 -3800
rect -21092 -4160 -20692 -4120
rect -20080 -3800 -19680 -3760
rect -20080 -4120 -20040 -3800
rect -19720 -4120 -19680 -3800
rect -20080 -4160 -19680 -4120
rect -19068 -3800 -18668 -3760
rect -19068 -4120 -19028 -3800
rect -18708 -4120 -18668 -3800
rect -19068 -4160 -18668 -4120
rect -18056 -3800 -17656 -3760
rect -18056 -4120 -18016 -3800
rect -17696 -4120 -17656 -3800
rect -18056 -4160 -17656 -4120
rect -17044 -3800 -16644 -3760
rect -17044 -4120 -17004 -3800
rect -16684 -4120 -16644 -3800
rect -17044 -4160 -16644 -4120
rect -16032 -3800 -15632 -3760
rect -16032 -4120 -15992 -3800
rect -15672 -4120 -15632 -3800
rect -16032 -4160 -15632 -4120
rect -15020 -3800 -14620 -3760
rect -15020 -4120 -14980 -3800
rect -14660 -4120 -14620 -3800
rect -15020 -4160 -14620 -4120
rect -14008 -3800 -13608 -3760
rect -14008 -4120 -13968 -3800
rect -13648 -4120 -13608 -3800
rect -14008 -4160 -13608 -4120
rect -12996 -3800 -12596 -3760
rect -12996 -4120 -12956 -3800
rect -12636 -4120 -12596 -3800
rect -12996 -4160 -12596 -4120
rect -11984 -3800 -11584 -3760
rect -11984 -4120 -11944 -3800
rect -11624 -4120 -11584 -3800
rect -11984 -4160 -11584 -4120
rect -10972 -3800 -10572 -3760
rect -10972 -4120 -10932 -3800
rect -10612 -4120 -10572 -3800
rect -10972 -4160 -10572 -4120
rect -9960 -3800 -9560 -3760
rect -9960 -4120 -9920 -3800
rect -9600 -4120 -9560 -3800
rect -9960 -4160 -9560 -4120
rect -8948 -3800 -8548 -3760
rect -8948 -4120 -8908 -3800
rect -8588 -4120 -8548 -3800
rect -8948 -4160 -8548 -4120
rect -7936 -3800 -7536 -3760
rect -7936 -4120 -7896 -3800
rect -7576 -4120 -7536 -3800
rect -7936 -4160 -7536 -4120
rect -6924 -3800 -6524 -3760
rect -6924 -4120 -6884 -3800
rect -6564 -4120 -6524 -3800
rect -6924 -4160 -6524 -4120
rect -5912 -3800 -5512 -3760
rect -5912 -4120 -5872 -3800
rect -5552 -4120 -5512 -3800
rect -5912 -4160 -5512 -4120
rect -4900 -3800 -4500 -3760
rect -4900 -4120 -4860 -3800
rect -4540 -4120 -4500 -3800
rect -4900 -4160 -4500 -4120
rect -3888 -3800 -3488 -3760
rect -3888 -4120 -3848 -3800
rect -3528 -4120 -3488 -3800
rect -3888 -4160 -3488 -4120
rect -2876 -3800 -2476 -3760
rect -2876 -4120 -2836 -3800
rect -2516 -4120 -2476 -3800
rect -2876 -4160 -2476 -4120
rect -1864 -3800 -1464 -3760
rect -1864 -4120 -1824 -3800
rect -1504 -4120 -1464 -3800
rect -1864 -4160 -1464 -4120
rect -852 -3800 -452 -3760
rect -852 -4120 -812 -3800
rect -492 -4120 -452 -3800
rect -852 -4160 -452 -4120
rect 160 -3800 560 -3760
rect 160 -4120 200 -3800
rect 520 -4120 560 -3800
rect 160 -4160 560 -4120
rect 1172 -3800 1572 -3760
rect 1172 -4120 1212 -3800
rect 1532 -4120 1572 -3800
rect 1172 -4160 1572 -4120
rect 2184 -3800 2584 -3760
rect 2184 -4120 2224 -3800
rect 2544 -4120 2584 -3800
rect 2184 -4160 2584 -4120
rect 3196 -3800 3596 -3760
rect 3196 -4120 3236 -3800
rect 3556 -4120 3596 -3800
rect 3196 -4160 3596 -4120
rect 4208 -3800 4608 -3760
rect 4208 -4120 4248 -3800
rect 4568 -4120 4608 -3800
rect 4208 -4160 4608 -4120
rect 5220 -3800 5620 -3760
rect 5220 -4120 5260 -3800
rect 5580 -4120 5620 -3800
rect 5220 -4160 5620 -4120
rect 6232 -3800 6632 -3760
rect 6232 -4120 6272 -3800
rect 6592 -4120 6632 -3800
rect 6232 -4160 6632 -4120
rect 7244 -3800 7644 -3760
rect 7244 -4120 7284 -3800
rect 7604 -4120 7644 -3800
rect 7244 -4160 7644 -4120
rect 8256 -3800 8656 -3760
rect 8256 -4120 8296 -3800
rect 8616 -4120 8656 -3800
rect 8256 -4160 8656 -4120
rect 9268 -3800 9668 -3760
rect 9268 -4120 9308 -3800
rect 9628 -4120 9668 -3800
rect 9268 -4160 9668 -4120
rect 10280 -3800 10680 -3760
rect 10280 -4120 10320 -3800
rect 10640 -4120 10680 -3800
rect 10280 -4160 10680 -4120
rect 11292 -3800 11692 -3760
rect 11292 -4120 11332 -3800
rect 11652 -4120 11692 -3800
rect 11292 -4160 11692 -4120
rect 12304 -3800 12704 -3760
rect 12304 -4120 12344 -3800
rect 12664 -4120 12704 -3800
rect 12304 -4160 12704 -4120
rect 13316 -3800 13716 -3760
rect 13316 -4120 13356 -3800
rect 13676 -4120 13716 -3800
rect 13316 -4160 13716 -4120
rect 14328 -3800 14728 -3760
rect 14328 -4120 14368 -3800
rect 14688 -4120 14728 -3800
rect 14328 -4160 14728 -4120
rect 15340 -3800 15740 -3760
rect 15340 -4120 15380 -3800
rect 15700 -4120 15740 -3800
rect 15340 -4160 15740 -4120
rect 16352 -3800 16752 -3760
rect 16352 -4120 16392 -3800
rect 16712 -4120 16752 -3800
rect 16352 -4160 16752 -4120
rect 17364 -3800 17764 -3760
rect 17364 -4120 17404 -3800
rect 17724 -4120 17764 -3800
rect 17364 -4160 17764 -4120
rect 18376 -3800 18776 -3760
rect 18376 -4120 18416 -3800
rect 18736 -4120 18776 -3800
rect 18376 -4160 18776 -4120
rect 19388 -3800 19788 -3760
rect 19388 -4120 19428 -3800
rect 19748 -4120 19788 -3800
rect 19388 -4160 19788 -4120
rect 20400 -3800 20800 -3760
rect 20400 -4120 20440 -3800
rect 20760 -4120 20800 -3800
rect 20400 -4160 20800 -4120
rect 21412 -3800 21812 -3760
rect 21412 -4120 21452 -3800
rect 21772 -4120 21812 -3800
rect 21412 -4160 21812 -4120
rect 22424 -3800 22824 -3760
rect 22424 -4120 22464 -3800
rect 22784 -4120 22824 -3800
rect 22424 -4160 22824 -4120
rect 23436 -3800 23836 -3760
rect 23436 -4120 23476 -3800
rect 23796 -4120 23836 -3800
rect 23436 -4160 23836 -4120
rect 24448 -3800 24848 -3760
rect 24448 -4120 24488 -3800
rect 24808 -4120 24848 -3800
rect 24448 -4160 24848 -4120
rect 25460 -3800 25860 -3760
rect 25460 -4120 25500 -3800
rect 25820 -4120 25860 -3800
rect 25460 -4160 25860 -4120
rect 26472 -3800 26872 -3760
rect 26472 -4120 26512 -3800
rect 26832 -4120 26872 -3800
rect 26472 -4160 26872 -4120
rect 27484 -3800 27884 -3760
rect 27484 -4120 27524 -3800
rect 27844 -4120 27884 -3800
rect 27484 -4160 27884 -4120
rect 28496 -3800 28896 -3760
rect 28496 -4120 28536 -3800
rect 28856 -4120 28896 -3800
rect 28496 -4160 28896 -4120
rect 29508 -3800 29908 -3760
rect 29508 -4120 29548 -3800
rect 29868 -4120 29908 -3800
rect 29508 -4160 29908 -4120
rect 30520 -3800 30920 -3760
rect 30520 -4120 30560 -3800
rect 30880 -4120 30920 -3800
rect 30520 -4160 30920 -4120
rect 31532 -3800 31932 -3760
rect 31532 -4120 31572 -3800
rect 31892 -4120 31932 -3800
rect 31532 -4160 31932 -4120
rect -32224 -4520 -31824 -4480
rect -32224 -4840 -32184 -4520
rect -31864 -4840 -31824 -4520
rect -32224 -4880 -31824 -4840
rect -31212 -4520 -30812 -4480
rect -31212 -4840 -31172 -4520
rect -30852 -4840 -30812 -4520
rect -31212 -4880 -30812 -4840
rect -30200 -4520 -29800 -4480
rect -30200 -4840 -30160 -4520
rect -29840 -4840 -29800 -4520
rect -30200 -4880 -29800 -4840
rect -29188 -4520 -28788 -4480
rect -29188 -4840 -29148 -4520
rect -28828 -4840 -28788 -4520
rect -29188 -4880 -28788 -4840
rect -28176 -4520 -27776 -4480
rect -28176 -4840 -28136 -4520
rect -27816 -4840 -27776 -4520
rect -28176 -4880 -27776 -4840
rect -27164 -4520 -26764 -4480
rect -27164 -4840 -27124 -4520
rect -26804 -4840 -26764 -4520
rect -27164 -4880 -26764 -4840
rect -26152 -4520 -25752 -4480
rect -26152 -4840 -26112 -4520
rect -25792 -4840 -25752 -4520
rect -26152 -4880 -25752 -4840
rect -25140 -4520 -24740 -4480
rect -25140 -4840 -25100 -4520
rect -24780 -4840 -24740 -4520
rect -25140 -4880 -24740 -4840
rect -24128 -4520 -23728 -4480
rect -24128 -4840 -24088 -4520
rect -23768 -4840 -23728 -4520
rect -24128 -4880 -23728 -4840
rect -23116 -4520 -22716 -4480
rect -23116 -4840 -23076 -4520
rect -22756 -4840 -22716 -4520
rect -23116 -4880 -22716 -4840
rect -22104 -4520 -21704 -4480
rect -22104 -4840 -22064 -4520
rect -21744 -4840 -21704 -4520
rect -22104 -4880 -21704 -4840
rect -21092 -4520 -20692 -4480
rect -21092 -4840 -21052 -4520
rect -20732 -4840 -20692 -4520
rect -21092 -4880 -20692 -4840
rect -20080 -4520 -19680 -4480
rect -20080 -4840 -20040 -4520
rect -19720 -4840 -19680 -4520
rect -20080 -4880 -19680 -4840
rect -19068 -4520 -18668 -4480
rect -19068 -4840 -19028 -4520
rect -18708 -4840 -18668 -4520
rect -19068 -4880 -18668 -4840
rect -18056 -4520 -17656 -4480
rect -18056 -4840 -18016 -4520
rect -17696 -4840 -17656 -4520
rect -18056 -4880 -17656 -4840
rect -17044 -4520 -16644 -4480
rect -17044 -4840 -17004 -4520
rect -16684 -4840 -16644 -4520
rect -17044 -4880 -16644 -4840
rect -16032 -4520 -15632 -4480
rect -16032 -4840 -15992 -4520
rect -15672 -4840 -15632 -4520
rect -16032 -4880 -15632 -4840
rect -15020 -4520 -14620 -4480
rect -15020 -4840 -14980 -4520
rect -14660 -4840 -14620 -4520
rect -15020 -4880 -14620 -4840
rect -14008 -4520 -13608 -4480
rect -14008 -4840 -13968 -4520
rect -13648 -4840 -13608 -4520
rect -14008 -4880 -13608 -4840
rect -12996 -4520 -12596 -4480
rect -12996 -4840 -12956 -4520
rect -12636 -4840 -12596 -4520
rect -12996 -4880 -12596 -4840
rect -11984 -4520 -11584 -4480
rect -11984 -4840 -11944 -4520
rect -11624 -4840 -11584 -4520
rect -11984 -4880 -11584 -4840
rect -10972 -4520 -10572 -4480
rect -10972 -4840 -10932 -4520
rect -10612 -4840 -10572 -4520
rect -10972 -4880 -10572 -4840
rect -9960 -4520 -9560 -4480
rect -9960 -4840 -9920 -4520
rect -9600 -4840 -9560 -4520
rect -9960 -4880 -9560 -4840
rect -8948 -4520 -8548 -4480
rect -8948 -4840 -8908 -4520
rect -8588 -4840 -8548 -4520
rect -8948 -4880 -8548 -4840
rect -7936 -4520 -7536 -4480
rect -7936 -4840 -7896 -4520
rect -7576 -4840 -7536 -4520
rect -7936 -4880 -7536 -4840
rect -6924 -4520 -6524 -4480
rect -6924 -4840 -6884 -4520
rect -6564 -4840 -6524 -4520
rect -6924 -4880 -6524 -4840
rect -5912 -4520 -5512 -4480
rect -5912 -4840 -5872 -4520
rect -5552 -4840 -5512 -4520
rect -5912 -4880 -5512 -4840
rect -4900 -4520 -4500 -4480
rect -4900 -4840 -4860 -4520
rect -4540 -4840 -4500 -4520
rect -4900 -4880 -4500 -4840
rect -3888 -4520 -3488 -4480
rect -3888 -4840 -3848 -4520
rect -3528 -4840 -3488 -4520
rect -3888 -4880 -3488 -4840
rect -2876 -4520 -2476 -4480
rect -2876 -4840 -2836 -4520
rect -2516 -4840 -2476 -4520
rect -2876 -4880 -2476 -4840
rect -1864 -4520 -1464 -4480
rect -1864 -4840 -1824 -4520
rect -1504 -4840 -1464 -4520
rect -1864 -4880 -1464 -4840
rect -852 -4520 -452 -4480
rect -852 -4840 -812 -4520
rect -492 -4840 -452 -4520
rect -852 -4880 -452 -4840
rect 160 -4520 560 -4480
rect 160 -4840 200 -4520
rect 520 -4840 560 -4520
rect 160 -4880 560 -4840
rect 1172 -4520 1572 -4480
rect 1172 -4840 1212 -4520
rect 1532 -4840 1572 -4520
rect 1172 -4880 1572 -4840
rect 2184 -4520 2584 -4480
rect 2184 -4840 2224 -4520
rect 2544 -4840 2584 -4520
rect 2184 -4880 2584 -4840
rect 3196 -4520 3596 -4480
rect 3196 -4840 3236 -4520
rect 3556 -4840 3596 -4520
rect 3196 -4880 3596 -4840
rect 4208 -4520 4608 -4480
rect 4208 -4840 4248 -4520
rect 4568 -4840 4608 -4520
rect 4208 -4880 4608 -4840
rect 5220 -4520 5620 -4480
rect 5220 -4840 5260 -4520
rect 5580 -4840 5620 -4520
rect 5220 -4880 5620 -4840
rect 6232 -4520 6632 -4480
rect 6232 -4840 6272 -4520
rect 6592 -4840 6632 -4520
rect 6232 -4880 6632 -4840
rect 7244 -4520 7644 -4480
rect 7244 -4840 7284 -4520
rect 7604 -4840 7644 -4520
rect 7244 -4880 7644 -4840
rect 8256 -4520 8656 -4480
rect 8256 -4840 8296 -4520
rect 8616 -4840 8656 -4520
rect 8256 -4880 8656 -4840
rect 9268 -4520 9668 -4480
rect 9268 -4840 9308 -4520
rect 9628 -4840 9668 -4520
rect 9268 -4880 9668 -4840
rect 10280 -4520 10680 -4480
rect 10280 -4840 10320 -4520
rect 10640 -4840 10680 -4520
rect 10280 -4880 10680 -4840
rect 11292 -4520 11692 -4480
rect 11292 -4840 11332 -4520
rect 11652 -4840 11692 -4520
rect 11292 -4880 11692 -4840
rect 12304 -4520 12704 -4480
rect 12304 -4840 12344 -4520
rect 12664 -4840 12704 -4520
rect 12304 -4880 12704 -4840
rect 13316 -4520 13716 -4480
rect 13316 -4840 13356 -4520
rect 13676 -4840 13716 -4520
rect 13316 -4880 13716 -4840
rect 14328 -4520 14728 -4480
rect 14328 -4840 14368 -4520
rect 14688 -4840 14728 -4520
rect 14328 -4880 14728 -4840
rect 15340 -4520 15740 -4480
rect 15340 -4840 15380 -4520
rect 15700 -4840 15740 -4520
rect 15340 -4880 15740 -4840
rect 16352 -4520 16752 -4480
rect 16352 -4840 16392 -4520
rect 16712 -4840 16752 -4520
rect 16352 -4880 16752 -4840
rect 17364 -4520 17764 -4480
rect 17364 -4840 17404 -4520
rect 17724 -4840 17764 -4520
rect 17364 -4880 17764 -4840
rect 18376 -4520 18776 -4480
rect 18376 -4840 18416 -4520
rect 18736 -4840 18776 -4520
rect 18376 -4880 18776 -4840
rect 19388 -4520 19788 -4480
rect 19388 -4840 19428 -4520
rect 19748 -4840 19788 -4520
rect 19388 -4880 19788 -4840
rect 20400 -4520 20800 -4480
rect 20400 -4840 20440 -4520
rect 20760 -4840 20800 -4520
rect 20400 -4880 20800 -4840
rect 21412 -4520 21812 -4480
rect 21412 -4840 21452 -4520
rect 21772 -4840 21812 -4520
rect 21412 -4880 21812 -4840
rect 22424 -4520 22824 -4480
rect 22424 -4840 22464 -4520
rect 22784 -4840 22824 -4520
rect 22424 -4880 22824 -4840
rect 23436 -4520 23836 -4480
rect 23436 -4840 23476 -4520
rect 23796 -4840 23836 -4520
rect 23436 -4880 23836 -4840
rect 24448 -4520 24848 -4480
rect 24448 -4840 24488 -4520
rect 24808 -4840 24848 -4520
rect 24448 -4880 24848 -4840
rect 25460 -4520 25860 -4480
rect 25460 -4840 25500 -4520
rect 25820 -4840 25860 -4520
rect 25460 -4880 25860 -4840
rect 26472 -4520 26872 -4480
rect 26472 -4840 26512 -4520
rect 26832 -4840 26872 -4520
rect 26472 -4880 26872 -4840
rect 27484 -4520 27884 -4480
rect 27484 -4840 27524 -4520
rect 27844 -4840 27884 -4520
rect 27484 -4880 27884 -4840
rect 28496 -4520 28896 -4480
rect 28496 -4840 28536 -4520
rect 28856 -4840 28896 -4520
rect 28496 -4880 28896 -4840
rect 29508 -4520 29908 -4480
rect 29508 -4840 29548 -4520
rect 29868 -4840 29908 -4520
rect 29508 -4880 29908 -4840
rect 30520 -4520 30920 -4480
rect 30520 -4840 30560 -4520
rect 30880 -4840 30920 -4520
rect 30520 -4880 30920 -4840
rect 31532 -4520 31932 -4480
rect 31532 -4840 31572 -4520
rect 31892 -4840 31932 -4520
rect 31532 -4880 31932 -4840
rect -32224 -5240 -31824 -5200
rect -32224 -5560 -32184 -5240
rect -31864 -5560 -31824 -5240
rect -32224 -5600 -31824 -5560
rect -31212 -5240 -30812 -5200
rect -31212 -5560 -31172 -5240
rect -30852 -5560 -30812 -5240
rect -31212 -5600 -30812 -5560
rect -30200 -5240 -29800 -5200
rect -30200 -5560 -30160 -5240
rect -29840 -5560 -29800 -5240
rect -30200 -5600 -29800 -5560
rect -29188 -5240 -28788 -5200
rect -29188 -5560 -29148 -5240
rect -28828 -5560 -28788 -5240
rect -29188 -5600 -28788 -5560
rect -28176 -5240 -27776 -5200
rect -28176 -5560 -28136 -5240
rect -27816 -5560 -27776 -5240
rect -28176 -5600 -27776 -5560
rect -27164 -5240 -26764 -5200
rect -27164 -5560 -27124 -5240
rect -26804 -5560 -26764 -5240
rect -27164 -5600 -26764 -5560
rect -26152 -5240 -25752 -5200
rect -26152 -5560 -26112 -5240
rect -25792 -5560 -25752 -5240
rect -26152 -5600 -25752 -5560
rect -25140 -5240 -24740 -5200
rect -25140 -5560 -25100 -5240
rect -24780 -5560 -24740 -5240
rect -25140 -5600 -24740 -5560
rect -24128 -5240 -23728 -5200
rect -24128 -5560 -24088 -5240
rect -23768 -5560 -23728 -5240
rect -24128 -5600 -23728 -5560
rect -23116 -5240 -22716 -5200
rect -23116 -5560 -23076 -5240
rect -22756 -5560 -22716 -5240
rect -23116 -5600 -22716 -5560
rect -22104 -5240 -21704 -5200
rect -22104 -5560 -22064 -5240
rect -21744 -5560 -21704 -5240
rect -22104 -5600 -21704 -5560
rect -21092 -5240 -20692 -5200
rect -21092 -5560 -21052 -5240
rect -20732 -5560 -20692 -5240
rect -21092 -5600 -20692 -5560
rect -20080 -5240 -19680 -5200
rect -20080 -5560 -20040 -5240
rect -19720 -5560 -19680 -5240
rect -20080 -5600 -19680 -5560
rect -19068 -5240 -18668 -5200
rect -19068 -5560 -19028 -5240
rect -18708 -5560 -18668 -5240
rect -19068 -5600 -18668 -5560
rect -18056 -5240 -17656 -5200
rect -18056 -5560 -18016 -5240
rect -17696 -5560 -17656 -5240
rect -18056 -5600 -17656 -5560
rect -17044 -5240 -16644 -5200
rect -17044 -5560 -17004 -5240
rect -16684 -5560 -16644 -5240
rect -17044 -5600 -16644 -5560
rect -16032 -5240 -15632 -5200
rect -16032 -5560 -15992 -5240
rect -15672 -5560 -15632 -5240
rect -16032 -5600 -15632 -5560
rect -15020 -5240 -14620 -5200
rect -15020 -5560 -14980 -5240
rect -14660 -5560 -14620 -5240
rect -15020 -5600 -14620 -5560
rect -14008 -5240 -13608 -5200
rect -14008 -5560 -13968 -5240
rect -13648 -5560 -13608 -5240
rect -14008 -5600 -13608 -5560
rect -12996 -5240 -12596 -5200
rect -12996 -5560 -12956 -5240
rect -12636 -5560 -12596 -5240
rect -12996 -5600 -12596 -5560
rect -11984 -5240 -11584 -5200
rect -11984 -5560 -11944 -5240
rect -11624 -5560 -11584 -5240
rect -11984 -5600 -11584 -5560
rect -10972 -5240 -10572 -5200
rect -10972 -5560 -10932 -5240
rect -10612 -5560 -10572 -5240
rect -10972 -5600 -10572 -5560
rect -9960 -5240 -9560 -5200
rect -9960 -5560 -9920 -5240
rect -9600 -5560 -9560 -5240
rect -9960 -5600 -9560 -5560
rect -8948 -5240 -8548 -5200
rect -8948 -5560 -8908 -5240
rect -8588 -5560 -8548 -5240
rect -8948 -5600 -8548 -5560
rect -7936 -5240 -7536 -5200
rect -7936 -5560 -7896 -5240
rect -7576 -5560 -7536 -5240
rect -7936 -5600 -7536 -5560
rect -6924 -5240 -6524 -5200
rect -6924 -5560 -6884 -5240
rect -6564 -5560 -6524 -5240
rect -6924 -5600 -6524 -5560
rect -5912 -5240 -5512 -5200
rect -5912 -5560 -5872 -5240
rect -5552 -5560 -5512 -5240
rect -5912 -5600 -5512 -5560
rect -4900 -5240 -4500 -5200
rect -4900 -5560 -4860 -5240
rect -4540 -5560 -4500 -5240
rect -4900 -5600 -4500 -5560
rect -3888 -5240 -3488 -5200
rect -3888 -5560 -3848 -5240
rect -3528 -5560 -3488 -5240
rect -3888 -5600 -3488 -5560
rect -2876 -5240 -2476 -5200
rect -2876 -5560 -2836 -5240
rect -2516 -5560 -2476 -5240
rect -2876 -5600 -2476 -5560
rect -1864 -5240 -1464 -5200
rect -1864 -5560 -1824 -5240
rect -1504 -5560 -1464 -5240
rect -1864 -5600 -1464 -5560
rect -852 -5240 -452 -5200
rect -852 -5560 -812 -5240
rect -492 -5560 -452 -5240
rect -852 -5600 -452 -5560
rect 160 -5240 560 -5200
rect 160 -5560 200 -5240
rect 520 -5560 560 -5240
rect 160 -5600 560 -5560
rect 1172 -5240 1572 -5200
rect 1172 -5560 1212 -5240
rect 1532 -5560 1572 -5240
rect 1172 -5600 1572 -5560
rect 2184 -5240 2584 -5200
rect 2184 -5560 2224 -5240
rect 2544 -5560 2584 -5240
rect 2184 -5600 2584 -5560
rect 3196 -5240 3596 -5200
rect 3196 -5560 3236 -5240
rect 3556 -5560 3596 -5240
rect 3196 -5600 3596 -5560
rect 4208 -5240 4608 -5200
rect 4208 -5560 4248 -5240
rect 4568 -5560 4608 -5240
rect 4208 -5600 4608 -5560
rect 5220 -5240 5620 -5200
rect 5220 -5560 5260 -5240
rect 5580 -5560 5620 -5240
rect 5220 -5600 5620 -5560
rect 6232 -5240 6632 -5200
rect 6232 -5560 6272 -5240
rect 6592 -5560 6632 -5240
rect 6232 -5600 6632 -5560
rect 7244 -5240 7644 -5200
rect 7244 -5560 7284 -5240
rect 7604 -5560 7644 -5240
rect 7244 -5600 7644 -5560
rect 8256 -5240 8656 -5200
rect 8256 -5560 8296 -5240
rect 8616 -5560 8656 -5240
rect 8256 -5600 8656 -5560
rect 9268 -5240 9668 -5200
rect 9268 -5560 9308 -5240
rect 9628 -5560 9668 -5240
rect 9268 -5600 9668 -5560
rect 10280 -5240 10680 -5200
rect 10280 -5560 10320 -5240
rect 10640 -5560 10680 -5240
rect 10280 -5600 10680 -5560
rect 11292 -5240 11692 -5200
rect 11292 -5560 11332 -5240
rect 11652 -5560 11692 -5240
rect 11292 -5600 11692 -5560
rect 12304 -5240 12704 -5200
rect 12304 -5560 12344 -5240
rect 12664 -5560 12704 -5240
rect 12304 -5600 12704 -5560
rect 13316 -5240 13716 -5200
rect 13316 -5560 13356 -5240
rect 13676 -5560 13716 -5240
rect 13316 -5600 13716 -5560
rect 14328 -5240 14728 -5200
rect 14328 -5560 14368 -5240
rect 14688 -5560 14728 -5240
rect 14328 -5600 14728 -5560
rect 15340 -5240 15740 -5200
rect 15340 -5560 15380 -5240
rect 15700 -5560 15740 -5240
rect 15340 -5600 15740 -5560
rect 16352 -5240 16752 -5200
rect 16352 -5560 16392 -5240
rect 16712 -5560 16752 -5240
rect 16352 -5600 16752 -5560
rect 17364 -5240 17764 -5200
rect 17364 -5560 17404 -5240
rect 17724 -5560 17764 -5240
rect 17364 -5600 17764 -5560
rect 18376 -5240 18776 -5200
rect 18376 -5560 18416 -5240
rect 18736 -5560 18776 -5240
rect 18376 -5600 18776 -5560
rect 19388 -5240 19788 -5200
rect 19388 -5560 19428 -5240
rect 19748 -5560 19788 -5240
rect 19388 -5600 19788 -5560
rect 20400 -5240 20800 -5200
rect 20400 -5560 20440 -5240
rect 20760 -5560 20800 -5240
rect 20400 -5600 20800 -5560
rect 21412 -5240 21812 -5200
rect 21412 -5560 21452 -5240
rect 21772 -5560 21812 -5240
rect 21412 -5600 21812 -5560
rect 22424 -5240 22824 -5200
rect 22424 -5560 22464 -5240
rect 22784 -5560 22824 -5240
rect 22424 -5600 22824 -5560
rect 23436 -5240 23836 -5200
rect 23436 -5560 23476 -5240
rect 23796 -5560 23836 -5240
rect 23436 -5600 23836 -5560
rect 24448 -5240 24848 -5200
rect 24448 -5560 24488 -5240
rect 24808 -5560 24848 -5240
rect 24448 -5600 24848 -5560
rect 25460 -5240 25860 -5200
rect 25460 -5560 25500 -5240
rect 25820 -5560 25860 -5240
rect 25460 -5600 25860 -5560
rect 26472 -5240 26872 -5200
rect 26472 -5560 26512 -5240
rect 26832 -5560 26872 -5240
rect 26472 -5600 26872 -5560
rect 27484 -5240 27884 -5200
rect 27484 -5560 27524 -5240
rect 27844 -5560 27884 -5240
rect 27484 -5600 27884 -5560
rect 28496 -5240 28896 -5200
rect 28496 -5560 28536 -5240
rect 28856 -5560 28896 -5240
rect 28496 -5600 28896 -5560
rect 29508 -5240 29908 -5200
rect 29508 -5560 29548 -5240
rect 29868 -5560 29908 -5240
rect 29508 -5600 29908 -5560
rect 30520 -5240 30920 -5200
rect 30520 -5560 30560 -5240
rect 30880 -5560 30920 -5240
rect 30520 -5600 30920 -5560
rect 31532 -5240 31932 -5200
rect 31532 -5560 31572 -5240
rect 31892 -5560 31932 -5240
rect 31532 -5600 31932 -5560
<< mimcapcontact >>
rect -32184 5240 -31864 5560
rect -31172 5240 -30852 5560
rect -30160 5240 -29840 5560
rect -29148 5240 -28828 5560
rect -28136 5240 -27816 5560
rect -27124 5240 -26804 5560
rect -26112 5240 -25792 5560
rect -25100 5240 -24780 5560
rect -24088 5240 -23768 5560
rect -23076 5240 -22756 5560
rect -22064 5240 -21744 5560
rect -21052 5240 -20732 5560
rect -20040 5240 -19720 5560
rect -19028 5240 -18708 5560
rect -18016 5240 -17696 5560
rect -17004 5240 -16684 5560
rect -15992 5240 -15672 5560
rect -14980 5240 -14660 5560
rect -13968 5240 -13648 5560
rect -12956 5240 -12636 5560
rect -11944 5240 -11624 5560
rect -10932 5240 -10612 5560
rect -9920 5240 -9600 5560
rect -8908 5240 -8588 5560
rect -7896 5240 -7576 5560
rect -6884 5240 -6564 5560
rect -5872 5240 -5552 5560
rect -4860 5240 -4540 5560
rect -3848 5240 -3528 5560
rect -2836 5240 -2516 5560
rect -1824 5240 -1504 5560
rect -812 5240 -492 5560
rect 200 5240 520 5560
rect 1212 5240 1532 5560
rect 2224 5240 2544 5560
rect 3236 5240 3556 5560
rect 4248 5240 4568 5560
rect 5260 5240 5580 5560
rect 6272 5240 6592 5560
rect 7284 5240 7604 5560
rect 8296 5240 8616 5560
rect 9308 5240 9628 5560
rect 10320 5240 10640 5560
rect 11332 5240 11652 5560
rect 12344 5240 12664 5560
rect 13356 5240 13676 5560
rect 14368 5240 14688 5560
rect 15380 5240 15700 5560
rect 16392 5240 16712 5560
rect 17404 5240 17724 5560
rect 18416 5240 18736 5560
rect 19428 5240 19748 5560
rect 20440 5240 20760 5560
rect 21452 5240 21772 5560
rect 22464 5240 22784 5560
rect 23476 5240 23796 5560
rect 24488 5240 24808 5560
rect 25500 5240 25820 5560
rect 26512 5240 26832 5560
rect 27524 5240 27844 5560
rect 28536 5240 28856 5560
rect 29548 5240 29868 5560
rect 30560 5240 30880 5560
rect 31572 5240 31892 5560
rect -32184 4520 -31864 4840
rect -31172 4520 -30852 4840
rect -30160 4520 -29840 4840
rect -29148 4520 -28828 4840
rect -28136 4520 -27816 4840
rect -27124 4520 -26804 4840
rect -26112 4520 -25792 4840
rect -25100 4520 -24780 4840
rect -24088 4520 -23768 4840
rect -23076 4520 -22756 4840
rect -22064 4520 -21744 4840
rect -21052 4520 -20732 4840
rect -20040 4520 -19720 4840
rect -19028 4520 -18708 4840
rect -18016 4520 -17696 4840
rect -17004 4520 -16684 4840
rect -15992 4520 -15672 4840
rect -14980 4520 -14660 4840
rect -13968 4520 -13648 4840
rect -12956 4520 -12636 4840
rect -11944 4520 -11624 4840
rect -10932 4520 -10612 4840
rect -9920 4520 -9600 4840
rect -8908 4520 -8588 4840
rect -7896 4520 -7576 4840
rect -6884 4520 -6564 4840
rect -5872 4520 -5552 4840
rect -4860 4520 -4540 4840
rect -3848 4520 -3528 4840
rect -2836 4520 -2516 4840
rect -1824 4520 -1504 4840
rect -812 4520 -492 4840
rect 200 4520 520 4840
rect 1212 4520 1532 4840
rect 2224 4520 2544 4840
rect 3236 4520 3556 4840
rect 4248 4520 4568 4840
rect 5260 4520 5580 4840
rect 6272 4520 6592 4840
rect 7284 4520 7604 4840
rect 8296 4520 8616 4840
rect 9308 4520 9628 4840
rect 10320 4520 10640 4840
rect 11332 4520 11652 4840
rect 12344 4520 12664 4840
rect 13356 4520 13676 4840
rect 14368 4520 14688 4840
rect 15380 4520 15700 4840
rect 16392 4520 16712 4840
rect 17404 4520 17724 4840
rect 18416 4520 18736 4840
rect 19428 4520 19748 4840
rect 20440 4520 20760 4840
rect 21452 4520 21772 4840
rect 22464 4520 22784 4840
rect 23476 4520 23796 4840
rect 24488 4520 24808 4840
rect 25500 4520 25820 4840
rect 26512 4520 26832 4840
rect 27524 4520 27844 4840
rect 28536 4520 28856 4840
rect 29548 4520 29868 4840
rect 30560 4520 30880 4840
rect 31572 4520 31892 4840
rect -32184 3800 -31864 4120
rect -31172 3800 -30852 4120
rect -30160 3800 -29840 4120
rect -29148 3800 -28828 4120
rect -28136 3800 -27816 4120
rect -27124 3800 -26804 4120
rect -26112 3800 -25792 4120
rect -25100 3800 -24780 4120
rect -24088 3800 -23768 4120
rect -23076 3800 -22756 4120
rect -22064 3800 -21744 4120
rect -21052 3800 -20732 4120
rect -20040 3800 -19720 4120
rect -19028 3800 -18708 4120
rect -18016 3800 -17696 4120
rect -17004 3800 -16684 4120
rect -15992 3800 -15672 4120
rect -14980 3800 -14660 4120
rect -13968 3800 -13648 4120
rect -12956 3800 -12636 4120
rect -11944 3800 -11624 4120
rect -10932 3800 -10612 4120
rect -9920 3800 -9600 4120
rect -8908 3800 -8588 4120
rect -7896 3800 -7576 4120
rect -6884 3800 -6564 4120
rect -5872 3800 -5552 4120
rect -4860 3800 -4540 4120
rect -3848 3800 -3528 4120
rect -2836 3800 -2516 4120
rect -1824 3800 -1504 4120
rect -812 3800 -492 4120
rect 200 3800 520 4120
rect 1212 3800 1532 4120
rect 2224 3800 2544 4120
rect 3236 3800 3556 4120
rect 4248 3800 4568 4120
rect 5260 3800 5580 4120
rect 6272 3800 6592 4120
rect 7284 3800 7604 4120
rect 8296 3800 8616 4120
rect 9308 3800 9628 4120
rect 10320 3800 10640 4120
rect 11332 3800 11652 4120
rect 12344 3800 12664 4120
rect 13356 3800 13676 4120
rect 14368 3800 14688 4120
rect 15380 3800 15700 4120
rect 16392 3800 16712 4120
rect 17404 3800 17724 4120
rect 18416 3800 18736 4120
rect 19428 3800 19748 4120
rect 20440 3800 20760 4120
rect 21452 3800 21772 4120
rect 22464 3800 22784 4120
rect 23476 3800 23796 4120
rect 24488 3800 24808 4120
rect 25500 3800 25820 4120
rect 26512 3800 26832 4120
rect 27524 3800 27844 4120
rect 28536 3800 28856 4120
rect 29548 3800 29868 4120
rect 30560 3800 30880 4120
rect 31572 3800 31892 4120
rect -32184 3080 -31864 3400
rect -31172 3080 -30852 3400
rect -30160 3080 -29840 3400
rect -29148 3080 -28828 3400
rect -28136 3080 -27816 3400
rect -27124 3080 -26804 3400
rect -26112 3080 -25792 3400
rect -25100 3080 -24780 3400
rect -24088 3080 -23768 3400
rect -23076 3080 -22756 3400
rect -22064 3080 -21744 3400
rect -21052 3080 -20732 3400
rect -20040 3080 -19720 3400
rect -19028 3080 -18708 3400
rect -18016 3080 -17696 3400
rect -17004 3080 -16684 3400
rect -15992 3080 -15672 3400
rect -14980 3080 -14660 3400
rect -13968 3080 -13648 3400
rect -12956 3080 -12636 3400
rect -11944 3080 -11624 3400
rect -10932 3080 -10612 3400
rect -9920 3080 -9600 3400
rect -8908 3080 -8588 3400
rect -7896 3080 -7576 3400
rect -6884 3080 -6564 3400
rect -5872 3080 -5552 3400
rect -4860 3080 -4540 3400
rect -3848 3080 -3528 3400
rect -2836 3080 -2516 3400
rect -1824 3080 -1504 3400
rect -812 3080 -492 3400
rect 200 3080 520 3400
rect 1212 3080 1532 3400
rect 2224 3080 2544 3400
rect 3236 3080 3556 3400
rect 4248 3080 4568 3400
rect 5260 3080 5580 3400
rect 6272 3080 6592 3400
rect 7284 3080 7604 3400
rect 8296 3080 8616 3400
rect 9308 3080 9628 3400
rect 10320 3080 10640 3400
rect 11332 3080 11652 3400
rect 12344 3080 12664 3400
rect 13356 3080 13676 3400
rect 14368 3080 14688 3400
rect 15380 3080 15700 3400
rect 16392 3080 16712 3400
rect 17404 3080 17724 3400
rect 18416 3080 18736 3400
rect 19428 3080 19748 3400
rect 20440 3080 20760 3400
rect 21452 3080 21772 3400
rect 22464 3080 22784 3400
rect 23476 3080 23796 3400
rect 24488 3080 24808 3400
rect 25500 3080 25820 3400
rect 26512 3080 26832 3400
rect 27524 3080 27844 3400
rect 28536 3080 28856 3400
rect 29548 3080 29868 3400
rect 30560 3080 30880 3400
rect 31572 3080 31892 3400
rect -32184 2360 -31864 2680
rect -31172 2360 -30852 2680
rect -30160 2360 -29840 2680
rect -29148 2360 -28828 2680
rect -28136 2360 -27816 2680
rect -27124 2360 -26804 2680
rect -26112 2360 -25792 2680
rect -25100 2360 -24780 2680
rect -24088 2360 -23768 2680
rect -23076 2360 -22756 2680
rect -22064 2360 -21744 2680
rect -21052 2360 -20732 2680
rect -20040 2360 -19720 2680
rect -19028 2360 -18708 2680
rect -18016 2360 -17696 2680
rect -17004 2360 -16684 2680
rect -15992 2360 -15672 2680
rect -14980 2360 -14660 2680
rect -13968 2360 -13648 2680
rect -12956 2360 -12636 2680
rect -11944 2360 -11624 2680
rect -10932 2360 -10612 2680
rect -9920 2360 -9600 2680
rect -8908 2360 -8588 2680
rect -7896 2360 -7576 2680
rect -6884 2360 -6564 2680
rect -5872 2360 -5552 2680
rect -4860 2360 -4540 2680
rect -3848 2360 -3528 2680
rect -2836 2360 -2516 2680
rect -1824 2360 -1504 2680
rect -812 2360 -492 2680
rect 200 2360 520 2680
rect 1212 2360 1532 2680
rect 2224 2360 2544 2680
rect 3236 2360 3556 2680
rect 4248 2360 4568 2680
rect 5260 2360 5580 2680
rect 6272 2360 6592 2680
rect 7284 2360 7604 2680
rect 8296 2360 8616 2680
rect 9308 2360 9628 2680
rect 10320 2360 10640 2680
rect 11332 2360 11652 2680
rect 12344 2360 12664 2680
rect 13356 2360 13676 2680
rect 14368 2360 14688 2680
rect 15380 2360 15700 2680
rect 16392 2360 16712 2680
rect 17404 2360 17724 2680
rect 18416 2360 18736 2680
rect 19428 2360 19748 2680
rect 20440 2360 20760 2680
rect 21452 2360 21772 2680
rect 22464 2360 22784 2680
rect 23476 2360 23796 2680
rect 24488 2360 24808 2680
rect 25500 2360 25820 2680
rect 26512 2360 26832 2680
rect 27524 2360 27844 2680
rect 28536 2360 28856 2680
rect 29548 2360 29868 2680
rect 30560 2360 30880 2680
rect 31572 2360 31892 2680
rect -32184 1640 -31864 1960
rect -31172 1640 -30852 1960
rect -30160 1640 -29840 1960
rect -29148 1640 -28828 1960
rect -28136 1640 -27816 1960
rect -27124 1640 -26804 1960
rect -26112 1640 -25792 1960
rect -25100 1640 -24780 1960
rect -24088 1640 -23768 1960
rect -23076 1640 -22756 1960
rect -22064 1640 -21744 1960
rect -21052 1640 -20732 1960
rect -20040 1640 -19720 1960
rect -19028 1640 -18708 1960
rect -18016 1640 -17696 1960
rect -17004 1640 -16684 1960
rect -15992 1640 -15672 1960
rect -14980 1640 -14660 1960
rect -13968 1640 -13648 1960
rect -12956 1640 -12636 1960
rect -11944 1640 -11624 1960
rect -10932 1640 -10612 1960
rect -9920 1640 -9600 1960
rect -8908 1640 -8588 1960
rect -7896 1640 -7576 1960
rect -6884 1640 -6564 1960
rect -5872 1640 -5552 1960
rect -4860 1640 -4540 1960
rect -3848 1640 -3528 1960
rect -2836 1640 -2516 1960
rect -1824 1640 -1504 1960
rect -812 1640 -492 1960
rect 200 1640 520 1960
rect 1212 1640 1532 1960
rect 2224 1640 2544 1960
rect 3236 1640 3556 1960
rect 4248 1640 4568 1960
rect 5260 1640 5580 1960
rect 6272 1640 6592 1960
rect 7284 1640 7604 1960
rect 8296 1640 8616 1960
rect 9308 1640 9628 1960
rect 10320 1640 10640 1960
rect 11332 1640 11652 1960
rect 12344 1640 12664 1960
rect 13356 1640 13676 1960
rect 14368 1640 14688 1960
rect 15380 1640 15700 1960
rect 16392 1640 16712 1960
rect 17404 1640 17724 1960
rect 18416 1640 18736 1960
rect 19428 1640 19748 1960
rect 20440 1640 20760 1960
rect 21452 1640 21772 1960
rect 22464 1640 22784 1960
rect 23476 1640 23796 1960
rect 24488 1640 24808 1960
rect 25500 1640 25820 1960
rect 26512 1640 26832 1960
rect 27524 1640 27844 1960
rect 28536 1640 28856 1960
rect 29548 1640 29868 1960
rect 30560 1640 30880 1960
rect 31572 1640 31892 1960
rect -32184 920 -31864 1240
rect -31172 920 -30852 1240
rect -30160 920 -29840 1240
rect -29148 920 -28828 1240
rect -28136 920 -27816 1240
rect -27124 920 -26804 1240
rect -26112 920 -25792 1240
rect -25100 920 -24780 1240
rect -24088 920 -23768 1240
rect -23076 920 -22756 1240
rect -22064 920 -21744 1240
rect -21052 920 -20732 1240
rect -20040 920 -19720 1240
rect -19028 920 -18708 1240
rect -18016 920 -17696 1240
rect -17004 920 -16684 1240
rect -15992 920 -15672 1240
rect -14980 920 -14660 1240
rect -13968 920 -13648 1240
rect -12956 920 -12636 1240
rect -11944 920 -11624 1240
rect -10932 920 -10612 1240
rect -9920 920 -9600 1240
rect -8908 920 -8588 1240
rect -7896 920 -7576 1240
rect -6884 920 -6564 1240
rect -5872 920 -5552 1240
rect -4860 920 -4540 1240
rect -3848 920 -3528 1240
rect -2836 920 -2516 1240
rect -1824 920 -1504 1240
rect -812 920 -492 1240
rect 200 920 520 1240
rect 1212 920 1532 1240
rect 2224 920 2544 1240
rect 3236 920 3556 1240
rect 4248 920 4568 1240
rect 5260 920 5580 1240
rect 6272 920 6592 1240
rect 7284 920 7604 1240
rect 8296 920 8616 1240
rect 9308 920 9628 1240
rect 10320 920 10640 1240
rect 11332 920 11652 1240
rect 12344 920 12664 1240
rect 13356 920 13676 1240
rect 14368 920 14688 1240
rect 15380 920 15700 1240
rect 16392 920 16712 1240
rect 17404 920 17724 1240
rect 18416 920 18736 1240
rect 19428 920 19748 1240
rect 20440 920 20760 1240
rect 21452 920 21772 1240
rect 22464 920 22784 1240
rect 23476 920 23796 1240
rect 24488 920 24808 1240
rect 25500 920 25820 1240
rect 26512 920 26832 1240
rect 27524 920 27844 1240
rect 28536 920 28856 1240
rect 29548 920 29868 1240
rect 30560 920 30880 1240
rect 31572 920 31892 1240
rect -32184 200 -31864 520
rect -31172 200 -30852 520
rect -30160 200 -29840 520
rect -29148 200 -28828 520
rect -28136 200 -27816 520
rect -27124 200 -26804 520
rect -26112 200 -25792 520
rect -25100 200 -24780 520
rect -24088 200 -23768 520
rect -23076 200 -22756 520
rect -22064 200 -21744 520
rect -21052 200 -20732 520
rect -20040 200 -19720 520
rect -19028 200 -18708 520
rect -18016 200 -17696 520
rect -17004 200 -16684 520
rect -15992 200 -15672 520
rect -14980 200 -14660 520
rect -13968 200 -13648 520
rect -12956 200 -12636 520
rect -11944 200 -11624 520
rect -10932 200 -10612 520
rect -9920 200 -9600 520
rect -8908 200 -8588 520
rect -7896 200 -7576 520
rect -6884 200 -6564 520
rect -5872 200 -5552 520
rect -4860 200 -4540 520
rect -3848 200 -3528 520
rect -2836 200 -2516 520
rect -1824 200 -1504 520
rect -812 200 -492 520
rect 200 200 520 520
rect 1212 200 1532 520
rect 2224 200 2544 520
rect 3236 200 3556 520
rect 4248 200 4568 520
rect 5260 200 5580 520
rect 6272 200 6592 520
rect 7284 200 7604 520
rect 8296 200 8616 520
rect 9308 200 9628 520
rect 10320 200 10640 520
rect 11332 200 11652 520
rect 12344 200 12664 520
rect 13356 200 13676 520
rect 14368 200 14688 520
rect 15380 200 15700 520
rect 16392 200 16712 520
rect 17404 200 17724 520
rect 18416 200 18736 520
rect 19428 200 19748 520
rect 20440 200 20760 520
rect 21452 200 21772 520
rect 22464 200 22784 520
rect 23476 200 23796 520
rect 24488 200 24808 520
rect 25500 200 25820 520
rect 26512 200 26832 520
rect 27524 200 27844 520
rect 28536 200 28856 520
rect 29548 200 29868 520
rect 30560 200 30880 520
rect 31572 200 31892 520
rect -32184 -520 -31864 -200
rect -31172 -520 -30852 -200
rect -30160 -520 -29840 -200
rect -29148 -520 -28828 -200
rect -28136 -520 -27816 -200
rect -27124 -520 -26804 -200
rect -26112 -520 -25792 -200
rect -25100 -520 -24780 -200
rect -24088 -520 -23768 -200
rect -23076 -520 -22756 -200
rect -22064 -520 -21744 -200
rect -21052 -520 -20732 -200
rect -20040 -520 -19720 -200
rect -19028 -520 -18708 -200
rect -18016 -520 -17696 -200
rect -17004 -520 -16684 -200
rect -15992 -520 -15672 -200
rect -14980 -520 -14660 -200
rect -13968 -520 -13648 -200
rect -12956 -520 -12636 -200
rect -11944 -520 -11624 -200
rect -10932 -520 -10612 -200
rect -9920 -520 -9600 -200
rect -8908 -520 -8588 -200
rect -7896 -520 -7576 -200
rect -6884 -520 -6564 -200
rect -5872 -520 -5552 -200
rect -4860 -520 -4540 -200
rect -3848 -520 -3528 -200
rect -2836 -520 -2516 -200
rect -1824 -520 -1504 -200
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect 1212 -520 1532 -200
rect 2224 -520 2544 -200
rect 3236 -520 3556 -200
rect 4248 -520 4568 -200
rect 5260 -520 5580 -200
rect 6272 -520 6592 -200
rect 7284 -520 7604 -200
rect 8296 -520 8616 -200
rect 9308 -520 9628 -200
rect 10320 -520 10640 -200
rect 11332 -520 11652 -200
rect 12344 -520 12664 -200
rect 13356 -520 13676 -200
rect 14368 -520 14688 -200
rect 15380 -520 15700 -200
rect 16392 -520 16712 -200
rect 17404 -520 17724 -200
rect 18416 -520 18736 -200
rect 19428 -520 19748 -200
rect 20440 -520 20760 -200
rect 21452 -520 21772 -200
rect 22464 -520 22784 -200
rect 23476 -520 23796 -200
rect 24488 -520 24808 -200
rect 25500 -520 25820 -200
rect 26512 -520 26832 -200
rect 27524 -520 27844 -200
rect 28536 -520 28856 -200
rect 29548 -520 29868 -200
rect 30560 -520 30880 -200
rect 31572 -520 31892 -200
rect -32184 -1240 -31864 -920
rect -31172 -1240 -30852 -920
rect -30160 -1240 -29840 -920
rect -29148 -1240 -28828 -920
rect -28136 -1240 -27816 -920
rect -27124 -1240 -26804 -920
rect -26112 -1240 -25792 -920
rect -25100 -1240 -24780 -920
rect -24088 -1240 -23768 -920
rect -23076 -1240 -22756 -920
rect -22064 -1240 -21744 -920
rect -21052 -1240 -20732 -920
rect -20040 -1240 -19720 -920
rect -19028 -1240 -18708 -920
rect -18016 -1240 -17696 -920
rect -17004 -1240 -16684 -920
rect -15992 -1240 -15672 -920
rect -14980 -1240 -14660 -920
rect -13968 -1240 -13648 -920
rect -12956 -1240 -12636 -920
rect -11944 -1240 -11624 -920
rect -10932 -1240 -10612 -920
rect -9920 -1240 -9600 -920
rect -8908 -1240 -8588 -920
rect -7896 -1240 -7576 -920
rect -6884 -1240 -6564 -920
rect -5872 -1240 -5552 -920
rect -4860 -1240 -4540 -920
rect -3848 -1240 -3528 -920
rect -2836 -1240 -2516 -920
rect -1824 -1240 -1504 -920
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect 1212 -1240 1532 -920
rect 2224 -1240 2544 -920
rect 3236 -1240 3556 -920
rect 4248 -1240 4568 -920
rect 5260 -1240 5580 -920
rect 6272 -1240 6592 -920
rect 7284 -1240 7604 -920
rect 8296 -1240 8616 -920
rect 9308 -1240 9628 -920
rect 10320 -1240 10640 -920
rect 11332 -1240 11652 -920
rect 12344 -1240 12664 -920
rect 13356 -1240 13676 -920
rect 14368 -1240 14688 -920
rect 15380 -1240 15700 -920
rect 16392 -1240 16712 -920
rect 17404 -1240 17724 -920
rect 18416 -1240 18736 -920
rect 19428 -1240 19748 -920
rect 20440 -1240 20760 -920
rect 21452 -1240 21772 -920
rect 22464 -1240 22784 -920
rect 23476 -1240 23796 -920
rect 24488 -1240 24808 -920
rect 25500 -1240 25820 -920
rect 26512 -1240 26832 -920
rect 27524 -1240 27844 -920
rect 28536 -1240 28856 -920
rect 29548 -1240 29868 -920
rect 30560 -1240 30880 -920
rect 31572 -1240 31892 -920
rect -32184 -1960 -31864 -1640
rect -31172 -1960 -30852 -1640
rect -30160 -1960 -29840 -1640
rect -29148 -1960 -28828 -1640
rect -28136 -1960 -27816 -1640
rect -27124 -1960 -26804 -1640
rect -26112 -1960 -25792 -1640
rect -25100 -1960 -24780 -1640
rect -24088 -1960 -23768 -1640
rect -23076 -1960 -22756 -1640
rect -22064 -1960 -21744 -1640
rect -21052 -1960 -20732 -1640
rect -20040 -1960 -19720 -1640
rect -19028 -1960 -18708 -1640
rect -18016 -1960 -17696 -1640
rect -17004 -1960 -16684 -1640
rect -15992 -1960 -15672 -1640
rect -14980 -1960 -14660 -1640
rect -13968 -1960 -13648 -1640
rect -12956 -1960 -12636 -1640
rect -11944 -1960 -11624 -1640
rect -10932 -1960 -10612 -1640
rect -9920 -1960 -9600 -1640
rect -8908 -1960 -8588 -1640
rect -7896 -1960 -7576 -1640
rect -6884 -1960 -6564 -1640
rect -5872 -1960 -5552 -1640
rect -4860 -1960 -4540 -1640
rect -3848 -1960 -3528 -1640
rect -2836 -1960 -2516 -1640
rect -1824 -1960 -1504 -1640
rect -812 -1960 -492 -1640
rect 200 -1960 520 -1640
rect 1212 -1960 1532 -1640
rect 2224 -1960 2544 -1640
rect 3236 -1960 3556 -1640
rect 4248 -1960 4568 -1640
rect 5260 -1960 5580 -1640
rect 6272 -1960 6592 -1640
rect 7284 -1960 7604 -1640
rect 8296 -1960 8616 -1640
rect 9308 -1960 9628 -1640
rect 10320 -1960 10640 -1640
rect 11332 -1960 11652 -1640
rect 12344 -1960 12664 -1640
rect 13356 -1960 13676 -1640
rect 14368 -1960 14688 -1640
rect 15380 -1960 15700 -1640
rect 16392 -1960 16712 -1640
rect 17404 -1960 17724 -1640
rect 18416 -1960 18736 -1640
rect 19428 -1960 19748 -1640
rect 20440 -1960 20760 -1640
rect 21452 -1960 21772 -1640
rect 22464 -1960 22784 -1640
rect 23476 -1960 23796 -1640
rect 24488 -1960 24808 -1640
rect 25500 -1960 25820 -1640
rect 26512 -1960 26832 -1640
rect 27524 -1960 27844 -1640
rect 28536 -1960 28856 -1640
rect 29548 -1960 29868 -1640
rect 30560 -1960 30880 -1640
rect 31572 -1960 31892 -1640
rect -32184 -2680 -31864 -2360
rect -31172 -2680 -30852 -2360
rect -30160 -2680 -29840 -2360
rect -29148 -2680 -28828 -2360
rect -28136 -2680 -27816 -2360
rect -27124 -2680 -26804 -2360
rect -26112 -2680 -25792 -2360
rect -25100 -2680 -24780 -2360
rect -24088 -2680 -23768 -2360
rect -23076 -2680 -22756 -2360
rect -22064 -2680 -21744 -2360
rect -21052 -2680 -20732 -2360
rect -20040 -2680 -19720 -2360
rect -19028 -2680 -18708 -2360
rect -18016 -2680 -17696 -2360
rect -17004 -2680 -16684 -2360
rect -15992 -2680 -15672 -2360
rect -14980 -2680 -14660 -2360
rect -13968 -2680 -13648 -2360
rect -12956 -2680 -12636 -2360
rect -11944 -2680 -11624 -2360
rect -10932 -2680 -10612 -2360
rect -9920 -2680 -9600 -2360
rect -8908 -2680 -8588 -2360
rect -7896 -2680 -7576 -2360
rect -6884 -2680 -6564 -2360
rect -5872 -2680 -5552 -2360
rect -4860 -2680 -4540 -2360
rect -3848 -2680 -3528 -2360
rect -2836 -2680 -2516 -2360
rect -1824 -2680 -1504 -2360
rect -812 -2680 -492 -2360
rect 200 -2680 520 -2360
rect 1212 -2680 1532 -2360
rect 2224 -2680 2544 -2360
rect 3236 -2680 3556 -2360
rect 4248 -2680 4568 -2360
rect 5260 -2680 5580 -2360
rect 6272 -2680 6592 -2360
rect 7284 -2680 7604 -2360
rect 8296 -2680 8616 -2360
rect 9308 -2680 9628 -2360
rect 10320 -2680 10640 -2360
rect 11332 -2680 11652 -2360
rect 12344 -2680 12664 -2360
rect 13356 -2680 13676 -2360
rect 14368 -2680 14688 -2360
rect 15380 -2680 15700 -2360
rect 16392 -2680 16712 -2360
rect 17404 -2680 17724 -2360
rect 18416 -2680 18736 -2360
rect 19428 -2680 19748 -2360
rect 20440 -2680 20760 -2360
rect 21452 -2680 21772 -2360
rect 22464 -2680 22784 -2360
rect 23476 -2680 23796 -2360
rect 24488 -2680 24808 -2360
rect 25500 -2680 25820 -2360
rect 26512 -2680 26832 -2360
rect 27524 -2680 27844 -2360
rect 28536 -2680 28856 -2360
rect 29548 -2680 29868 -2360
rect 30560 -2680 30880 -2360
rect 31572 -2680 31892 -2360
rect -32184 -3400 -31864 -3080
rect -31172 -3400 -30852 -3080
rect -30160 -3400 -29840 -3080
rect -29148 -3400 -28828 -3080
rect -28136 -3400 -27816 -3080
rect -27124 -3400 -26804 -3080
rect -26112 -3400 -25792 -3080
rect -25100 -3400 -24780 -3080
rect -24088 -3400 -23768 -3080
rect -23076 -3400 -22756 -3080
rect -22064 -3400 -21744 -3080
rect -21052 -3400 -20732 -3080
rect -20040 -3400 -19720 -3080
rect -19028 -3400 -18708 -3080
rect -18016 -3400 -17696 -3080
rect -17004 -3400 -16684 -3080
rect -15992 -3400 -15672 -3080
rect -14980 -3400 -14660 -3080
rect -13968 -3400 -13648 -3080
rect -12956 -3400 -12636 -3080
rect -11944 -3400 -11624 -3080
rect -10932 -3400 -10612 -3080
rect -9920 -3400 -9600 -3080
rect -8908 -3400 -8588 -3080
rect -7896 -3400 -7576 -3080
rect -6884 -3400 -6564 -3080
rect -5872 -3400 -5552 -3080
rect -4860 -3400 -4540 -3080
rect -3848 -3400 -3528 -3080
rect -2836 -3400 -2516 -3080
rect -1824 -3400 -1504 -3080
rect -812 -3400 -492 -3080
rect 200 -3400 520 -3080
rect 1212 -3400 1532 -3080
rect 2224 -3400 2544 -3080
rect 3236 -3400 3556 -3080
rect 4248 -3400 4568 -3080
rect 5260 -3400 5580 -3080
rect 6272 -3400 6592 -3080
rect 7284 -3400 7604 -3080
rect 8296 -3400 8616 -3080
rect 9308 -3400 9628 -3080
rect 10320 -3400 10640 -3080
rect 11332 -3400 11652 -3080
rect 12344 -3400 12664 -3080
rect 13356 -3400 13676 -3080
rect 14368 -3400 14688 -3080
rect 15380 -3400 15700 -3080
rect 16392 -3400 16712 -3080
rect 17404 -3400 17724 -3080
rect 18416 -3400 18736 -3080
rect 19428 -3400 19748 -3080
rect 20440 -3400 20760 -3080
rect 21452 -3400 21772 -3080
rect 22464 -3400 22784 -3080
rect 23476 -3400 23796 -3080
rect 24488 -3400 24808 -3080
rect 25500 -3400 25820 -3080
rect 26512 -3400 26832 -3080
rect 27524 -3400 27844 -3080
rect 28536 -3400 28856 -3080
rect 29548 -3400 29868 -3080
rect 30560 -3400 30880 -3080
rect 31572 -3400 31892 -3080
rect -32184 -4120 -31864 -3800
rect -31172 -4120 -30852 -3800
rect -30160 -4120 -29840 -3800
rect -29148 -4120 -28828 -3800
rect -28136 -4120 -27816 -3800
rect -27124 -4120 -26804 -3800
rect -26112 -4120 -25792 -3800
rect -25100 -4120 -24780 -3800
rect -24088 -4120 -23768 -3800
rect -23076 -4120 -22756 -3800
rect -22064 -4120 -21744 -3800
rect -21052 -4120 -20732 -3800
rect -20040 -4120 -19720 -3800
rect -19028 -4120 -18708 -3800
rect -18016 -4120 -17696 -3800
rect -17004 -4120 -16684 -3800
rect -15992 -4120 -15672 -3800
rect -14980 -4120 -14660 -3800
rect -13968 -4120 -13648 -3800
rect -12956 -4120 -12636 -3800
rect -11944 -4120 -11624 -3800
rect -10932 -4120 -10612 -3800
rect -9920 -4120 -9600 -3800
rect -8908 -4120 -8588 -3800
rect -7896 -4120 -7576 -3800
rect -6884 -4120 -6564 -3800
rect -5872 -4120 -5552 -3800
rect -4860 -4120 -4540 -3800
rect -3848 -4120 -3528 -3800
rect -2836 -4120 -2516 -3800
rect -1824 -4120 -1504 -3800
rect -812 -4120 -492 -3800
rect 200 -4120 520 -3800
rect 1212 -4120 1532 -3800
rect 2224 -4120 2544 -3800
rect 3236 -4120 3556 -3800
rect 4248 -4120 4568 -3800
rect 5260 -4120 5580 -3800
rect 6272 -4120 6592 -3800
rect 7284 -4120 7604 -3800
rect 8296 -4120 8616 -3800
rect 9308 -4120 9628 -3800
rect 10320 -4120 10640 -3800
rect 11332 -4120 11652 -3800
rect 12344 -4120 12664 -3800
rect 13356 -4120 13676 -3800
rect 14368 -4120 14688 -3800
rect 15380 -4120 15700 -3800
rect 16392 -4120 16712 -3800
rect 17404 -4120 17724 -3800
rect 18416 -4120 18736 -3800
rect 19428 -4120 19748 -3800
rect 20440 -4120 20760 -3800
rect 21452 -4120 21772 -3800
rect 22464 -4120 22784 -3800
rect 23476 -4120 23796 -3800
rect 24488 -4120 24808 -3800
rect 25500 -4120 25820 -3800
rect 26512 -4120 26832 -3800
rect 27524 -4120 27844 -3800
rect 28536 -4120 28856 -3800
rect 29548 -4120 29868 -3800
rect 30560 -4120 30880 -3800
rect 31572 -4120 31892 -3800
rect -32184 -4840 -31864 -4520
rect -31172 -4840 -30852 -4520
rect -30160 -4840 -29840 -4520
rect -29148 -4840 -28828 -4520
rect -28136 -4840 -27816 -4520
rect -27124 -4840 -26804 -4520
rect -26112 -4840 -25792 -4520
rect -25100 -4840 -24780 -4520
rect -24088 -4840 -23768 -4520
rect -23076 -4840 -22756 -4520
rect -22064 -4840 -21744 -4520
rect -21052 -4840 -20732 -4520
rect -20040 -4840 -19720 -4520
rect -19028 -4840 -18708 -4520
rect -18016 -4840 -17696 -4520
rect -17004 -4840 -16684 -4520
rect -15992 -4840 -15672 -4520
rect -14980 -4840 -14660 -4520
rect -13968 -4840 -13648 -4520
rect -12956 -4840 -12636 -4520
rect -11944 -4840 -11624 -4520
rect -10932 -4840 -10612 -4520
rect -9920 -4840 -9600 -4520
rect -8908 -4840 -8588 -4520
rect -7896 -4840 -7576 -4520
rect -6884 -4840 -6564 -4520
rect -5872 -4840 -5552 -4520
rect -4860 -4840 -4540 -4520
rect -3848 -4840 -3528 -4520
rect -2836 -4840 -2516 -4520
rect -1824 -4840 -1504 -4520
rect -812 -4840 -492 -4520
rect 200 -4840 520 -4520
rect 1212 -4840 1532 -4520
rect 2224 -4840 2544 -4520
rect 3236 -4840 3556 -4520
rect 4248 -4840 4568 -4520
rect 5260 -4840 5580 -4520
rect 6272 -4840 6592 -4520
rect 7284 -4840 7604 -4520
rect 8296 -4840 8616 -4520
rect 9308 -4840 9628 -4520
rect 10320 -4840 10640 -4520
rect 11332 -4840 11652 -4520
rect 12344 -4840 12664 -4520
rect 13356 -4840 13676 -4520
rect 14368 -4840 14688 -4520
rect 15380 -4840 15700 -4520
rect 16392 -4840 16712 -4520
rect 17404 -4840 17724 -4520
rect 18416 -4840 18736 -4520
rect 19428 -4840 19748 -4520
rect 20440 -4840 20760 -4520
rect 21452 -4840 21772 -4520
rect 22464 -4840 22784 -4520
rect 23476 -4840 23796 -4520
rect 24488 -4840 24808 -4520
rect 25500 -4840 25820 -4520
rect 26512 -4840 26832 -4520
rect 27524 -4840 27844 -4520
rect 28536 -4840 28856 -4520
rect 29548 -4840 29868 -4520
rect 30560 -4840 30880 -4520
rect 31572 -4840 31892 -4520
rect -32184 -5560 -31864 -5240
rect -31172 -5560 -30852 -5240
rect -30160 -5560 -29840 -5240
rect -29148 -5560 -28828 -5240
rect -28136 -5560 -27816 -5240
rect -27124 -5560 -26804 -5240
rect -26112 -5560 -25792 -5240
rect -25100 -5560 -24780 -5240
rect -24088 -5560 -23768 -5240
rect -23076 -5560 -22756 -5240
rect -22064 -5560 -21744 -5240
rect -21052 -5560 -20732 -5240
rect -20040 -5560 -19720 -5240
rect -19028 -5560 -18708 -5240
rect -18016 -5560 -17696 -5240
rect -17004 -5560 -16684 -5240
rect -15992 -5560 -15672 -5240
rect -14980 -5560 -14660 -5240
rect -13968 -5560 -13648 -5240
rect -12956 -5560 -12636 -5240
rect -11944 -5560 -11624 -5240
rect -10932 -5560 -10612 -5240
rect -9920 -5560 -9600 -5240
rect -8908 -5560 -8588 -5240
rect -7896 -5560 -7576 -5240
rect -6884 -5560 -6564 -5240
rect -5872 -5560 -5552 -5240
rect -4860 -5560 -4540 -5240
rect -3848 -5560 -3528 -5240
rect -2836 -5560 -2516 -5240
rect -1824 -5560 -1504 -5240
rect -812 -5560 -492 -5240
rect 200 -5560 520 -5240
rect 1212 -5560 1532 -5240
rect 2224 -5560 2544 -5240
rect 3236 -5560 3556 -5240
rect 4248 -5560 4568 -5240
rect 5260 -5560 5580 -5240
rect 6272 -5560 6592 -5240
rect 7284 -5560 7604 -5240
rect 8296 -5560 8616 -5240
rect 9308 -5560 9628 -5240
rect 10320 -5560 10640 -5240
rect 11332 -5560 11652 -5240
rect 12344 -5560 12664 -5240
rect 13356 -5560 13676 -5240
rect 14368 -5560 14688 -5240
rect 15380 -5560 15700 -5240
rect 16392 -5560 16712 -5240
rect 17404 -5560 17724 -5240
rect 18416 -5560 18736 -5240
rect 19428 -5560 19748 -5240
rect 20440 -5560 20760 -5240
rect 21452 -5560 21772 -5240
rect 22464 -5560 22784 -5240
rect 23476 -5560 23796 -5240
rect 24488 -5560 24808 -5240
rect 25500 -5560 25820 -5240
rect 26512 -5560 26832 -5240
rect 27524 -5560 27844 -5240
rect 28536 -5560 28856 -5240
rect 29548 -5560 29868 -5240
rect 30560 -5560 30880 -5240
rect 31572 -5560 31892 -5240
<< metal4 >>
rect -32076 5561 -31972 5760
rect -31596 5612 -31492 5760
rect -32185 5560 -31863 5561
rect -32185 5240 -32184 5560
rect -31864 5240 -31863 5560
rect -32185 5239 -31863 5240
rect -32076 4841 -31972 5239
rect -31596 5188 -31576 5612
rect -31512 5188 -31492 5612
rect -31064 5561 -30960 5760
rect -30584 5612 -30480 5760
rect -31173 5560 -30851 5561
rect -31173 5240 -31172 5560
rect -30852 5240 -30851 5560
rect -31173 5239 -30851 5240
rect -31596 4892 -31492 5188
rect -32185 4840 -31863 4841
rect -32185 4520 -32184 4840
rect -31864 4520 -31863 4840
rect -32185 4519 -31863 4520
rect -32076 4121 -31972 4519
rect -31596 4468 -31576 4892
rect -31512 4468 -31492 4892
rect -31064 4841 -30960 5239
rect -30584 5188 -30564 5612
rect -30500 5188 -30480 5612
rect -30052 5561 -29948 5760
rect -29572 5612 -29468 5760
rect -30161 5560 -29839 5561
rect -30161 5240 -30160 5560
rect -29840 5240 -29839 5560
rect -30161 5239 -29839 5240
rect -30584 4892 -30480 5188
rect -31173 4840 -30851 4841
rect -31173 4520 -31172 4840
rect -30852 4520 -30851 4840
rect -31173 4519 -30851 4520
rect -31596 4172 -31492 4468
rect -32185 4120 -31863 4121
rect -32185 3800 -32184 4120
rect -31864 3800 -31863 4120
rect -32185 3799 -31863 3800
rect -32076 3401 -31972 3799
rect -31596 3748 -31576 4172
rect -31512 3748 -31492 4172
rect -31064 4121 -30960 4519
rect -30584 4468 -30564 4892
rect -30500 4468 -30480 4892
rect -30052 4841 -29948 5239
rect -29572 5188 -29552 5612
rect -29488 5188 -29468 5612
rect -29040 5561 -28936 5760
rect -28560 5612 -28456 5760
rect -29149 5560 -28827 5561
rect -29149 5240 -29148 5560
rect -28828 5240 -28827 5560
rect -29149 5239 -28827 5240
rect -29572 4892 -29468 5188
rect -30161 4840 -29839 4841
rect -30161 4520 -30160 4840
rect -29840 4520 -29839 4840
rect -30161 4519 -29839 4520
rect -30584 4172 -30480 4468
rect -31173 4120 -30851 4121
rect -31173 3800 -31172 4120
rect -30852 3800 -30851 4120
rect -31173 3799 -30851 3800
rect -31596 3452 -31492 3748
rect -32185 3400 -31863 3401
rect -32185 3080 -32184 3400
rect -31864 3080 -31863 3400
rect -32185 3079 -31863 3080
rect -32076 2681 -31972 3079
rect -31596 3028 -31576 3452
rect -31512 3028 -31492 3452
rect -31064 3401 -30960 3799
rect -30584 3748 -30564 4172
rect -30500 3748 -30480 4172
rect -30052 4121 -29948 4519
rect -29572 4468 -29552 4892
rect -29488 4468 -29468 4892
rect -29040 4841 -28936 5239
rect -28560 5188 -28540 5612
rect -28476 5188 -28456 5612
rect -28028 5561 -27924 5760
rect -27548 5612 -27444 5760
rect -28137 5560 -27815 5561
rect -28137 5240 -28136 5560
rect -27816 5240 -27815 5560
rect -28137 5239 -27815 5240
rect -28560 4892 -28456 5188
rect -29149 4840 -28827 4841
rect -29149 4520 -29148 4840
rect -28828 4520 -28827 4840
rect -29149 4519 -28827 4520
rect -29572 4172 -29468 4468
rect -30161 4120 -29839 4121
rect -30161 3800 -30160 4120
rect -29840 3800 -29839 4120
rect -30161 3799 -29839 3800
rect -30584 3452 -30480 3748
rect -31173 3400 -30851 3401
rect -31173 3080 -31172 3400
rect -30852 3080 -30851 3400
rect -31173 3079 -30851 3080
rect -31596 2732 -31492 3028
rect -32185 2680 -31863 2681
rect -32185 2360 -32184 2680
rect -31864 2360 -31863 2680
rect -32185 2359 -31863 2360
rect -32076 1961 -31972 2359
rect -31596 2308 -31576 2732
rect -31512 2308 -31492 2732
rect -31064 2681 -30960 3079
rect -30584 3028 -30564 3452
rect -30500 3028 -30480 3452
rect -30052 3401 -29948 3799
rect -29572 3748 -29552 4172
rect -29488 3748 -29468 4172
rect -29040 4121 -28936 4519
rect -28560 4468 -28540 4892
rect -28476 4468 -28456 4892
rect -28028 4841 -27924 5239
rect -27548 5188 -27528 5612
rect -27464 5188 -27444 5612
rect -27016 5561 -26912 5760
rect -26536 5612 -26432 5760
rect -27125 5560 -26803 5561
rect -27125 5240 -27124 5560
rect -26804 5240 -26803 5560
rect -27125 5239 -26803 5240
rect -27548 4892 -27444 5188
rect -28137 4840 -27815 4841
rect -28137 4520 -28136 4840
rect -27816 4520 -27815 4840
rect -28137 4519 -27815 4520
rect -28560 4172 -28456 4468
rect -29149 4120 -28827 4121
rect -29149 3800 -29148 4120
rect -28828 3800 -28827 4120
rect -29149 3799 -28827 3800
rect -29572 3452 -29468 3748
rect -30161 3400 -29839 3401
rect -30161 3080 -30160 3400
rect -29840 3080 -29839 3400
rect -30161 3079 -29839 3080
rect -30584 2732 -30480 3028
rect -31173 2680 -30851 2681
rect -31173 2360 -31172 2680
rect -30852 2360 -30851 2680
rect -31173 2359 -30851 2360
rect -31596 2012 -31492 2308
rect -32185 1960 -31863 1961
rect -32185 1640 -32184 1960
rect -31864 1640 -31863 1960
rect -32185 1639 -31863 1640
rect -32076 1241 -31972 1639
rect -31596 1588 -31576 2012
rect -31512 1588 -31492 2012
rect -31064 1961 -30960 2359
rect -30584 2308 -30564 2732
rect -30500 2308 -30480 2732
rect -30052 2681 -29948 3079
rect -29572 3028 -29552 3452
rect -29488 3028 -29468 3452
rect -29040 3401 -28936 3799
rect -28560 3748 -28540 4172
rect -28476 3748 -28456 4172
rect -28028 4121 -27924 4519
rect -27548 4468 -27528 4892
rect -27464 4468 -27444 4892
rect -27016 4841 -26912 5239
rect -26536 5188 -26516 5612
rect -26452 5188 -26432 5612
rect -26004 5561 -25900 5760
rect -25524 5612 -25420 5760
rect -26113 5560 -25791 5561
rect -26113 5240 -26112 5560
rect -25792 5240 -25791 5560
rect -26113 5239 -25791 5240
rect -26536 4892 -26432 5188
rect -27125 4840 -26803 4841
rect -27125 4520 -27124 4840
rect -26804 4520 -26803 4840
rect -27125 4519 -26803 4520
rect -27548 4172 -27444 4468
rect -28137 4120 -27815 4121
rect -28137 3800 -28136 4120
rect -27816 3800 -27815 4120
rect -28137 3799 -27815 3800
rect -28560 3452 -28456 3748
rect -29149 3400 -28827 3401
rect -29149 3080 -29148 3400
rect -28828 3080 -28827 3400
rect -29149 3079 -28827 3080
rect -29572 2732 -29468 3028
rect -30161 2680 -29839 2681
rect -30161 2360 -30160 2680
rect -29840 2360 -29839 2680
rect -30161 2359 -29839 2360
rect -30584 2012 -30480 2308
rect -31173 1960 -30851 1961
rect -31173 1640 -31172 1960
rect -30852 1640 -30851 1960
rect -31173 1639 -30851 1640
rect -31596 1292 -31492 1588
rect -32185 1240 -31863 1241
rect -32185 920 -32184 1240
rect -31864 920 -31863 1240
rect -32185 919 -31863 920
rect -32076 521 -31972 919
rect -31596 868 -31576 1292
rect -31512 868 -31492 1292
rect -31064 1241 -30960 1639
rect -30584 1588 -30564 2012
rect -30500 1588 -30480 2012
rect -30052 1961 -29948 2359
rect -29572 2308 -29552 2732
rect -29488 2308 -29468 2732
rect -29040 2681 -28936 3079
rect -28560 3028 -28540 3452
rect -28476 3028 -28456 3452
rect -28028 3401 -27924 3799
rect -27548 3748 -27528 4172
rect -27464 3748 -27444 4172
rect -27016 4121 -26912 4519
rect -26536 4468 -26516 4892
rect -26452 4468 -26432 4892
rect -26004 4841 -25900 5239
rect -25524 5188 -25504 5612
rect -25440 5188 -25420 5612
rect -24992 5561 -24888 5760
rect -24512 5612 -24408 5760
rect -25101 5560 -24779 5561
rect -25101 5240 -25100 5560
rect -24780 5240 -24779 5560
rect -25101 5239 -24779 5240
rect -25524 4892 -25420 5188
rect -26113 4840 -25791 4841
rect -26113 4520 -26112 4840
rect -25792 4520 -25791 4840
rect -26113 4519 -25791 4520
rect -26536 4172 -26432 4468
rect -27125 4120 -26803 4121
rect -27125 3800 -27124 4120
rect -26804 3800 -26803 4120
rect -27125 3799 -26803 3800
rect -27548 3452 -27444 3748
rect -28137 3400 -27815 3401
rect -28137 3080 -28136 3400
rect -27816 3080 -27815 3400
rect -28137 3079 -27815 3080
rect -28560 2732 -28456 3028
rect -29149 2680 -28827 2681
rect -29149 2360 -29148 2680
rect -28828 2360 -28827 2680
rect -29149 2359 -28827 2360
rect -29572 2012 -29468 2308
rect -30161 1960 -29839 1961
rect -30161 1640 -30160 1960
rect -29840 1640 -29839 1960
rect -30161 1639 -29839 1640
rect -30584 1292 -30480 1588
rect -31173 1240 -30851 1241
rect -31173 920 -31172 1240
rect -30852 920 -30851 1240
rect -31173 919 -30851 920
rect -31596 572 -31492 868
rect -32185 520 -31863 521
rect -32185 200 -32184 520
rect -31864 200 -31863 520
rect -32185 199 -31863 200
rect -32076 -199 -31972 199
rect -31596 148 -31576 572
rect -31512 148 -31492 572
rect -31064 521 -30960 919
rect -30584 868 -30564 1292
rect -30500 868 -30480 1292
rect -30052 1241 -29948 1639
rect -29572 1588 -29552 2012
rect -29488 1588 -29468 2012
rect -29040 1961 -28936 2359
rect -28560 2308 -28540 2732
rect -28476 2308 -28456 2732
rect -28028 2681 -27924 3079
rect -27548 3028 -27528 3452
rect -27464 3028 -27444 3452
rect -27016 3401 -26912 3799
rect -26536 3748 -26516 4172
rect -26452 3748 -26432 4172
rect -26004 4121 -25900 4519
rect -25524 4468 -25504 4892
rect -25440 4468 -25420 4892
rect -24992 4841 -24888 5239
rect -24512 5188 -24492 5612
rect -24428 5188 -24408 5612
rect -23980 5561 -23876 5760
rect -23500 5612 -23396 5760
rect -24089 5560 -23767 5561
rect -24089 5240 -24088 5560
rect -23768 5240 -23767 5560
rect -24089 5239 -23767 5240
rect -24512 4892 -24408 5188
rect -25101 4840 -24779 4841
rect -25101 4520 -25100 4840
rect -24780 4520 -24779 4840
rect -25101 4519 -24779 4520
rect -25524 4172 -25420 4468
rect -26113 4120 -25791 4121
rect -26113 3800 -26112 4120
rect -25792 3800 -25791 4120
rect -26113 3799 -25791 3800
rect -26536 3452 -26432 3748
rect -27125 3400 -26803 3401
rect -27125 3080 -27124 3400
rect -26804 3080 -26803 3400
rect -27125 3079 -26803 3080
rect -27548 2732 -27444 3028
rect -28137 2680 -27815 2681
rect -28137 2360 -28136 2680
rect -27816 2360 -27815 2680
rect -28137 2359 -27815 2360
rect -28560 2012 -28456 2308
rect -29149 1960 -28827 1961
rect -29149 1640 -29148 1960
rect -28828 1640 -28827 1960
rect -29149 1639 -28827 1640
rect -29572 1292 -29468 1588
rect -30161 1240 -29839 1241
rect -30161 920 -30160 1240
rect -29840 920 -29839 1240
rect -30161 919 -29839 920
rect -30584 572 -30480 868
rect -31173 520 -30851 521
rect -31173 200 -31172 520
rect -30852 200 -30851 520
rect -31173 199 -30851 200
rect -31596 -148 -31492 148
rect -32185 -200 -31863 -199
rect -32185 -520 -32184 -200
rect -31864 -520 -31863 -200
rect -32185 -521 -31863 -520
rect -32076 -919 -31972 -521
rect -31596 -572 -31576 -148
rect -31512 -572 -31492 -148
rect -31064 -199 -30960 199
rect -30584 148 -30564 572
rect -30500 148 -30480 572
rect -30052 521 -29948 919
rect -29572 868 -29552 1292
rect -29488 868 -29468 1292
rect -29040 1241 -28936 1639
rect -28560 1588 -28540 2012
rect -28476 1588 -28456 2012
rect -28028 1961 -27924 2359
rect -27548 2308 -27528 2732
rect -27464 2308 -27444 2732
rect -27016 2681 -26912 3079
rect -26536 3028 -26516 3452
rect -26452 3028 -26432 3452
rect -26004 3401 -25900 3799
rect -25524 3748 -25504 4172
rect -25440 3748 -25420 4172
rect -24992 4121 -24888 4519
rect -24512 4468 -24492 4892
rect -24428 4468 -24408 4892
rect -23980 4841 -23876 5239
rect -23500 5188 -23480 5612
rect -23416 5188 -23396 5612
rect -22968 5561 -22864 5760
rect -22488 5612 -22384 5760
rect -23077 5560 -22755 5561
rect -23077 5240 -23076 5560
rect -22756 5240 -22755 5560
rect -23077 5239 -22755 5240
rect -23500 4892 -23396 5188
rect -24089 4840 -23767 4841
rect -24089 4520 -24088 4840
rect -23768 4520 -23767 4840
rect -24089 4519 -23767 4520
rect -24512 4172 -24408 4468
rect -25101 4120 -24779 4121
rect -25101 3800 -25100 4120
rect -24780 3800 -24779 4120
rect -25101 3799 -24779 3800
rect -25524 3452 -25420 3748
rect -26113 3400 -25791 3401
rect -26113 3080 -26112 3400
rect -25792 3080 -25791 3400
rect -26113 3079 -25791 3080
rect -26536 2732 -26432 3028
rect -27125 2680 -26803 2681
rect -27125 2360 -27124 2680
rect -26804 2360 -26803 2680
rect -27125 2359 -26803 2360
rect -27548 2012 -27444 2308
rect -28137 1960 -27815 1961
rect -28137 1640 -28136 1960
rect -27816 1640 -27815 1960
rect -28137 1639 -27815 1640
rect -28560 1292 -28456 1588
rect -29149 1240 -28827 1241
rect -29149 920 -29148 1240
rect -28828 920 -28827 1240
rect -29149 919 -28827 920
rect -29572 572 -29468 868
rect -30161 520 -29839 521
rect -30161 200 -30160 520
rect -29840 200 -29839 520
rect -30161 199 -29839 200
rect -30584 -148 -30480 148
rect -31173 -200 -30851 -199
rect -31173 -520 -31172 -200
rect -30852 -520 -30851 -200
rect -31173 -521 -30851 -520
rect -31596 -868 -31492 -572
rect -32185 -920 -31863 -919
rect -32185 -1240 -32184 -920
rect -31864 -1240 -31863 -920
rect -32185 -1241 -31863 -1240
rect -32076 -1639 -31972 -1241
rect -31596 -1292 -31576 -868
rect -31512 -1292 -31492 -868
rect -31064 -919 -30960 -521
rect -30584 -572 -30564 -148
rect -30500 -572 -30480 -148
rect -30052 -199 -29948 199
rect -29572 148 -29552 572
rect -29488 148 -29468 572
rect -29040 521 -28936 919
rect -28560 868 -28540 1292
rect -28476 868 -28456 1292
rect -28028 1241 -27924 1639
rect -27548 1588 -27528 2012
rect -27464 1588 -27444 2012
rect -27016 1961 -26912 2359
rect -26536 2308 -26516 2732
rect -26452 2308 -26432 2732
rect -26004 2681 -25900 3079
rect -25524 3028 -25504 3452
rect -25440 3028 -25420 3452
rect -24992 3401 -24888 3799
rect -24512 3748 -24492 4172
rect -24428 3748 -24408 4172
rect -23980 4121 -23876 4519
rect -23500 4468 -23480 4892
rect -23416 4468 -23396 4892
rect -22968 4841 -22864 5239
rect -22488 5188 -22468 5612
rect -22404 5188 -22384 5612
rect -21956 5561 -21852 5760
rect -21476 5612 -21372 5760
rect -22065 5560 -21743 5561
rect -22065 5240 -22064 5560
rect -21744 5240 -21743 5560
rect -22065 5239 -21743 5240
rect -22488 4892 -22384 5188
rect -23077 4840 -22755 4841
rect -23077 4520 -23076 4840
rect -22756 4520 -22755 4840
rect -23077 4519 -22755 4520
rect -23500 4172 -23396 4468
rect -24089 4120 -23767 4121
rect -24089 3800 -24088 4120
rect -23768 3800 -23767 4120
rect -24089 3799 -23767 3800
rect -24512 3452 -24408 3748
rect -25101 3400 -24779 3401
rect -25101 3080 -25100 3400
rect -24780 3080 -24779 3400
rect -25101 3079 -24779 3080
rect -25524 2732 -25420 3028
rect -26113 2680 -25791 2681
rect -26113 2360 -26112 2680
rect -25792 2360 -25791 2680
rect -26113 2359 -25791 2360
rect -26536 2012 -26432 2308
rect -27125 1960 -26803 1961
rect -27125 1640 -27124 1960
rect -26804 1640 -26803 1960
rect -27125 1639 -26803 1640
rect -27548 1292 -27444 1588
rect -28137 1240 -27815 1241
rect -28137 920 -28136 1240
rect -27816 920 -27815 1240
rect -28137 919 -27815 920
rect -28560 572 -28456 868
rect -29149 520 -28827 521
rect -29149 200 -29148 520
rect -28828 200 -28827 520
rect -29149 199 -28827 200
rect -29572 -148 -29468 148
rect -30161 -200 -29839 -199
rect -30161 -520 -30160 -200
rect -29840 -520 -29839 -200
rect -30161 -521 -29839 -520
rect -30584 -868 -30480 -572
rect -31173 -920 -30851 -919
rect -31173 -1240 -31172 -920
rect -30852 -1240 -30851 -920
rect -31173 -1241 -30851 -1240
rect -31596 -1588 -31492 -1292
rect -32185 -1640 -31863 -1639
rect -32185 -1960 -32184 -1640
rect -31864 -1960 -31863 -1640
rect -32185 -1961 -31863 -1960
rect -32076 -2359 -31972 -1961
rect -31596 -2012 -31576 -1588
rect -31512 -2012 -31492 -1588
rect -31064 -1639 -30960 -1241
rect -30584 -1292 -30564 -868
rect -30500 -1292 -30480 -868
rect -30052 -919 -29948 -521
rect -29572 -572 -29552 -148
rect -29488 -572 -29468 -148
rect -29040 -199 -28936 199
rect -28560 148 -28540 572
rect -28476 148 -28456 572
rect -28028 521 -27924 919
rect -27548 868 -27528 1292
rect -27464 868 -27444 1292
rect -27016 1241 -26912 1639
rect -26536 1588 -26516 2012
rect -26452 1588 -26432 2012
rect -26004 1961 -25900 2359
rect -25524 2308 -25504 2732
rect -25440 2308 -25420 2732
rect -24992 2681 -24888 3079
rect -24512 3028 -24492 3452
rect -24428 3028 -24408 3452
rect -23980 3401 -23876 3799
rect -23500 3748 -23480 4172
rect -23416 3748 -23396 4172
rect -22968 4121 -22864 4519
rect -22488 4468 -22468 4892
rect -22404 4468 -22384 4892
rect -21956 4841 -21852 5239
rect -21476 5188 -21456 5612
rect -21392 5188 -21372 5612
rect -20944 5561 -20840 5760
rect -20464 5612 -20360 5760
rect -21053 5560 -20731 5561
rect -21053 5240 -21052 5560
rect -20732 5240 -20731 5560
rect -21053 5239 -20731 5240
rect -21476 4892 -21372 5188
rect -22065 4840 -21743 4841
rect -22065 4520 -22064 4840
rect -21744 4520 -21743 4840
rect -22065 4519 -21743 4520
rect -22488 4172 -22384 4468
rect -23077 4120 -22755 4121
rect -23077 3800 -23076 4120
rect -22756 3800 -22755 4120
rect -23077 3799 -22755 3800
rect -23500 3452 -23396 3748
rect -24089 3400 -23767 3401
rect -24089 3080 -24088 3400
rect -23768 3080 -23767 3400
rect -24089 3079 -23767 3080
rect -24512 2732 -24408 3028
rect -25101 2680 -24779 2681
rect -25101 2360 -25100 2680
rect -24780 2360 -24779 2680
rect -25101 2359 -24779 2360
rect -25524 2012 -25420 2308
rect -26113 1960 -25791 1961
rect -26113 1640 -26112 1960
rect -25792 1640 -25791 1960
rect -26113 1639 -25791 1640
rect -26536 1292 -26432 1588
rect -27125 1240 -26803 1241
rect -27125 920 -27124 1240
rect -26804 920 -26803 1240
rect -27125 919 -26803 920
rect -27548 572 -27444 868
rect -28137 520 -27815 521
rect -28137 200 -28136 520
rect -27816 200 -27815 520
rect -28137 199 -27815 200
rect -28560 -148 -28456 148
rect -29149 -200 -28827 -199
rect -29149 -520 -29148 -200
rect -28828 -520 -28827 -200
rect -29149 -521 -28827 -520
rect -29572 -868 -29468 -572
rect -30161 -920 -29839 -919
rect -30161 -1240 -30160 -920
rect -29840 -1240 -29839 -920
rect -30161 -1241 -29839 -1240
rect -30584 -1588 -30480 -1292
rect -31173 -1640 -30851 -1639
rect -31173 -1960 -31172 -1640
rect -30852 -1960 -30851 -1640
rect -31173 -1961 -30851 -1960
rect -31596 -2308 -31492 -2012
rect -32185 -2360 -31863 -2359
rect -32185 -2680 -32184 -2360
rect -31864 -2680 -31863 -2360
rect -32185 -2681 -31863 -2680
rect -32076 -3079 -31972 -2681
rect -31596 -2732 -31576 -2308
rect -31512 -2732 -31492 -2308
rect -31064 -2359 -30960 -1961
rect -30584 -2012 -30564 -1588
rect -30500 -2012 -30480 -1588
rect -30052 -1639 -29948 -1241
rect -29572 -1292 -29552 -868
rect -29488 -1292 -29468 -868
rect -29040 -919 -28936 -521
rect -28560 -572 -28540 -148
rect -28476 -572 -28456 -148
rect -28028 -199 -27924 199
rect -27548 148 -27528 572
rect -27464 148 -27444 572
rect -27016 521 -26912 919
rect -26536 868 -26516 1292
rect -26452 868 -26432 1292
rect -26004 1241 -25900 1639
rect -25524 1588 -25504 2012
rect -25440 1588 -25420 2012
rect -24992 1961 -24888 2359
rect -24512 2308 -24492 2732
rect -24428 2308 -24408 2732
rect -23980 2681 -23876 3079
rect -23500 3028 -23480 3452
rect -23416 3028 -23396 3452
rect -22968 3401 -22864 3799
rect -22488 3748 -22468 4172
rect -22404 3748 -22384 4172
rect -21956 4121 -21852 4519
rect -21476 4468 -21456 4892
rect -21392 4468 -21372 4892
rect -20944 4841 -20840 5239
rect -20464 5188 -20444 5612
rect -20380 5188 -20360 5612
rect -19932 5561 -19828 5760
rect -19452 5612 -19348 5760
rect -20041 5560 -19719 5561
rect -20041 5240 -20040 5560
rect -19720 5240 -19719 5560
rect -20041 5239 -19719 5240
rect -20464 4892 -20360 5188
rect -21053 4840 -20731 4841
rect -21053 4520 -21052 4840
rect -20732 4520 -20731 4840
rect -21053 4519 -20731 4520
rect -21476 4172 -21372 4468
rect -22065 4120 -21743 4121
rect -22065 3800 -22064 4120
rect -21744 3800 -21743 4120
rect -22065 3799 -21743 3800
rect -22488 3452 -22384 3748
rect -23077 3400 -22755 3401
rect -23077 3080 -23076 3400
rect -22756 3080 -22755 3400
rect -23077 3079 -22755 3080
rect -23500 2732 -23396 3028
rect -24089 2680 -23767 2681
rect -24089 2360 -24088 2680
rect -23768 2360 -23767 2680
rect -24089 2359 -23767 2360
rect -24512 2012 -24408 2308
rect -25101 1960 -24779 1961
rect -25101 1640 -25100 1960
rect -24780 1640 -24779 1960
rect -25101 1639 -24779 1640
rect -25524 1292 -25420 1588
rect -26113 1240 -25791 1241
rect -26113 920 -26112 1240
rect -25792 920 -25791 1240
rect -26113 919 -25791 920
rect -26536 572 -26432 868
rect -27125 520 -26803 521
rect -27125 200 -27124 520
rect -26804 200 -26803 520
rect -27125 199 -26803 200
rect -27548 -148 -27444 148
rect -28137 -200 -27815 -199
rect -28137 -520 -28136 -200
rect -27816 -520 -27815 -200
rect -28137 -521 -27815 -520
rect -28560 -868 -28456 -572
rect -29149 -920 -28827 -919
rect -29149 -1240 -29148 -920
rect -28828 -1240 -28827 -920
rect -29149 -1241 -28827 -1240
rect -29572 -1588 -29468 -1292
rect -30161 -1640 -29839 -1639
rect -30161 -1960 -30160 -1640
rect -29840 -1960 -29839 -1640
rect -30161 -1961 -29839 -1960
rect -30584 -2308 -30480 -2012
rect -31173 -2360 -30851 -2359
rect -31173 -2680 -31172 -2360
rect -30852 -2680 -30851 -2360
rect -31173 -2681 -30851 -2680
rect -31596 -3028 -31492 -2732
rect -32185 -3080 -31863 -3079
rect -32185 -3400 -32184 -3080
rect -31864 -3400 -31863 -3080
rect -32185 -3401 -31863 -3400
rect -32076 -3799 -31972 -3401
rect -31596 -3452 -31576 -3028
rect -31512 -3452 -31492 -3028
rect -31064 -3079 -30960 -2681
rect -30584 -2732 -30564 -2308
rect -30500 -2732 -30480 -2308
rect -30052 -2359 -29948 -1961
rect -29572 -2012 -29552 -1588
rect -29488 -2012 -29468 -1588
rect -29040 -1639 -28936 -1241
rect -28560 -1292 -28540 -868
rect -28476 -1292 -28456 -868
rect -28028 -919 -27924 -521
rect -27548 -572 -27528 -148
rect -27464 -572 -27444 -148
rect -27016 -199 -26912 199
rect -26536 148 -26516 572
rect -26452 148 -26432 572
rect -26004 521 -25900 919
rect -25524 868 -25504 1292
rect -25440 868 -25420 1292
rect -24992 1241 -24888 1639
rect -24512 1588 -24492 2012
rect -24428 1588 -24408 2012
rect -23980 1961 -23876 2359
rect -23500 2308 -23480 2732
rect -23416 2308 -23396 2732
rect -22968 2681 -22864 3079
rect -22488 3028 -22468 3452
rect -22404 3028 -22384 3452
rect -21956 3401 -21852 3799
rect -21476 3748 -21456 4172
rect -21392 3748 -21372 4172
rect -20944 4121 -20840 4519
rect -20464 4468 -20444 4892
rect -20380 4468 -20360 4892
rect -19932 4841 -19828 5239
rect -19452 5188 -19432 5612
rect -19368 5188 -19348 5612
rect -18920 5561 -18816 5760
rect -18440 5612 -18336 5760
rect -19029 5560 -18707 5561
rect -19029 5240 -19028 5560
rect -18708 5240 -18707 5560
rect -19029 5239 -18707 5240
rect -19452 4892 -19348 5188
rect -20041 4840 -19719 4841
rect -20041 4520 -20040 4840
rect -19720 4520 -19719 4840
rect -20041 4519 -19719 4520
rect -20464 4172 -20360 4468
rect -21053 4120 -20731 4121
rect -21053 3800 -21052 4120
rect -20732 3800 -20731 4120
rect -21053 3799 -20731 3800
rect -21476 3452 -21372 3748
rect -22065 3400 -21743 3401
rect -22065 3080 -22064 3400
rect -21744 3080 -21743 3400
rect -22065 3079 -21743 3080
rect -22488 2732 -22384 3028
rect -23077 2680 -22755 2681
rect -23077 2360 -23076 2680
rect -22756 2360 -22755 2680
rect -23077 2359 -22755 2360
rect -23500 2012 -23396 2308
rect -24089 1960 -23767 1961
rect -24089 1640 -24088 1960
rect -23768 1640 -23767 1960
rect -24089 1639 -23767 1640
rect -24512 1292 -24408 1588
rect -25101 1240 -24779 1241
rect -25101 920 -25100 1240
rect -24780 920 -24779 1240
rect -25101 919 -24779 920
rect -25524 572 -25420 868
rect -26113 520 -25791 521
rect -26113 200 -26112 520
rect -25792 200 -25791 520
rect -26113 199 -25791 200
rect -26536 -148 -26432 148
rect -27125 -200 -26803 -199
rect -27125 -520 -27124 -200
rect -26804 -520 -26803 -200
rect -27125 -521 -26803 -520
rect -27548 -868 -27444 -572
rect -28137 -920 -27815 -919
rect -28137 -1240 -28136 -920
rect -27816 -1240 -27815 -920
rect -28137 -1241 -27815 -1240
rect -28560 -1588 -28456 -1292
rect -29149 -1640 -28827 -1639
rect -29149 -1960 -29148 -1640
rect -28828 -1960 -28827 -1640
rect -29149 -1961 -28827 -1960
rect -29572 -2308 -29468 -2012
rect -30161 -2360 -29839 -2359
rect -30161 -2680 -30160 -2360
rect -29840 -2680 -29839 -2360
rect -30161 -2681 -29839 -2680
rect -30584 -3028 -30480 -2732
rect -31173 -3080 -30851 -3079
rect -31173 -3400 -31172 -3080
rect -30852 -3400 -30851 -3080
rect -31173 -3401 -30851 -3400
rect -31596 -3748 -31492 -3452
rect -32185 -3800 -31863 -3799
rect -32185 -4120 -32184 -3800
rect -31864 -4120 -31863 -3800
rect -32185 -4121 -31863 -4120
rect -32076 -4519 -31972 -4121
rect -31596 -4172 -31576 -3748
rect -31512 -4172 -31492 -3748
rect -31064 -3799 -30960 -3401
rect -30584 -3452 -30564 -3028
rect -30500 -3452 -30480 -3028
rect -30052 -3079 -29948 -2681
rect -29572 -2732 -29552 -2308
rect -29488 -2732 -29468 -2308
rect -29040 -2359 -28936 -1961
rect -28560 -2012 -28540 -1588
rect -28476 -2012 -28456 -1588
rect -28028 -1639 -27924 -1241
rect -27548 -1292 -27528 -868
rect -27464 -1292 -27444 -868
rect -27016 -919 -26912 -521
rect -26536 -572 -26516 -148
rect -26452 -572 -26432 -148
rect -26004 -199 -25900 199
rect -25524 148 -25504 572
rect -25440 148 -25420 572
rect -24992 521 -24888 919
rect -24512 868 -24492 1292
rect -24428 868 -24408 1292
rect -23980 1241 -23876 1639
rect -23500 1588 -23480 2012
rect -23416 1588 -23396 2012
rect -22968 1961 -22864 2359
rect -22488 2308 -22468 2732
rect -22404 2308 -22384 2732
rect -21956 2681 -21852 3079
rect -21476 3028 -21456 3452
rect -21392 3028 -21372 3452
rect -20944 3401 -20840 3799
rect -20464 3748 -20444 4172
rect -20380 3748 -20360 4172
rect -19932 4121 -19828 4519
rect -19452 4468 -19432 4892
rect -19368 4468 -19348 4892
rect -18920 4841 -18816 5239
rect -18440 5188 -18420 5612
rect -18356 5188 -18336 5612
rect -17908 5561 -17804 5760
rect -17428 5612 -17324 5760
rect -18017 5560 -17695 5561
rect -18017 5240 -18016 5560
rect -17696 5240 -17695 5560
rect -18017 5239 -17695 5240
rect -18440 4892 -18336 5188
rect -19029 4840 -18707 4841
rect -19029 4520 -19028 4840
rect -18708 4520 -18707 4840
rect -19029 4519 -18707 4520
rect -19452 4172 -19348 4468
rect -20041 4120 -19719 4121
rect -20041 3800 -20040 4120
rect -19720 3800 -19719 4120
rect -20041 3799 -19719 3800
rect -20464 3452 -20360 3748
rect -21053 3400 -20731 3401
rect -21053 3080 -21052 3400
rect -20732 3080 -20731 3400
rect -21053 3079 -20731 3080
rect -21476 2732 -21372 3028
rect -22065 2680 -21743 2681
rect -22065 2360 -22064 2680
rect -21744 2360 -21743 2680
rect -22065 2359 -21743 2360
rect -22488 2012 -22384 2308
rect -23077 1960 -22755 1961
rect -23077 1640 -23076 1960
rect -22756 1640 -22755 1960
rect -23077 1639 -22755 1640
rect -23500 1292 -23396 1588
rect -24089 1240 -23767 1241
rect -24089 920 -24088 1240
rect -23768 920 -23767 1240
rect -24089 919 -23767 920
rect -24512 572 -24408 868
rect -25101 520 -24779 521
rect -25101 200 -25100 520
rect -24780 200 -24779 520
rect -25101 199 -24779 200
rect -25524 -148 -25420 148
rect -26113 -200 -25791 -199
rect -26113 -520 -26112 -200
rect -25792 -520 -25791 -200
rect -26113 -521 -25791 -520
rect -26536 -868 -26432 -572
rect -27125 -920 -26803 -919
rect -27125 -1240 -27124 -920
rect -26804 -1240 -26803 -920
rect -27125 -1241 -26803 -1240
rect -27548 -1588 -27444 -1292
rect -28137 -1640 -27815 -1639
rect -28137 -1960 -28136 -1640
rect -27816 -1960 -27815 -1640
rect -28137 -1961 -27815 -1960
rect -28560 -2308 -28456 -2012
rect -29149 -2360 -28827 -2359
rect -29149 -2680 -29148 -2360
rect -28828 -2680 -28827 -2360
rect -29149 -2681 -28827 -2680
rect -29572 -3028 -29468 -2732
rect -30161 -3080 -29839 -3079
rect -30161 -3400 -30160 -3080
rect -29840 -3400 -29839 -3080
rect -30161 -3401 -29839 -3400
rect -30584 -3748 -30480 -3452
rect -31173 -3800 -30851 -3799
rect -31173 -4120 -31172 -3800
rect -30852 -4120 -30851 -3800
rect -31173 -4121 -30851 -4120
rect -31596 -4468 -31492 -4172
rect -32185 -4520 -31863 -4519
rect -32185 -4840 -32184 -4520
rect -31864 -4840 -31863 -4520
rect -32185 -4841 -31863 -4840
rect -32076 -5239 -31972 -4841
rect -31596 -4892 -31576 -4468
rect -31512 -4892 -31492 -4468
rect -31064 -4519 -30960 -4121
rect -30584 -4172 -30564 -3748
rect -30500 -4172 -30480 -3748
rect -30052 -3799 -29948 -3401
rect -29572 -3452 -29552 -3028
rect -29488 -3452 -29468 -3028
rect -29040 -3079 -28936 -2681
rect -28560 -2732 -28540 -2308
rect -28476 -2732 -28456 -2308
rect -28028 -2359 -27924 -1961
rect -27548 -2012 -27528 -1588
rect -27464 -2012 -27444 -1588
rect -27016 -1639 -26912 -1241
rect -26536 -1292 -26516 -868
rect -26452 -1292 -26432 -868
rect -26004 -919 -25900 -521
rect -25524 -572 -25504 -148
rect -25440 -572 -25420 -148
rect -24992 -199 -24888 199
rect -24512 148 -24492 572
rect -24428 148 -24408 572
rect -23980 521 -23876 919
rect -23500 868 -23480 1292
rect -23416 868 -23396 1292
rect -22968 1241 -22864 1639
rect -22488 1588 -22468 2012
rect -22404 1588 -22384 2012
rect -21956 1961 -21852 2359
rect -21476 2308 -21456 2732
rect -21392 2308 -21372 2732
rect -20944 2681 -20840 3079
rect -20464 3028 -20444 3452
rect -20380 3028 -20360 3452
rect -19932 3401 -19828 3799
rect -19452 3748 -19432 4172
rect -19368 3748 -19348 4172
rect -18920 4121 -18816 4519
rect -18440 4468 -18420 4892
rect -18356 4468 -18336 4892
rect -17908 4841 -17804 5239
rect -17428 5188 -17408 5612
rect -17344 5188 -17324 5612
rect -16896 5561 -16792 5760
rect -16416 5612 -16312 5760
rect -17005 5560 -16683 5561
rect -17005 5240 -17004 5560
rect -16684 5240 -16683 5560
rect -17005 5239 -16683 5240
rect -17428 4892 -17324 5188
rect -18017 4840 -17695 4841
rect -18017 4520 -18016 4840
rect -17696 4520 -17695 4840
rect -18017 4519 -17695 4520
rect -18440 4172 -18336 4468
rect -19029 4120 -18707 4121
rect -19029 3800 -19028 4120
rect -18708 3800 -18707 4120
rect -19029 3799 -18707 3800
rect -19452 3452 -19348 3748
rect -20041 3400 -19719 3401
rect -20041 3080 -20040 3400
rect -19720 3080 -19719 3400
rect -20041 3079 -19719 3080
rect -20464 2732 -20360 3028
rect -21053 2680 -20731 2681
rect -21053 2360 -21052 2680
rect -20732 2360 -20731 2680
rect -21053 2359 -20731 2360
rect -21476 2012 -21372 2308
rect -22065 1960 -21743 1961
rect -22065 1640 -22064 1960
rect -21744 1640 -21743 1960
rect -22065 1639 -21743 1640
rect -22488 1292 -22384 1588
rect -23077 1240 -22755 1241
rect -23077 920 -23076 1240
rect -22756 920 -22755 1240
rect -23077 919 -22755 920
rect -23500 572 -23396 868
rect -24089 520 -23767 521
rect -24089 200 -24088 520
rect -23768 200 -23767 520
rect -24089 199 -23767 200
rect -24512 -148 -24408 148
rect -25101 -200 -24779 -199
rect -25101 -520 -25100 -200
rect -24780 -520 -24779 -200
rect -25101 -521 -24779 -520
rect -25524 -868 -25420 -572
rect -26113 -920 -25791 -919
rect -26113 -1240 -26112 -920
rect -25792 -1240 -25791 -920
rect -26113 -1241 -25791 -1240
rect -26536 -1588 -26432 -1292
rect -27125 -1640 -26803 -1639
rect -27125 -1960 -27124 -1640
rect -26804 -1960 -26803 -1640
rect -27125 -1961 -26803 -1960
rect -27548 -2308 -27444 -2012
rect -28137 -2360 -27815 -2359
rect -28137 -2680 -28136 -2360
rect -27816 -2680 -27815 -2360
rect -28137 -2681 -27815 -2680
rect -28560 -3028 -28456 -2732
rect -29149 -3080 -28827 -3079
rect -29149 -3400 -29148 -3080
rect -28828 -3400 -28827 -3080
rect -29149 -3401 -28827 -3400
rect -29572 -3748 -29468 -3452
rect -30161 -3800 -29839 -3799
rect -30161 -4120 -30160 -3800
rect -29840 -4120 -29839 -3800
rect -30161 -4121 -29839 -4120
rect -30584 -4468 -30480 -4172
rect -31173 -4520 -30851 -4519
rect -31173 -4840 -31172 -4520
rect -30852 -4840 -30851 -4520
rect -31173 -4841 -30851 -4840
rect -31596 -5188 -31492 -4892
rect -32185 -5240 -31863 -5239
rect -32185 -5560 -32184 -5240
rect -31864 -5560 -31863 -5240
rect -32185 -5561 -31863 -5560
rect -32076 -5760 -31972 -5561
rect -31596 -5612 -31576 -5188
rect -31512 -5612 -31492 -5188
rect -31064 -5239 -30960 -4841
rect -30584 -4892 -30564 -4468
rect -30500 -4892 -30480 -4468
rect -30052 -4519 -29948 -4121
rect -29572 -4172 -29552 -3748
rect -29488 -4172 -29468 -3748
rect -29040 -3799 -28936 -3401
rect -28560 -3452 -28540 -3028
rect -28476 -3452 -28456 -3028
rect -28028 -3079 -27924 -2681
rect -27548 -2732 -27528 -2308
rect -27464 -2732 -27444 -2308
rect -27016 -2359 -26912 -1961
rect -26536 -2012 -26516 -1588
rect -26452 -2012 -26432 -1588
rect -26004 -1639 -25900 -1241
rect -25524 -1292 -25504 -868
rect -25440 -1292 -25420 -868
rect -24992 -919 -24888 -521
rect -24512 -572 -24492 -148
rect -24428 -572 -24408 -148
rect -23980 -199 -23876 199
rect -23500 148 -23480 572
rect -23416 148 -23396 572
rect -22968 521 -22864 919
rect -22488 868 -22468 1292
rect -22404 868 -22384 1292
rect -21956 1241 -21852 1639
rect -21476 1588 -21456 2012
rect -21392 1588 -21372 2012
rect -20944 1961 -20840 2359
rect -20464 2308 -20444 2732
rect -20380 2308 -20360 2732
rect -19932 2681 -19828 3079
rect -19452 3028 -19432 3452
rect -19368 3028 -19348 3452
rect -18920 3401 -18816 3799
rect -18440 3748 -18420 4172
rect -18356 3748 -18336 4172
rect -17908 4121 -17804 4519
rect -17428 4468 -17408 4892
rect -17344 4468 -17324 4892
rect -16896 4841 -16792 5239
rect -16416 5188 -16396 5612
rect -16332 5188 -16312 5612
rect -15884 5561 -15780 5760
rect -15404 5612 -15300 5760
rect -15993 5560 -15671 5561
rect -15993 5240 -15992 5560
rect -15672 5240 -15671 5560
rect -15993 5239 -15671 5240
rect -16416 4892 -16312 5188
rect -17005 4840 -16683 4841
rect -17005 4520 -17004 4840
rect -16684 4520 -16683 4840
rect -17005 4519 -16683 4520
rect -17428 4172 -17324 4468
rect -18017 4120 -17695 4121
rect -18017 3800 -18016 4120
rect -17696 3800 -17695 4120
rect -18017 3799 -17695 3800
rect -18440 3452 -18336 3748
rect -19029 3400 -18707 3401
rect -19029 3080 -19028 3400
rect -18708 3080 -18707 3400
rect -19029 3079 -18707 3080
rect -19452 2732 -19348 3028
rect -20041 2680 -19719 2681
rect -20041 2360 -20040 2680
rect -19720 2360 -19719 2680
rect -20041 2359 -19719 2360
rect -20464 2012 -20360 2308
rect -21053 1960 -20731 1961
rect -21053 1640 -21052 1960
rect -20732 1640 -20731 1960
rect -21053 1639 -20731 1640
rect -21476 1292 -21372 1588
rect -22065 1240 -21743 1241
rect -22065 920 -22064 1240
rect -21744 920 -21743 1240
rect -22065 919 -21743 920
rect -22488 572 -22384 868
rect -23077 520 -22755 521
rect -23077 200 -23076 520
rect -22756 200 -22755 520
rect -23077 199 -22755 200
rect -23500 -148 -23396 148
rect -24089 -200 -23767 -199
rect -24089 -520 -24088 -200
rect -23768 -520 -23767 -200
rect -24089 -521 -23767 -520
rect -24512 -868 -24408 -572
rect -25101 -920 -24779 -919
rect -25101 -1240 -25100 -920
rect -24780 -1240 -24779 -920
rect -25101 -1241 -24779 -1240
rect -25524 -1588 -25420 -1292
rect -26113 -1640 -25791 -1639
rect -26113 -1960 -26112 -1640
rect -25792 -1960 -25791 -1640
rect -26113 -1961 -25791 -1960
rect -26536 -2308 -26432 -2012
rect -27125 -2360 -26803 -2359
rect -27125 -2680 -27124 -2360
rect -26804 -2680 -26803 -2360
rect -27125 -2681 -26803 -2680
rect -27548 -3028 -27444 -2732
rect -28137 -3080 -27815 -3079
rect -28137 -3400 -28136 -3080
rect -27816 -3400 -27815 -3080
rect -28137 -3401 -27815 -3400
rect -28560 -3748 -28456 -3452
rect -29149 -3800 -28827 -3799
rect -29149 -4120 -29148 -3800
rect -28828 -4120 -28827 -3800
rect -29149 -4121 -28827 -4120
rect -29572 -4468 -29468 -4172
rect -30161 -4520 -29839 -4519
rect -30161 -4840 -30160 -4520
rect -29840 -4840 -29839 -4520
rect -30161 -4841 -29839 -4840
rect -30584 -5188 -30480 -4892
rect -31173 -5240 -30851 -5239
rect -31173 -5560 -31172 -5240
rect -30852 -5560 -30851 -5240
rect -31173 -5561 -30851 -5560
rect -31596 -5760 -31492 -5612
rect -31064 -5760 -30960 -5561
rect -30584 -5612 -30564 -5188
rect -30500 -5612 -30480 -5188
rect -30052 -5239 -29948 -4841
rect -29572 -4892 -29552 -4468
rect -29488 -4892 -29468 -4468
rect -29040 -4519 -28936 -4121
rect -28560 -4172 -28540 -3748
rect -28476 -4172 -28456 -3748
rect -28028 -3799 -27924 -3401
rect -27548 -3452 -27528 -3028
rect -27464 -3452 -27444 -3028
rect -27016 -3079 -26912 -2681
rect -26536 -2732 -26516 -2308
rect -26452 -2732 -26432 -2308
rect -26004 -2359 -25900 -1961
rect -25524 -2012 -25504 -1588
rect -25440 -2012 -25420 -1588
rect -24992 -1639 -24888 -1241
rect -24512 -1292 -24492 -868
rect -24428 -1292 -24408 -868
rect -23980 -919 -23876 -521
rect -23500 -572 -23480 -148
rect -23416 -572 -23396 -148
rect -22968 -199 -22864 199
rect -22488 148 -22468 572
rect -22404 148 -22384 572
rect -21956 521 -21852 919
rect -21476 868 -21456 1292
rect -21392 868 -21372 1292
rect -20944 1241 -20840 1639
rect -20464 1588 -20444 2012
rect -20380 1588 -20360 2012
rect -19932 1961 -19828 2359
rect -19452 2308 -19432 2732
rect -19368 2308 -19348 2732
rect -18920 2681 -18816 3079
rect -18440 3028 -18420 3452
rect -18356 3028 -18336 3452
rect -17908 3401 -17804 3799
rect -17428 3748 -17408 4172
rect -17344 3748 -17324 4172
rect -16896 4121 -16792 4519
rect -16416 4468 -16396 4892
rect -16332 4468 -16312 4892
rect -15884 4841 -15780 5239
rect -15404 5188 -15384 5612
rect -15320 5188 -15300 5612
rect -14872 5561 -14768 5760
rect -14392 5612 -14288 5760
rect -14981 5560 -14659 5561
rect -14981 5240 -14980 5560
rect -14660 5240 -14659 5560
rect -14981 5239 -14659 5240
rect -15404 4892 -15300 5188
rect -15993 4840 -15671 4841
rect -15993 4520 -15992 4840
rect -15672 4520 -15671 4840
rect -15993 4519 -15671 4520
rect -16416 4172 -16312 4468
rect -17005 4120 -16683 4121
rect -17005 3800 -17004 4120
rect -16684 3800 -16683 4120
rect -17005 3799 -16683 3800
rect -17428 3452 -17324 3748
rect -18017 3400 -17695 3401
rect -18017 3080 -18016 3400
rect -17696 3080 -17695 3400
rect -18017 3079 -17695 3080
rect -18440 2732 -18336 3028
rect -19029 2680 -18707 2681
rect -19029 2360 -19028 2680
rect -18708 2360 -18707 2680
rect -19029 2359 -18707 2360
rect -19452 2012 -19348 2308
rect -20041 1960 -19719 1961
rect -20041 1640 -20040 1960
rect -19720 1640 -19719 1960
rect -20041 1639 -19719 1640
rect -20464 1292 -20360 1588
rect -21053 1240 -20731 1241
rect -21053 920 -21052 1240
rect -20732 920 -20731 1240
rect -21053 919 -20731 920
rect -21476 572 -21372 868
rect -22065 520 -21743 521
rect -22065 200 -22064 520
rect -21744 200 -21743 520
rect -22065 199 -21743 200
rect -22488 -148 -22384 148
rect -23077 -200 -22755 -199
rect -23077 -520 -23076 -200
rect -22756 -520 -22755 -200
rect -23077 -521 -22755 -520
rect -23500 -868 -23396 -572
rect -24089 -920 -23767 -919
rect -24089 -1240 -24088 -920
rect -23768 -1240 -23767 -920
rect -24089 -1241 -23767 -1240
rect -24512 -1588 -24408 -1292
rect -25101 -1640 -24779 -1639
rect -25101 -1960 -25100 -1640
rect -24780 -1960 -24779 -1640
rect -25101 -1961 -24779 -1960
rect -25524 -2308 -25420 -2012
rect -26113 -2360 -25791 -2359
rect -26113 -2680 -26112 -2360
rect -25792 -2680 -25791 -2360
rect -26113 -2681 -25791 -2680
rect -26536 -3028 -26432 -2732
rect -27125 -3080 -26803 -3079
rect -27125 -3400 -27124 -3080
rect -26804 -3400 -26803 -3080
rect -27125 -3401 -26803 -3400
rect -27548 -3748 -27444 -3452
rect -28137 -3800 -27815 -3799
rect -28137 -4120 -28136 -3800
rect -27816 -4120 -27815 -3800
rect -28137 -4121 -27815 -4120
rect -28560 -4468 -28456 -4172
rect -29149 -4520 -28827 -4519
rect -29149 -4840 -29148 -4520
rect -28828 -4840 -28827 -4520
rect -29149 -4841 -28827 -4840
rect -29572 -5188 -29468 -4892
rect -30161 -5240 -29839 -5239
rect -30161 -5560 -30160 -5240
rect -29840 -5560 -29839 -5240
rect -30161 -5561 -29839 -5560
rect -30584 -5760 -30480 -5612
rect -30052 -5760 -29948 -5561
rect -29572 -5612 -29552 -5188
rect -29488 -5612 -29468 -5188
rect -29040 -5239 -28936 -4841
rect -28560 -4892 -28540 -4468
rect -28476 -4892 -28456 -4468
rect -28028 -4519 -27924 -4121
rect -27548 -4172 -27528 -3748
rect -27464 -4172 -27444 -3748
rect -27016 -3799 -26912 -3401
rect -26536 -3452 -26516 -3028
rect -26452 -3452 -26432 -3028
rect -26004 -3079 -25900 -2681
rect -25524 -2732 -25504 -2308
rect -25440 -2732 -25420 -2308
rect -24992 -2359 -24888 -1961
rect -24512 -2012 -24492 -1588
rect -24428 -2012 -24408 -1588
rect -23980 -1639 -23876 -1241
rect -23500 -1292 -23480 -868
rect -23416 -1292 -23396 -868
rect -22968 -919 -22864 -521
rect -22488 -572 -22468 -148
rect -22404 -572 -22384 -148
rect -21956 -199 -21852 199
rect -21476 148 -21456 572
rect -21392 148 -21372 572
rect -20944 521 -20840 919
rect -20464 868 -20444 1292
rect -20380 868 -20360 1292
rect -19932 1241 -19828 1639
rect -19452 1588 -19432 2012
rect -19368 1588 -19348 2012
rect -18920 1961 -18816 2359
rect -18440 2308 -18420 2732
rect -18356 2308 -18336 2732
rect -17908 2681 -17804 3079
rect -17428 3028 -17408 3452
rect -17344 3028 -17324 3452
rect -16896 3401 -16792 3799
rect -16416 3748 -16396 4172
rect -16332 3748 -16312 4172
rect -15884 4121 -15780 4519
rect -15404 4468 -15384 4892
rect -15320 4468 -15300 4892
rect -14872 4841 -14768 5239
rect -14392 5188 -14372 5612
rect -14308 5188 -14288 5612
rect -13860 5561 -13756 5760
rect -13380 5612 -13276 5760
rect -13969 5560 -13647 5561
rect -13969 5240 -13968 5560
rect -13648 5240 -13647 5560
rect -13969 5239 -13647 5240
rect -14392 4892 -14288 5188
rect -14981 4840 -14659 4841
rect -14981 4520 -14980 4840
rect -14660 4520 -14659 4840
rect -14981 4519 -14659 4520
rect -15404 4172 -15300 4468
rect -15993 4120 -15671 4121
rect -15993 3800 -15992 4120
rect -15672 3800 -15671 4120
rect -15993 3799 -15671 3800
rect -16416 3452 -16312 3748
rect -17005 3400 -16683 3401
rect -17005 3080 -17004 3400
rect -16684 3080 -16683 3400
rect -17005 3079 -16683 3080
rect -17428 2732 -17324 3028
rect -18017 2680 -17695 2681
rect -18017 2360 -18016 2680
rect -17696 2360 -17695 2680
rect -18017 2359 -17695 2360
rect -18440 2012 -18336 2308
rect -19029 1960 -18707 1961
rect -19029 1640 -19028 1960
rect -18708 1640 -18707 1960
rect -19029 1639 -18707 1640
rect -19452 1292 -19348 1588
rect -20041 1240 -19719 1241
rect -20041 920 -20040 1240
rect -19720 920 -19719 1240
rect -20041 919 -19719 920
rect -20464 572 -20360 868
rect -21053 520 -20731 521
rect -21053 200 -21052 520
rect -20732 200 -20731 520
rect -21053 199 -20731 200
rect -21476 -148 -21372 148
rect -22065 -200 -21743 -199
rect -22065 -520 -22064 -200
rect -21744 -520 -21743 -200
rect -22065 -521 -21743 -520
rect -22488 -868 -22384 -572
rect -23077 -920 -22755 -919
rect -23077 -1240 -23076 -920
rect -22756 -1240 -22755 -920
rect -23077 -1241 -22755 -1240
rect -23500 -1588 -23396 -1292
rect -24089 -1640 -23767 -1639
rect -24089 -1960 -24088 -1640
rect -23768 -1960 -23767 -1640
rect -24089 -1961 -23767 -1960
rect -24512 -2308 -24408 -2012
rect -25101 -2360 -24779 -2359
rect -25101 -2680 -25100 -2360
rect -24780 -2680 -24779 -2360
rect -25101 -2681 -24779 -2680
rect -25524 -3028 -25420 -2732
rect -26113 -3080 -25791 -3079
rect -26113 -3400 -26112 -3080
rect -25792 -3400 -25791 -3080
rect -26113 -3401 -25791 -3400
rect -26536 -3748 -26432 -3452
rect -27125 -3800 -26803 -3799
rect -27125 -4120 -27124 -3800
rect -26804 -4120 -26803 -3800
rect -27125 -4121 -26803 -4120
rect -27548 -4468 -27444 -4172
rect -28137 -4520 -27815 -4519
rect -28137 -4840 -28136 -4520
rect -27816 -4840 -27815 -4520
rect -28137 -4841 -27815 -4840
rect -28560 -5188 -28456 -4892
rect -29149 -5240 -28827 -5239
rect -29149 -5560 -29148 -5240
rect -28828 -5560 -28827 -5240
rect -29149 -5561 -28827 -5560
rect -29572 -5760 -29468 -5612
rect -29040 -5760 -28936 -5561
rect -28560 -5612 -28540 -5188
rect -28476 -5612 -28456 -5188
rect -28028 -5239 -27924 -4841
rect -27548 -4892 -27528 -4468
rect -27464 -4892 -27444 -4468
rect -27016 -4519 -26912 -4121
rect -26536 -4172 -26516 -3748
rect -26452 -4172 -26432 -3748
rect -26004 -3799 -25900 -3401
rect -25524 -3452 -25504 -3028
rect -25440 -3452 -25420 -3028
rect -24992 -3079 -24888 -2681
rect -24512 -2732 -24492 -2308
rect -24428 -2732 -24408 -2308
rect -23980 -2359 -23876 -1961
rect -23500 -2012 -23480 -1588
rect -23416 -2012 -23396 -1588
rect -22968 -1639 -22864 -1241
rect -22488 -1292 -22468 -868
rect -22404 -1292 -22384 -868
rect -21956 -919 -21852 -521
rect -21476 -572 -21456 -148
rect -21392 -572 -21372 -148
rect -20944 -199 -20840 199
rect -20464 148 -20444 572
rect -20380 148 -20360 572
rect -19932 521 -19828 919
rect -19452 868 -19432 1292
rect -19368 868 -19348 1292
rect -18920 1241 -18816 1639
rect -18440 1588 -18420 2012
rect -18356 1588 -18336 2012
rect -17908 1961 -17804 2359
rect -17428 2308 -17408 2732
rect -17344 2308 -17324 2732
rect -16896 2681 -16792 3079
rect -16416 3028 -16396 3452
rect -16332 3028 -16312 3452
rect -15884 3401 -15780 3799
rect -15404 3748 -15384 4172
rect -15320 3748 -15300 4172
rect -14872 4121 -14768 4519
rect -14392 4468 -14372 4892
rect -14308 4468 -14288 4892
rect -13860 4841 -13756 5239
rect -13380 5188 -13360 5612
rect -13296 5188 -13276 5612
rect -12848 5561 -12744 5760
rect -12368 5612 -12264 5760
rect -12957 5560 -12635 5561
rect -12957 5240 -12956 5560
rect -12636 5240 -12635 5560
rect -12957 5239 -12635 5240
rect -13380 4892 -13276 5188
rect -13969 4840 -13647 4841
rect -13969 4520 -13968 4840
rect -13648 4520 -13647 4840
rect -13969 4519 -13647 4520
rect -14392 4172 -14288 4468
rect -14981 4120 -14659 4121
rect -14981 3800 -14980 4120
rect -14660 3800 -14659 4120
rect -14981 3799 -14659 3800
rect -15404 3452 -15300 3748
rect -15993 3400 -15671 3401
rect -15993 3080 -15992 3400
rect -15672 3080 -15671 3400
rect -15993 3079 -15671 3080
rect -16416 2732 -16312 3028
rect -17005 2680 -16683 2681
rect -17005 2360 -17004 2680
rect -16684 2360 -16683 2680
rect -17005 2359 -16683 2360
rect -17428 2012 -17324 2308
rect -18017 1960 -17695 1961
rect -18017 1640 -18016 1960
rect -17696 1640 -17695 1960
rect -18017 1639 -17695 1640
rect -18440 1292 -18336 1588
rect -19029 1240 -18707 1241
rect -19029 920 -19028 1240
rect -18708 920 -18707 1240
rect -19029 919 -18707 920
rect -19452 572 -19348 868
rect -20041 520 -19719 521
rect -20041 200 -20040 520
rect -19720 200 -19719 520
rect -20041 199 -19719 200
rect -20464 -148 -20360 148
rect -21053 -200 -20731 -199
rect -21053 -520 -21052 -200
rect -20732 -520 -20731 -200
rect -21053 -521 -20731 -520
rect -21476 -868 -21372 -572
rect -22065 -920 -21743 -919
rect -22065 -1240 -22064 -920
rect -21744 -1240 -21743 -920
rect -22065 -1241 -21743 -1240
rect -22488 -1588 -22384 -1292
rect -23077 -1640 -22755 -1639
rect -23077 -1960 -23076 -1640
rect -22756 -1960 -22755 -1640
rect -23077 -1961 -22755 -1960
rect -23500 -2308 -23396 -2012
rect -24089 -2360 -23767 -2359
rect -24089 -2680 -24088 -2360
rect -23768 -2680 -23767 -2360
rect -24089 -2681 -23767 -2680
rect -24512 -3028 -24408 -2732
rect -25101 -3080 -24779 -3079
rect -25101 -3400 -25100 -3080
rect -24780 -3400 -24779 -3080
rect -25101 -3401 -24779 -3400
rect -25524 -3748 -25420 -3452
rect -26113 -3800 -25791 -3799
rect -26113 -4120 -26112 -3800
rect -25792 -4120 -25791 -3800
rect -26113 -4121 -25791 -4120
rect -26536 -4468 -26432 -4172
rect -27125 -4520 -26803 -4519
rect -27125 -4840 -27124 -4520
rect -26804 -4840 -26803 -4520
rect -27125 -4841 -26803 -4840
rect -27548 -5188 -27444 -4892
rect -28137 -5240 -27815 -5239
rect -28137 -5560 -28136 -5240
rect -27816 -5560 -27815 -5240
rect -28137 -5561 -27815 -5560
rect -28560 -5760 -28456 -5612
rect -28028 -5760 -27924 -5561
rect -27548 -5612 -27528 -5188
rect -27464 -5612 -27444 -5188
rect -27016 -5239 -26912 -4841
rect -26536 -4892 -26516 -4468
rect -26452 -4892 -26432 -4468
rect -26004 -4519 -25900 -4121
rect -25524 -4172 -25504 -3748
rect -25440 -4172 -25420 -3748
rect -24992 -3799 -24888 -3401
rect -24512 -3452 -24492 -3028
rect -24428 -3452 -24408 -3028
rect -23980 -3079 -23876 -2681
rect -23500 -2732 -23480 -2308
rect -23416 -2732 -23396 -2308
rect -22968 -2359 -22864 -1961
rect -22488 -2012 -22468 -1588
rect -22404 -2012 -22384 -1588
rect -21956 -1639 -21852 -1241
rect -21476 -1292 -21456 -868
rect -21392 -1292 -21372 -868
rect -20944 -919 -20840 -521
rect -20464 -572 -20444 -148
rect -20380 -572 -20360 -148
rect -19932 -199 -19828 199
rect -19452 148 -19432 572
rect -19368 148 -19348 572
rect -18920 521 -18816 919
rect -18440 868 -18420 1292
rect -18356 868 -18336 1292
rect -17908 1241 -17804 1639
rect -17428 1588 -17408 2012
rect -17344 1588 -17324 2012
rect -16896 1961 -16792 2359
rect -16416 2308 -16396 2732
rect -16332 2308 -16312 2732
rect -15884 2681 -15780 3079
rect -15404 3028 -15384 3452
rect -15320 3028 -15300 3452
rect -14872 3401 -14768 3799
rect -14392 3748 -14372 4172
rect -14308 3748 -14288 4172
rect -13860 4121 -13756 4519
rect -13380 4468 -13360 4892
rect -13296 4468 -13276 4892
rect -12848 4841 -12744 5239
rect -12368 5188 -12348 5612
rect -12284 5188 -12264 5612
rect -11836 5561 -11732 5760
rect -11356 5612 -11252 5760
rect -11945 5560 -11623 5561
rect -11945 5240 -11944 5560
rect -11624 5240 -11623 5560
rect -11945 5239 -11623 5240
rect -12368 4892 -12264 5188
rect -12957 4840 -12635 4841
rect -12957 4520 -12956 4840
rect -12636 4520 -12635 4840
rect -12957 4519 -12635 4520
rect -13380 4172 -13276 4468
rect -13969 4120 -13647 4121
rect -13969 3800 -13968 4120
rect -13648 3800 -13647 4120
rect -13969 3799 -13647 3800
rect -14392 3452 -14288 3748
rect -14981 3400 -14659 3401
rect -14981 3080 -14980 3400
rect -14660 3080 -14659 3400
rect -14981 3079 -14659 3080
rect -15404 2732 -15300 3028
rect -15993 2680 -15671 2681
rect -15993 2360 -15992 2680
rect -15672 2360 -15671 2680
rect -15993 2359 -15671 2360
rect -16416 2012 -16312 2308
rect -17005 1960 -16683 1961
rect -17005 1640 -17004 1960
rect -16684 1640 -16683 1960
rect -17005 1639 -16683 1640
rect -17428 1292 -17324 1588
rect -18017 1240 -17695 1241
rect -18017 920 -18016 1240
rect -17696 920 -17695 1240
rect -18017 919 -17695 920
rect -18440 572 -18336 868
rect -19029 520 -18707 521
rect -19029 200 -19028 520
rect -18708 200 -18707 520
rect -19029 199 -18707 200
rect -19452 -148 -19348 148
rect -20041 -200 -19719 -199
rect -20041 -520 -20040 -200
rect -19720 -520 -19719 -200
rect -20041 -521 -19719 -520
rect -20464 -868 -20360 -572
rect -21053 -920 -20731 -919
rect -21053 -1240 -21052 -920
rect -20732 -1240 -20731 -920
rect -21053 -1241 -20731 -1240
rect -21476 -1588 -21372 -1292
rect -22065 -1640 -21743 -1639
rect -22065 -1960 -22064 -1640
rect -21744 -1960 -21743 -1640
rect -22065 -1961 -21743 -1960
rect -22488 -2308 -22384 -2012
rect -23077 -2360 -22755 -2359
rect -23077 -2680 -23076 -2360
rect -22756 -2680 -22755 -2360
rect -23077 -2681 -22755 -2680
rect -23500 -3028 -23396 -2732
rect -24089 -3080 -23767 -3079
rect -24089 -3400 -24088 -3080
rect -23768 -3400 -23767 -3080
rect -24089 -3401 -23767 -3400
rect -24512 -3748 -24408 -3452
rect -25101 -3800 -24779 -3799
rect -25101 -4120 -25100 -3800
rect -24780 -4120 -24779 -3800
rect -25101 -4121 -24779 -4120
rect -25524 -4468 -25420 -4172
rect -26113 -4520 -25791 -4519
rect -26113 -4840 -26112 -4520
rect -25792 -4840 -25791 -4520
rect -26113 -4841 -25791 -4840
rect -26536 -5188 -26432 -4892
rect -27125 -5240 -26803 -5239
rect -27125 -5560 -27124 -5240
rect -26804 -5560 -26803 -5240
rect -27125 -5561 -26803 -5560
rect -27548 -5760 -27444 -5612
rect -27016 -5760 -26912 -5561
rect -26536 -5612 -26516 -5188
rect -26452 -5612 -26432 -5188
rect -26004 -5239 -25900 -4841
rect -25524 -4892 -25504 -4468
rect -25440 -4892 -25420 -4468
rect -24992 -4519 -24888 -4121
rect -24512 -4172 -24492 -3748
rect -24428 -4172 -24408 -3748
rect -23980 -3799 -23876 -3401
rect -23500 -3452 -23480 -3028
rect -23416 -3452 -23396 -3028
rect -22968 -3079 -22864 -2681
rect -22488 -2732 -22468 -2308
rect -22404 -2732 -22384 -2308
rect -21956 -2359 -21852 -1961
rect -21476 -2012 -21456 -1588
rect -21392 -2012 -21372 -1588
rect -20944 -1639 -20840 -1241
rect -20464 -1292 -20444 -868
rect -20380 -1292 -20360 -868
rect -19932 -919 -19828 -521
rect -19452 -572 -19432 -148
rect -19368 -572 -19348 -148
rect -18920 -199 -18816 199
rect -18440 148 -18420 572
rect -18356 148 -18336 572
rect -17908 521 -17804 919
rect -17428 868 -17408 1292
rect -17344 868 -17324 1292
rect -16896 1241 -16792 1639
rect -16416 1588 -16396 2012
rect -16332 1588 -16312 2012
rect -15884 1961 -15780 2359
rect -15404 2308 -15384 2732
rect -15320 2308 -15300 2732
rect -14872 2681 -14768 3079
rect -14392 3028 -14372 3452
rect -14308 3028 -14288 3452
rect -13860 3401 -13756 3799
rect -13380 3748 -13360 4172
rect -13296 3748 -13276 4172
rect -12848 4121 -12744 4519
rect -12368 4468 -12348 4892
rect -12284 4468 -12264 4892
rect -11836 4841 -11732 5239
rect -11356 5188 -11336 5612
rect -11272 5188 -11252 5612
rect -10824 5561 -10720 5760
rect -10344 5612 -10240 5760
rect -10933 5560 -10611 5561
rect -10933 5240 -10932 5560
rect -10612 5240 -10611 5560
rect -10933 5239 -10611 5240
rect -11356 4892 -11252 5188
rect -11945 4840 -11623 4841
rect -11945 4520 -11944 4840
rect -11624 4520 -11623 4840
rect -11945 4519 -11623 4520
rect -12368 4172 -12264 4468
rect -12957 4120 -12635 4121
rect -12957 3800 -12956 4120
rect -12636 3800 -12635 4120
rect -12957 3799 -12635 3800
rect -13380 3452 -13276 3748
rect -13969 3400 -13647 3401
rect -13969 3080 -13968 3400
rect -13648 3080 -13647 3400
rect -13969 3079 -13647 3080
rect -14392 2732 -14288 3028
rect -14981 2680 -14659 2681
rect -14981 2360 -14980 2680
rect -14660 2360 -14659 2680
rect -14981 2359 -14659 2360
rect -15404 2012 -15300 2308
rect -15993 1960 -15671 1961
rect -15993 1640 -15992 1960
rect -15672 1640 -15671 1960
rect -15993 1639 -15671 1640
rect -16416 1292 -16312 1588
rect -17005 1240 -16683 1241
rect -17005 920 -17004 1240
rect -16684 920 -16683 1240
rect -17005 919 -16683 920
rect -17428 572 -17324 868
rect -18017 520 -17695 521
rect -18017 200 -18016 520
rect -17696 200 -17695 520
rect -18017 199 -17695 200
rect -18440 -148 -18336 148
rect -19029 -200 -18707 -199
rect -19029 -520 -19028 -200
rect -18708 -520 -18707 -200
rect -19029 -521 -18707 -520
rect -19452 -868 -19348 -572
rect -20041 -920 -19719 -919
rect -20041 -1240 -20040 -920
rect -19720 -1240 -19719 -920
rect -20041 -1241 -19719 -1240
rect -20464 -1588 -20360 -1292
rect -21053 -1640 -20731 -1639
rect -21053 -1960 -21052 -1640
rect -20732 -1960 -20731 -1640
rect -21053 -1961 -20731 -1960
rect -21476 -2308 -21372 -2012
rect -22065 -2360 -21743 -2359
rect -22065 -2680 -22064 -2360
rect -21744 -2680 -21743 -2360
rect -22065 -2681 -21743 -2680
rect -22488 -3028 -22384 -2732
rect -23077 -3080 -22755 -3079
rect -23077 -3400 -23076 -3080
rect -22756 -3400 -22755 -3080
rect -23077 -3401 -22755 -3400
rect -23500 -3748 -23396 -3452
rect -24089 -3800 -23767 -3799
rect -24089 -4120 -24088 -3800
rect -23768 -4120 -23767 -3800
rect -24089 -4121 -23767 -4120
rect -24512 -4468 -24408 -4172
rect -25101 -4520 -24779 -4519
rect -25101 -4840 -25100 -4520
rect -24780 -4840 -24779 -4520
rect -25101 -4841 -24779 -4840
rect -25524 -5188 -25420 -4892
rect -26113 -5240 -25791 -5239
rect -26113 -5560 -26112 -5240
rect -25792 -5560 -25791 -5240
rect -26113 -5561 -25791 -5560
rect -26536 -5760 -26432 -5612
rect -26004 -5760 -25900 -5561
rect -25524 -5612 -25504 -5188
rect -25440 -5612 -25420 -5188
rect -24992 -5239 -24888 -4841
rect -24512 -4892 -24492 -4468
rect -24428 -4892 -24408 -4468
rect -23980 -4519 -23876 -4121
rect -23500 -4172 -23480 -3748
rect -23416 -4172 -23396 -3748
rect -22968 -3799 -22864 -3401
rect -22488 -3452 -22468 -3028
rect -22404 -3452 -22384 -3028
rect -21956 -3079 -21852 -2681
rect -21476 -2732 -21456 -2308
rect -21392 -2732 -21372 -2308
rect -20944 -2359 -20840 -1961
rect -20464 -2012 -20444 -1588
rect -20380 -2012 -20360 -1588
rect -19932 -1639 -19828 -1241
rect -19452 -1292 -19432 -868
rect -19368 -1292 -19348 -868
rect -18920 -919 -18816 -521
rect -18440 -572 -18420 -148
rect -18356 -572 -18336 -148
rect -17908 -199 -17804 199
rect -17428 148 -17408 572
rect -17344 148 -17324 572
rect -16896 521 -16792 919
rect -16416 868 -16396 1292
rect -16332 868 -16312 1292
rect -15884 1241 -15780 1639
rect -15404 1588 -15384 2012
rect -15320 1588 -15300 2012
rect -14872 1961 -14768 2359
rect -14392 2308 -14372 2732
rect -14308 2308 -14288 2732
rect -13860 2681 -13756 3079
rect -13380 3028 -13360 3452
rect -13296 3028 -13276 3452
rect -12848 3401 -12744 3799
rect -12368 3748 -12348 4172
rect -12284 3748 -12264 4172
rect -11836 4121 -11732 4519
rect -11356 4468 -11336 4892
rect -11272 4468 -11252 4892
rect -10824 4841 -10720 5239
rect -10344 5188 -10324 5612
rect -10260 5188 -10240 5612
rect -9812 5561 -9708 5760
rect -9332 5612 -9228 5760
rect -9921 5560 -9599 5561
rect -9921 5240 -9920 5560
rect -9600 5240 -9599 5560
rect -9921 5239 -9599 5240
rect -10344 4892 -10240 5188
rect -10933 4840 -10611 4841
rect -10933 4520 -10932 4840
rect -10612 4520 -10611 4840
rect -10933 4519 -10611 4520
rect -11356 4172 -11252 4468
rect -11945 4120 -11623 4121
rect -11945 3800 -11944 4120
rect -11624 3800 -11623 4120
rect -11945 3799 -11623 3800
rect -12368 3452 -12264 3748
rect -12957 3400 -12635 3401
rect -12957 3080 -12956 3400
rect -12636 3080 -12635 3400
rect -12957 3079 -12635 3080
rect -13380 2732 -13276 3028
rect -13969 2680 -13647 2681
rect -13969 2360 -13968 2680
rect -13648 2360 -13647 2680
rect -13969 2359 -13647 2360
rect -14392 2012 -14288 2308
rect -14981 1960 -14659 1961
rect -14981 1640 -14980 1960
rect -14660 1640 -14659 1960
rect -14981 1639 -14659 1640
rect -15404 1292 -15300 1588
rect -15993 1240 -15671 1241
rect -15993 920 -15992 1240
rect -15672 920 -15671 1240
rect -15993 919 -15671 920
rect -16416 572 -16312 868
rect -17005 520 -16683 521
rect -17005 200 -17004 520
rect -16684 200 -16683 520
rect -17005 199 -16683 200
rect -17428 -148 -17324 148
rect -18017 -200 -17695 -199
rect -18017 -520 -18016 -200
rect -17696 -520 -17695 -200
rect -18017 -521 -17695 -520
rect -18440 -868 -18336 -572
rect -19029 -920 -18707 -919
rect -19029 -1240 -19028 -920
rect -18708 -1240 -18707 -920
rect -19029 -1241 -18707 -1240
rect -19452 -1588 -19348 -1292
rect -20041 -1640 -19719 -1639
rect -20041 -1960 -20040 -1640
rect -19720 -1960 -19719 -1640
rect -20041 -1961 -19719 -1960
rect -20464 -2308 -20360 -2012
rect -21053 -2360 -20731 -2359
rect -21053 -2680 -21052 -2360
rect -20732 -2680 -20731 -2360
rect -21053 -2681 -20731 -2680
rect -21476 -3028 -21372 -2732
rect -22065 -3080 -21743 -3079
rect -22065 -3400 -22064 -3080
rect -21744 -3400 -21743 -3080
rect -22065 -3401 -21743 -3400
rect -22488 -3748 -22384 -3452
rect -23077 -3800 -22755 -3799
rect -23077 -4120 -23076 -3800
rect -22756 -4120 -22755 -3800
rect -23077 -4121 -22755 -4120
rect -23500 -4468 -23396 -4172
rect -24089 -4520 -23767 -4519
rect -24089 -4840 -24088 -4520
rect -23768 -4840 -23767 -4520
rect -24089 -4841 -23767 -4840
rect -24512 -5188 -24408 -4892
rect -25101 -5240 -24779 -5239
rect -25101 -5560 -25100 -5240
rect -24780 -5560 -24779 -5240
rect -25101 -5561 -24779 -5560
rect -25524 -5760 -25420 -5612
rect -24992 -5760 -24888 -5561
rect -24512 -5612 -24492 -5188
rect -24428 -5612 -24408 -5188
rect -23980 -5239 -23876 -4841
rect -23500 -4892 -23480 -4468
rect -23416 -4892 -23396 -4468
rect -22968 -4519 -22864 -4121
rect -22488 -4172 -22468 -3748
rect -22404 -4172 -22384 -3748
rect -21956 -3799 -21852 -3401
rect -21476 -3452 -21456 -3028
rect -21392 -3452 -21372 -3028
rect -20944 -3079 -20840 -2681
rect -20464 -2732 -20444 -2308
rect -20380 -2732 -20360 -2308
rect -19932 -2359 -19828 -1961
rect -19452 -2012 -19432 -1588
rect -19368 -2012 -19348 -1588
rect -18920 -1639 -18816 -1241
rect -18440 -1292 -18420 -868
rect -18356 -1292 -18336 -868
rect -17908 -919 -17804 -521
rect -17428 -572 -17408 -148
rect -17344 -572 -17324 -148
rect -16896 -199 -16792 199
rect -16416 148 -16396 572
rect -16332 148 -16312 572
rect -15884 521 -15780 919
rect -15404 868 -15384 1292
rect -15320 868 -15300 1292
rect -14872 1241 -14768 1639
rect -14392 1588 -14372 2012
rect -14308 1588 -14288 2012
rect -13860 1961 -13756 2359
rect -13380 2308 -13360 2732
rect -13296 2308 -13276 2732
rect -12848 2681 -12744 3079
rect -12368 3028 -12348 3452
rect -12284 3028 -12264 3452
rect -11836 3401 -11732 3799
rect -11356 3748 -11336 4172
rect -11272 3748 -11252 4172
rect -10824 4121 -10720 4519
rect -10344 4468 -10324 4892
rect -10260 4468 -10240 4892
rect -9812 4841 -9708 5239
rect -9332 5188 -9312 5612
rect -9248 5188 -9228 5612
rect -8800 5561 -8696 5760
rect -8320 5612 -8216 5760
rect -8909 5560 -8587 5561
rect -8909 5240 -8908 5560
rect -8588 5240 -8587 5560
rect -8909 5239 -8587 5240
rect -9332 4892 -9228 5188
rect -9921 4840 -9599 4841
rect -9921 4520 -9920 4840
rect -9600 4520 -9599 4840
rect -9921 4519 -9599 4520
rect -10344 4172 -10240 4468
rect -10933 4120 -10611 4121
rect -10933 3800 -10932 4120
rect -10612 3800 -10611 4120
rect -10933 3799 -10611 3800
rect -11356 3452 -11252 3748
rect -11945 3400 -11623 3401
rect -11945 3080 -11944 3400
rect -11624 3080 -11623 3400
rect -11945 3079 -11623 3080
rect -12368 2732 -12264 3028
rect -12957 2680 -12635 2681
rect -12957 2360 -12956 2680
rect -12636 2360 -12635 2680
rect -12957 2359 -12635 2360
rect -13380 2012 -13276 2308
rect -13969 1960 -13647 1961
rect -13969 1640 -13968 1960
rect -13648 1640 -13647 1960
rect -13969 1639 -13647 1640
rect -14392 1292 -14288 1588
rect -14981 1240 -14659 1241
rect -14981 920 -14980 1240
rect -14660 920 -14659 1240
rect -14981 919 -14659 920
rect -15404 572 -15300 868
rect -15993 520 -15671 521
rect -15993 200 -15992 520
rect -15672 200 -15671 520
rect -15993 199 -15671 200
rect -16416 -148 -16312 148
rect -17005 -200 -16683 -199
rect -17005 -520 -17004 -200
rect -16684 -520 -16683 -200
rect -17005 -521 -16683 -520
rect -17428 -868 -17324 -572
rect -18017 -920 -17695 -919
rect -18017 -1240 -18016 -920
rect -17696 -1240 -17695 -920
rect -18017 -1241 -17695 -1240
rect -18440 -1588 -18336 -1292
rect -19029 -1640 -18707 -1639
rect -19029 -1960 -19028 -1640
rect -18708 -1960 -18707 -1640
rect -19029 -1961 -18707 -1960
rect -19452 -2308 -19348 -2012
rect -20041 -2360 -19719 -2359
rect -20041 -2680 -20040 -2360
rect -19720 -2680 -19719 -2360
rect -20041 -2681 -19719 -2680
rect -20464 -3028 -20360 -2732
rect -21053 -3080 -20731 -3079
rect -21053 -3400 -21052 -3080
rect -20732 -3400 -20731 -3080
rect -21053 -3401 -20731 -3400
rect -21476 -3748 -21372 -3452
rect -22065 -3800 -21743 -3799
rect -22065 -4120 -22064 -3800
rect -21744 -4120 -21743 -3800
rect -22065 -4121 -21743 -4120
rect -22488 -4468 -22384 -4172
rect -23077 -4520 -22755 -4519
rect -23077 -4840 -23076 -4520
rect -22756 -4840 -22755 -4520
rect -23077 -4841 -22755 -4840
rect -23500 -5188 -23396 -4892
rect -24089 -5240 -23767 -5239
rect -24089 -5560 -24088 -5240
rect -23768 -5560 -23767 -5240
rect -24089 -5561 -23767 -5560
rect -24512 -5760 -24408 -5612
rect -23980 -5760 -23876 -5561
rect -23500 -5612 -23480 -5188
rect -23416 -5612 -23396 -5188
rect -22968 -5239 -22864 -4841
rect -22488 -4892 -22468 -4468
rect -22404 -4892 -22384 -4468
rect -21956 -4519 -21852 -4121
rect -21476 -4172 -21456 -3748
rect -21392 -4172 -21372 -3748
rect -20944 -3799 -20840 -3401
rect -20464 -3452 -20444 -3028
rect -20380 -3452 -20360 -3028
rect -19932 -3079 -19828 -2681
rect -19452 -2732 -19432 -2308
rect -19368 -2732 -19348 -2308
rect -18920 -2359 -18816 -1961
rect -18440 -2012 -18420 -1588
rect -18356 -2012 -18336 -1588
rect -17908 -1639 -17804 -1241
rect -17428 -1292 -17408 -868
rect -17344 -1292 -17324 -868
rect -16896 -919 -16792 -521
rect -16416 -572 -16396 -148
rect -16332 -572 -16312 -148
rect -15884 -199 -15780 199
rect -15404 148 -15384 572
rect -15320 148 -15300 572
rect -14872 521 -14768 919
rect -14392 868 -14372 1292
rect -14308 868 -14288 1292
rect -13860 1241 -13756 1639
rect -13380 1588 -13360 2012
rect -13296 1588 -13276 2012
rect -12848 1961 -12744 2359
rect -12368 2308 -12348 2732
rect -12284 2308 -12264 2732
rect -11836 2681 -11732 3079
rect -11356 3028 -11336 3452
rect -11272 3028 -11252 3452
rect -10824 3401 -10720 3799
rect -10344 3748 -10324 4172
rect -10260 3748 -10240 4172
rect -9812 4121 -9708 4519
rect -9332 4468 -9312 4892
rect -9248 4468 -9228 4892
rect -8800 4841 -8696 5239
rect -8320 5188 -8300 5612
rect -8236 5188 -8216 5612
rect -7788 5561 -7684 5760
rect -7308 5612 -7204 5760
rect -7897 5560 -7575 5561
rect -7897 5240 -7896 5560
rect -7576 5240 -7575 5560
rect -7897 5239 -7575 5240
rect -8320 4892 -8216 5188
rect -8909 4840 -8587 4841
rect -8909 4520 -8908 4840
rect -8588 4520 -8587 4840
rect -8909 4519 -8587 4520
rect -9332 4172 -9228 4468
rect -9921 4120 -9599 4121
rect -9921 3800 -9920 4120
rect -9600 3800 -9599 4120
rect -9921 3799 -9599 3800
rect -10344 3452 -10240 3748
rect -10933 3400 -10611 3401
rect -10933 3080 -10932 3400
rect -10612 3080 -10611 3400
rect -10933 3079 -10611 3080
rect -11356 2732 -11252 3028
rect -11945 2680 -11623 2681
rect -11945 2360 -11944 2680
rect -11624 2360 -11623 2680
rect -11945 2359 -11623 2360
rect -12368 2012 -12264 2308
rect -12957 1960 -12635 1961
rect -12957 1640 -12956 1960
rect -12636 1640 -12635 1960
rect -12957 1639 -12635 1640
rect -13380 1292 -13276 1588
rect -13969 1240 -13647 1241
rect -13969 920 -13968 1240
rect -13648 920 -13647 1240
rect -13969 919 -13647 920
rect -14392 572 -14288 868
rect -14981 520 -14659 521
rect -14981 200 -14980 520
rect -14660 200 -14659 520
rect -14981 199 -14659 200
rect -15404 -148 -15300 148
rect -15993 -200 -15671 -199
rect -15993 -520 -15992 -200
rect -15672 -520 -15671 -200
rect -15993 -521 -15671 -520
rect -16416 -868 -16312 -572
rect -17005 -920 -16683 -919
rect -17005 -1240 -17004 -920
rect -16684 -1240 -16683 -920
rect -17005 -1241 -16683 -1240
rect -17428 -1588 -17324 -1292
rect -18017 -1640 -17695 -1639
rect -18017 -1960 -18016 -1640
rect -17696 -1960 -17695 -1640
rect -18017 -1961 -17695 -1960
rect -18440 -2308 -18336 -2012
rect -19029 -2360 -18707 -2359
rect -19029 -2680 -19028 -2360
rect -18708 -2680 -18707 -2360
rect -19029 -2681 -18707 -2680
rect -19452 -3028 -19348 -2732
rect -20041 -3080 -19719 -3079
rect -20041 -3400 -20040 -3080
rect -19720 -3400 -19719 -3080
rect -20041 -3401 -19719 -3400
rect -20464 -3748 -20360 -3452
rect -21053 -3800 -20731 -3799
rect -21053 -4120 -21052 -3800
rect -20732 -4120 -20731 -3800
rect -21053 -4121 -20731 -4120
rect -21476 -4468 -21372 -4172
rect -22065 -4520 -21743 -4519
rect -22065 -4840 -22064 -4520
rect -21744 -4840 -21743 -4520
rect -22065 -4841 -21743 -4840
rect -22488 -5188 -22384 -4892
rect -23077 -5240 -22755 -5239
rect -23077 -5560 -23076 -5240
rect -22756 -5560 -22755 -5240
rect -23077 -5561 -22755 -5560
rect -23500 -5760 -23396 -5612
rect -22968 -5760 -22864 -5561
rect -22488 -5612 -22468 -5188
rect -22404 -5612 -22384 -5188
rect -21956 -5239 -21852 -4841
rect -21476 -4892 -21456 -4468
rect -21392 -4892 -21372 -4468
rect -20944 -4519 -20840 -4121
rect -20464 -4172 -20444 -3748
rect -20380 -4172 -20360 -3748
rect -19932 -3799 -19828 -3401
rect -19452 -3452 -19432 -3028
rect -19368 -3452 -19348 -3028
rect -18920 -3079 -18816 -2681
rect -18440 -2732 -18420 -2308
rect -18356 -2732 -18336 -2308
rect -17908 -2359 -17804 -1961
rect -17428 -2012 -17408 -1588
rect -17344 -2012 -17324 -1588
rect -16896 -1639 -16792 -1241
rect -16416 -1292 -16396 -868
rect -16332 -1292 -16312 -868
rect -15884 -919 -15780 -521
rect -15404 -572 -15384 -148
rect -15320 -572 -15300 -148
rect -14872 -199 -14768 199
rect -14392 148 -14372 572
rect -14308 148 -14288 572
rect -13860 521 -13756 919
rect -13380 868 -13360 1292
rect -13296 868 -13276 1292
rect -12848 1241 -12744 1639
rect -12368 1588 -12348 2012
rect -12284 1588 -12264 2012
rect -11836 1961 -11732 2359
rect -11356 2308 -11336 2732
rect -11272 2308 -11252 2732
rect -10824 2681 -10720 3079
rect -10344 3028 -10324 3452
rect -10260 3028 -10240 3452
rect -9812 3401 -9708 3799
rect -9332 3748 -9312 4172
rect -9248 3748 -9228 4172
rect -8800 4121 -8696 4519
rect -8320 4468 -8300 4892
rect -8236 4468 -8216 4892
rect -7788 4841 -7684 5239
rect -7308 5188 -7288 5612
rect -7224 5188 -7204 5612
rect -6776 5561 -6672 5760
rect -6296 5612 -6192 5760
rect -6885 5560 -6563 5561
rect -6885 5240 -6884 5560
rect -6564 5240 -6563 5560
rect -6885 5239 -6563 5240
rect -7308 4892 -7204 5188
rect -7897 4840 -7575 4841
rect -7897 4520 -7896 4840
rect -7576 4520 -7575 4840
rect -7897 4519 -7575 4520
rect -8320 4172 -8216 4468
rect -8909 4120 -8587 4121
rect -8909 3800 -8908 4120
rect -8588 3800 -8587 4120
rect -8909 3799 -8587 3800
rect -9332 3452 -9228 3748
rect -9921 3400 -9599 3401
rect -9921 3080 -9920 3400
rect -9600 3080 -9599 3400
rect -9921 3079 -9599 3080
rect -10344 2732 -10240 3028
rect -10933 2680 -10611 2681
rect -10933 2360 -10932 2680
rect -10612 2360 -10611 2680
rect -10933 2359 -10611 2360
rect -11356 2012 -11252 2308
rect -11945 1960 -11623 1961
rect -11945 1640 -11944 1960
rect -11624 1640 -11623 1960
rect -11945 1639 -11623 1640
rect -12368 1292 -12264 1588
rect -12957 1240 -12635 1241
rect -12957 920 -12956 1240
rect -12636 920 -12635 1240
rect -12957 919 -12635 920
rect -13380 572 -13276 868
rect -13969 520 -13647 521
rect -13969 200 -13968 520
rect -13648 200 -13647 520
rect -13969 199 -13647 200
rect -14392 -148 -14288 148
rect -14981 -200 -14659 -199
rect -14981 -520 -14980 -200
rect -14660 -520 -14659 -200
rect -14981 -521 -14659 -520
rect -15404 -868 -15300 -572
rect -15993 -920 -15671 -919
rect -15993 -1240 -15992 -920
rect -15672 -1240 -15671 -920
rect -15993 -1241 -15671 -1240
rect -16416 -1588 -16312 -1292
rect -17005 -1640 -16683 -1639
rect -17005 -1960 -17004 -1640
rect -16684 -1960 -16683 -1640
rect -17005 -1961 -16683 -1960
rect -17428 -2308 -17324 -2012
rect -18017 -2360 -17695 -2359
rect -18017 -2680 -18016 -2360
rect -17696 -2680 -17695 -2360
rect -18017 -2681 -17695 -2680
rect -18440 -3028 -18336 -2732
rect -19029 -3080 -18707 -3079
rect -19029 -3400 -19028 -3080
rect -18708 -3400 -18707 -3080
rect -19029 -3401 -18707 -3400
rect -19452 -3748 -19348 -3452
rect -20041 -3800 -19719 -3799
rect -20041 -4120 -20040 -3800
rect -19720 -4120 -19719 -3800
rect -20041 -4121 -19719 -4120
rect -20464 -4468 -20360 -4172
rect -21053 -4520 -20731 -4519
rect -21053 -4840 -21052 -4520
rect -20732 -4840 -20731 -4520
rect -21053 -4841 -20731 -4840
rect -21476 -5188 -21372 -4892
rect -22065 -5240 -21743 -5239
rect -22065 -5560 -22064 -5240
rect -21744 -5560 -21743 -5240
rect -22065 -5561 -21743 -5560
rect -22488 -5760 -22384 -5612
rect -21956 -5760 -21852 -5561
rect -21476 -5612 -21456 -5188
rect -21392 -5612 -21372 -5188
rect -20944 -5239 -20840 -4841
rect -20464 -4892 -20444 -4468
rect -20380 -4892 -20360 -4468
rect -19932 -4519 -19828 -4121
rect -19452 -4172 -19432 -3748
rect -19368 -4172 -19348 -3748
rect -18920 -3799 -18816 -3401
rect -18440 -3452 -18420 -3028
rect -18356 -3452 -18336 -3028
rect -17908 -3079 -17804 -2681
rect -17428 -2732 -17408 -2308
rect -17344 -2732 -17324 -2308
rect -16896 -2359 -16792 -1961
rect -16416 -2012 -16396 -1588
rect -16332 -2012 -16312 -1588
rect -15884 -1639 -15780 -1241
rect -15404 -1292 -15384 -868
rect -15320 -1292 -15300 -868
rect -14872 -919 -14768 -521
rect -14392 -572 -14372 -148
rect -14308 -572 -14288 -148
rect -13860 -199 -13756 199
rect -13380 148 -13360 572
rect -13296 148 -13276 572
rect -12848 521 -12744 919
rect -12368 868 -12348 1292
rect -12284 868 -12264 1292
rect -11836 1241 -11732 1639
rect -11356 1588 -11336 2012
rect -11272 1588 -11252 2012
rect -10824 1961 -10720 2359
rect -10344 2308 -10324 2732
rect -10260 2308 -10240 2732
rect -9812 2681 -9708 3079
rect -9332 3028 -9312 3452
rect -9248 3028 -9228 3452
rect -8800 3401 -8696 3799
rect -8320 3748 -8300 4172
rect -8236 3748 -8216 4172
rect -7788 4121 -7684 4519
rect -7308 4468 -7288 4892
rect -7224 4468 -7204 4892
rect -6776 4841 -6672 5239
rect -6296 5188 -6276 5612
rect -6212 5188 -6192 5612
rect -5764 5561 -5660 5760
rect -5284 5612 -5180 5760
rect -5873 5560 -5551 5561
rect -5873 5240 -5872 5560
rect -5552 5240 -5551 5560
rect -5873 5239 -5551 5240
rect -6296 4892 -6192 5188
rect -6885 4840 -6563 4841
rect -6885 4520 -6884 4840
rect -6564 4520 -6563 4840
rect -6885 4519 -6563 4520
rect -7308 4172 -7204 4468
rect -7897 4120 -7575 4121
rect -7897 3800 -7896 4120
rect -7576 3800 -7575 4120
rect -7897 3799 -7575 3800
rect -8320 3452 -8216 3748
rect -8909 3400 -8587 3401
rect -8909 3080 -8908 3400
rect -8588 3080 -8587 3400
rect -8909 3079 -8587 3080
rect -9332 2732 -9228 3028
rect -9921 2680 -9599 2681
rect -9921 2360 -9920 2680
rect -9600 2360 -9599 2680
rect -9921 2359 -9599 2360
rect -10344 2012 -10240 2308
rect -10933 1960 -10611 1961
rect -10933 1640 -10932 1960
rect -10612 1640 -10611 1960
rect -10933 1639 -10611 1640
rect -11356 1292 -11252 1588
rect -11945 1240 -11623 1241
rect -11945 920 -11944 1240
rect -11624 920 -11623 1240
rect -11945 919 -11623 920
rect -12368 572 -12264 868
rect -12957 520 -12635 521
rect -12957 200 -12956 520
rect -12636 200 -12635 520
rect -12957 199 -12635 200
rect -13380 -148 -13276 148
rect -13969 -200 -13647 -199
rect -13969 -520 -13968 -200
rect -13648 -520 -13647 -200
rect -13969 -521 -13647 -520
rect -14392 -868 -14288 -572
rect -14981 -920 -14659 -919
rect -14981 -1240 -14980 -920
rect -14660 -1240 -14659 -920
rect -14981 -1241 -14659 -1240
rect -15404 -1588 -15300 -1292
rect -15993 -1640 -15671 -1639
rect -15993 -1960 -15992 -1640
rect -15672 -1960 -15671 -1640
rect -15993 -1961 -15671 -1960
rect -16416 -2308 -16312 -2012
rect -17005 -2360 -16683 -2359
rect -17005 -2680 -17004 -2360
rect -16684 -2680 -16683 -2360
rect -17005 -2681 -16683 -2680
rect -17428 -3028 -17324 -2732
rect -18017 -3080 -17695 -3079
rect -18017 -3400 -18016 -3080
rect -17696 -3400 -17695 -3080
rect -18017 -3401 -17695 -3400
rect -18440 -3748 -18336 -3452
rect -19029 -3800 -18707 -3799
rect -19029 -4120 -19028 -3800
rect -18708 -4120 -18707 -3800
rect -19029 -4121 -18707 -4120
rect -19452 -4468 -19348 -4172
rect -20041 -4520 -19719 -4519
rect -20041 -4840 -20040 -4520
rect -19720 -4840 -19719 -4520
rect -20041 -4841 -19719 -4840
rect -20464 -5188 -20360 -4892
rect -21053 -5240 -20731 -5239
rect -21053 -5560 -21052 -5240
rect -20732 -5560 -20731 -5240
rect -21053 -5561 -20731 -5560
rect -21476 -5760 -21372 -5612
rect -20944 -5760 -20840 -5561
rect -20464 -5612 -20444 -5188
rect -20380 -5612 -20360 -5188
rect -19932 -5239 -19828 -4841
rect -19452 -4892 -19432 -4468
rect -19368 -4892 -19348 -4468
rect -18920 -4519 -18816 -4121
rect -18440 -4172 -18420 -3748
rect -18356 -4172 -18336 -3748
rect -17908 -3799 -17804 -3401
rect -17428 -3452 -17408 -3028
rect -17344 -3452 -17324 -3028
rect -16896 -3079 -16792 -2681
rect -16416 -2732 -16396 -2308
rect -16332 -2732 -16312 -2308
rect -15884 -2359 -15780 -1961
rect -15404 -2012 -15384 -1588
rect -15320 -2012 -15300 -1588
rect -14872 -1639 -14768 -1241
rect -14392 -1292 -14372 -868
rect -14308 -1292 -14288 -868
rect -13860 -919 -13756 -521
rect -13380 -572 -13360 -148
rect -13296 -572 -13276 -148
rect -12848 -199 -12744 199
rect -12368 148 -12348 572
rect -12284 148 -12264 572
rect -11836 521 -11732 919
rect -11356 868 -11336 1292
rect -11272 868 -11252 1292
rect -10824 1241 -10720 1639
rect -10344 1588 -10324 2012
rect -10260 1588 -10240 2012
rect -9812 1961 -9708 2359
rect -9332 2308 -9312 2732
rect -9248 2308 -9228 2732
rect -8800 2681 -8696 3079
rect -8320 3028 -8300 3452
rect -8236 3028 -8216 3452
rect -7788 3401 -7684 3799
rect -7308 3748 -7288 4172
rect -7224 3748 -7204 4172
rect -6776 4121 -6672 4519
rect -6296 4468 -6276 4892
rect -6212 4468 -6192 4892
rect -5764 4841 -5660 5239
rect -5284 5188 -5264 5612
rect -5200 5188 -5180 5612
rect -4752 5561 -4648 5760
rect -4272 5612 -4168 5760
rect -4861 5560 -4539 5561
rect -4861 5240 -4860 5560
rect -4540 5240 -4539 5560
rect -4861 5239 -4539 5240
rect -5284 4892 -5180 5188
rect -5873 4840 -5551 4841
rect -5873 4520 -5872 4840
rect -5552 4520 -5551 4840
rect -5873 4519 -5551 4520
rect -6296 4172 -6192 4468
rect -6885 4120 -6563 4121
rect -6885 3800 -6884 4120
rect -6564 3800 -6563 4120
rect -6885 3799 -6563 3800
rect -7308 3452 -7204 3748
rect -7897 3400 -7575 3401
rect -7897 3080 -7896 3400
rect -7576 3080 -7575 3400
rect -7897 3079 -7575 3080
rect -8320 2732 -8216 3028
rect -8909 2680 -8587 2681
rect -8909 2360 -8908 2680
rect -8588 2360 -8587 2680
rect -8909 2359 -8587 2360
rect -9332 2012 -9228 2308
rect -9921 1960 -9599 1961
rect -9921 1640 -9920 1960
rect -9600 1640 -9599 1960
rect -9921 1639 -9599 1640
rect -10344 1292 -10240 1588
rect -10933 1240 -10611 1241
rect -10933 920 -10932 1240
rect -10612 920 -10611 1240
rect -10933 919 -10611 920
rect -11356 572 -11252 868
rect -11945 520 -11623 521
rect -11945 200 -11944 520
rect -11624 200 -11623 520
rect -11945 199 -11623 200
rect -12368 -148 -12264 148
rect -12957 -200 -12635 -199
rect -12957 -520 -12956 -200
rect -12636 -520 -12635 -200
rect -12957 -521 -12635 -520
rect -13380 -868 -13276 -572
rect -13969 -920 -13647 -919
rect -13969 -1240 -13968 -920
rect -13648 -1240 -13647 -920
rect -13969 -1241 -13647 -1240
rect -14392 -1588 -14288 -1292
rect -14981 -1640 -14659 -1639
rect -14981 -1960 -14980 -1640
rect -14660 -1960 -14659 -1640
rect -14981 -1961 -14659 -1960
rect -15404 -2308 -15300 -2012
rect -15993 -2360 -15671 -2359
rect -15993 -2680 -15992 -2360
rect -15672 -2680 -15671 -2360
rect -15993 -2681 -15671 -2680
rect -16416 -3028 -16312 -2732
rect -17005 -3080 -16683 -3079
rect -17005 -3400 -17004 -3080
rect -16684 -3400 -16683 -3080
rect -17005 -3401 -16683 -3400
rect -17428 -3748 -17324 -3452
rect -18017 -3800 -17695 -3799
rect -18017 -4120 -18016 -3800
rect -17696 -4120 -17695 -3800
rect -18017 -4121 -17695 -4120
rect -18440 -4468 -18336 -4172
rect -19029 -4520 -18707 -4519
rect -19029 -4840 -19028 -4520
rect -18708 -4840 -18707 -4520
rect -19029 -4841 -18707 -4840
rect -19452 -5188 -19348 -4892
rect -20041 -5240 -19719 -5239
rect -20041 -5560 -20040 -5240
rect -19720 -5560 -19719 -5240
rect -20041 -5561 -19719 -5560
rect -20464 -5760 -20360 -5612
rect -19932 -5760 -19828 -5561
rect -19452 -5612 -19432 -5188
rect -19368 -5612 -19348 -5188
rect -18920 -5239 -18816 -4841
rect -18440 -4892 -18420 -4468
rect -18356 -4892 -18336 -4468
rect -17908 -4519 -17804 -4121
rect -17428 -4172 -17408 -3748
rect -17344 -4172 -17324 -3748
rect -16896 -3799 -16792 -3401
rect -16416 -3452 -16396 -3028
rect -16332 -3452 -16312 -3028
rect -15884 -3079 -15780 -2681
rect -15404 -2732 -15384 -2308
rect -15320 -2732 -15300 -2308
rect -14872 -2359 -14768 -1961
rect -14392 -2012 -14372 -1588
rect -14308 -2012 -14288 -1588
rect -13860 -1639 -13756 -1241
rect -13380 -1292 -13360 -868
rect -13296 -1292 -13276 -868
rect -12848 -919 -12744 -521
rect -12368 -572 -12348 -148
rect -12284 -572 -12264 -148
rect -11836 -199 -11732 199
rect -11356 148 -11336 572
rect -11272 148 -11252 572
rect -10824 521 -10720 919
rect -10344 868 -10324 1292
rect -10260 868 -10240 1292
rect -9812 1241 -9708 1639
rect -9332 1588 -9312 2012
rect -9248 1588 -9228 2012
rect -8800 1961 -8696 2359
rect -8320 2308 -8300 2732
rect -8236 2308 -8216 2732
rect -7788 2681 -7684 3079
rect -7308 3028 -7288 3452
rect -7224 3028 -7204 3452
rect -6776 3401 -6672 3799
rect -6296 3748 -6276 4172
rect -6212 3748 -6192 4172
rect -5764 4121 -5660 4519
rect -5284 4468 -5264 4892
rect -5200 4468 -5180 4892
rect -4752 4841 -4648 5239
rect -4272 5188 -4252 5612
rect -4188 5188 -4168 5612
rect -3740 5561 -3636 5760
rect -3260 5612 -3156 5760
rect -3849 5560 -3527 5561
rect -3849 5240 -3848 5560
rect -3528 5240 -3527 5560
rect -3849 5239 -3527 5240
rect -4272 4892 -4168 5188
rect -4861 4840 -4539 4841
rect -4861 4520 -4860 4840
rect -4540 4520 -4539 4840
rect -4861 4519 -4539 4520
rect -5284 4172 -5180 4468
rect -5873 4120 -5551 4121
rect -5873 3800 -5872 4120
rect -5552 3800 -5551 4120
rect -5873 3799 -5551 3800
rect -6296 3452 -6192 3748
rect -6885 3400 -6563 3401
rect -6885 3080 -6884 3400
rect -6564 3080 -6563 3400
rect -6885 3079 -6563 3080
rect -7308 2732 -7204 3028
rect -7897 2680 -7575 2681
rect -7897 2360 -7896 2680
rect -7576 2360 -7575 2680
rect -7897 2359 -7575 2360
rect -8320 2012 -8216 2308
rect -8909 1960 -8587 1961
rect -8909 1640 -8908 1960
rect -8588 1640 -8587 1960
rect -8909 1639 -8587 1640
rect -9332 1292 -9228 1588
rect -9921 1240 -9599 1241
rect -9921 920 -9920 1240
rect -9600 920 -9599 1240
rect -9921 919 -9599 920
rect -10344 572 -10240 868
rect -10933 520 -10611 521
rect -10933 200 -10932 520
rect -10612 200 -10611 520
rect -10933 199 -10611 200
rect -11356 -148 -11252 148
rect -11945 -200 -11623 -199
rect -11945 -520 -11944 -200
rect -11624 -520 -11623 -200
rect -11945 -521 -11623 -520
rect -12368 -868 -12264 -572
rect -12957 -920 -12635 -919
rect -12957 -1240 -12956 -920
rect -12636 -1240 -12635 -920
rect -12957 -1241 -12635 -1240
rect -13380 -1588 -13276 -1292
rect -13969 -1640 -13647 -1639
rect -13969 -1960 -13968 -1640
rect -13648 -1960 -13647 -1640
rect -13969 -1961 -13647 -1960
rect -14392 -2308 -14288 -2012
rect -14981 -2360 -14659 -2359
rect -14981 -2680 -14980 -2360
rect -14660 -2680 -14659 -2360
rect -14981 -2681 -14659 -2680
rect -15404 -3028 -15300 -2732
rect -15993 -3080 -15671 -3079
rect -15993 -3400 -15992 -3080
rect -15672 -3400 -15671 -3080
rect -15993 -3401 -15671 -3400
rect -16416 -3748 -16312 -3452
rect -17005 -3800 -16683 -3799
rect -17005 -4120 -17004 -3800
rect -16684 -4120 -16683 -3800
rect -17005 -4121 -16683 -4120
rect -17428 -4468 -17324 -4172
rect -18017 -4520 -17695 -4519
rect -18017 -4840 -18016 -4520
rect -17696 -4840 -17695 -4520
rect -18017 -4841 -17695 -4840
rect -18440 -5188 -18336 -4892
rect -19029 -5240 -18707 -5239
rect -19029 -5560 -19028 -5240
rect -18708 -5560 -18707 -5240
rect -19029 -5561 -18707 -5560
rect -19452 -5760 -19348 -5612
rect -18920 -5760 -18816 -5561
rect -18440 -5612 -18420 -5188
rect -18356 -5612 -18336 -5188
rect -17908 -5239 -17804 -4841
rect -17428 -4892 -17408 -4468
rect -17344 -4892 -17324 -4468
rect -16896 -4519 -16792 -4121
rect -16416 -4172 -16396 -3748
rect -16332 -4172 -16312 -3748
rect -15884 -3799 -15780 -3401
rect -15404 -3452 -15384 -3028
rect -15320 -3452 -15300 -3028
rect -14872 -3079 -14768 -2681
rect -14392 -2732 -14372 -2308
rect -14308 -2732 -14288 -2308
rect -13860 -2359 -13756 -1961
rect -13380 -2012 -13360 -1588
rect -13296 -2012 -13276 -1588
rect -12848 -1639 -12744 -1241
rect -12368 -1292 -12348 -868
rect -12284 -1292 -12264 -868
rect -11836 -919 -11732 -521
rect -11356 -572 -11336 -148
rect -11272 -572 -11252 -148
rect -10824 -199 -10720 199
rect -10344 148 -10324 572
rect -10260 148 -10240 572
rect -9812 521 -9708 919
rect -9332 868 -9312 1292
rect -9248 868 -9228 1292
rect -8800 1241 -8696 1639
rect -8320 1588 -8300 2012
rect -8236 1588 -8216 2012
rect -7788 1961 -7684 2359
rect -7308 2308 -7288 2732
rect -7224 2308 -7204 2732
rect -6776 2681 -6672 3079
rect -6296 3028 -6276 3452
rect -6212 3028 -6192 3452
rect -5764 3401 -5660 3799
rect -5284 3748 -5264 4172
rect -5200 3748 -5180 4172
rect -4752 4121 -4648 4519
rect -4272 4468 -4252 4892
rect -4188 4468 -4168 4892
rect -3740 4841 -3636 5239
rect -3260 5188 -3240 5612
rect -3176 5188 -3156 5612
rect -2728 5561 -2624 5760
rect -2248 5612 -2144 5760
rect -2837 5560 -2515 5561
rect -2837 5240 -2836 5560
rect -2516 5240 -2515 5560
rect -2837 5239 -2515 5240
rect -3260 4892 -3156 5188
rect -3849 4840 -3527 4841
rect -3849 4520 -3848 4840
rect -3528 4520 -3527 4840
rect -3849 4519 -3527 4520
rect -4272 4172 -4168 4468
rect -4861 4120 -4539 4121
rect -4861 3800 -4860 4120
rect -4540 3800 -4539 4120
rect -4861 3799 -4539 3800
rect -5284 3452 -5180 3748
rect -5873 3400 -5551 3401
rect -5873 3080 -5872 3400
rect -5552 3080 -5551 3400
rect -5873 3079 -5551 3080
rect -6296 2732 -6192 3028
rect -6885 2680 -6563 2681
rect -6885 2360 -6884 2680
rect -6564 2360 -6563 2680
rect -6885 2359 -6563 2360
rect -7308 2012 -7204 2308
rect -7897 1960 -7575 1961
rect -7897 1640 -7896 1960
rect -7576 1640 -7575 1960
rect -7897 1639 -7575 1640
rect -8320 1292 -8216 1588
rect -8909 1240 -8587 1241
rect -8909 920 -8908 1240
rect -8588 920 -8587 1240
rect -8909 919 -8587 920
rect -9332 572 -9228 868
rect -9921 520 -9599 521
rect -9921 200 -9920 520
rect -9600 200 -9599 520
rect -9921 199 -9599 200
rect -10344 -148 -10240 148
rect -10933 -200 -10611 -199
rect -10933 -520 -10932 -200
rect -10612 -520 -10611 -200
rect -10933 -521 -10611 -520
rect -11356 -868 -11252 -572
rect -11945 -920 -11623 -919
rect -11945 -1240 -11944 -920
rect -11624 -1240 -11623 -920
rect -11945 -1241 -11623 -1240
rect -12368 -1588 -12264 -1292
rect -12957 -1640 -12635 -1639
rect -12957 -1960 -12956 -1640
rect -12636 -1960 -12635 -1640
rect -12957 -1961 -12635 -1960
rect -13380 -2308 -13276 -2012
rect -13969 -2360 -13647 -2359
rect -13969 -2680 -13968 -2360
rect -13648 -2680 -13647 -2360
rect -13969 -2681 -13647 -2680
rect -14392 -3028 -14288 -2732
rect -14981 -3080 -14659 -3079
rect -14981 -3400 -14980 -3080
rect -14660 -3400 -14659 -3080
rect -14981 -3401 -14659 -3400
rect -15404 -3748 -15300 -3452
rect -15993 -3800 -15671 -3799
rect -15993 -4120 -15992 -3800
rect -15672 -4120 -15671 -3800
rect -15993 -4121 -15671 -4120
rect -16416 -4468 -16312 -4172
rect -17005 -4520 -16683 -4519
rect -17005 -4840 -17004 -4520
rect -16684 -4840 -16683 -4520
rect -17005 -4841 -16683 -4840
rect -17428 -5188 -17324 -4892
rect -18017 -5240 -17695 -5239
rect -18017 -5560 -18016 -5240
rect -17696 -5560 -17695 -5240
rect -18017 -5561 -17695 -5560
rect -18440 -5760 -18336 -5612
rect -17908 -5760 -17804 -5561
rect -17428 -5612 -17408 -5188
rect -17344 -5612 -17324 -5188
rect -16896 -5239 -16792 -4841
rect -16416 -4892 -16396 -4468
rect -16332 -4892 -16312 -4468
rect -15884 -4519 -15780 -4121
rect -15404 -4172 -15384 -3748
rect -15320 -4172 -15300 -3748
rect -14872 -3799 -14768 -3401
rect -14392 -3452 -14372 -3028
rect -14308 -3452 -14288 -3028
rect -13860 -3079 -13756 -2681
rect -13380 -2732 -13360 -2308
rect -13296 -2732 -13276 -2308
rect -12848 -2359 -12744 -1961
rect -12368 -2012 -12348 -1588
rect -12284 -2012 -12264 -1588
rect -11836 -1639 -11732 -1241
rect -11356 -1292 -11336 -868
rect -11272 -1292 -11252 -868
rect -10824 -919 -10720 -521
rect -10344 -572 -10324 -148
rect -10260 -572 -10240 -148
rect -9812 -199 -9708 199
rect -9332 148 -9312 572
rect -9248 148 -9228 572
rect -8800 521 -8696 919
rect -8320 868 -8300 1292
rect -8236 868 -8216 1292
rect -7788 1241 -7684 1639
rect -7308 1588 -7288 2012
rect -7224 1588 -7204 2012
rect -6776 1961 -6672 2359
rect -6296 2308 -6276 2732
rect -6212 2308 -6192 2732
rect -5764 2681 -5660 3079
rect -5284 3028 -5264 3452
rect -5200 3028 -5180 3452
rect -4752 3401 -4648 3799
rect -4272 3748 -4252 4172
rect -4188 3748 -4168 4172
rect -3740 4121 -3636 4519
rect -3260 4468 -3240 4892
rect -3176 4468 -3156 4892
rect -2728 4841 -2624 5239
rect -2248 5188 -2228 5612
rect -2164 5188 -2144 5612
rect -1716 5561 -1612 5760
rect -1236 5612 -1132 5760
rect -1825 5560 -1503 5561
rect -1825 5240 -1824 5560
rect -1504 5240 -1503 5560
rect -1825 5239 -1503 5240
rect -2248 4892 -2144 5188
rect -2837 4840 -2515 4841
rect -2837 4520 -2836 4840
rect -2516 4520 -2515 4840
rect -2837 4519 -2515 4520
rect -3260 4172 -3156 4468
rect -3849 4120 -3527 4121
rect -3849 3800 -3848 4120
rect -3528 3800 -3527 4120
rect -3849 3799 -3527 3800
rect -4272 3452 -4168 3748
rect -4861 3400 -4539 3401
rect -4861 3080 -4860 3400
rect -4540 3080 -4539 3400
rect -4861 3079 -4539 3080
rect -5284 2732 -5180 3028
rect -5873 2680 -5551 2681
rect -5873 2360 -5872 2680
rect -5552 2360 -5551 2680
rect -5873 2359 -5551 2360
rect -6296 2012 -6192 2308
rect -6885 1960 -6563 1961
rect -6885 1640 -6884 1960
rect -6564 1640 -6563 1960
rect -6885 1639 -6563 1640
rect -7308 1292 -7204 1588
rect -7897 1240 -7575 1241
rect -7897 920 -7896 1240
rect -7576 920 -7575 1240
rect -7897 919 -7575 920
rect -8320 572 -8216 868
rect -8909 520 -8587 521
rect -8909 200 -8908 520
rect -8588 200 -8587 520
rect -8909 199 -8587 200
rect -9332 -148 -9228 148
rect -9921 -200 -9599 -199
rect -9921 -520 -9920 -200
rect -9600 -520 -9599 -200
rect -9921 -521 -9599 -520
rect -10344 -868 -10240 -572
rect -10933 -920 -10611 -919
rect -10933 -1240 -10932 -920
rect -10612 -1240 -10611 -920
rect -10933 -1241 -10611 -1240
rect -11356 -1588 -11252 -1292
rect -11945 -1640 -11623 -1639
rect -11945 -1960 -11944 -1640
rect -11624 -1960 -11623 -1640
rect -11945 -1961 -11623 -1960
rect -12368 -2308 -12264 -2012
rect -12957 -2360 -12635 -2359
rect -12957 -2680 -12956 -2360
rect -12636 -2680 -12635 -2360
rect -12957 -2681 -12635 -2680
rect -13380 -3028 -13276 -2732
rect -13969 -3080 -13647 -3079
rect -13969 -3400 -13968 -3080
rect -13648 -3400 -13647 -3080
rect -13969 -3401 -13647 -3400
rect -14392 -3748 -14288 -3452
rect -14981 -3800 -14659 -3799
rect -14981 -4120 -14980 -3800
rect -14660 -4120 -14659 -3800
rect -14981 -4121 -14659 -4120
rect -15404 -4468 -15300 -4172
rect -15993 -4520 -15671 -4519
rect -15993 -4840 -15992 -4520
rect -15672 -4840 -15671 -4520
rect -15993 -4841 -15671 -4840
rect -16416 -5188 -16312 -4892
rect -17005 -5240 -16683 -5239
rect -17005 -5560 -17004 -5240
rect -16684 -5560 -16683 -5240
rect -17005 -5561 -16683 -5560
rect -17428 -5760 -17324 -5612
rect -16896 -5760 -16792 -5561
rect -16416 -5612 -16396 -5188
rect -16332 -5612 -16312 -5188
rect -15884 -5239 -15780 -4841
rect -15404 -4892 -15384 -4468
rect -15320 -4892 -15300 -4468
rect -14872 -4519 -14768 -4121
rect -14392 -4172 -14372 -3748
rect -14308 -4172 -14288 -3748
rect -13860 -3799 -13756 -3401
rect -13380 -3452 -13360 -3028
rect -13296 -3452 -13276 -3028
rect -12848 -3079 -12744 -2681
rect -12368 -2732 -12348 -2308
rect -12284 -2732 -12264 -2308
rect -11836 -2359 -11732 -1961
rect -11356 -2012 -11336 -1588
rect -11272 -2012 -11252 -1588
rect -10824 -1639 -10720 -1241
rect -10344 -1292 -10324 -868
rect -10260 -1292 -10240 -868
rect -9812 -919 -9708 -521
rect -9332 -572 -9312 -148
rect -9248 -572 -9228 -148
rect -8800 -199 -8696 199
rect -8320 148 -8300 572
rect -8236 148 -8216 572
rect -7788 521 -7684 919
rect -7308 868 -7288 1292
rect -7224 868 -7204 1292
rect -6776 1241 -6672 1639
rect -6296 1588 -6276 2012
rect -6212 1588 -6192 2012
rect -5764 1961 -5660 2359
rect -5284 2308 -5264 2732
rect -5200 2308 -5180 2732
rect -4752 2681 -4648 3079
rect -4272 3028 -4252 3452
rect -4188 3028 -4168 3452
rect -3740 3401 -3636 3799
rect -3260 3748 -3240 4172
rect -3176 3748 -3156 4172
rect -2728 4121 -2624 4519
rect -2248 4468 -2228 4892
rect -2164 4468 -2144 4892
rect -1716 4841 -1612 5239
rect -1236 5188 -1216 5612
rect -1152 5188 -1132 5612
rect -704 5561 -600 5760
rect -224 5612 -120 5760
rect -813 5560 -491 5561
rect -813 5240 -812 5560
rect -492 5240 -491 5560
rect -813 5239 -491 5240
rect -1236 4892 -1132 5188
rect -1825 4840 -1503 4841
rect -1825 4520 -1824 4840
rect -1504 4520 -1503 4840
rect -1825 4519 -1503 4520
rect -2248 4172 -2144 4468
rect -2837 4120 -2515 4121
rect -2837 3800 -2836 4120
rect -2516 3800 -2515 4120
rect -2837 3799 -2515 3800
rect -3260 3452 -3156 3748
rect -3849 3400 -3527 3401
rect -3849 3080 -3848 3400
rect -3528 3080 -3527 3400
rect -3849 3079 -3527 3080
rect -4272 2732 -4168 3028
rect -4861 2680 -4539 2681
rect -4861 2360 -4860 2680
rect -4540 2360 -4539 2680
rect -4861 2359 -4539 2360
rect -5284 2012 -5180 2308
rect -5873 1960 -5551 1961
rect -5873 1640 -5872 1960
rect -5552 1640 -5551 1960
rect -5873 1639 -5551 1640
rect -6296 1292 -6192 1588
rect -6885 1240 -6563 1241
rect -6885 920 -6884 1240
rect -6564 920 -6563 1240
rect -6885 919 -6563 920
rect -7308 572 -7204 868
rect -7897 520 -7575 521
rect -7897 200 -7896 520
rect -7576 200 -7575 520
rect -7897 199 -7575 200
rect -8320 -148 -8216 148
rect -8909 -200 -8587 -199
rect -8909 -520 -8908 -200
rect -8588 -520 -8587 -200
rect -8909 -521 -8587 -520
rect -9332 -868 -9228 -572
rect -9921 -920 -9599 -919
rect -9921 -1240 -9920 -920
rect -9600 -1240 -9599 -920
rect -9921 -1241 -9599 -1240
rect -10344 -1588 -10240 -1292
rect -10933 -1640 -10611 -1639
rect -10933 -1960 -10932 -1640
rect -10612 -1960 -10611 -1640
rect -10933 -1961 -10611 -1960
rect -11356 -2308 -11252 -2012
rect -11945 -2360 -11623 -2359
rect -11945 -2680 -11944 -2360
rect -11624 -2680 -11623 -2360
rect -11945 -2681 -11623 -2680
rect -12368 -3028 -12264 -2732
rect -12957 -3080 -12635 -3079
rect -12957 -3400 -12956 -3080
rect -12636 -3400 -12635 -3080
rect -12957 -3401 -12635 -3400
rect -13380 -3748 -13276 -3452
rect -13969 -3800 -13647 -3799
rect -13969 -4120 -13968 -3800
rect -13648 -4120 -13647 -3800
rect -13969 -4121 -13647 -4120
rect -14392 -4468 -14288 -4172
rect -14981 -4520 -14659 -4519
rect -14981 -4840 -14980 -4520
rect -14660 -4840 -14659 -4520
rect -14981 -4841 -14659 -4840
rect -15404 -5188 -15300 -4892
rect -15993 -5240 -15671 -5239
rect -15993 -5560 -15992 -5240
rect -15672 -5560 -15671 -5240
rect -15993 -5561 -15671 -5560
rect -16416 -5760 -16312 -5612
rect -15884 -5760 -15780 -5561
rect -15404 -5612 -15384 -5188
rect -15320 -5612 -15300 -5188
rect -14872 -5239 -14768 -4841
rect -14392 -4892 -14372 -4468
rect -14308 -4892 -14288 -4468
rect -13860 -4519 -13756 -4121
rect -13380 -4172 -13360 -3748
rect -13296 -4172 -13276 -3748
rect -12848 -3799 -12744 -3401
rect -12368 -3452 -12348 -3028
rect -12284 -3452 -12264 -3028
rect -11836 -3079 -11732 -2681
rect -11356 -2732 -11336 -2308
rect -11272 -2732 -11252 -2308
rect -10824 -2359 -10720 -1961
rect -10344 -2012 -10324 -1588
rect -10260 -2012 -10240 -1588
rect -9812 -1639 -9708 -1241
rect -9332 -1292 -9312 -868
rect -9248 -1292 -9228 -868
rect -8800 -919 -8696 -521
rect -8320 -572 -8300 -148
rect -8236 -572 -8216 -148
rect -7788 -199 -7684 199
rect -7308 148 -7288 572
rect -7224 148 -7204 572
rect -6776 521 -6672 919
rect -6296 868 -6276 1292
rect -6212 868 -6192 1292
rect -5764 1241 -5660 1639
rect -5284 1588 -5264 2012
rect -5200 1588 -5180 2012
rect -4752 1961 -4648 2359
rect -4272 2308 -4252 2732
rect -4188 2308 -4168 2732
rect -3740 2681 -3636 3079
rect -3260 3028 -3240 3452
rect -3176 3028 -3156 3452
rect -2728 3401 -2624 3799
rect -2248 3748 -2228 4172
rect -2164 3748 -2144 4172
rect -1716 4121 -1612 4519
rect -1236 4468 -1216 4892
rect -1152 4468 -1132 4892
rect -704 4841 -600 5239
rect -224 5188 -204 5612
rect -140 5188 -120 5612
rect 308 5561 412 5760
rect 788 5612 892 5760
rect 199 5560 521 5561
rect 199 5240 200 5560
rect 520 5240 521 5560
rect 199 5239 521 5240
rect -224 4892 -120 5188
rect -813 4840 -491 4841
rect -813 4520 -812 4840
rect -492 4520 -491 4840
rect -813 4519 -491 4520
rect -1236 4172 -1132 4468
rect -1825 4120 -1503 4121
rect -1825 3800 -1824 4120
rect -1504 3800 -1503 4120
rect -1825 3799 -1503 3800
rect -2248 3452 -2144 3748
rect -2837 3400 -2515 3401
rect -2837 3080 -2836 3400
rect -2516 3080 -2515 3400
rect -2837 3079 -2515 3080
rect -3260 2732 -3156 3028
rect -3849 2680 -3527 2681
rect -3849 2360 -3848 2680
rect -3528 2360 -3527 2680
rect -3849 2359 -3527 2360
rect -4272 2012 -4168 2308
rect -4861 1960 -4539 1961
rect -4861 1640 -4860 1960
rect -4540 1640 -4539 1960
rect -4861 1639 -4539 1640
rect -5284 1292 -5180 1588
rect -5873 1240 -5551 1241
rect -5873 920 -5872 1240
rect -5552 920 -5551 1240
rect -5873 919 -5551 920
rect -6296 572 -6192 868
rect -6885 520 -6563 521
rect -6885 200 -6884 520
rect -6564 200 -6563 520
rect -6885 199 -6563 200
rect -7308 -148 -7204 148
rect -7897 -200 -7575 -199
rect -7897 -520 -7896 -200
rect -7576 -520 -7575 -200
rect -7897 -521 -7575 -520
rect -8320 -868 -8216 -572
rect -8909 -920 -8587 -919
rect -8909 -1240 -8908 -920
rect -8588 -1240 -8587 -920
rect -8909 -1241 -8587 -1240
rect -9332 -1588 -9228 -1292
rect -9921 -1640 -9599 -1639
rect -9921 -1960 -9920 -1640
rect -9600 -1960 -9599 -1640
rect -9921 -1961 -9599 -1960
rect -10344 -2308 -10240 -2012
rect -10933 -2360 -10611 -2359
rect -10933 -2680 -10932 -2360
rect -10612 -2680 -10611 -2360
rect -10933 -2681 -10611 -2680
rect -11356 -3028 -11252 -2732
rect -11945 -3080 -11623 -3079
rect -11945 -3400 -11944 -3080
rect -11624 -3400 -11623 -3080
rect -11945 -3401 -11623 -3400
rect -12368 -3748 -12264 -3452
rect -12957 -3800 -12635 -3799
rect -12957 -4120 -12956 -3800
rect -12636 -4120 -12635 -3800
rect -12957 -4121 -12635 -4120
rect -13380 -4468 -13276 -4172
rect -13969 -4520 -13647 -4519
rect -13969 -4840 -13968 -4520
rect -13648 -4840 -13647 -4520
rect -13969 -4841 -13647 -4840
rect -14392 -5188 -14288 -4892
rect -14981 -5240 -14659 -5239
rect -14981 -5560 -14980 -5240
rect -14660 -5560 -14659 -5240
rect -14981 -5561 -14659 -5560
rect -15404 -5760 -15300 -5612
rect -14872 -5760 -14768 -5561
rect -14392 -5612 -14372 -5188
rect -14308 -5612 -14288 -5188
rect -13860 -5239 -13756 -4841
rect -13380 -4892 -13360 -4468
rect -13296 -4892 -13276 -4468
rect -12848 -4519 -12744 -4121
rect -12368 -4172 -12348 -3748
rect -12284 -4172 -12264 -3748
rect -11836 -3799 -11732 -3401
rect -11356 -3452 -11336 -3028
rect -11272 -3452 -11252 -3028
rect -10824 -3079 -10720 -2681
rect -10344 -2732 -10324 -2308
rect -10260 -2732 -10240 -2308
rect -9812 -2359 -9708 -1961
rect -9332 -2012 -9312 -1588
rect -9248 -2012 -9228 -1588
rect -8800 -1639 -8696 -1241
rect -8320 -1292 -8300 -868
rect -8236 -1292 -8216 -868
rect -7788 -919 -7684 -521
rect -7308 -572 -7288 -148
rect -7224 -572 -7204 -148
rect -6776 -199 -6672 199
rect -6296 148 -6276 572
rect -6212 148 -6192 572
rect -5764 521 -5660 919
rect -5284 868 -5264 1292
rect -5200 868 -5180 1292
rect -4752 1241 -4648 1639
rect -4272 1588 -4252 2012
rect -4188 1588 -4168 2012
rect -3740 1961 -3636 2359
rect -3260 2308 -3240 2732
rect -3176 2308 -3156 2732
rect -2728 2681 -2624 3079
rect -2248 3028 -2228 3452
rect -2164 3028 -2144 3452
rect -1716 3401 -1612 3799
rect -1236 3748 -1216 4172
rect -1152 3748 -1132 4172
rect -704 4121 -600 4519
rect -224 4468 -204 4892
rect -140 4468 -120 4892
rect 308 4841 412 5239
rect 788 5188 808 5612
rect 872 5188 892 5612
rect 1320 5561 1424 5760
rect 1800 5612 1904 5760
rect 1211 5560 1533 5561
rect 1211 5240 1212 5560
rect 1532 5240 1533 5560
rect 1211 5239 1533 5240
rect 788 4892 892 5188
rect 199 4840 521 4841
rect 199 4520 200 4840
rect 520 4520 521 4840
rect 199 4519 521 4520
rect -224 4172 -120 4468
rect -813 4120 -491 4121
rect -813 3800 -812 4120
rect -492 3800 -491 4120
rect -813 3799 -491 3800
rect -1236 3452 -1132 3748
rect -1825 3400 -1503 3401
rect -1825 3080 -1824 3400
rect -1504 3080 -1503 3400
rect -1825 3079 -1503 3080
rect -2248 2732 -2144 3028
rect -2837 2680 -2515 2681
rect -2837 2360 -2836 2680
rect -2516 2360 -2515 2680
rect -2837 2359 -2515 2360
rect -3260 2012 -3156 2308
rect -3849 1960 -3527 1961
rect -3849 1640 -3848 1960
rect -3528 1640 -3527 1960
rect -3849 1639 -3527 1640
rect -4272 1292 -4168 1588
rect -4861 1240 -4539 1241
rect -4861 920 -4860 1240
rect -4540 920 -4539 1240
rect -4861 919 -4539 920
rect -5284 572 -5180 868
rect -5873 520 -5551 521
rect -5873 200 -5872 520
rect -5552 200 -5551 520
rect -5873 199 -5551 200
rect -6296 -148 -6192 148
rect -6885 -200 -6563 -199
rect -6885 -520 -6884 -200
rect -6564 -520 -6563 -200
rect -6885 -521 -6563 -520
rect -7308 -868 -7204 -572
rect -7897 -920 -7575 -919
rect -7897 -1240 -7896 -920
rect -7576 -1240 -7575 -920
rect -7897 -1241 -7575 -1240
rect -8320 -1588 -8216 -1292
rect -8909 -1640 -8587 -1639
rect -8909 -1960 -8908 -1640
rect -8588 -1960 -8587 -1640
rect -8909 -1961 -8587 -1960
rect -9332 -2308 -9228 -2012
rect -9921 -2360 -9599 -2359
rect -9921 -2680 -9920 -2360
rect -9600 -2680 -9599 -2360
rect -9921 -2681 -9599 -2680
rect -10344 -3028 -10240 -2732
rect -10933 -3080 -10611 -3079
rect -10933 -3400 -10932 -3080
rect -10612 -3400 -10611 -3080
rect -10933 -3401 -10611 -3400
rect -11356 -3748 -11252 -3452
rect -11945 -3800 -11623 -3799
rect -11945 -4120 -11944 -3800
rect -11624 -4120 -11623 -3800
rect -11945 -4121 -11623 -4120
rect -12368 -4468 -12264 -4172
rect -12957 -4520 -12635 -4519
rect -12957 -4840 -12956 -4520
rect -12636 -4840 -12635 -4520
rect -12957 -4841 -12635 -4840
rect -13380 -5188 -13276 -4892
rect -13969 -5240 -13647 -5239
rect -13969 -5560 -13968 -5240
rect -13648 -5560 -13647 -5240
rect -13969 -5561 -13647 -5560
rect -14392 -5760 -14288 -5612
rect -13860 -5760 -13756 -5561
rect -13380 -5612 -13360 -5188
rect -13296 -5612 -13276 -5188
rect -12848 -5239 -12744 -4841
rect -12368 -4892 -12348 -4468
rect -12284 -4892 -12264 -4468
rect -11836 -4519 -11732 -4121
rect -11356 -4172 -11336 -3748
rect -11272 -4172 -11252 -3748
rect -10824 -3799 -10720 -3401
rect -10344 -3452 -10324 -3028
rect -10260 -3452 -10240 -3028
rect -9812 -3079 -9708 -2681
rect -9332 -2732 -9312 -2308
rect -9248 -2732 -9228 -2308
rect -8800 -2359 -8696 -1961
rect -8320 -2012 -8300 -1588
rect -8236 -2012 -8216 -1588
rect -7788 -1639 -7684 -1241
rect -7308 -1292 -7288 -868
rect -7224 -1292 -7204 -868
rect -6776 -919 -6672 -521
rect -6296 -572 -6276 -148
rect -6212 -572 -6192 -148
rect -5764 -199 -5660 199
rect -5284 148 -5264 572
rect -5200 148 -5180 572
rect -4752 521 -4648 919
rect -4272 868 -4252 1292
rect -4188 868 -4168 1292
rect -3740 1241 -3636 1639
rect -3260 1588 -3240 2012
rect -3176 1588 -3156 2012
rect -2728 1961 -2624 2359
rect -2248 2308 -2228 2732
rect -2164 2308 -2144 2732
rect -1716 2681 -1612 3079
rect -1236 3028 -1216 3452
rect -1152 3028 -1132 3452
rect -704 3401 -600 3799
rect -224 3748 -204 4172
rect -140 3748 -120 4172
rect 308 4121 412 4519
rect 788 4468 808 4892
rect 872 4468 892 4892
rect 1320 4841 1424 5239
rect 1800 5188 1820 5612
rect 1884 5188 1904 5612
rect 2332 5561 2436 5760
rect 2812 5612 2916 5760
rect 2223 5560 2545 5561
rect 2223 5240 2224 5560
rect 2544 5240 2545 5560
rect 2223 5239 2545 5240
rect 1800 4892 1904 5188
rect 1211 4840 1533 4841
rect 1211 4520 1212 4840
rect 1532 4520 1533 4840
rect 1211 4519 1533 4520
rect 788 4172 892 4468
rect 199 4120 521 4121
rect 199 3800 200 4120
rect 520 3800 521 4120
rect 199 3799 521 3800
rect -224 3452 -120 3748
rect -813 3400 -491 3401
rect -813 3080 -812 3400
rect -492 3080 -491 3400
rect -813 3079 -491 3080
rect -1236 2732 -1132 3028
rect -1825 2680 -1503 2681
rect -1825 2360 -1824 2680
rect -1504 2360 -1503 2680
rect -1825 2359 -1503 2360
rect -2248 2012 -2144 2308
rect -2837 1960 -2515 1961
rect -2837 1640 -2836 1960
rect -2516 1640 -2515 1960
rect -2837 1639 -2515 1640
rect -3260 1292 -3156 1588
rect -3849 1240 -3527 1241
rect -3849 920 -3848 1240
rect -3528 920 -3527 1240
rect -3849 919 -3527 920
rect -4272 572 -4168 868
rect -4861 520 -4539 521
rect -4861 200 -4860 520
rect -4540 200 -4539 520
rect -4861 199 -4539 200
rect -5284 -148 -5180 148
rect -5873 -200 -5551 -199
rect -5873 -520 -5872 -200
rect -5552 -520 -5551 -200
rect -5873 -521 -5551 -520
rect -6296 -868 -6192 -572
rect -6885 -920 -6563 -919
rect -6885 -1240 -6884 -920
rect -6564 -1240 -6563 -920
rect -6885 -1241 -6563 -1240
rect -7308 -1588 -7204 -1292
rect -7897 -1640 -7575 -1639
rect -7897 -1960 -7896 -1640
rect -7576 -1960 -7575 -1640
rect -7897 -1961 -7575 -1960
rect -8320 -2308 -8216 -2012
rect -8909 -2360 -8587 -2359
rect -8909 -2680 -8908 -2360
rect -8588 -2680 -8587 -2360
rect -8909 -2681 -8587 -2680
rect -9332 -3028 -9228 -2732
rect -9921 -3080 -9599 -3079
rect -9921 -3400 -9920 -3080
rect -9600 -3400 -9599 -3080
rect -9921 -3401 -9599 -3400
rect -10344 -3748 -10240 -3452
rect -10933 -3800 -10611 -3799
rect -10933 -4120 -10932 -3800
rect -10612 -4120 -10611 -3800
rect -10933 -4121 -10611 -4120
rect -11356 -4468 -11252 -4172
rect -11945 -4520 -11623 -4519
rect -11945 -4840 -11944 -4520
rect -11624 -4840 -11623 -4520
rect -11945 -4841 -11623 -4840
rect -12368 -5188 -12264 -4892
rect -12957 -5240 -12635 -5239
rect -12957 -5560 -12956 -5240
rect -12636 -5560 -12635 -5240
rect -12957 -5561 -12635 -5560
rect -13380 -5760 -13276 -5612
rect -12848 -5760 -12744 -5561
rect -12368 -5612 -12348 -5188
rect -12284 -5612 -12264 -5188
rect -11836 -5239 -11732 -4841
rect -11356 -4892 -11336 -4468
rect -11272 -4892 -11252 -4468
rect -10824 -4519 -10720 -4121
rect -10344 -4172 -10324 -3748
rect -10260 -4172 -10240 -3748
rect -9812 -3799 -9708 -3401
rect -9332 -3452 -9312 -3028
rect -9248 -3452 -9228 -3028
rect -8800 -3079 -8696 -2681
rect -8320 -2732 -8300 -2308
rect -8236 -2732 -8216 -2308
rect -7788 -2359 -7684 -1961
rect -7308 -2012 -7288 -1588
rect -7224 -2012 -7204 -1588
rect -6776 -1639 -6672 -1241
rect -6296 -1292 -6276 -868
rect -6212 -1292 -6192 -868
rect -5764 -919 -5660 -521
rect -5284 -572 -5264 -148
rect -5200 -572 -5180 -148
rect -4752 -199 -4648 199
rect -4272 148 -4252 572
rect -4188 148 -4168 572
rect -3740 521 -3636 919
rect -3260 868 -3240 1292
rect -3176 868 -3156 1292
rect -2728 1241 -2624 1639
rect -2248 1588 -2228 2012
rect -2164 1588 -2144 2012
rect -1716 1961 -1612 2359
rect -1236 2308 -1216 2732
rect -1152 2308 -1132 2732
rect -704 2681 -600 3079
rect -224 3028 -204 3452
rect -140 3028 -120 3452
rect 308 3401 412 3799
rect 788 3748 808 4172
rect 872 3748 892 4172
rect 1320 4121 1424 4519
rect 1800 4468 1820 4892
rect 1884 4468 1904 4892
rect 2332 4841 2436 5239
rect 2812 5188 2832 5612
rect 2896 5188 2916 5612
rect 3344 5561 3448 5760
rect 3824 5612 3928 5760
rect 3235 5560 3557 5561
rect 3235 5240 3236 5560
rect 3556 5240 3557 5560
rect 3235 5239 3557 5240
rect 2812 4892 2916 5188
rect 2223 4840 2545 4841
rect 2223 4520 2224 4840
rect 2544 4520 2545 4840
rect 2223 4519 2545 4520
rect 1800 4172 1904 4468
rect 1211 4120 1533 4121
rect 1211 3800 1212 4120
rect 1532 3800 1533 4120
rect 1211 3799 1533 3800
rect 788 3452 892 3748
rect 199 3400 521 3401
rect 199 3080 200 3400
rect 520 3080 521 3400
rect 199 3079 521 3080
rect -224 2732 -120 3028
rect -813 2680 -491 2681
rect -813 2360 -812 2680
rect -492 2360 -491 2680
rect -813 2359 -491 2360
rect -1236 2012 -1132 2308
rect -1825 1960 -1503 1961
rect -1825 1640 -1824 1960
rect -1504 1640 -1503 1960
rect -1825 1639 -1503 1640
rect -2248 1292 -2144 1588
rect -2837 1240 -2515 1241
rect -2837 920 -2836 1240
rect -2516 920 -2515 1240
rect -2837 919 -2515 920
rect -3260 572 -3156 868
rect -3849 520 -3527 521
rect -3849 200 -3848 520
rect -3528 200 -3527 520
rect -3849 199 -3527 200
rect -4272 -148 -4168 148
rect -4861 -200 -4539 -199
rect -4861 -520 -4860 -200
rect -4540 -520 -4539 -200
rect -4861 -521 -4539 -520
rect -5284 -868 -5180 -572
rect -5873 -920 -5551 -919
rect -5873 -1240 -5872 -920
rect -5552 -1240 -5551 -920
rect -5873 -1241 -5551 -1240
rect -6296 -1588 -6192 -1292
rect -6885 -1640 -6563 -1639
rect -6885 -1960 -6884 -1640
rect -6564 -1960 -6563 -1640
rect -6885 -1961 -6563 -1960
rect -7308 -2308 -7204 -2012
rect -7897 -2360 -7575 -2359
rect -7897 -2680 -7896 -2360
rect -7576 -2680 -7575 -2360
rect -7897 -2681 -7575 -2680
rect -8320 -3028 -8216 -2732
rect -8909 -3080 -8587 -3079
rect -8909 -3400 -8908 -3080
rect -8588 -3400 -8587 -3080
rect -8909 -3401 -8587 -3400
rect -9332 -3748 -9228 -3452
rect -9921 -3800 -9599 -3799
rect -9921 -4120 -9920 -3800
rect -9600 -4120 -9599 -3800
rect -9921 -4121 -9599 -4120
rect -10344 -4468 -10240 -4172
rect -10933 -4520 -10611 -4519
rect -10933 -4840 -10932 -4520
rect -10612 -4840 -10611 -4520
rect -10933 -4841 -10611 -4840
rect -11356 -5188 -11252 -4892
rect -11945 -5240 -11623 -5239
rect -11945 -5560 -11944 -5240
rect -11624 -5560 -11623 -5240
rect -11945 -5561 -11623 -5560
rect -12368 -5760 -12264 -5612
rect -11836 -5760 -11732 -5561
rect -11356 -5612 -11336 -5188
rect -11272 -5612 -11252 -5188
rect -10824 -5239 -10720 -4841
rect -10344 -4892 -10324 -4468
rect -10260 -4892 -10240 -4468
rect -9812 -4519 -9708 -4121
rect -9332 -4172 -9312 -3748
rect -9248 -4172 -9228 -3748
rect -8800 -3799 -8696 -3401
rect -8320 -3452 -8300 -3028
rect -8236 -3452 -8216 -3028
rect -7788 -3079 -7684 -2681
rect -7308 -2732 -7288 -2308
rect -7224 -2732 -7204 -2308
rect -6776 -2359 -6672 -1961
rect -6296 -2012 -6276 -1588
rect -6212 -2012 -6192 -1588
rect -5764 -1639 -5660 -1241
rect -5284 -1292 -5264 -868
rect -5200 -1292 -5180 -868
rect -4752 -919 -4648 -521
rect -4272 -572 -4252 -148
rect -4188 -572 -4168 -148
rect -3740 -199 -3636 199
rect -3260 148 -3240 572
rect -3176 148 -3156 572
rect -2728 521 -2624 919
rect -2248 868 -2228 1292
rect -2164 868 -2144 1292
rect -1716 1241 -1612 1639
rect -1236 1588 -1216 2012
rect -1152 1588 -1132 2012
rect -704 1961 -600 2359
rect -224 2308 -204 2732
rect -140 2308 -120 2732
rect 308 2681 412 3079
rect 788 3028 808 3452
rect 872 3028 892 3452
rect 1320 3401 1424 3799
rect 1800 3748 1820 4172
rect 1884 3748 1904 4172
rect 2332 4121 2436 4519
rect 2812 4468 2832 4892
rect 2896 4468 2916 4892
rect 3344 4841 3448 5239
rect 3824 5188 3844 5612
rect 3908 5188 3928 5612
rect 4356 5561 4460 5760
rect 4836 5612 4940 5760
rect 4247 5560 4569 5561
rect 4247 5240 4248 5560
rect 4568 5240 4569 5560
rect 4247 5239 4569 5240
rect 3824 4892 3928 5188
rect 3235 4840 3557 4841
rect 3235 4520 3236 4840
rect 3556 4520 3557 4840
rect 3235 4519 3557 4520
rect 2812 4172 2916 4468
rect 2223 4120 2545 4121
rect 2223 3800 2224 4120
rect 2544 3800 2545 4120
rect 2223 3799 2545 3800
rect 1800 3452 1904 3748
rect 1211 3400 1533 3401
rect 1211 3080 1212 3400
rect 1532 3080 1533 3400
rect 1211 3079 1533 3080
rect 788 2732 892 3028
rect 199 2680 521 2681
rect 199 2360 200 2680
rect 520 2360 521 2680
rect 199 2359 521 2360
rect -224 2012 -120 2308
rect -813 1960 -491 1961
rect -813 1640 -812 1960
rect -492 1640 -491 1960
rect -813 1639 -491 1640
rect -1236 1292 -1132 1588
rect -1825 1240 -1503 1241
rect -1825 920 -1824 1240
rect -1504 920 -1503 1240
rect -1825 919 -1503 920
rect -2248 572 -2144 868
rect -2837 520 -2515 521
rect -2837 200 -2836 520
rect -2516 200 -2515 520
rect -2837 199 -2515 200
rect -3260 -148 -3156 148
rect -3849 -200 -3527 -199
rect -3849 -520 -3848 -200
rect -3528 -520 -3527 -200
rect -3849 -521 -3527 -520
rect -4272 -868 -4168 -572
rect -4861 -920 -4539 -919
rect -4861 -1240 -4860 -920
rect -4540 -1240 -4539 -920
rect -4861 -1241 -4539 -1240
rect -5284 -1588 -5180 -1292
rect -5873 -1640 -5551 -1639
rect -5873 -1960 -5872 -1640
rect -5552 -1960 -5551 -1640
rect -5873 -1961 -5551 -1960
rect -6296 -2308 -6192 -2012
rect -6885 -2360 -6563 -2359
rect -6885 -2680 -6884 -2360
rect -6564 -2680 -6563 -2360
rect -6885 -2681 -6563 -2680
rect -7308 -3028 -7204 -2732
rect -7897 -3080 -7575 -3079
rect -7897 -3400 -7896 -3080
rect -7576 -3400 -7575 -3080
rect -7897 -3401 -7575 -3400
rect -8320 -3748 -8216 -3452
rect -8909 -3800 -8587 -3799
rect -8909 -4120 -8908 -3800
rect -8588 -4120 -8587 -3800
rect -8909 -4121 -8587 -4120
rect -9332 -4468 -9228 -4172
rect -9921 -4520 -9599 -4519
rect -9921 -4840 -9920 -4520
rect -9600 -4840 -9599 -4520
rect -9921 -4841 -9599 -4840
rect -10344 -5188 -10240 -4892
rect -10933 -5240 -10611 -5239
rect -10933 -5560 -10932 -5240
rect -10612 -5560 -10611 -5240
rect -10933 -5561 -10611 -5560
rect -11356 -5760 -11252 -5612
rect -10824 -5760 -10720 -5561
rect -10344 -5612 -10324 -5188
rect -10260 -5612 -10240 -5188
rect -9812 -5239 -9708 -4841
rect -9332 -4892 -9312 -4468
rect -9248 -4892 -9228 -4468
rect -8800 -4519 -8696 -4121
rect -8320 -4172 -8300 -3748
rect -8236 -4172 -8216 -3748
rect -7788 -3799 -7684 -3401
rect -7308 -3452 -7288 -3028
rect -7224 -3452 -7204 -3028
rect -6776 -3079 -6672 -2681
rect -6296 -2732 -6276 -2308
rect -6212 -2732 -6192 -2308
rect -5764 -2359 -5660 -1961
rect -5284 -2012 -5264 -1588
rect -5200 -2012 -5180 -1588
rect -4752 -1639 -4648 -1241
rect -4272 -1292 -4252 -868
rect -4188 -1292 -4168 -868
rect -3740 -919 -3636 -521
rect -3260 -572 -3240 -148
rect -3176 -572 -3156 -148
rect -2728 -199 -2624 199
rect -2248 148 -2228 572
rect -2164 148 -2144 572
rect -1716 521 -1612 919
rect -1236 868 -1216 1292
rect -1152 868 -1132 1292
rect -704 1241 -600 1639
rect -224 1588 -204 2012
rect -140 1588 -120 2012
rect 308 1961 412 2359
rect 788 2308 808 2732
rect 872 2308 892 2732
rect 1320 2681 1424 3079
rect 1800 3028 1820 3452
rect 1884 3028 1904 3452
rect 2332 3401 2436 3799
rect 2812 3748 2832 4172
rect 2896 3748 2916 4172
rect 3344 4121 3448 4519
rect 3824 4468 3844 4892
rect 3908 4468 3928 4892
rect 4356 4841 4460 5239
rect 4836 5188 4856 5612
rect 4920 5188 4940 5612
rect 5368 5561 5472 5760
rect 5848 5612 5952 5760
rect 5259 5560 5581 5561
rect 5259 5240 5260 5560
rect 5580 5240 5581 5560
rect 5259 5239 5581 5240
rect 4836 4892 4940 5188
rect 4247 4840 4569 4841
rect 4247 4520 4248 4840
rect 4568 4520 4569 4840
rect 4247 4519 4569 4520
rect 3824 4172 3928 4468
rect 3235 4120 3557 4121
rect 3235 3800 3236 4120
rect 3556 3800 3557 4120
rect 3235 3799 3557 3800
rect 2812 3452 2916 3748
rect 2223 3400 2545 3401
rect 2223 3080 2224 3400
rect 2544 3080 2545 3400
rect 2223 3079 2545 3080
rect 1800 2732 1904 3028
rect 1211 2680 1533 2681
rect 1211 2360 1212 2680
rect 1532 2360 1533 2680
rect 1211 2359 1533 2360
rect 788 2012 892 2308
rect 199 1960 521 1961
rect 199 1640 200 1960
rect 520 1640 521 1960
rect 199 1639 521 1640
rect -224 1292 -120 1588
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -1236 572 -1132 868
rect -1825 520 -1503 521
rect -1825 200 -1824 520
rect -1504 200 -1503 520
rect -1825 199 -1503 200
rect -2248 -148 -2144 148
rect -2837 -200 -2515 -199
rect -2837 -520 -2836 -200
rect -2516 -520 -2515 -200
rect -2837 -521 -2515 -520
rect -3260 -868 -3156 -572
rect -3849 -920 -3527 -919
rect -3849 -1240 -3848 -920
rect -3528 -1240 -3527 -920
rect -3849 -1241 -3527 -1240
rect -4272 -1588 -4168 -1292
rect -4861 -1640 -4539 -1639
rect -4861 -1960 -4860 -1640
rect -4540 -1960 -4539 -1640
rect -4861 -1961 -4539 -1960
rect -5284 -2308 -5180 -2012
rect -5873 -2360 -5551 -2359
rect -5873 -2680 -5872 -2360
rect -5552 -2680 -5551 -2360
rect -5873 -2681 -5551 -2680
rect -6296 -3028 -6192 -2732
rect -6885 -3080 -6563 -3079
rect -6885 -3400 -6884 -3080
rect -6564 -3400 -6563 -3080
rect -6885 -3401 -6563 -3400
rect -7308 -3748 -7204 -3452
rect -7897 -3800 -7575 -3799
rect -7897 -4120 -7896 -3800
rect -7576 -4120 -7575 -3800
rect -7897 -4121 -7575 -4120
rect -8320 -4468 -8216 -4172
rect -8909 -4520 -8587 -4519
rect -8909 -4840 -8908 -4520
rect -8588 -4840 -8587 -4520
rect -8909 -4841 -8587 -4840
rect -9332 -5188 -9228 -4892
rect -9921 -5240 -9599 -5239
rect -9921 -5560 -9920 -5240
rect -9600 -5560 -9599 -5240
rect -9921 -5561 -9599 -5560
rect -10344 -5760 -10240 -5612
rect -9812 -5760 -9708 -5561
rect -9332 -5612 -9312 -5188
rect -9248 -5612 -9228 -5188
rect -8800 -5239 -8696 -4841
rect -8320 -4892 -8300 -4468
rect -8236 -4892 -8216 -4468
rect -7788 -4519 -7684 -4121
rect -7308 -4172 -7288 -3748
rect -7224 -4172 -7204 -3748
rect -6776 -3799 -6672 -3401
rect -6296 -3452 -6276 -3028
rect -6212 -3452 -6192 -3028
rect -5764 -3079 -5660 -2681
rect -5284 -2732 -5264 -2308
rect -5200 -2732 -5180 -2308
rect -4752 -2359 -4648 -1961
rect -4272 -2012 -4252 -1588
rect -4188 -2012 -4168 -1588
rect -3740 -1639 -3636 -1241
rect -3260 -1292 -3240 -868
rect -3176 -1292 -3156 -868
rect -2728 -919 -2624 -521
rect -2248 -572 -2228 -148
rect -2164 -572 -2144 -148
rect -1716 -199 -1612 199
rect -1236 148 -1216 572
rect -1152 148 -1132 572
rect -704 521 -600 919
rect -224 868 -204 1292
rect -140 868 -120 1292
rect 308 1241 412 1639
rect 788 1588 808 2012
rect 872 1588 892 2012
rect 1320 1961 1424 2359
rect 1800 2308 1820 2732
rect 1884 2308 1904 2732
rect 2332 2681 2436 3079
rect 2812 3028 2832 3452
rect 2896 3028 2916 3452
rect 3344 3401 3448 3799
rect 3824 3748 3844 4172
rect 3908 3748 3928 4172
rect 4356 4121 4460 4519
rect 4836 4468 4856 4892
rect 4920 4468 4940 4892
rect 5368 4841 5472 5239
rect 5848 5188 5868 5612
rect 5932 5188 5952 5612
rect 6380 5561 6484 5760
rect 6860 5612 6964 5760
rect 6271 5560 6593 5561
rect 6271 5240 6272 5560
rect 6592 5240 6593 5560
rect 6271 5239 6593 5240
rect 5848 4892 5952 5188
rect 5259 4840 5581 4841
rect 5259 4520 5260 4840
rect 5580 4520 5581 4840
rect 5259 4519 5581 4520
rect 4836 4172 4940 4468
rect 4247 4120 4569 4121
rect 4247 3800 4248 4120
rect 4568 3800 4569 4120
rect 4247 3799 4569 3800
rect 3824 3452 3928 3748
rect 3235 3400 3557 3401
rect 3235 3080 3236 3400
rect 3556 3080 3557 3400
rect 3235 3079 3557 3080
rect 2812 2732 2916 3028
rect 2223 2680 2545 2681
rect 2223 2360 2224 2680
rect 2544 2360 2545 2680
rect 2223 2359 2545 2360
rect 1800 2012 1904 2308
rect 1211 1960 1533 1961
rect 1211 1640 1212 1960
rect 1532 1640 1533 1960
rect 1211 1639 1533 1640
rect 788 1292 892 1588
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -224 572 -120 868
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -1236 -148 -1132 148
rect -1825 -200 -1503 -199
rect -1825 -520 -1824 -200
rect -1504 -520 -1503 -200
rect -1825 -521 -1503 -520
rect -2248 -868 -2144 -572
rect -2837 -920 -2515 -919
rect -2837 -1240 -2836 -920
rect -2516 -1240 -2515 -920
rect -2837 -1241 -2515 -1240
rect -3260 -1588 -3156 -1292
rect -3849 -1640 -3527 -1639
rect -3849 -1960 -3848 -1640
rect -3528 -1960 -3527 -1640
rect -3849 -1961 -3527 -1960
rect -4272 -2308 -4168 -2012
rect -4861 -2360 -4539 -2359
rect -4861 -2680 -4860 -2360
rect -4540 -2680 -4539 -2360
rect -4861 -2681 -4539 -2680
rect -5284 -3028 -5180 -2732
rect -5873 -3080 -5551 -3079
rect -5873 -3400 -5872 -3080
rect -5552 -3400 -5551 -3080
rect -5873 -3401 -5551 -3400
rect -6296 -3748 -6192 -3452
rect -6885 -3800 -6563 -3799
rect -6885 -4120 -6884 -3800
rect -6564 -4120 -6563 -3800
rect -6885 -4121 -6563 -4120
rect -7308 -4468 -7204 -4172
rect -7897 -4520 -7575 -4519
rect -7897 -4840 -7896 -4520
rect -7576 -4840 -7575 -4520
rect -7897 -4841 -7575 -4840
rect -8320 -5188 -8216 -4892
rect -8909 -5240 -8587 -5239
rect -8909 -5560 -8908 -5240
rect -8588 -5560 -8587 -5240
rect -8909 -5561 -8587 -5560
rect -9332 -5760 -9228 -5612
rect -8800 -5760 -8696 -5561
rect -8320 -5612 -8300 -5188
rect -8236 -5612 -8216 -5188
rect -7788 -5239 -7684 -4841
rect -7308 -4892 -7288 -4468
rect -7224 -4892 -7204 -4468
rect -6776 -4519 -6672 -4121
rect -6296 -4172 -6276 -3748
rect -6212 -4172 -6192 -3748
rect -5764 -3799 -5660 -3401
rect -5284 -3452 -5264 -3028
rect -5200 -3452 -5180 -3028
rect -4752 -3079 -4648 -2681
rect -4272 -2732 -4252 -2308
rect -4188 -2732 -4168 -2308
rect -3740 -2359 -3636 -1961
rect -3260 -2012 -3240 -1588
rect -3176 -2012 -3156 -1588
rect -2728 -1639 -2624 -1241
rect -2248 -1292 -2228 -868
rect -2164 -1292 -2144 -868
rect -1716 -919 -1612 -521
rect -1236 -572 -1216 -148
rect -1152 -572 -1132 -148
rect -704 -199 -600 199
rect -224 148 -204 572
rect -140 148 -120 572
rect 308 521 412 919
rect 788 868 808 1292
rect 872 868 892 1292
rect 1320 1241 1424 1639
rect 1800 1588 1820 2012
rect 1884 1588 1904 2012
rect 2332 1961 2436 2359
rect 2812 2308 2832 2732
rect 2896 2308 2916 2732
rect 3344 2681 3448 3079
rect 3824 3028 3844 3452
rect 3908 3028 3928 3452
rect 4356 3401 4460 3799
rect 4836 3748 4856 4172
rect 4920 3748 4940 4172
rect 5368 4121 5472 4519
rect 5848 4468 5868 4892
rect 5932 4468 5952 4892
rect 6380 4841 6484 5239
rect 6860 5188 6880 5612
rect 6944 5188 6964 5612
rect 7392 5561 7496 5760
rect 7872 5612 7976 5760
rect 7283 5560 7605 5561
rect 7283 5240 7284 5560
rect 7604 5240 7605 5560
rect 7283 5239 7605 5240
rect 6860 4892 6964 5188
rect 6271 4840 6593 4841
rect 6271 4520 6272 4840
rect 6592 4520 6593 4840
rect 6271 4519 6593 4520
rect 5848 4172 5952 4468
rect 5259 4120 5581 4121
rect 5259 3800 5260 4120
rect 5580 3800 5581 4120
rect 5259 3799 5581 3800
rect 4836 3452 4940 3748
rect 4247 3400 4569 3401
rect 4247 3080 4248 3400
rect 4568 3080 4569 3400
rect 4247 3079 4569 3080
rect 3824 2732 3928 3028
rect 3235 2680 3557 2681
rect 3235 2360 3236 2680
rect 3556 2360 3557 2680
rect 3235 2359 3557 2360
rect 2812 2012 2916 2308
rect 2223 1960 2545 1961
rect 2223 1640 2224 1960
rect 2544 1640 2545 1960
rect 2223 1639 2545 1640
rect 1800 1292 1904 1588
rect 1211 1240 1533 1241
rect 1211 920 1212 1240
rect 1532 920 1533 1240
rect 1211 919 1533 920
rect 788 572 892 868
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -1236 -868 -1132 -572
rect -1825 -920 -1503 -919
rect -1825 -1240 -1824 -920
rect -1504 -1240 -1503 -920
rect -1825 -1241 -1503 -1240
rect -2248 -1588 -2144 -1292
rect -2837 -1640 -2515 -1639
rect -2837 -1960 -2836 -1640
rect -2516 -1960 -2515 -1640
rect -2837 -1961 -2515 -1960
rect -3260 -2308 -3156 -2012
rect -3849 -2360 -3527 -2359
rect -3849 -2680 -3848 -2360
rect -3528 -2680 -3527 -2360
rect -3849 -2681 -3527 -2680
rect -4272 -3028 -4168 -2732
rect -4861 -3080 -4539 -3079
rect -4861 -3400 -4860 -3080
rect -4540 -3400 -4539 -3080
rect -4861 -3401 -4539 -3400
rect -5284 -3748 -5180 -3452
rect -5873 -3800 -5551 -3799
rect -5873 -4120 -5872 -3800
rect -5552 -4120 -5551 -3800
rect -5873 -4121 -5551 -4120
rect -6296 -4468 -6192 -4172
rect -6885 -4520 -6563 -4519
rect -6885 -4840 -6884 -4520
rect -6564 -4840 -6563 -4520
rect -6885 -4841 -6563 -4840
rect -7308 -5188 -7204 -4892
rect -7897 -5240 -7575 -5239
rect -7897 -5560 -7896 -5240
rect -7576 -5560 -7575 -5240
rect -7897 -5561 -7575 -5560
rect -8320 -5760 -8216 -5612
rect -7788 -5760 -7684 -5561
rect -7308 -5612 -7288 -5188
rect -7224 -5612 -7204 -5188
rect -6776 -5239 -6672 -4841
rect -6296 -4892 -6276 -4468
rect -6212 -4892 -6192 -4468
rect -5764 -4519 -5660 -4121
rect -5284 -4172 -5264 -3748
rect -5200 -4172 -5180 -3748
rect -4752 -3799 -4648 -3401
rect -4272 -3452 -4252 -3028
rect -4188 -3452 -4168 -3028
rect -3740 -3079 -3636 -2681
rect -3260 -2732 -3240 -2308
rect -3176 -2732 -3156 -2308
rect -2728 -2359 -2624 -1961
rect -2248 -2012 -2228 -1588
rect -2164 -2012 -2144 -1588
rect -1716 -1639 -1612 -1241
rect -1236 -1292 -1216 -868
rect -1152 -1292 -1132 -868
rect -704 -919 -600 -521
rect -224 -572 -204 -148
rect -140 -572 -120 -148
rect 308 -199 412 199
rect 788 148 808 572
rect 872 148 892 572
rect 1320 521 1424 919
rect 1800 868 1820 1292
rect 1884 868 1904 1292
rect 2332 1241 2436 1639
rect 2812 1588 2832 2012
rect 2896 1588 2916 2012
rect 3344 1961 3448 2359
rect 3824 2308 3844 2732
rect 3908 2308 3928 2732
rect 4356 2681 4460 3079
rect 4836 3028 4856 3452
rect 4920 3028 4940 3452
rect 5368 3401 5472 3799
rect 5848 3748 5868 4172
rect 5932 3748 5952 4172
rect 6380 4121 6484 4519
rect 6860 4468 6880 4892
rect 6944 4468 6964 4892
rect 7392 4841 7496 5239
rect 7872 5188 7892 5612
rect 7956 5188 7976 5612
rect 8404 5561 8508 5760
rect 8884 5612 8988 5760
rect 8295 5560 8617 5561
rect 8295 5240 8296 5560
rect 8616 5240 8617 5560
rect 8295 5239 8617 5240
rect 7872 4892 7976 5188
rect 7283 4840 7605 4841
rect 7283 4520 7284 4840
rect 7604 4520 7605 4840
rect 7283 4519 7605 4520
rect 6860 4172 6964 4468
rect 6271 4120 6593 4121
rect 6271 3800 6272 4120
rect 6592 3800 6593 4120
rect 6271 3799 6593 3800
rect 5848 3452 5952 3748
rect 5259 3400 5581 3401
rect 5259 3080 5260 3400
rect 5580 3080 5581 3400
rect 5259 3079 5581 3080
rect 4836 2732 4940 3028
rect 4247 2680 4569 2681
rect 4247 2360 4248 2680
rect 4568 2360 4569 2680
rect 4247 2359 4569 2360
rect 3824 2012 3928 2308
rect 3235 1960 3557 1961
rect 3235 1640 3236 1960
rect 3556 1640 3557 1960
rect 3235 1639 3557 1640
rect 2812 1292 2916 1588
rect 2223 1240 2545 1241
rect 2223 920 2224 1240
rect 2544 920 2545 1240
rect 2223 919 2545 920
rect 1800 572 1904 868
rect 1211 520 1533 521
rect 1211 200 1212 520
rect 1532 200 1533 520
rect 1211 199 1533 200
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -224 -868 -120 -572
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -1236 -1588 -1132 -1292
rect -1825 -1640 -1503 -1639
rect -1825 -1960 -1824 -1640
rect -1504 -1960 -1503 -1640
rect -1825 -1961 -1503 -1960
rect -2248 -2308 -2144 -2012
rect -2837 -2360 -2515 -2359
rect -2837 -2680 -2836 -2360
rect -2516 -2680 -2515 -2360
rect -2837 -2681 -2515 -2680
rect -3260 -3028 -3156 -2732
rect -3849 -3080 -3527 -3079
rect -3849 -3400 -3848 -3080
rect -3528 -3400 -3527 -3080
rect -3849 -3401 -3527 -3400
rect -4272 -3748 -4168 -3452
rect -4861 -3800 -4539 -3799
rect -4861 -4120 -4860 -3800
rect -4540 -4120 -4539 -3800
rect -4861 -4121 -4539 -4120
rect -5284 -4468 -5180 -4172
rect -5873 -4520 -5551 -4519
rect -5873 -4840 -5872 -4520
rect -5552 -4840 -5551 -4520
rect -5873 -4841 -5551 -4840
rect -6296 -5188 -6192 -4892
rect -6885 -5240 -6563 -5239
rect -6885 -5560 -6884 -5240
rect -6564 -5560 -6563 -5240
rect -6885 -5561 -6563 -5560
rect -7308 -5760 -7204 -5612
rect -6776 -5760 -6672 -5561
rect -6296 -5612 -6276 -5188
rect -6212 -5612 -6192 -5188
rect -5764 -5239 -5660 -4841
rect -5284 -4892 -5264 -4468
rect -5200 -4892 -5180 -4468
rect -4752 -4519 -4648 -4121
rect -4272 -4172 -4252 -3748
rect -4188 -4172 -4168 -3748
rect -3740 -3799 -3636 -3401
rect -3260 -3452 -3240 -3028
rect -3176 -3452 -3156 -3028
rect -2728 -3079 -2624 -2681
rect -2248 -2732 -2228 -2308
rect -2164 -2732 -2144 -2308
rect -1716 -2359 -1612 -1961
rect -1236 -2012 -1216 -1588
rect -1152 -2012 -1132 -1588
rect -704 -1639 -600 -1241
rect -224 -1292 -204 -868
rect -140 -1292 -120 -868
rect 308 -919 412 -521
rect 788 -572 808 -148
rect 872 -572 892 -148
rect 1320 -199 1424 199
rect 1800 148 1820 572
rect 1884 148 1904 572
rect 2332 521 2436 919
rect 2812 868 2832 1292
rect 2896 868 2916 1292
rect 3344 1241 3448 1639
rect 3824 1588 3844 2012
rect 3908 1588 3928 2012
rect 4356 1961 4460 2359
rect 4836 2308 4856 2732
rect 4920 2308 4940 2732
rect 5368 2681 5472 3079
rect 5848 3028 5868 3452
rect 5932 3028 5952 3452
rect 6380 3401 6484 3799
rect 6860 3748 6880 4172
rect 6944 3748 6964 4172
rect 7392 4121 7496 4519
rect 7872 4468 7892 4892
rect 7956 4468 7976 4892
rect 8404 4841 8508 5239
rect 8884 5188 8904 5612
rect 8968 5188 8988 5612
rect 9416 5561 9520 5760
rect 9896 5612 10000 5760
rect 9307 5560 9629 5561
rect 9307 5240 9308 5560
rect 9628 5240 9629 5560
rect 9307 5239 9629 5240
rect 8884 4892 8988 5188
rect 8295 4840 8617 4841
rect 8295 4520 8296 4840
rect 8616 4520 8617 4840
rect 8295 4519 8617 4520
rect 7872 4172 7976 4468
rect 7283 4120 7605 4121
rect 7283 3800 7284 4120
rect 7604 3800 7605 4120
rect 7283 3799 7605 3800
rect 6860 3452 6964 3748
rect 6271 3400 6593 3401
rect 6271 3080 6272 3400
rect 6592 3080 6593 3400
rect 6271 3079 6593 3080
rect 5848 2732 5952 3028
rect 5259 2680 5581 2681
rect 5259 2360 5260 2680
rect 5580 2360 5581 2680
rect 5259 2359 5581 2360
rect 4836 2012 4940 2308
rect 4247 1960 4569 1961
rect 4247 1640 4248 1960
rect 4568 1640 4569 1960
rect 4247 1639 4569 1640
rect 3824 1292 3928 1588
rect 3235 1240 3557 1241
rect 3235 920 3236 1240
rect 3556 920 3557 1240
rect 3235 919 3557 920
rect 2812 572 2916 868
rect 2223 520 2545 521
rect 2223 200 2224 520
rect 2544 200 2545 520
rect 2223 199 2545 200
rect 1800 -148 1904 148
rect 1211 -200 1533 -199
rect 1211 -520 1212 -200
rect 1532 -520 1533 -200
rect 1211 -521 1533 -520
rect 788 -868 892 -572
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -224 -1588 -120 -1292
rect -813 -1640 -491 -1639
rect -813 -1960 -812 -1640
rect -492 -1960 -491 -1640
rect -813 -1961 -491 -1960
rect -1236 -2308 -1132 -2012
rect -1825 -2360 -1503 -2359
rect -1825 -2680 -1824 -2360
rect -1504 -2680 -1503 -2360
rect -1825 -2681 -1503 -2680
rect -2248 -3028 -2144 -2732
rect -2837 -3080 -2515 -3079
rect -2837 -3400 -2836 -3080
rect -2516 -3400 -2515 -3080
rect -2837 -3401 -2515 -3400
rect -3260 -3748 -3156 -3452
rect -3849 -3800 -3527 -3799
rect -3849 -4120 -3848 -3800
rect -3528 -4120 -3527 -3800
rect -3849 -4121 -3527 -4120
rect -4272 -4468 -4168 -4172
rect -4861 -4520 -4539 -4519
rect -4861 -4840 -4860 -4520
rect -4540 -4840 -4539 -4520
rect -4861 -4841 -4539 -4840
rect -5284 -5188 -5180 -4892
rect -5873 -5240 -5551 -5239
rect -5873 -5560 -5872 -5240
rect -5552 -5560 -5551 -5240
rect -5873 -5561 -5551 -5560
rect -6296 -5760 -6192 -5612
rect -5764 -5760 -5660 -5561
rect -5284 -5612 -5264 -5188
rect -5200 -5612 -5180 -5188
rect -4752 -5239 -4648 -4841
rect -4272 -4892 -4252 -4468
rect -4188 -4892 -4168 -4468
rect -3740 -4519 -3636 -4121
rect -3260 -4172 -3240 -3748
rect -3176 -4172 -3156 -3748
rect -2728 -3799 -2624 -3401
rect -2248 -3452 -2228 -3028
rect -2164 -3452 -2144 -3028
rect -1716 -3079 -1612 -2681
rect -1236 -2732 -1216 -2308
rect -1152 -2732 -1132 -2308
rect -704 -2359 -600 -1961
rect -224 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect 308 -1639 412 -1241
rect 788 -1292 808 -868
rect 872 -1292 892 -868
rect 1320 -919 1424 -521
rect 1800 -572 1820 -148
rect 1884 -572 1904 -148
rect 2332 -199 2436 199
rect 2812 148 2832 572
rect 2896 148 2916 572
rect 3344 521 3448 919
rect 3824 868 3844 1292
rect 3908 868 3928 1292
rect 4356 1241 4460 1639
rect 4836 1588 4856 2012
rect 4920 1588 4940 2012
rect 5368 1961 5472 2359
rect 5848 2308 5868 2732
rect 5932 2308 5952 2732
rect 6380 2681 6484 3079
rect 6860 3028 6880 3452
rect 6944 3028 6964 3452
rect 7392 3401 7496 3799
rect 7872 3748 7892 4172
rect 7956 3748 7976 4172
rect 8404 4121 8508 4519
rect 8884 4468 8904 4892
rect 8968 4468 8988 4892
rect 9416 4841 9520 5239
rect 9896 5188 9916 5612
rect 9980 5188 10000 5612
rect 10428 5561 10532 5760
rect 10908 5612 11012 5760
rect 10319 5560 10641 5561
rect 10319 5240 10320 5560
rect 10640 5240 10641 5560
rect 10319 5239 10641 5240
rect 9896 4892 10000 5188
rect 9307 4840 9629 4841
rect 9307 4520 9308 4840
rect 9628 4520 9629 4840
rect 9307 4519 9629 4520
rect 8884 4172 8988 4468
rect 8295 4120 8617 4121
rect 8295 3800 8296 4120
rect 8616 3800 8617 4120
rect 8295 3799 8617 3800
rect 7872 3452 7976 3748
rect 7283 3400 7605 3401
rect 7283 3080 7284 3400
rect 7604 3080 7605 3400
rect 7283 3079 7605 3080
rect 6860 2732 6964 3028
rect 6271 2680 6593 2681
rect 6271 2360 6272 2680
rect 6592 2360 6593 2680
rect 6271 2359 6593 2360
rect 5848 2012 5952 2308
rect 5259 1960 5581 1961
rect 5259 1640 5260 1960
rect 5580 1640 5581 1960
rect 5259 1639 5581 1640
rect 4836 1292 4940 1588
rect 4247 1240 4569 1241
rect 4247 920 4248 1240
rect 4568 920 4569 1240
rect 4247 919 4569 920
rect 3824 572 3928 868
rect 3235 520 3557 521
rect 3235 200 3236 520
rect 3556 200 3557 520
rect 3235 199 3557 200
rect 2812 -148 2916 148
rect 2223 -200 2545 -199
rect 2223 -520 2224 -200
rect 2544 -520 2545 -200
rect 2223 -521 2545 -520
rect 1800 -868 1904 -572
rect 1211 -920 1533 -919
rect 1211 -1240 1212 -920
rect 1532 -1240 1533 -920
rect 1211 -1241 1533 -1240
rect 788 -1588 892 -1292
rect 199 -1640 521 -1639
rect 199 -1960 200 -1640
rect 520 -1960 521 -1640
rect 199 -1961 521 -1960
rect -224 -2308 -120 -2012
rect -813 -2360 -491 -2359
rect -813 -2680 -812 -2360
rect -492 -2680 -491 -2360
rect -813 -2681 -491 -2680
rect -1236 -3028 -1132 -2732
rect -1825 -3080 -1503 -3079
rect -1825 -3400 -1824 -3080
rect -1504 -3400 -1503 -3080
rect -1825 -3401 -1503 -3400
rect -2248 -3748 -2144 -3452
rect -2837 -3800 -2515 -3799
rect -2837 -4120 -2836 -3800
rect -2516 -4120 -2515 -3800
rect -2837 -4121 -2515 -4120
rect -3260 -4468 -3156 -4172
rect -3849 -4520 -3527 -4519
rect -3849 -4840 -3848 -4520
rect -3528 -4840 -3527 -4520
rect -3849 -4841 -3527 -4840
rect -4272 -5188 -4168 -4892
rect -4861 -5240 -4539 -5239
rect -4861 -5560 -4860 -5240
rect -4540 -5560 -4539 -5240
rect -4861 -5561 -4539 -5560
rect -5284 -5760 -5180 -5612
rect -4752 -5760 -4648 -5561
rect -4272 -5612 -4252 -5188
rect -4188 -5612 -4168 -5188
rect -3740 -5239 -3636 -4841
rect -3260 -4892 -3240 -4468
rect -3176 -4892 -3156 -4468
rect -2728 -4519 -2624 -4121
rect -2248 -4172 -2228 -3748
rect -2164 -4172 -2144 -3748
rect -1716 -3799 -1612 -3401
rect -1236 -3452 -1216 -3028
rect -1152 -3452 -1132 -3028
rect -704 -3079 -600 -2681
rect -224 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect 308 -2359 412 -1961
rect 788 -2012 808 -1588
rect 872 -2012 892 -1588
rect 1320 -1639 1424 -1241
rect 1800 -1292 1820 -868
rect 1884 -1292 1904 -868
rect 2332 -919 2436 -521
rect 2812 -572 2832 -148
rect 2896 -572 2916 -148
rect 3344 -199 3448 199
rect 3824 148 3844 572
rect 3908 148 3928 572
rect 4356 521 4460 919
rect 4836 868 4856 1292
rect 4920 868 4940 1292
rect 5368 1241 5472 1639
rect 5848 1588 5868 2012
rect 5932 1588 5952 2012
rect 6380 1961 6484 2359
rect 6860 2308 6880 2732
rect 6944 2308 6964 2732
rect 7392 2681 7496 3079
rect 7872 3028 7892 3452
rect 7956 3028 7976 3452
rect 8404 3401 8508 3799
rect 8884 3748 8904 4172
rect 8968 3748 8988 4172
rect 9416 4121 9520 4519
rect 9896 4468 9916 4892
rect 9980 4468 10000 4892
rect 10428 4841 10532 5239
rect 10908 5188 10928 5612
rect 10992 5188 11012 5612
rect 11440 5561 11544 5760
rect 11920 5612 12024 5760
rect 11331 5560 11653 5561
rect 11331 5240 11332 5560
rect 11652 5240 11653 5560
rect 11331 5239 11653 5240
rect 10908 4892 11012 5188
rect 10319 4840 10641 4841
rect 10319 4520 10320 4840
rect 10640 4520 10641 4840
rect 10319 4519 10641 4520
rect 9896 4172 10000 4468
rect 9307 4120 9629 4121
rect 9307 3800 9308 4120
rect 9628 3800 9629 4120
rect 9307 3799 9629 3800
rect 8884 3452 8988 3748
rect 8295 3400 8617 3401
rect 8295 3080 8296 3400
rect 8616 3080 8617 3400
rect 8295 3079 8617 3080
rect 7872 2732 7976 3028
rect 7283 2680 7605 2681
rect 7283 2360 7284 2680
rect 7604 2360 7605 2680
rect 7283 2359 7605 2360
rect 6860 2012 6964 2308
rect 6271 1960 6593 1961
rect 6271 1640 6272 1960
rect 6592 1640 6593 1960
rect 6271 1639 6593 1640
rect 5848 1292 5952 1588
rect 5259 1240 5581 1241
rect 5259 920 5260 1240
rect 5580 920 5581 1240
rect 5259 919 5581 920
rect 4836 572 4940 868
rect 4247 520 4569 521
rect 4247 200 4248 520
rect 4568 200 4569 520
rect 4247 199 4569 200
rect 3824 -148 3928 148
rect 3235 -200 3557 -199
rect 3235 -520 3236 -200
rect 3556 -520 3557 -200
rect 3235 -521 3557 -520
rect 2812 -868 2916 -572
rect 2223 -920 2545 -919
rect 2223 -1240 2224 -920
rect 2544 -1240 2545 -920
rect 2223 -1241 2545 -1240
rect 1800 -1588 1904 -1292
rect 1211 -1640 1533 -1639
rect 1211 -1960 1212 -1640
rect 1532 -1960 1533 -1640
rect 1211 -1961 1533 -1960
rect 788 -2308 892 -2012
rect 199 -2360 521 -2359
rect 199 -2680 200 -2360
rect 520 -2680 521 -2360
rect 199 -2681 521 -2680
rect -224 -3028 -120 -2732
rect -813 -3080 -491 -3079
rect -813 -3400 -812 -3080
rect -492 -3400 -491 -3080
rect -813 -3401 -491 -3400
rect -1236 -3748 -1132 -3452
rect -1825 -3800 -1503 -3799
rect -1825 -4120 -1824 -3800
rect -1504 -4120 -1503 -3800
rect -1825 -4121 -1503 -4120
rect -2248 -4468 -2144 -4172
rect -2837 -4520 -2515 -4519
rect -2837 -4840 -2836 -4520
rect -2516 -4840 -2515 -4520
rect -2837 -4841 -2515 -4840
rect -3260 -5188 -3156 -4892
rect -3849 -5240 -3527 -5239
rect -3849 -5560 -3848 -5240
rect -3528 -5560 -3527 -5240
rect -3849 -5561 -3527 -5560
rect -4272 -5760 -4168 -5612
rect -3740 -5760 -3636 -5561
rect -3260 -5612 -3240 -5188
rect -3176 -5612 -3156 -5188
rect -2728 -5239 -2624 -4841
rect -2248 -4892 -2228 -4468
rect -2164 -4892 -2144 -4468
rect -1716 -4519 -1612 -4121
rect -1236 -4172 -1216 -3748
rect -1152 -4172 -1132 -3748
rect -704 -3799 -600 -3401
rect -224 -3452 -204 -3028
rect -140 -3452 -120 -3028
rect 308 -3079 412 -2681
rect 788 -2732 808 -2308
rect 872 -2732 892 -2308
rect 1320 -2359 1424 -1961
rect 1800 -2012 1820 -1588
rect 1884 -2012 1904 -1588
rect 2332 -1639 2436 -1241
rect 2812 -1292 2832 -868
rect 2896 -1292 2916 -868
rect 3344 -919 3448 -521
rect 3824 -572 3844 -148
rect 3908 -572 3928 -148
rect 4356 -199 4460 199
rect 4836 148 4856 572
rect 4920 148 4940 572
rect 5368 521 5472 919
rect 5848 868 5868 1292
rect 5932 868 5952 1292
rect 6380 1241 6484 1639
rect 6860 1588 6880 2012
rect 6944 1588 6964 2012
rect 7392 1961 7496 2359
rect 7872 2308 7892 2732
rect 7956 2308 7976 2732
rect 8404 2681 8508 3079
rect 8884 3028 8904 3452
rect 8968 3028 8988 3452
rect 9416 3401 9520 3799
rect 9896 3748 9916 4172
rect 9980 3748 10000 4172
rect 10428 4121 10532 4519
rect 10908 4468 10928 4892
rect 10992 4468 11012 4892
rect 11440 4841 11544 5239
rect 11920 5188 11940 5612
rect 12004 5188 12024 5612
rect 12452 5561 12556 5760
rect 12932 5612 13036 5760
rect 12343 5560 12665 5561
rect 12343 5240 12344 5560
rect 12664 5240 12665 5560
rect 12343 5239 12665 5240
rect 11920 4892 12024 5188
rect 11331 4840 11653 4841
rect 11331 4520 11332 4840
rect 11652 4520 11653 4840
rect 11331 4519 11653 4520
rect 10908 4172 11012 4468
rect 10319 4120 10641 4121
rect 10319 3800 10320 4120
rect 10640 3800 10641 4120
rect 10319 3799 10641 3800
rect 9896 3452 10000 3748
rect 9307 3400 9629 3401
rect 9307 3080 9308 3400
rect 9628 3080 9629 3400
rect 9307 3079 9629 3080
rect 8884 2732 8988 3028
rect 8295 2680 8617 2681
rect 8295 2360 8296 2680
rect 8616 2360 8617 2680
rect 8295 2359 8617 2360
rect 7872 2012 7976 2308
rect 7283 1960 7605 1961
rect 7283 1640 7284 1960
rect 7604 1640 7605 1960
rect 7283 1639 7605 1640
rect 6860 1292 6964 1588
rect 6271 1240 6593 1241
rect 6271 920 6272 1240
rect 6592 920 6593 1240
rect 6271 919 6593 920
rect 5848 572 5952 868
rect 5259 520 5581 521
rect 5259 200 5260 520
rect 5580 200 5581 520
rect 5259 199 5581 200
rect 4836 -148 4940 148
rect 4247 -200 4569 -199
rect 4247 -520 4248 -200
rect 4568 -520 4569 -200
rect 4247 -521 4569 -520
rect 3824 -868 3928 -572
rect 3235 -920 3557 -919
rect 3235 -1240 3236 -920
rect 3556 -1240 3557 -920
rect 3235 -1241 3557 -1240
rect 2812 -1588 2916 -1292
rect 2223 -1640 2545 -1639
rect 2223 -1960 2224 -1640
rect 2544 -1960 2545 -1640
rect 2223 -1961 2545 -1960
rect 1800 -2308 1904 -2012
rect 1211 -2360 1533 -2359
rect 1211 -2680 1212 -2360
rect 1532 -2680 1533 -2360
rect 1211 -2681 1533 -2680
rect 788 -3028 892 -2732
rect 199 -3080 521 -3079
rect 199 -3400 200 -3080
rect 520 -3400 521 -3080
rect 199 -3401 521 -3400
rect -224 -3748 -120 -3452
rect -813 -3800 -491 -3799
rect -813 -4120 -812 -3800
rect -492 -4120 -491 -3800
rect -813 -4121 -491 -4120
rect -1236 -4468 -1132 -4172
rect -1825 -4520 -1503 -4519
rect -1825 -4840 -1824 -4520
rect -1504 -4840 -1503 -4520
rect -1825 -4841 -1503 -4840
rect -2248 -5188 -2144 -4892
rect -2837 -5240 -2515 -5239
rect -2837 -5560 -2836 -5240
rect -2516 -5560 -2515 -5240
rect -2837 -5561 -2515 -5560
rect -3260 -5760 -3156 -5612
rect -2728 -5760 -2624 -5561
rect -2248 -5612 -2228 -5188
rect -2164 -5612 -2144 -5188
rect -1716 -5239 -1612 -4841
rect -1236 -4892 -1216 -4468
rect -1152 -4892 -1132 -4468
rect -704 -4519 -600 -4121
rect -224 -4172 -204 -3748
rect -140 -4172 -120 -3748
rect 308 -3799 412 -3401
rect 788 -3452 808 -3028
rect 872 -3452 892 -3028
rect 1320 -3079 1424 -2681
rect 1800 -2732 1820 -2308
rect 1884 -2732 1904 -2308
rect 2332 -2359 2436 -1961
rect 2812 -2012 2832 -1588
rect 2896 -2012 2916 -1588
rect 3344 -1639 3448 -1241
rect 3824 -1292 3844 -868
rect 3908 -1292 3928 -868
rect 4356 -919 4460 -521
rect 4836 -572 4856 -148
rect 4920 -572 4940 -148
rect 5368 -199 5472 199
rect 5848 148 5868 572
rect 5932 148 5952 572
rect 6380 521 6484 919
rect 6860 868 6880 1292
rect 6944 868 6964 1292
rect 7392 1241 7496 1639
rect 7872 1588 7892 2012
rect 7956 1588 7976 2012
rect 8404 1961 8508 2359
rect 8884 2308 8904 2732
rect 8968 2308 8988 2732
rect 9416 2681 9520 3079
rect 9896 3028 9916 3452
rect 9980 3028 10000 3452
rect 10428 3401 10532 3799
rect 10908 3748 10928 4172
rect 10992 3748 11012 4172
rect 11440 4121 11544 4519
rect 11920 4468 11940 4892
rect 12004 4468 12024 4892
rect 12452 4841 12556 5239
rect 12932 5188 12952 5612
rect 13016 5188 13036 5612
rect 13464 5561 13568 5760
rect 13944 5612 14048 5760
rect 13355 5560 13677 5561
rect 13355 5240 13356 5560
rect 13676 5240 13677 5560
rect 13355 5239 13677 5240
rect 12932 4892 13036 5188
rect 12343 4840 12665 4841
rect 12343 4520 12344 4840
rect 12664 4520 12665 4840
rect 12343 4519 12665 4520
rect 11920 4172 12024 4468
rect 11331 4120 11653 4121
rect 11331 3800 11332 4120
rect 11652 3800 11653 4120
rect 11331 3799 11653 3800
rect 10908 3452 11012 3748
rect 10319 3400 10641 3401
rect 10319 3080 10320 3400
rect 10640 3080 10641 3400
rect 10319 3079 10641 3080
rect 9896 2732 10000 3028
rect 9307 2680 9629 2681
rect 9307 2360 9308 2680
rect 9628 2360 9629 2680
rect 9307 2359 9629 2360
rect 8884 2012 8988 2308
rect 8295 1960 8617 1961
rect 8295 1640 8296 1960
rect 8616 1640 8617 1960
rect 8295 1639 8617 1640
rect 7872 1292 7976 1588
rect 7283 1240 7605 1241
rect 7283 920 7284 1240
rect 7604 920 7605 1240
rect 7283 919 7605 920
rect 6860 572 6964 868
rect 6271 520 6593 521
rect 6271 200 6272 520
rect 6592 200 6593 520
rect 6271 199 6593 200
rect 5848 -148 5952 148
rect 5259 -200 5581 -199
rect 5259 -520 5260 -200
rect 5580 -520 5581 -200
rect 5259 -521 5581 -520
rect 4836 -868 4940 -572
rect 4247 -920 4569 -919
rect 4247 -1240 4248 -920
rect 4568 -1240 4569 -920
rect 4247 -1241 4569 -1240
rect 3824 -1588 3928 -1292
rect 3235 -1640 3557 -1639
rect 3235 -1960 3236 -1640
rect 3556 -1960 3557 -1640
rect 3235 -1961 3557 -1960
rect 2812 -2308 2916 -2012
rect 2223 -2360 2545 -2359
rect 2223 -2680 2224 -2360
rect 2544 -2680 2545 -2360
rect 2223 -2681 2545 -2680
rect 1800 -3028 1904 -2732
rect 1211 -3080 1533 -3079
rect 1211 -3400 1212 -3080
rect 1532 -3400 1533 -3080
rect 1211 -3401 1533 -3400
rect 788 -3748 892 -3452
rect 199 -3800 521 -3799
rect 199 -4120 200 -3800
rect 520 -4120 521 -3800
rect 199 -4121 521 -4120
rect -224 -4468 -120 -4172
rect -813 -4520 -491 -4519
rect -813 -4840 -812 -4520
rect -492 -4840 -491 -4520
rect -813 -4841 -491 -4840
rect -1236 -5188 -1132 -4892
rect -1825 -5240 -1503 -5239
rect -1825 -5560 -1824 -5240
rect -1504 -5560 -1503 -5240
rect -1825 -5561 -1503 -5560
rect -2248 -5760 -2144 -5612
rect -1716 -5760 -1612 -5561
rect -1236 -5612 -1216 -5188
rect -1152 -5612 -1132 -5188
rect -704 -5239 -600 -4841
rect -224 -4892 -204 -4468
rect -140 -4892 -120 -4468
rect 308 -4519 412 -4121
rect 788 -4172 808 -3748
rect 872 -4172 892 -3748
rect 1320 -3799 1424 -3401
rect 1800 -3452 1820 -3028
rect 1884 -3452 1904 -3028
rect 2332 -3079 2436 -2681
rect 2812 -2732 2832 -2308
rect 2896 -2732 2916 -2308
rect 3344 -2359 3448 -1961
rect 3824 -2012 3844 -1588
rect 3908 -2012 3928 -1588
rect 4356 -1639 4460 -1241
rect 4836 -1292 4856 -868
rect 4920 -1292 4940 -868
rect 5368 -919 5472 -521
rect 5848 -572 5868 -148
rect 5932 -572 5952 -148
rect 6380 -199 6484 199
rect 6860 148 6880 572
rect 6944 148 6964 572
rect 7392 521 7496 919
rect 7872 868 7892 1292
rect 7956 868 7976 1292
rect 8404 1241 8508 1639
rect 8884 1588 8904 2012
rect 8968 1588 8988 2012
rect 9416 1961 9520 2359
rect 9896 2308 9916 2732
rect 9980 2308 10000 2732
rect 10428 2681 10532 3079
rect 10908 3028 10928 3452
rect 10992 3028 11012 3452
rect 11440 3401 11544 3799
rect 11920 3748 11940 4172
rect 12004 3748 12024 4172
rect 12452 4121 12556 4519
rect 12932 4468 12952 4892
rect 13016 4468 13036 4892
rect 13464 4841 13568 5239
rect 13944 5188 13964 5612
rect 14028 5188 14048 5612
rect 14476 5561 14580 5760
rect 14956 5612 15060 5760
rect 14367 5560 14689 5561
rect 14367 5240 14368 5560
rect 14688 5240 14689 5560
rect 14367 5239 14689 5240
rect 13944 4892 14048 5188
rect 13355 4840 13677 4841
rect 13355 4520 13356 4840
rect 13676 4520 13677 4840
rect 13355 4519 13677 4520
rect 12932 4172 13036 4468
rect 12343 4120 12665 4121
rect 12343 3800 12344 4120
rect 12664 3800 12665 4120
rect 12343 3799 12665 3800
rect 11920 3452 12024 3748
rect 11331 3400 11653 3401
rect 11331 3080 11332 3400
rect 11652 3080 11653 3400
rect 11331 3079 11653 3080
rect 10908 2732 11012 3028
rect 10319 2680 10641 2681
rect 10319 2360 10320 2680
rect 10640 2360 10641 2680
rect 10319 2359 10641 2360
rect 9896 2012 10000 2308
rect 9307 1960 9629 1961
rect 9307 1640 9308 1960
rect 9628 1640 9629 1960
rect 9307 1639 9629 1640
rect 8884 1292 8988 1588
rect 8295 1240 8617 1241
rect 8295 920 8296 1240
rect 8616 920 8617 1240
rect 8295 919 8617 920
rect 7872 572 7976 868
rect 7283 520 7605 521
rect 7283 200 7284 520
rect 7604 200 7605 520
rect 7283 199 7605 200
rect 6860 -148 6964 148
rect 6271 -200 6593 -199
rect 6271 -520 6272 -200
rect 6592 -520 6593 -200
rect 6271 -521 6593 -520
rect 5848 -868 5952 -572
rect 5259 -920 5581 -919
rect 5259 -1240 5260 -920
rect 5580 -1240 5581 -920
rect 5259 -1241 5581 -1240
rect 4836 -1588 4940 -1292
rect 4247 -1640 4569 -1639
rect 4247 -1960 4248 -1640
rect 4568 -1960 4569 -1640
rect 4247 -1961 4569 -1960
rect 3824 -2308 3928 -2012
rect 3235 -2360 3557 -2359
rect 3235 -2680 3236 -2360
rect 3556 -2680 3557 -2360
rect 3235 -2681 3557 -2680
rect 2812 -3028 2916 -2732
rect 2223 -3080 2545 -3079
rect 2223 -3400 2224 -3080
rect 2544 -3400 2545 -3080
rect 2223 -3401 2545 -3400
rect 1800 -3748 1904 -3452
rect 1211 -3800 1533 -3799
rect 1211 -4120 1212 -3800
rect 1532 -4120 1533 -3800
rect 1211 -4121 1533 -4120
rect 788 -4468 892 -4172
rect 199 -4520 521 -4519
rect 199 -4840 200 -4520
rect 520 -4840 521 -4520
rect 199 -4841 521 -4840
rect -224 -5188 -120 -4892
rect -813 -5240 -491 -5239
rect -813 -5560 -812 -5240
rect -492 -5560 -491 -5240
rect -813 -5561 -491 -5560
rect -1236 -5760 -1132 -5612
rect -704 -5760 -600 -5561
rect -224 -5612 -204 -5188
rect -140 -5612 -120 -5188
rect 308 -5239 412 -4841
rect 788 -4892 808 -4468
rect 872 -4892 892 -4468
rect 1320 -4519 1424 -4121
rect 1800 -4172 1820 -3748
rect 1884 -4172 1904 -3748
rect 2332 -3799 2436 -3401
rect 2812 -3452 2832 -3028
rect 2896 -3452 2916 -3028
rect 3344 -3079 3448 -2681
rect 3824 -2732 3844 -2308
rect 3908 -2732 3928 -2308
rect 4356 -2359 4460 -1961
rect 4836 -2012 4856 -1588
rect 4920 -2012 4940 -1588
rect 5368 -1639 5472 -1241
rect 5848 -1292 5868 -868
rect 5932 -1292 5952 -868
rect 6380 -919 6484 -521
rect 6860 -572 6880 -148
rect 6944 -572 6964 -148
rect 7392 -199 7496 199
rect 7872 148 7892 572
rect 7956 148 7976 572
rect 8404 521 8508 919
rect 8884 868 8904 1292
rect 8968 868 8988 1292
rect 9416 1241 9520 1639
rect 9896 1588 9916 2012
rect 9980 1588 10000 2012
rect 10428 1961 10532 2359
rect 10908 2308 10928 2732
rect 10992 2308 11012 2732
rect 11440 2681 11544 3079
rect 11920 3028 11940 3452
rect 12004 3028 12024 3452
rect 12452 3401 12556 3799
rect 12932 3748 12952 4172
rect 13016 3748 13036 4172
rect 13464 4121 13568 4519
rect 13944 4468 13964 4892
rect 14028 4468 14048 4892
rect 14476 4841 14580 5239
rect 14956 5188 14976 5612
rect 15040 5188 15060 5612
rect 15488 5561 15592 5760
rect 15968 5612 16072 5760
rect 15379 5560 15701 5561
rect 15379 5240 15380 5560
rect 15700 5240 15701 5560
rect 15379 5239 15701 5240
rect 14956 4892 15060 5188
rect 14367 4840 14689 4841
rect 14367 4520 14368 4840
rect 14688 4520 14689 4840
rect 14367 4519 14689 4520
rect 13944 4172 14048 4468
rect 13355 4120 13677 4121
rect 13355 3800 13356 4120
rect 13676 3800 13677 4120
rect 13355 3799 13677 3800
rect 12932 3452 13036 3748
rect 12343 3400 12665 3401
rect 12343 3080 12344 3400
rect 12664 3080 12665 3400
rect 12343 3079 12665 3080
rect 11920 2732 12024 3028
rect 11331 2680 11653 2681
rect 11331 2360 11332 2680
rect 11652 2360 11653 2680
rect 11331 2359 11653 2360
rect 10908 2012 11012 2308
rect 10319 1960 10641 1961
rect 10319 1640 10320 1960
rect 10640 1640 10641 1960
rect 10319 1639 10641 1640
rect 9896 1292 10000 1588
rect 9307 1240 9629 1241
rect 9307 920 9308 1240
rect 9628 920 9629 1240
rect 9307 919 9629 920
rect 8884 572 8988 868
rect 8295 520 8617 521
rect 8295 200 8296 520
rect 8616 200 8617 520
rect 8295 199 8617 200
rect 7872 -148 7976 148
rect 7283 -200 7605 -199
rect 7283 -520 7284 -200
rect 7604 -520 7605 -200
rect 7283 -521 7605 -520
rect 6860 -868 6964 -572
rect 6271 -920 6593 -919
rect 6271 -1240 6272 -920
rect 6592 -1240 6593 -920
rect 6271 -1241 6593 -1240
rect 5848 -1588 5952 -1292
rect 5259 -1640 5581 -1639
rect 5259 -1960 5260 -1640
rect 5580 -1960 5581 -1640
rect 5259 -1961 5581 -1960
rect 4836 -2308 4940 -2012
rect 4247 -2360 4569 -2359
rect 4247 -2680 4248 -2360
rect 4568 -2680 4569 -2360
rect 4247 -2681 4569 -2680
rect 3824 -3028 3928 -2732
rect 3235 -3080 3557 -3079
rect 3235 -3400 3236 -3080
rect 3556 -3400 3557 -3080
rect 3235 -3401 3557 -3400
rect 2812 -3748 2916 -3452
rect 2223 -3800 2545 -3799
rect 2223 -4120 2224 -3800
rect 2544 -4120 2545 -3800
rect 2223 -4121 2545 -4120
rect 1800 -4468 1904 -4172
rect 1211 -4520 1533 -4519
rect 1211 -4840 1212 -4520
rect 1532 -4840 1533 -4520
rect 1211 -4841 1533 -4840
rect 788 -5188 892 -4892
rect 199 -5240 521 -5239
rect 199 -5560 200 -5240
rect 520 -5560 521 -5240
rect 199 -5561 521 -5560
rect -224 -5760 -120 -5612
rect 308 -5760 412 -5561
rect 788 -5612 808 -5188
rect 872 -5612 892 -5188
rect 1320 -5239 1424 -4841
rect 1800 -4892 1820 -4468
rect 1884 -4892 1904 -4468
rect 2332 -4519 2436 -4121
rect 2812 -4172 2832 -3748
rect 2896 -4172 2916 -3748
rect 3344 -3799 3448 -3401
rect 3824 -3452 3844 -3028
rect 3908 -3452 3928 -3028
rect 4356 -3079 4460 -2681
rect 4836 -2732 4856 -2308
rect 4920 -2732 4940 -2308
rect 5368 -2359 5472 -1961
rect 5848 -2012 5868 -1588
rect 5932 -2012 5952 -1588
rect 6380 -1639 6484 -1241
rect 6860 -1292 6880 -868
rect 6944 -1292 6964 -868
rect 7392 -919 7496 -521
rect 7872 -572 7892 -148
rect 7956 -572 7976 -148
rect 8404 -199 8508 199
rect 8884 148 8904 572
rect 8968 148 8988 572
rect 9416 521 9520 919
rect 9896 868 9916 1292
rect 9980 868 10000 1292
rect 10428 1241 10532 1639
rect 10908 1588 10928 2012
rect 10992 1588 11012 2012
rect 11440 1961 11544 2359
rect 11920 2308 11940 2732
rect 12004 2308 12024 2732
rect 12452 2681 12556 3079
rect 12932 3028 12952 3452
rect 13016 3028 13036 3452
rect 13464 3401 13568 3799
rect 13944 3748 13964 4172
rect 14028 3748 14048 4172
rect 14476 4121 14580 4519
rect 14956 4468 14976 4892
rect 15040 4468 15060 4892
rect 15488 4841 15592 5239
rect 15968 5188 15988 5612
rect 16052 5188 16072 5612
rect 16500 5561 16604 5760
rect 16980 5612 17084 5760
rect 16391 5560 16713 5561
rect 16391 5240 16392 5560
rect 16712 5240 16713 5560
rect 16391 5239 16713 5240
rect 15968 4892 16072 5188
rect 15379 4840 15701 4841
rect 15379 4520 15380 4840
rect 15700 4520 15701 4840
rect 15379 4519 15701 4520
rect 14956 4172 15060 4468
rect 14367 4120 14689 4121
rect 14367 3800 14368 4120
rect 14688 3800 14689 4120
rect 14367 3799 14689 3800
rect 13944 3452 14048 3748
rect 13355 3400 13677 3401
rect 13355 3080 13356 3400
rect 13676 3080 13677 3400
rect 13355 3079 13677 3080
rect 12932 2732 13036 3028
rect 12343 2680 12665 2681
rect 12343 2360 12344 2680
rect 12664 2360 12665 2680
rect 12343 2359 12665 2360
rect 11920 2012 12024 2308
rect 11331 1960 11653 1961
rect 11331 1640 11332 1960
rect 11652 1640 11653 1960
rect 11331 1639 11653 1640
rect 10908 1292 11012 1588
rect 10319 1240 10641 1241
rect 10319 920 10320 1240
rect 10640 920 10641 1240
rect 10319 919 10641 920
rect 9896 572 10000 868
rect 9307 520 9629 521
rect 9307 200 9308 520
rect 9628 200 9629 520
rect 9307 199 9629 200
rect 8884 -148 8988 148
rect 8295 -200 8617 -199
rect 8295 -520 8296 -200
rect 8616 -520 8617 -200
rect 8295 -521 8617 -520
rect 7872 -868 7976 -572
rect 7283 -920 7605 -919
rect 7283 -1240 7284 -920
rect 7604 -1240 7605 -920
rect 7283 -1241 7605 -1240
rect 6860 -1588 6964 -1292
rect 6271 -1640 6593 -1639
rect 6271 -1960 6272 -1640
rect 6592 -1960 6593 -1640
rect 6271 -1961 6593 -1960
rect 5848 -2308 5952 -2012
rect 5259 -2360 5581 -2359
rect 5259 -2680 5260 -2360
rect 5580 -2680 5581 -2360
rect 5259 -2681 5581 -2680
rect 4836 -3028 4940 -2732
rect 4247 -3080 4569 -3079
rect 4247 -3400 4248 -3080
rect 4568 -3400 4569 -3080
rect 4247 -3401 4569 -3400
rect 3824 -3748 3928 -3452
rect 3235 -3800 3557 -3799
rect 3235 -4120 3236 -3800
rect 3556 -4120 3557 -3800
rect 3235 -4121 3557 -4120
rect 2812 -4468 2916 -4172
rect 2223 -4520 2545 -4519
rect 2223 -4840 2224 -4520
rect 2544 -4840 2545 -4520
rect 2223 -4841 2545 -4840
rect 1800 -5188 1904 -4892
rect 1211 -5240 1533 -5239
rect 1211 -5560 1212 -5240
rect 1532 -5560 1533 -5240
rect 1211 -5561 1533 -5560
rect 788 -5760 892 -5612
rect 1320 -5760 1424 -5561
rect 1800 -5612 1820 -5188
rect 1884 -5612 1904 -5188
rect 2332 -5239 2436 -4841
rect 2812 -4892 2832 -4468
rect 2896 -4892 2916 -4468
rect 3344 -4519 3448 -4121
rect 3824 -4172 3844 -3748
rect 3908 -4172 3928 -3748
rect 4356 -3799 4460 -3401
rect 4836 -3452 4856 -3028
rect 4920 -3452 4940 -3028
rect 5368 -3079 5472 -2681
rect 5848 -2732 5868 -2308
rect 5932 -2732 5952 -2308
rect 6380 -2359 6484 -1961
rect 6860 -2012 6880 -1588
rect 6944 -2012 6964 -1588
rect 7392 -1639 7496 -1241
rect 7872 -1292 7892 -868
rect 7956 -1292 7976 -868
rect 8404 -919 8508 -521
rect 8884 -572 8904 -148
rect 8968 -572 8988 -148
rect 9416 -199 9520 199
rect 9896 148 9916 572
rect 9980 148 10000 572
rect 10428 521 10532 919
rect 10908 868 10928 1292
rect 10992 868 11012 1292
rect 11440 1241 11544 1639
rect 11920 1588 11940 2012
rect 12004 1588 12024 2012
rect 12452 1961 12556 2359
rect 12932 2308 12952 2732
rect 13016 2308 13036 2732
rect 13464 2681 13568 3079
rect 13944 3028 13964 3452
rect 14028 3028 14048 3452
rect 14476 3401 14580 3799
rect 14956 3748 14976 4172
rect 15040 3748 15060 4172
rect 15488 4121 15592 4519
rect 15968 4468 15988 4892
rect 16052 4468 16072 4892
rect 16500 4841 16604 5239
rect 16980 5188 17000 5612
rect 17064 5188 17084 5612
rect 17512 5561 17616 5760
rect 17992 5612 18096 5760
rect 17403 5560 17725 5561
rect 17403 5240 17404 5560
rect 17724 5240 17725 5560
rect 17403 5239 17725 5240
rect 16980 4892 17084 5188
rect 16391 4840 16713 4841
rect 16391 4520 16392 4840
rect 16712 4520 16713 4840
rect 16391 4519 16713 4520
rect 15968 4172 16072 4468
rect 15379 4120 15701 4121
rect 15379 3800 15380 4120
rect 15700 3800 15701 4120
rect 15379 3799 15701 3800
rect 14956 3452 15060 3748
rect 14367 3400 14689 3401
rect 14367 3080 14368 3400
rect 14688 3080 14689 3400
rect 14367 3079 14689 3080
rect 13944 2732 14048 3028
rect 13355 2680 13677 2681
rect 13355 2360 13356 2680
rect 13676 2360 13677 2680
rect 13355 2359 13677 2360
rect 12932 2012 13036 2308
rect 12343 1960 12665 1961
rect 12343 1640 12344 1960
rect 12664 1640 12665 1960
rect 12343 1639 12665 1640
rect 11920 1292 12024 1588
rect 11331 1240 11653 1241
rect 11331 920 11332 1240
rect 11652 920 11653 1240
rect 11331 919 11653 920
rect 10908 572 11012 868
rect 10319 520 10641 521
rect 10319 200 10320 520
rect 10640 200 10641 520
rect 10319 199 10641 200
rect 9896 -148 10000 148
rect 9307 -200 9629 -199
rect 9307 -520 9308 -200
rect 9628 -520 9629 -200
rect 9307 -521 9629 -520
rect 8884 -868 8988 -572
rect 8295 -920 8617 -919
rect 8295 -1240 8296 -920
rect 8616 -1240 8617 -920
rect 8295 -1241 8617 -1240
rect 7872 -1588 7976 -1292
rect 7283 -1640 7605 -1639
rect 7283 -1960 7284 -1640
rect 7604 -1960 7605 -1640
rect 7283 -1961 7605 -1960
rect 6860 -2308 6964 -2012
rect 6271 -2360 6593 -2359
rect 6271 -2680 6272 -2360
rect 6592 -2680 6593 -2360
rect 6271 -2681 6593 -2680
rect 5848 -3028 5952 -2732
rect 5259 -3080 5581 -3079
rect 5259 -3400 5260 -3080
rect 5580 -3400 5581 -3080
rect 5259 -3401 5581 -3400
rect 4836 -3748 4940 -3452
rect 4247 -3800 4569 -3799
rect 4247 -4120 4248 -3800
rect 4568 -4120 4569 -3800
rect 4247 -4121 4569 -4120
rect 3824 -4468 3928 -4172
rect 3235 -4520 3557 -4519
rect 3235 -4840 3236 -4520
rect 3556 -4840 3557 -4520
rect 3235 -4841 3557 -4840
rect 2812 -5188 2916 -4892
rect 2223 -5240 2545 -5239
rect 2223 -5560 2224 -5240
rect 2544 -5560 2545 -5240
rect 2223 -5561 2545 -5560
rect 1800 -5760 1904 -5612
rect 2332 -5760 2436 -5561
rect 2812 -5612 2832 -5188
rect 2896 -5612 2916 -5188
rect 3344 -5239 3448 -4841
rect 3824 -4892 3844 -4468
rect 3908 -4892 3928 -4468
rect 4356 -4519 4460 -4121
rect 4836 -4172 4856 -3748
rect 4920 -4172 4940 -3748
rect 5368 -3799 5472 -3401
rect 5848 -3452 5868 -3028
rect 5932 -3452 5952 -3028
rect 6380 -3079 6484 -2681
rect 6860 -2732 6880 -2308
rect 6944 -2732 6964 -2308
rect 7392 -2359 7496 -1961
rect 7872 -2012 7892 -1588
rect 7956 -2012 7976 -1588
rect 8404 -1639 8508 -1241
rect 8884 -1292 8904 -868
rect 8968 -1292 8988 -868
rect 9416 -919 9520 -521
rect 9896 -572 9916 -148
rect 9980 -572 10000 -148
rect 10428 -199 10532 199
rect 10908 148 10928 572
rect 10992 148 11012 572
rect 11440 521 11544 919
rect 11920 868 11940 1292
rect 12004 868 12024 1292
rect 12452 1241 12556 1639
rect 12932 1588 12952 2012
rect 13016 1588 13036 2012
rect 13464 1961 13568 2359
rect 13944 2308 13964 2732
rect 14028 2308 14048 2732
rect 14476 2681 14580 3079
rect 14956 3028 14976 3452
rect 15040 3028 15060 3452
rect 15488 3401 15592 3799
rect 15968 3748 15988 4172
rect 16052 3748 16072 4172
rect 16500 4121 16604 4519
rect 16980 4468 17000 4892
rect 17064 4468 17084 4892
rect 17512 4841 17616 5239
rect 17992 5188 18012 5612
rect 18076 5188 18096 5612
rect 18524 5561 18628 5760
rect 19004 5612 19108 5760
rect 18415 5560 18737 5561
rect 18415 5240 18416 5560
rect 18736 5240 18737 5560
rect 18415 5239 18737 5240
rect 17992 4892 18096 5188
rect 17403 4840 17725 4841
rect 17403 4520 17404 4840
rect 17724 4520 17725 4840
rect 17403 4519 17725 4520
rect 16980 4172 17084 4468
rect 16391 4120 16713 4121
rect 16391 3800 16392 4120
rect 16712 3800 16713 4120
rect 16391 3799 16713 3800
rect 15968 3452 16072 3748
rect 15379 3400 15701 3401
rect 15379 3080 15380 3400
rect 15700 3080 15701 3400
rect 15379 3079 15701 3080
rect 14956 2732 15060 3028
rect 14367 2680 14689 2681
rect 14367 2360 14368 2680
rect 14688 2360 14689 2680
rect 14367 2359 14689 2360
rect 13944 2012 14048 2308
rect 13355 1960 13677 1961
rect 13355 1640 13356 1960
rect 13676 1640 13677 1960
rect 13355 1639 13677 1640
rect 12932 1292 13036 1588
rect 12343 1240 12665 1241
rect 12343 920 12344 1240
rect 12664 920 12665 1240
rect 12343 919 12665 920
rect 11920 572 12024 868
rect 11331 520 11653 521
rect 11331 200 11332 520
rect 11652 200 11653 520
rect 11331 199 11653 200
rect 10908 -148 11012 148
rect 10319 -200 10641 -199
rect 10319 -520 10320 -200
rect 10640 -520 10641 -200
rect 10319 -521 10641 -520
rect 9896 -868 10000 -572
rect 9307 -920 9629 -919
rect 9307 -1240 9308 -920
rect 9628 -1240 9629 -920
rect 9307 -1241 9629 -1240
rect 8884 -1588 8988 -1292
rect 8295 -1640 8617 -1639
rect 8295 -1960 8296 -1640
rect 8616 -1960 8617 -1640
rect 8295 -1961 8617 -1960
rect 7872 -2308 7976 -2012
rect 7283 -2360 7605 -2359
rect 7283 -2680 7284 -2360
rect 7604 -2680 7605 -2360
rect 7283 -2681 7605 -2680
rect 6860 -3028 6964 -2732
rect 6271 -3080 6593 -3079
rect 6271 -3400 6272 -3080
rect 6592 -3400 6593 -3080
rect 6271 -3401 6593 -3400
rect 5848 -3748 5952 -3452
rect 5259 -3800 5581 -3799
rect 5259 -4120 5260 -3800
rect 5580 -4120 5581 -3800
rect 5259 -4121 5581 -4120
rect 4836 -4468 4940 -4172
rect 4247 -4520 4569 -4519
rect 4247 -4840 4248 -4520
rect 4568 -4840 4569 -4520
rect 4247 -4841 4569 -4840
rect 3824 -5188 3928 -4892
rect 3235 -5240 3557 -5239
rect 3235 -5560 3236 -5240
rect 3556 -5560 3557 -5240
rect 3235 -5561 3557 -5560
rect 2812 -5760 2916 -5612
rect 3344 -5760 3448 -5561
rect 3824 -5612 3844 -5188
rect 3908 -5612 3928 -5188
rect 4356 -5239 4460 -4841
rect 4836 -4892 4856 -4468
rect 4920 -4892 4940 -4468
rect 5368 -4519 5472 -4121
rect 5848 -4172 5868 -3748
rect 5932 -4172 5952 -3748
rect 6380 -3799 6484 -3401
rect 6860 -3452 6880 -3028
rect 6944 -3452 6964 -3028
rect 7392 -3079 7496 -2681
rect 7872 -2732 7892 -2308
rect 7956 -2732 7976 -2308
rect 8404 -2359 8508 -1961
rect 8884 -2012 8904 -1588
rect 8968 -2012 8988 -1588
rect 9416 -1639 9520 -1241
rect 9896 -1292 9916 -868
rect 9980 -1292 10000 -868
rect 10428 -919 10532 -521
rect 10908 -572 10928 -148
rect 10992 -572 11012 -148
rect 11440 -199 11544 199
rect 11920 148 11940 572
rect 12004 148 12024 572
rect 12452 521 12556 919
rect 12932 868 12952 1292
rect 13016 868 13036 1292
rect 13464 1241 13568 1639
rect 13944 1588 13964 2012
rect 14028 1588 14048 2012
rect 14476 1961 14580 2359
rect 14956 2308 14976 2732
rect 15040 2308 15060 2732
rect 15488 2681 15592 3079
rect 15968 3028 15988 3452
rect 16052 3028 16072 3452
rect 16500 3401 16604 3799
rect 16980 3748 17000 4172
rect 17064 3748 17084 4172
rect 17512 4121 17616 4519
rect 17992 4468 18012 4892
rect 18076 4468 18096 4892
rect 18524 4841 18628 5239
rect 19004 5188 19024 5612
rect 19088 5188 19108 5612
rect 19536 5561 19640 5760
rect 20016 5612 20120 5760
rect 19427 5560 19749 5561
rect 19427 5240 19428 5560
rect 19748 5240 19749 5560
rect 19427 5239 19749 5240
rect 19004 4892 19108 5188
rect 18415 4840 18737 4841
rect 18415 4520 18416 4840
rect 18736 4520 18737 4840
rect 18415 4519 18737 4520
rect 17992 4172 18096 4468
rect 17403 4120 17725 4121
rect 17403 3800 17404 4120
rect 17724 3800 17725 4120
rect 17403 3799 17725 3800
rect 16980 3452 17084 3748
rect 16391 3400 16713 3401
rect 16391 3080 16392 3400
rect 16712 3080 16713 3400
rect 16391 3079 16713 3080
rect 15968 2732 16072 3028
rect 15379 2680 15701 2681
rect 15379 2360 15380 2680
rect 15700 2360 15701 2680
rect 15379 2359 15701 2360
rect 14956 2012 15060 2308
rect 14367 1960 14689 1961
rect 14367 1640 14368 1960
rect 14688 1640 14689 1960
rect 14367 1639 14689 1640
rect 13944 1292 14048 1588
rect 13355 1240 13677 1241
rect 13355 920 13356 1240
rect 13676 920 13677 1240
rect 13355 919 13677 920
rect 12932 572 13036 868
rect 12343 520 12665 521
rect 12343 200 12344 520
rect 12664 200 12665 520
rect 12343 199 12665 200
rect 11920 -148 12024 148
rect 11331 -200 11653 -199
rect 11331 -520 11332 -200
rect 11652 -520 11653 -200
rect 11331 -521 11653 -520
rect 10908 -868 11012 -572
rect 10319 -920 10641 -919
rect 10319 -1240 10320 -920
rect 10640 -1240 10641 -920
rect 10319 -1241 10641 -1240
rect 9896 -1588 10000 -1292
rect 9307 -1640 9629 -1639
rect 9307 -1960 9308 -1640
rect 9628 -1960 9629 -1640
rect 9307 -1961 9629 -1960
rect 8884 -2308 8988 -2012
rect 8295 -2360 8617 -2359
rect 8295 -2680 8296 -2360
rect 8616 -2680 8617 -2360
rect 8295 -2681 8617 -2680
rect 7872 -3028 7976 -2732
rect 7283 -3080 7605 -3079
rect 7283 -3400 7284 -3080
rect 7604 -3400 7605 -3080
rect 7283 -3401 7605 -3400
rect 6860 -3748 6964 -3452
rect 6271 -3800 6593 -3799
rect 6271 -4120 6272 -3800
rect 6592 -4120 6593 -3800
rect 6271 -4121 6593 -4120
rect 5848 -4468 5952 -4172
rect 5259 -4520 5581 -4519
rect 5259 -4840 5260 -4520
rect 5580 -4840 5581 -4520
rect 5259 -4841 5581 -4840
rect 4836 -5188 4940 -4892
rect 4247 -5240 4569 -5239
rect 4247 -5560 4248 -5240
rect 4568 -5560 4569 -5240
rect 4247 -5561 4569 -5560
rect 3824 -5760 3928 -5612
rect 4356 -5760 4460 -5561
rect 4836 -5612 4856 -5188
rect 4920 -5612 4940 -5188
rect 5368 -5239 5472 -4841
rect 5848 -4892 5868 -4468
rect 5932 -4892 5952 -4468
rect 6380 -4519 6484 -4121
rect 6860 -4172 6880 -3748
rect 6944 -4172 6964 -3748
rect 7392 -3799 7496 -3401
rect 7872 -3452 7892 -3028
rect 7956 -3452 7976 -3028
rect 8404 -3079 8508 -2681
rect 8884 -2732 8904 -2308
rect 8968 -2732 8988 -2308
rect 9416 -2359 9520 -1961
rect 9896 -2012 9916 -1588
rect 9980 -2012 10000 -1588
rect 10428 -1639 10532 -1241
rect 10908 -1292 10928 -868
rect 10992 -1292 11012 -868
rect 11440 -919 11544 -521
rect 11920 -572 11940 -148
rect 12004 -572 12024 -148
rect 12452 -199 12556 199
rect 12932 148 12952 572
rect 13016 148 13036 572
rect 13464 521 13568 919
rect 13944 868 13964 1292
rect 14028 868 14048 1292
rect 14476 1241 14580 1639
rect 14956 1588 14976 2012
rect 15040 1588 15060 2012
rect 15488 1961 15592 2359
rect 15968 2308 15988 2732
rect 16052 2308 16072 2732
rect 16500 2681 16604 3079
rect 16980 3028 17000 3452
rect 17064 3028 17084 3452
rect 17512 3401 17616 3799
rect 17992 3748 18012 4172
rect 18076 3748 18096 4172
rect 18524 4121 18628 4519
rect 19004 4468 19024 4892
rect 19088 4468 19108 4892
rect 19536 4841 19640 5239
rect 20016 5188 20036 5612
rect 20100 5188 20120 5612
rect 20548 5561 20652 5760
rect 21028 5612 21132 5760
rect 20439 5560 20761 5561
rect 20439 5240 20440 5560
rect 20760 5240 20761 5560
rect 20439 5239 20761 5240
rect 20016 4892 20120 5188
rect 19427 4840 19749 4841
rect 19427 4520 19428 4840
rect 19748 4520 19749 4840
rect 19427 4519 19749 4520
rect 19004 4172 19108 4468
rect 18415 4120 18737 4121
rect 18415 3800 18416 4120
rect 18736 3800 18737 4120
rect 18415 3799 18737 3800
rect 17992 3452 18096 3748
rect 17403 3400 17725 3401
rect 17403 3080 17404 3400
rect 17724 3080 17725 3400
rect 17403 3079 17725 3080
rect 16980 2732 17084 3028
rect 16391 2680 16713 2681
rect 16391 2360 16392 2680
rect 16712 2360 16713 2680
rect 16391 2359 16713 2360
rect 15968 2012 16072 2308
rect 15379 1960 15701 1961
rect 15379 1640 15380 1960
rect 15700 1640 15701 1960
rect 15379 1639 15701 1640
rect 14956 1292 15060 1588
rect 14367 1240 14689 1241
rect 14367 920 14368 1240
rect 14688 920 14689 1240
rect 14367 919 14689 920
rect 13944 572 14048 868
rect 13355 520 13677 521
rect 13355 200 13356 520
rect 13676 200 13677 520
rect 13355 199 13677 200
rect 12932 -148 13036 148
rect 12343 -200 12665 -199
rect 12343 -520 12344 -200
rect 12664 -520 12665 -200
rect 12343 -521 12665 -520
rect 11920 -868 12024 -572
rect 11331 -920 11653 -919
rect 11331 -1240 11332 -920
rect 11652 -1240 11653 -920
rect 11331 -1241 11653 -1240
rect 10908 -1588 11012 -1292
rect 10319 -1640 10641 -1639
rect 10319 -1960 10320 -1640
rect 10640 -1960 10641 -1640
rect 10319 -1961 10641 -1960
rect 9896 -2308 10000 -2012
rect 9307 -2360 9629 -2359
rect 9307 -2680 9308 -2360
rect 9628 -2680 9629 -2360
rect 9307 -2681 9629 -2680
rect 8884 -3028 8988 -2732
rect 8295 -3080 8617 -3079
rect 8295 -3400 8296 -3080
rect 8616 -3400 8617 -3080
rect 8295 -3401 8617 -3400
rect 7872 -3748 7976 -3452
rect 7283 -3800 7605 -3799
rect 7283 -4120 7284 -3800
rect 7604 -4120 7605 -3800
rect 7283 -4121 7605 -4120
rect 6860 -4468 6964 -4172
rect 6271 -4520 6593 -4519
rect 6271 -4840 6272 -4520
rect 6592 -4840 6593 -4520
rect 6271 -4841 6593 -4840
rect 5848 -5188 5952 -4892
rect 5259 -5240 5581 -5239
rect 5259 -5560 5260 -5240
rect 5580 -5560 5581 -5240
rect 5259 -5561 5581 -5560
rect 4836 -5760 4940 -5612
rect 5368 -5760 5472 -5561
rect 5848 -5612 5868 -5188
rect 5932 -5612 5952 -5188
rect 6380 -5239 6484 -4841
rect 6860 -4892 6880 -4468
rect 6944 -4892 6964 -4468
rect 7392 -4519 7496 -4121
rect 7872 -4172 7892 -3748
rect 7956 -4172 7976 -3748
rect 8404 -3799 8508 -3401
rect 8884 -3452 8904 -3028
rect 8968 -3452 8988 -3028
rect 9416 -3079 9520 -2681
rect 9896 -2732 9916 -2308
rect 9980 -2732 10000 -2308
rect 10428 -2359 10532 -1961
rect 10908 -2012 10928 -1588
rect 10992 -2012 11012 -1588
rect 11440 -1639 11544 -1241
rect 11920 -1292 11940 -868
rect 12004 -1292 12024 -868
rect 12452 -919 12556 -521
rect 12932 -572 12952 -148
rect 13016 -572 13036 -148
rect 13464 -199 13568 199
rect 13944 148 13964 572
rect 14028 148 14048 572
rect 14476 521 14580 919
rect 14956 868 14976 1292
rect 15040 868 15060 1292
rect 15488 1241 15592 1639
rect 15968 1588 15988 2012
rect 16052 1588 16072 2012
rect 16500 1961 16604 2359
rect 16980 2308 17000 2732
rect 17064 2308 17084 2732
rect 17512 2681 17616 3079
rect 17992 3028 18012 3452
rect 18076 3028 18096 3452
rect 18524 3401 18628 3799
rect 19004 3748 19024 4172
rect 19088 3748 19108 4172
rect 19536 4121 19640 4519
rect 20016 4468 20036 4892
rect 20100 4468 20120 4892
rect 20548 4841 20652 5239
rect 21028 5188 21048 5612
rect 21112 5188 21132 5612
rect 21560 5561 21664 5760
rect 22040 5612 22144 5760
rect 21451 5560 21773 5561
rect 21451 5240 21452 5560
rect 21772 5240 21773 5560
rect 21451 5239 21773 5240
rect 21028 4892 21132 5188
rect 20439 4840 20761 4841
rect 20439 4520 20440 4840
rect 20760 4520 20761 4840
rect 20439 4519 20761 4520
rect 20016 4172 20120 4468
rect 19427 4120 19749 4121
rect 19427 3800 19428 4120
rect 19748 3800 19749 4120
rect 19427 3799 19749 3800
rect 19004 3452 19108 3748
rect 18415 3400 18737 3401
rect 18415 3080 18416 3400
rect 18736 3080 18737 3400
rect 18415 3079 18737 3080
rect 17992 2732 18096 3028
rect 17403 2680 17725 2681
rect 17403 2360 17404 2680
rect 17724 2360 17725 2680
rect 17403 2359 17725 2360
rect 16980 2012 17084 2308
rect 16391 1960 16713 1961
rect 16391 1640 16392 1960
rect 16712 1640 16713 1960
rect 16391 1639 16713 1640
rect 15968 1292 16072 1588
rect 15379 1240 15701 1241
rect 15379 920 15380 1240
rect 15700 920 15701 1240
rect 15379 919 15701 920
rect 14956 572 15060 868
rect 14367 520 14689 521
rect 14367 200 14368 520
rect 14688 200 14689 520
rect 14367 199 14689 200
rect 13944 -148 14048 148
rect 13355 -200 13677 -199
rect 13355 -520 13356 -200
rect 13676 -520 13677 -200
rect 13355 -521 13677 -520
rect 12932 -868 13036 -572
rect 12343 -920 12665 -919
rect 12343 -1240 12344 -920
rect 12664 -1240 12665 -920
rect 12343 -1241 12665 -1240
rect 11920 -1588 12024 -1292
rect 11331 -1640 11653 -1639
rect 11331 -1960 11332 -1640
rect 11652 -1960 11653 -1640
rect 11331 -1961 11653 -1960
rect 10908 -2308 11012 -2012
rect 10319 -2360 10641 -2359
rect 10319 -2680 10320 -2360
rect 10640 -2680 10641 -2360
rect 10319 -2681 10641 -2680
rect 9896 -3028 10000 -2732
rect 9307 -3080 9629 -3079
rect 9307 -3400 9308 -3080
rect 9628 -3400 9629 -3080
rect 9307 -3401 9629 -3400
rect 8884 -3748 8988 -3452
rect 8295 -3800 8617 -3799
rect 8295 -4120 8296 -3800
rect 8616 -4120 8617 -3800
rect 8295 -4121 8617 -4120
rect 7872 -4468 7976 -4172
rect 7283 -4520 7605 -4519
rect 7283 -4840 7284 -4520
rect 7604 -4840 7605 -4520
rect 7283 -4841 7605 -4840
rect 6860 -5188 6964 -4892
rect 6271 -5240 6593 -5239
rect 6271 -5560 6272 -5240
rect 6592 -5560 6593 -5240
rect 6271 -5561 6593 -5560
rect 5848 -5760 5952 -5612
rect 6380 -5760 6484 -5561
rect 6860 -5612 6880 -5188
rect 6944 -5612 6964 -5188
rect 7392 -5239 7496 -4841
rect 7872 -4892 7892 -4468
rect 7956 -4892 7976 -4468
rect 8404 -4519 8508 -4121
rect 8884 -4172 8904 -3748
rect 8968 -4172 8988 -3748
rect 9416 -3799 9520 -3401
rect 9896 -3452 9916 -3028
rect 9980 -3452 10000 -3028
rect 10428 -3079 10532 -2681
rect 10908 -2732 10928 -2308
rect 10992 -2732 11012 -2308
rect 11440 -2359 11544 -1961
rect 11920 -2012 11940 -1588
rect 12004 -2012 12024 -1588
rect 12452 -1639 12556 -1241
rect 12932 -1292 12952 -868
rect 13016 -1292 13036 -868
rect 13464 -919 13568 -521
rect 13944 -572 13964 -148
rect 14028 -572 14048 -148
rect 14476 -199 14580 199
rect 14956 148 14976 572
rect 15040 148 15060 572
rect 15488 521 15592 919
rect 15968 868 15988 1292
rect 16052 868 16072 1292
rect 16500 1241 16604 1639
rect 16980 1588 17000 2012
rect 17064 1588 17084 2012
rect 17512 1961 17616 2359
rect 17992 2308 18012 2732
rect 18076 2308 18096 2732
rect 18524 2681 18628 3079
rect 19004 3028 19024 3452
rect 19088 3028 19108 3452
rect 19536 3401 19640 3799
rect 20016 3748 20036 4172
rect 20100 3748 20120 4172
rect 20548 4121 20652 4519
rect 21028 4468 21048 4892
rect 21112 4468 21132 4892
rect 21560 4841 21664 5239
rect 22040 5188 22060 5612
rect 22124 5188 22144 5612
rect 22572 5561 22676 5760
rect 23052 5612 23156 5760
rect 22463 5560 22785 5561
rect 22463 5240 22464 5560
rect 22784 5240 22785 5560
rect 22463 5239 22785 5240
rect 22040 4892 22144 5188
rect 21451 4840 21773 4841
rect 21451 4520 21452 4840
rect 21772 4520 21773 4840
rect 21451 4519 21773 4520
rect 21028 4172 21132 4468
rect 20439 4120 20761 4121
rect 20439 3800 20440 4120
rect 20760 3800 20761 4120
rect 20439 3799 20761 3800
rect 20016 3452 20120 3748
rect 19427 3400 19749 3401
rect 19427 3080 19428 3400
rect 19748 3080 19749 3400
rect 19427 3079 19749 3080
rect 19004 2732 19108 3028
rect 18415 2680 18737 2681
rect 18415 2360 18416 2680
rect 18736 2360 18737 2680
rect 18415 2359 18737 2360
rect 17992 2012 18096 2308
rect 17403 1960 17725 1961
rect 17403 1640 17404 1960
rect 17724 1640 17725 1960
rect 17403 1639 17725 1640
rect 16980 1292 17084 1588
rect 16391 1240 16713 1241
rect 16391 920 16392 1240
rect 16712 920 16713 1240
rect 16391 919 16713 920
rect 15968 572 16072 868
rect 15379 520 15701 521
rect 15379 200 15380 520
rect 15700 200 15701 520
rect 15379 199 15701 200
rect 14956 -148 15060 148
rect 14367 -200 14689 -199
rect 14367 -520 14368 -200
rect 14688 -520 14689 -200
rect 14367 -521 14689 -520
rect 13944 -868 14048 -572
rect 13355 -920 13677 -919
rect 13355 -1240 13356 -920
rect 13676 -1240 13677 -920
rect 13355 -1241 13677 -1240
rect 12932 -1588 13036 -1292
rect 12343 -1640 12665 -1639
rect 12343 -1960 12344 -1640
rect 12664 -1960 12665 -1640
rect 12343 -1961 12665 -1960
rect 11920 -2308 12024 -2012
rect 11331 -2360 11653 -2359
rect 11331 -2680 11332 -2360
rect 11652 -2680 11653 -2360
rect 11331 -2681 11653 -2680
rect 10908 -3028 11012 -2732
rect 10319 -3080 10641 -3079
rect 10319 -3400 10320 -3080
rect 10640 -3400 10641 -3080
rect 10319 -3401 10641 -3400
rect 9896 -3748 10000 -3452
rect 9307 -3800 9629 -3799
rect 9307 -4120 9308 -3800
rect 9628 -4120 9629 -3800
rect 9307 -4121 9629 -4120
rect 8884 -4468 8988 -4172
rect 8295 -4520 8617 -4519
rect 8295 -4840 8296 -4520
rect 8616 -4840 8617 -4520
rect 8295 -4841 8617 -4840
rect 7872 -5188 7976 -4892
rect 7283 -5240 7605 -5239
rect 7283 -5560 7284 -5240
rect 7604 -5560 7605 -5240
rect 7283 -5561 7605 -5560
rect 6860 -5760 6964 -5612
rect 7392 -5760 7496 -5561
rect 7872 -5612 7892 -5188
rect 7956 -5612 7976 -5188
rect 8404 -5239 8508 -4841
rect 8884 -4892 8904 -4468
rect 8968 -4892 8988 -4468
rect 9416 -4519 9520 -4121
rect 9896 -4172 9916 -3748
rect 9980 -4172 10000 -3748
rect 10428 -3799 10532 -3401
rect 10908 -3452 10928 -3028
rect 10992 -3452 11012 -3028
rect 11440 -3079 11544 -2681
rect 11920 -2732 11940 -2308
rect 12004 -2732 12024 -2308
rect 12452 -2359 12556 -1961
rect 12932 -2012 12952 -1588
rect 13016 -2012 13036 -1588
rect 13464 -1639 13568 -1241
rect 13944 -1292 13964 -868
rect 14028 -1292 14048 -868
rect 14476 -919 14580 -521
rect 14956 -572 14976 -148
rect 15040 -572 15060 -148
rect 15488 -199 15592 199
rect 15968 148 15988 572
rect 16052 148 16072 572
rect 16500 521 16604 919
rect 16980 868 17000 1292
rect 17064 868 17084 1292
rect 17512 1241 17616 1639
rect 17992 1588 18012 2012
rect 18076 1588 18096 2012
rect 18524 1961 18628 2359
rect 19004 2308 19024 2732
rect 19088 2308 19108 2732
rect 19536 2681 19640 3079
rect 20016 3028 20036 3452
rect 20100 3028 20120 3452
rect 20548 3401 20652 3799
rect 21028 3748 21048 4172
rect 21112 3748 21132 4172
rect 21560 4121 21664 4519
rect 22040 4468 22060 4892
rect 22124 4468 22144 4892
rect 22572 4841 22676 5239
rect 23052 5188 23072 5612
rect 23136 5188 23156 5612
rect 23584 5561 23688 5760
rect 24064 5612 24168 5760
rect 23475 5560 23797 5561
rect 23475 5240 23476 5560
rect 23796 5240 23797 5560
rect 23475 5239 23797 5240
rect 23052 4892 23156 5188
rect 22463 4840 22785 4841
rect 22463 4520 22464 4840
rect 22784 4520 22785 4840
rect 22463 4519 22785 4520
rect 22040 4172 22144 4468
rect 21451 4120 21773 4121
rect 21451 3800 21452 4120
rect 21772 3800 21773 4120
rect 21451 3799 21773 3800
rect 21028 3452 21132 3748
rect 20439 3400 20761 3401
rect 20439 3080 20440 3400
rect 20760 3080 20761 3400
rect 20439 3079 20761 3080
rect 20016 2732 20120 3028
rect 19427 2680 19749 2681
rect 19427 2360 19428 2680
rect 19748 2360 19749 2680
rect 19427 2359 19749 2360
rect 19004 2012 19108 2308
rect 18415 1960 18737 1961
rect 18415 1640 18416 1960
rect 18736 1640 18737 1960
rect 18415 1639 18737 1640
rect 17992 1292 18096 1588
rect 17403 1240 17725 1241
rect 17403 920 17404 1240
rect 17724 920 17725 1240
rect 17403 919 17725 920
rect 16980 572 17084 868
rect 16391 520 16713 521
rect 16391 200 16392 520
rect 16712 200 16713 520
rect 16391 199 16713 200
rect 15968 -148 16072 148
rect 15379 -200 15701 -199
rect 15379 -520 15380 -200
rect 15700 -520 15701 -200
rect 15379 -521 15701 -520
rect 14956 -868 15060 -572
rect 14367 -920 14689 -919
rect 14367 -1240 14368 -920
rect 14688 -1240 14689 -920
rect 14367 -1241 14689 -1240
rect 13944 -1588 14048 -1292
rect 13355 -1640 13677 -1639
rect 13355 -1960 13356 -1640
rect 13676 -1960 13677 -1640
rect 13355 -1961 13677 -1960
rect 12932 -2308 13036 -2012
rect 12343 -2360 12665 -2359
rect 12343 -2680 12344 -2360
rect 12664 -2680 12665 -2360
rect 12343 -2681 12665 -2680
rect 11920 -3028 12024 -2732
rect 11331 -3080 11653 -3079
rect 11331 -3400 11332 -3080
rect 11652 -3400 11653 -3080
rect 11331 -3401 11653 -3400
rect 10908 -3748 11012 -3452
rect 10319 -3800 10641 -3799
rect 10319 -4120 10320 -3800
rect 10640 -4120 10641 -3800
rect 10319 -4121 10641 -4120
rect 9896 -4468 10000 -4172
rect 9307 -4520 9629 -4519
rect 9307 -4840 9308 -4520
rect 9628 -4840 9629 -4520
rect 9307 -4841 9629 -4840
rect 8884 -5188 8988 -4892
rect 8295 -5240 8617 -5239
rect 8295 -5560 8296 -5240
rect 8616 -5560 8617 -5240
rect 8295 -5561 8617 -5560
rect 7872 -5760 7976 -5612
rect 8404 -5760 8508 -5561
rect 8884 -5612 8904 -5188
rect 8968 -5612 8988 -5188
rect 9416 -5239 9520 -4841
rect 9896 -4892 9916 -4468
rect 9980 -4892 10000 -4468
rect 10428 -4519 10532 -4121
rect 10908 -4172 10928 -3748
rect 10992 -4172 11012 -3748
rect 11440 -3799 11544 -3401
rect 11920 -3452 11940 -3028
rect 12004 -3452 12024 -3028
rect 12452 -3079 12556 -2681
rect 12932 -2732 12952 -2308
rect 13016 -2732 13036 -2308
rect 13464 -2359 13568 -1961
rect 13944 -2012 13964 -1588
rect 14028 -2012 14048 -1588
rect 14476 -1639 14580 -1241
rect 14956 -1292 14976 -868
rect 15040 -1292 15060 -868
rect 15488 -919 15592 -521
rect 15968 -572 15988 -148
rect 16052 -572 16072 -148
rect 16500 -199 16604 199
rect 16980 148 17000 572
rect 17064 148 17084 572
rect 17512 521 17616 919
rect 17992 868 18012 1292
rect 18076 868 18096 1292
rect 18524 1241 18628 1639
rect 19004 1588 19024 2012
rect 19088 1588 19108 2012
rect 19536 1961 19640 2359
rect 20016 2308 20036 2732
rect 20100 2308 20120 2732
rect 20548 2681 20652 3079
rect 21028 3028 21048 3452
rect 21112 3028 21132 3452
rect 21560 3401 21664 3799
rect 22040 3748 22060 4172
rect 22124 3748 22144 4172
rect 22572 4121 22676 4519
rect 23052 4468 23072 4892
rect 23136 4468 23156 4892
rect 23584 4841 23688 5239
rect 24064 5188 24084 5612
rect 24148 5188 24168 5612
rect 24596 5561 24700 5760
rect 25076 5612 25180 5760
rect 24487 5560 24809 5561
rect 24487 5240 24488 5560
rect 24808 5240 24809 5560
rect 24487 5239 24809 5240
rect 24064 4892 24168 5188
rect 23475 4840 23797 4841
rect 23475 4520 23476 4840
rect 23796 4520 23797 4840
rect 23475 4519 23797 4520
rect 23052 4172 23156 4468
rect 22463 4120 22785 4121
rect 22463 3800 22464 4120
rect 22784 3800 22785 4120
rect 22463 3799 22785 3800
rect 22040 3452 22144 3748
rect 21451 3400 21773 3401
rect 21451 3080 21452 3400
rect 21772 3080 21773 3400
rect 21451 3079 21773 3080
rect 21028 2732 21132 3028
rect 20439 2680 20761 2681
rect 20439 2360 20440 2680
rect 20760 2360 20761 2680
rect 20439 2359 20761 2360
rect 20016 2012 20120 2308
rect 19427 1960 19749 1961
rect 19427 1640 19428 1960
rect 19748 1640 19749 1960
rect 19427 1639 19749 1640
rect 19004 1292 19108 1588
rect 18415 1240 18737 1241
rect 18415 920 18416 1240
rect 18736 920 18737 1240
rect 18415 919 18737 920
rect 17992 572 18096 868
rect 17403 520 17725 521
rect 17403 200 17404 520
rect 17724 200 17725 520
rect 17403 199 17725 200
rect 16980 -148 17084 148
rect 16391 -200 16713 -199
rect 16391 -520 16392 -200
rect 16712 -520 16713 -200
rect 16391 -521 16713 -520
rect 15968 -868 16072 -572
rect 15379 -920 15701 -919
rect 15379 -1240 15380 -920
rect 15700 -1240 15701 -920
rect 15379 -1241 15701 -1240
rect 14956 -1588 15060 -1292
rect 14367 -1640 14689 -1639
rect 14367 -1960 14368 -1640
rect 14688 -1960 14689 -1640
rect 14367 -1961 14689 -1960
rect 13944 -2308 14048 -2012
rect 13355 -2360 13677 -2359
rect 13355 -2680 13356 -2360
rect 13676 -2680 13677 -2360
rect 13355 -2681 13677 -2680
rect 12932 -3028 13036 -2732
rect 12343 -3080 12665 -3079
rect 12343 -3400 12344 -3080
rect 12664 -3400 12665 -3080
rect 12343 -3401 12665 -3400
rect 11920 -3748 12024 -3452
rect 11331 -3800 11653 -3799
rect 11331 -4120 11332 -3800
rect 11652 -4120 11653 -3800
rect 11331 -4121 11653 -4120
rect 10908 -4468 11012 -4172
rect 10319 -4520 10641 -4519
rect 10319 -4840 10320 -4520
rect 10640 -4840 10641 -4520
rect 10319 -4841 10641 -4840
rect 9896 -5188 10000 -4892
rect 9307 -5240 9629 -5239
rect 9307 -5560 9308 -5240
rect 9628 -5560 9629 -5240
rect 9307 -5561 9629 -5560
rect 8884 -5760 8988 -5612
rect 9416 -5760 9520 -5561
rect 9896 -5612 9916 -5188
rect 9980 -5612 10000 -5188
rect 10428 -5239 10532 -4841
rect 10908 -4892 10928 -4468
rect 10992 -4892 11012 -4468
rect 11440 -4519 11544 -4121
rect 11920 -4172 11940 -3748
rect 12004 -4172 12024 -3748
rect 12452 -3799 12556 -3401
rect 12932 -3452 12952 -3028
rect 13016 -3452 13036 -3028
rect 13464 -3079 13568 -2681
rect 13944 -2732 13964 -2308
rect 14028 -2732 14048 -2308
rect 14476 -2359 14580 -1961
rect 14956 -2012 14976 -1588
rect 15040 -2012 15060 -1588
rect 15488 -1639 15592 -1241
rect 15968 -1292 15988 -868
rect 16052 -1292 16072 -868
rect 16500 -919 16604 -521
rect 16980 -572 17000 -148
rect 17064 -572 17084 -148
rect 17512 -199 17616 199
rect 17992 148 18012 572
rect 18076 148 18096 572
rect 18524 521 18628 919
rect 19004 868 19024 1292
rect 19088 868 19108 1292
rect 19536 1241 19640 1639
rect 20016 1588 20036 2012
rect 20100 1588 20120 2012
rect 20548 1961 20652 2359
rect 21028 2308 21048 2732
rect 21112 2308 21132 2732
rect 21560 2681 21664 3079
rect 22040 3028 22060 3452
rect 22124 3028 22144 3452
rect 22572 3401 22676 3799
rect 23052 3748 23072 4172
rect 23136 3748 23156 4172
rect 23584 4121 23688 4519
rect 24064 4468 24084 4892
rect 24148 4468 24168 4892
rect 24596 4841 24700 5239
rect 25076 5188 25096 5612
rect 25160 5188 25180 5612
rect 25608 5561 25712 5760
rect 26088 5612 26192 5760
rect 25499 5560 25821 5561
rect 25499 5240 25500 5560
rect 25820 5240 25821 5560
rect 25499 5239 25821 5240
rect 25076 4892 25180 5188
rect 24487 4840 24809 4841
rect 24487 4520 24488 4840
rect 24808 4520 24809 4840
rect 24487 4519 24809 4520
rect 24064 4172 24168 4468
rect 23475 4120 23797 4121
rect 23475 3800 23476 4120
rect 23796 3800 23797 4120
rect 23475 3799 23797 3800
rect 23052 3452 23156 3748
rect 22463 3400 22785 3401
rect 22463 3080 22464 3400
rect 22784 3080 22785 3400
rect 22463 3079 22785 3080
rect 22040 2732 22144 3028
rect 21451 2680 21773 2681
rect 21451 2360 21452 2680
rect 21772 2360 21773 2680
rect 21451 2359 21773 2360
rect 21028 2012 21132 2308
rect 20439 1960 20761 1961
rect 20439 1640 20440 1960
rect 20760 1640 20761 1960
rect 20439 1639 20761 1640
rect 20016 1292 20120 1588
rect 19427 1240 19749 1241
rect 19427 920 19428 1240
rect 19748 920 19749 1240
rect 19427 919 19749 920
rect 19004 572 19108 868
rect 18415 520 18737 521
rect 18415 200 18416 520
rect 18736 200 18737 520
rect 18415 199 18737 200
rect 17992 -148 18096 148
rect 17403 -200 17725 -199
rect 17403 -520 17404 -200
rect 17724 -520 17725 -200
rect 17403 -521 17725 -520
rect 16980 -868 17084 -572
rect 16391 -920 16713 -919
rect 16391 -1240 16392 -920
rect 16712 -1240 16713 -920
rect 16391 -1241 16713 -1240
rect 15968 -1588 16072 -1292
rect 15379 -1640 15701 -1639
rect 15379 -1960 15380 -1640
rect 15700 -1960 15701 -1640
rect 15379 -1961 15701 -1960
rect 14956 -2308 15060 -2012
rect 14367 -2360 14689 -2359
rect 14367 -2680 14368 -2360
rect 14688 -2680 14689 -2360
rect 14367 -2681 14689 -2680
rect 13944 -3028 14048 -2732
rect 13355 -3080 13677 -3079
rect 13355 -3400 13356 -3080
rect 13676 -3400 13677 -3080
rect 13355 -3401 13677 -3400
rect 12932 -3748 13036 -3452
rect 12343 -3800 12665 -3799
rect 12343 -4120 12344 -3800
rect 12664 -4120 12665 -3800
rect 12343 -4121 12665 -4120
rect 11920 -4468 12024 -4172
rect 11331 -4520 11653 -4519
rect 11331 -4840 11332 -4520
rect 11652 -4840 11653 -4520
rect 11331 -4841 11653 -4840
rect 10908 -5188 11012 -4892
rect 10319 -5240 10641 -5239
rect 10319 -5560 10320 -5240
rect 10640 -5560 10641 -5240
rect 10319 -5561 10641 -5560
rect 9896 -5760 10000 -5612
rect 10428 -5760 10532 -5561
rect 10908 -5612 10928 -5188
rect 10992 -5612 11012 -5188
rect 11440 -5239 11544 -4841
rect 11920 -4892 11940 -4468
rect 12004 -4892 12024 -4468
rect 12452 -4519 12556 -4121
rect 12932 -4172 12952 -3748
rect 13016 -4172 13036 -3748
rect 13464 -3799 13568 -3401
rect 13944 -3452 13964 -3028
rect 14028 -3452 14048 -3028
rect 14476 -3079 14580 -2681
rect 14956 -2732 14976 -2308
rect 15040 -2732 15060 -2308
rect 15488 -2359 15592 -1961
rect 15968 -2012 15988 -1588
rect 16052 -2012 16072 -1588
rect 16500 -1639 16604 -1241
rect 16980 -1292 17000 -868
rect 17064 -1292 17084 -868
rect 17512 -919 17616 -521
rect 17992 -572 18012 -148
rect 18076 -572 18096 -148
rect 18524 -199 18628 199
rect 19004 148 19024 572
rect 19088 148 19108 572
rect 19536 521 19640 919
rect 20016 868 20036 1292
rect 20100 868 20120 1292
rect 20548 1241 20652 1639
rect 21028 1588 21048 2012
rect 21112 1588 21132 2012
rect 21560 1961 21664 2359
rect 22040 2308 22060 2732
rect 22124 2308 22144 2732
rect 22572 2681 22676 3079
rect 23052 3028 23072 3452
rect 23136 3028 23156 3452
rect 23584 3401 23688 3799
rect 24064 3748 24084 4172
rect 24148 3748 24168 4172
rect 24596 4121 24700 4519
rect 25076 4468 25096 4892
rect 25160 4468 25180 4892
rect 25608 4841 25712 5239
rect 26088 5188 26108 5612
rect 26172 5188 26192 5612
rect 26620 5561 26724 5760
rect 27100 5612 27204 5760
rect 26511 5560 26833 5561
rect 26511 5240 26512 5560
rect 26832 5240 26833 5560
rect 26511 5239 26833 5240
rect 26088 4892 26192 5188
rect 25499 4840 25821 4841
rect 25499 4520 25500 4840
rect 25820 4520 25821 4840
rect 25499 4519 25821 4520
rect 25076 4172 25180 4468
rect 24487 4120 24809 4121
rect 24487 3800 24488 4120
rect 24808 3800 24809 4120
rect 24487 3799 24809 3800
rect 24064 3452 24168 3748
rect 23475 3400 23797 3401
rect 23475 3080 23476 3400
rect 23796 3080 23797 3400
rect 23475 3079 23797 3080
rect 23052 2732 23156 3028
rect 22463 2680 22785 2681
rect 22463 2360 22464 2680
rect 22784 2360 22785 2680
rect 22463 2359 22785 2360
rect 22040 2012 22144 2308
rect 21451 1960 21773 1961
rect 21451 1640 21452 1960
rect 21772 1640 21773 1960
rect 21451 1639 21773 1640
rect 21028 1292 21132 1588
rect 20439 1240 20761 1241
rect 20439 920 20440 1240
rect 20760 920 20761 1240
rect 20439 919 20761 920
rect 20016 572 20120 868
rect 19427 520 19749 521
rect 19427 200 19428 520
rect 19748 200 19749 520
rect 19427 199 19749 200
rect 19004 -148 19108 148
rect 18415 -200 18737 -199
rect 18415 -520 18416 -200
rect 18736 -520 18737 -200
rect 18415 -521 18737 -520
rect 17992 -868 18096 -572
rect 17403 -920 17725 -919
rect 17403 -1240 17404 -920
rect 17724 -1240 17725 -920
rect 17403 -1241 17725 -1240
rect 16980 -1588 17084 -1292
rect 16391 -1640 16713 -1639
rect 16391 -1960 16392 -1640
rect 16712 -1960 16713 -1640
rect 16391 -1961 16713 -1960
rect 15968 -2308 16072 -2012
rect 15379 -2360 15701 -2359
rect 15379 -2680 15380 -2360
rect 15700 -2680 15701 -2360
rect 15379 -2681 15701 -2680
rect 14956 -3028 15060 -2732
rect 14367 -3080 14689 -3079
rect 14367 -3400 14368 -3080
rect 14688 -3400 14689 -3080
rect 14367 -3401 14689 -3400
rect 13944 -3748 14048 -3452
rect 13355 -3800 13677 -3799
rect 13355 -4120 13356 -3800
rect 13676 -4120 13677 -3800
rect 13355 -4121 13677 -4120
rect 12932 -4468 13036 -4172
rect 12343 -4520 12665 -4519
rect 12343 -4840 12344 -4520
rect 12664 -4840 12665 -4520
rect 12343 -4841 12665 -4840
rect 11920 -5188 12024 -4892
rect 11331 -5240 11653 -5239
rect 11331 -5560 11332 -5240
rect 11652 -5560 11653 -5240
rect 11331 -5561 11653 -5560
rect 10908 -5760 11012 -5612
rect 11440 -5760 11544 -5561
rect 11920 -5612 11940 -5188
rect 12004 -5612 12024 -5188
rect 12452 -5239 12556 -4841
rect 12932 -4892 12952 -4468
rect 13016 -4892 13036 -4468
rect 13464 -4519 13568 -4121
rect 13944 -4172 13964 -3748
rect 14028 -4172 14048 -3748
rect 14476 -3799 14580 -3401
rect 14956 -3452 14976 -3028
rect 15040 -3452 15060 -3028
rect 15488 -3079 15592 -2681
rect 15968 -2732 15988 -2308
rect 16052 -2732 16072 -2308
rect 16500 -2359 16604 -1961
rect 16980 -2012 17000 -1588
rect 17064 -2012 17084 -1588
rect 17512 -1639 17616 -1241
rect 17992 -1292 18012 -868
rect 18076 -1292 18096 -868
rect 18524 -919 18628 -521
rect 19004 -572 19024 -148
rect 19088 -572 19108 -148
rect 19536 -199 19640 199
rect 20016 148 20036 572
rect 20100 148 20120 572
rect 20548 521 20652 919
rect 21028 868 21048 1292
rect 21112 868 21132 1292
rect 21560 1241 21664 1639
rect 22040 1588 22060 2012
rect 22124 1588 22144 2012
rect 22572 1961 22676 2359
rect 23052 2308 23072 2732
rect 23136 2308 23156 2732
rect 23584 2681 23688 3079
rect 24064 3028 24084 3452
rect 24148 3028 24168 3452
rect 24596 3401 24700 3799
rect 25076 3748 25096 4172
rect 25160 3748 25180 4172
rect 25608 4121 25712 4519
rect 26088 4468 26108 4892
rect 26172 4468 26192 4892
rect 26620 4841 26724 5239
rect 27100 5188 27120 5612
rect 27184 5188 27204 5612
rect 27632 5561 27736 5760
rect 28112 5612 28216 5760
rect 27523 5560 27845 5561
rect 27523 5240 27524 5560
rect 27844 5240 27845 5560
rect 27523 5239 27845 5240
rect 27100 4892 27204 5188
rect 26511 4840 26833 4841
rect 26511 4520 26512 4840
rect 26832 4520 26833 4840
rect 26511 4519 26833 4520
rect 26088 4172 26192 4468
rect 25499 4120 25821 4121
rect 25499 3800 25500 4120
rect 25820 3800 25821 4120
rect 25499 3799 25821 3800
rect 25076 3452 25180 3748
rect 24487 3400 24809 3401
rect 24487 3080 24488 3400
rect 24808 3080 24809 3400
rect 24487 3079 24809 3080
rect 24064 2732 24168 3028
rect 23475 2680 23797 2681
rect 23475 2360 23476 2680
rect 23796 2360 23797 2680
rect 23475 2359 23797 2360
rect 23052 2012 23156 2308
rect 22463 1960 22785 1961
rect 22463 1640 22464 1960
rect 22784 1640 22785 1960
rect 22463 1639 22785 1640
rect 22040 1292 22144 1588
rect 21451 1240 21773 1241
rect 21451 920 21452 1240
rect 21772 920 21773 1240
rect 21451 919 21773 920
rect 21028 572 21132 868
rect 20439 520 20761 521
rect 20439 200 20440 520
rect 20760 200 20761 520
rect 20439 199 20761 200
rect 20016 -148 20120 148
rect 19427 -200 19749 -199
rect 19427 -520 19428 -200
rect 19748 -520 19749 -200
rect 19427 -521 19749 -520
rect 19004 -868 19108 -572
rect 18415 -920 18737 -919
rect 18415 -1240 18416 -920
rect 18736 -1240 18737 -920
rect 18415 -1241 18737 -1240
rect 17992 -1588 18096 -1292
rect 17403 -1640 17725 -1639
rect 17403 -1960 17404 -1640
rect 17724 -1960 17725 -1640
rect 17403 -1961 17725 -1960
rect 16980 -2308 17084 -2012
rect 16391 -2360 16713 -2359
rect 16391 -2680 16392 -2360
rect 16712 -2680 16713 -2360
rect 16391 -2681 16713 -2680
rect 15968 -3028 16072 -2732
rect 15379 -3080 15701 -3079
rect 15379 -3400 15380 -3080
rect 15700 -3400 15701 -3080
rect 15379 -3401 15701 -3400
rect 14956 -3748 15060 -3452
rect 14367 -3800 14689 -3799
rect 14367 -4120 14368 -3800
rect 14688 -4120 14689 -3800
rect 14367 -4121 14689 -4120
rect 13944 -4468 14048 -4172
rect 13355 -4520 13677 -4519
rect 13355 -4840 13356 -4520
rect 13676 -4840 13677 -4520
rect 13355 -4841 13677 -4840
rect 12932 -5188 13036 -4892
rect 12343 -5240 12665 -5239
rect 12343 -5560 12344 -5240
rect 12664 -5560 12665 -5240
rect 12343 -5561 12665 -5560
rect 11920 -5760 12024 -5612
rect 12452 -5760 12556 -5561
rect 12932 -5612 12952 -5188
rect 13016 -5612 13036 -5188
rect 13464 -5239 13568 -4841
rect 13944 -4892 13964 -4468
rect 14028 -4892 14048 -4468
rect 14476 -4519 14580 -4121
rect 14956 -4172 14976 -3748
rect 15040 -4172 15060 -3748
rect 15488 -3799 15592 -3401
rect 15968 -3452 15988 -3028
rect 16052 -3452 16072 -3028
rect 16500 -3079 16604 -2681
rect 16980 -2732 17000 -2308
rect 17064 -2732 17084 -2308
rect 17512 -2359 17616 -1961
rect 17992 -2012 18012 -1588
rect 18076 -2012 18096 -1588
rect 18524 -1639 18628 -1241
rect 19004 -1292 19024 -868
rect 19088 -1292 19108 -868
rect 19536 -919 19640 -521
rect 20016 -572 20036 -148
rect 20100 -572 20120 -148
rect 20548 -199 20652 199
rect 21028 148 21048 572
rect 21112 148 21132 572
rect 21560 521 21664 919
rect 22040 868 22060 1292
rect 22124 868 22144 1292
rect 22572 1241 22676 1639
rect 23052 1588 23072 2012
rect 23136 1588 23156 2012
rect 23584 1961 23688 2359
rect 24064 2308 24084 2732
rect 24148 2308 24168 2732
rect 24596 2681 24700 3079
rect 25076 3028 25096 3452
rect 25160 3028 25180 3452
rect 25608 3401 25712 3799
rect 26088 3748 26108 4172
rect 26172 3748 26192 4172
rect 26620 4121 26724 4519
rect 27100 4468 27120 4892
rect 27184 4468 27204 4892
rect 27632 4841 27736 5239
rect 28112 5188 28132 5612
rect 28196 5188 28216 5612
rect 28644 5561 28748 5760
rect 29124 5612 29228 5760
rect 28535 5560 28857 5561
rect 28535 5240 28536 5560
rect 28856 5240 28857 5560
rect 28535 5239 28857 5240
rect 28112 4892 28216 5188
rect 27523 4840 27845 4841
rect 27523 4520 27524 4840
rect 27844 4520 27845 4840
rect 27523 4519 27845 4520
rect 27100 4172 27204 4468
rect 26511 4120 26833 4121
rect 26511 3800 26512 4120
rect 26832 3800 26833 4120
rect 26511 3799 26833 3800
rect 26088 3452 26192 3748
rect 25499 3400 25821 3401
rect 25499 3080 25500 3400
rect 25820 3080 25821 3400
rect 25499 3079 25821 3080
rect 25076 2732 25180 3028
rect 24487 2680 24809 2681
rect 24487 2360 24488 2680
rect 24808 2360 24809 2680
rect 24487 2359 24809 2360
rect 24064 2012 24168 2308
rect 23475 1960 23797 1961
rect 23475 1640 23476 1960
rect 23796 1640 23797 1960
rect 23475 1639 23797 1640
rect 23052 1292 23156 1588
rect 22463 1240 22785 1241
rect 22463 920 22464 1240
rect 22784 920 22785 1240
rect 22463 919 22785 920
rect 22040 572 22144 868
rect 21451 520 21773 521
rect 21451 200 21452 520
rect 21772 200 21773 520
rect 21451 199 21773 200
rect 21028 -148 21132 148
rect 20439 -200 20761 -199
rect 20439 -520 20440 -200
rect 20760 -520 20761 -200
rect 20439 -521 20761 -520
rect 20016 -868 20120 -572
rect 19427 -920 19749 -919
rect 19427 -1240 19428 -920
rect 19748 -1240 19749 -920
rect 19427 -1241 19749 -1240
rect 19004 -1588 19108 -1292
rect 18415 -1640 18737 -1639
rect 18415 -1960 18416 -1640
rect 18736 -1960 18737 -1640
rect 18415 -1961 18737 -1960
rect 17992 -2308 18096 -2012
rect 17403 -2360 17725 -2359
rect 17403 -2680 17404 -2360
rect 17724 -2680 17725 -2360
rect 17403 -2681 17725 -2680
rect 16980 -3028 17084 -2732
rect 16391 -3080 16713 -3079
rect 16391 -3400 16392 -3080
rect 16712 -3400 16713 -3080
rect 16391 -3401 16713 -3400
rect 15968 -3748 16072 -3452
rect 15379 -3800 15701 -3799
rect 15379 -4120 15380 -3800
rect 15700 -4120 15701 -3800
rect 15379 -4121 15701 -4120
rect 14956 -4468 15060 -4172
rect 14367 -4520 14689 -4519
rect 14367 -4840 14368 -4520
rect 14688 -4840 14689 -4520
rect 14367 -4841 14689 -4840
rect 13944 -5188 14048 -4892
rect 13355 -5240 13677 -5239
rect 13355 -5560 13356 -5240
rect 13676 -5560 13677 -5240
rect 13355 -5561 13677 -5560
rect 12932 -5760 13036 -5612
rect 13464 -5760 13568 -5561
rect 13944 -5612 13964 -5188
rect 14028 -5612 14048 -5188
rect 14476 -5239 14580 -4841
rect 14956 -4892 14976 -4468
rect 15040 -4892 15060 -4468
rect 15488 -4519 15592 -4121
rect 15968 -4172 15988 -3748
rect 16052 -4172 16072 -3748
rect 16500 -3799 16604 -3401
rect 16980 -3452 17000 -3028
rect 17064 -3452 17084 -3028
rect 17512 -3079 17616 -2681
rect 17992 -2732 18012 -2308
rect 18076 -2732 18096 -2308
rect 18524 -2359 18628 -1961
rect 19004 -2012 19024 -1588
rect 19088 -2012 19108 -1588
rect 19536 -1639 19640 -1241
rect 20016 -1292 20036 -868
rect 20100 -1292 20120 -868
rect 20548 -919 20652 -521
rect 21028 -572 21048 -148
rect 21112 -572 21132 -148
rect 21560 -199 21664 199
rect 22040 148 22060 572
rect 22124 148 22144 572
rect 22572 521 22676 919
rect 23052 868 23072 1292
rect 23136 868 23156 1292
rect 23584 1241 23688 1639
rect 24064 1588 24084 2012
rect 24148 1588 24168 2012
rect 24596 1961 24700 2359
rect 25076 2308 25096 2732
rect 25160 2308 25180 2732
rect 25608 2681 25712 3079
rect 26088 3028 26108 3452
rect 26172 3028 26192 3452
rect 26620 3401 26724 3799
rect 27100 3748 27120 4172
rect 27184 3748 27204 4172
rect 27632 4121 27736 4519
rect 28112 4468 28132 4892
rect 28196 4468 28216 4892
rect 28644 4841 28748 5239
rect 29124 5188 29144 5612
rect 29208 5188 29228 5612
rect 29656 5561 29760 5760
rect 30136 5612 30240 5760
rect 29547 5560 29869 5561
rect 29547 5240 29548 5560
rect 29868 5240 29869 5560
rect 29547 5239 29869 5240
rect 29124 4892 29228 5188
rect 28535 4840 28857 4841
rect 28535 4520 28536 4840
rect 28856 4520 28857 4840
rect 28535 4519 28857 4520
rect 28112 4172 28216 4468
rect 27523 4120 27845 4121
rect 27523 3800 27524 4120
rect 27844 3800 27845 4120
rect 27523 3799 27845 3800
rect 27100 3452 27204 3748
rect 26511 3400 26833 3401
rect 26511 3080 26512 3400
rect 26832 3080 26833 3400
rect 26511 3079 26833 3080
rect 26088 2732 26192 3028
rect 25499 2680 25821 2681
rect 25499 2360 25500 2680
rect 25820 2360 25821 2680
rect 25499 2359 25821 2360
rect 25076 2012 25180 2308
rect 24487 1960 24809 1961
rect 24487 1640 24488 1960
rect 24808 1640 24809 1960
rect 24487 1639 24809 1640
rect 24064 1292 24168 1588
rect 23475 1240 23797 1241
rect 23475 920 23476 1240
rect 23796 920 23797 1240
rect 23475 919 23797 920
rect 23052 572 23156 868
rect 22463 520 22785 521
rect 22463 200 22464 520
rect 22784 200 22785 520
rect 22463 199 22785 200
rect 22040 -148 22144 148
rect 21451 -200 21773 -199
rect 21451 -520 21452 -200
rect 21772 -520 21773 -200
rect 21451 -521 21773 -520
rect 21028 -868 21132 -572
rect 20439 -920 20761 -919
rect 20439 -1240 20440 -920
rect 20760 -1240 20761 -920
rect 20439 -1241 20761 -1240
rect 20016 -1588 20120 -1292
rect 19427 -1640 19749 -1639
rect 19427 -1960 19428 -1640
rect 19748 -1960 19749 -1640
rect 19427 -1961 19749 -1960
rect 19004 -2308 19108 -2012
rect 18415 -2360 18737 -2359
rect 18415 -2680 18416 -2360
rect 18736 -2680 18737 -2360
rect 18415 -2681 18737 -2680
rect 17992 -3028 18096 -2732
rect 17403 -3080 17725 -3079
rect 17403 -3400 17404 -3080
rect 17724 -3400 17725 -3080
rect 17403 -3401 17725 -3400
rect 16980 -3748 17084 -3452
rect 16391 -3800 16713 -3799
rect 16391 -4120 16392 -3800
rect 16712 -4120 16713 -3800
rect 16391 -4121 16713 -4120
rect 15968 -4468 16072 -4172
rect 15379 -4520 15701 -4519
rect 15379 -4840 15380 -4520
rect 15700 -4840 15701 -4520
rect 15379 -4841 15701 -4840
rect 14956 -5188 15060 -4892
rect 14367 -5240 14689 -5239
rect 14367 -5560 14368 -5240
rect 14688 -5560 14689 -5240
rect 14367 -5561 14689 -5560
rect 13944 -5760 14048 -5612
rect 14476 -5760 14580 -5561
rect 14956 -5612 14976 -5188
rect 15040 -5612 15060 -5188
rect 15488 -5239 15592 -4841
rect 15968 -4892 15988 -4468
rect 16052 -4892 16072 -4468
rect 16500 -4519 16604 -4121
rect 16980 -4172 17000 -3748
rect 17064 -4172 17084 -3748
rect 17512 -3799 17616 -3401
rect 17992 -3452 18012 -3028
rect 18076 -3452 18096 -3028
rect 18524 -3079 18628 -2681
rect 19004 -2732 19024 -2308
rect 19088 -2732 19108 -2308
rect 19536 -2359 19640 -1961
rect 20016 -2012 20036 -1588
rect 20100 -2012 20120 -1588
rect 20548 -1639 20652 -1241
rect 21028 -1292 21048 -868
rect 21112 -1292 21132 -868
rect 21560 -919 21664 -521
rect 22040 -572 22060 -148
rect 22124 -572 22144 -148
rect 22572 -199 22676 199
rect 23052 148 23072 572
rect 23136 148 23156 572
rect 23584 521 23688 919
rect 24064 868 24084 1292
rect 24148 868 24168 1292
rect 24596 1241 24700 1639
rect 25076 1588 25096 2012
rect 25160 1588 25180 2012
rect 25608 1961 25712 2359
rect 26088 2308 26108 2732
rect 26172 2308 26192 2732
rect 26620 2681 26724 3079
rect 27100 3028 27120 3452
rect 27184 3028 27204 3452
rect 27632 3401 27736 3799
rect 28112 3748 28132 4172
rect 28196 3748 28216 4172
rect 28644 4121 28748 4519
rect 29124 4468 29144 4892
rect 29208 4468 29228 4892
rect 29656 4841 29760 5239
rect 30136 5188 30156 5612
rect 30220 5188 30240 5612
rect 30668 5561 30772 5760
rect 31148 5612 31252 5760
rect 30559 5560 30881 5561
rect 30559 5240 30560 5560
rect 30880 5240 30881 5560
rect 30559 5239 30881 5240
rect 30136 4892 30240 5188
rect 29547 4840 29869 4841
rect 29547 4520 29548 4840
rect 29868 4520 29869 4840
rect 29547 4519 29869 4520
rect 29124 4172 29228 4468
rect 28535 4120 28857 4121
rect 28535 3800 28536 4120
rect 28856 3800 28857 4120
rect 28535 3799 28857 3800
rect 28112 3452 28216 3748
rect 27523 3400 27845 3401
rect 27523 3080 27524 3400
rect 27844 3080 27845 3400
rect 27523 3079 27845 3080
rect 27100 2732 27204 3028
rect 26511 2680 26833 2681
rect 26511 2360 26512 2680
rect 26832 2360 26833 2680
rect 26511 2359 26833 2360
rect 26088 2012 26192 2308
rect 25499 1960 25821 1961
rect 25499 1640 25500 1960
rect 25820 1640 25821 1960
rect 25499 1639 25821 1640
rect 25076 1292 25180 1588
rect 24487 1240 24809 1241
rect 24487 920 24488 1240
rect 24808 920 24809 1240
rect 24487 919 24809 920
rect 24064 572 24168 868
rect 23475 520 23797 521
rect 23475 200 23476 520
rect 23796 200 23797 520
rect 23475 199 23797 200
rect 23052 -148 23156 148
rect 22463 -200 22785 -199
rect 22463 -520 22464 -200
rect 22784 -520 22785 -200
rect 22463 -521 22785 -520
rect 22040 -868 22144 -572
rect 21451 -920 21773 -919
rect 21451 -1240 21452 -920
rect 21772 -1240 21773 -920
rect 21451 -1241 21773 -1240
rect 21028 -1588 21132 -1292
rect 20439 -1640 20761 -1639
rect 20439 -1960 20440 -1640
rect 20760 -1960 20761 -1640
rect 20439 -1961 20761 -1960
rect 20016 -2308 20120 -2012
rect 19427 -2360 19749 -2359
rect 19427 -2680 19428 -2360
rect 19748 -2680 19749 -2360
rect 19427 -2681 19749 -2680
rect 19004 -3028 19108 -2732
rect 18415 -3080 18737 -3079
rect 18415 -3400 18416 -3080
rect 18736 -3400 18737 -3080
rect 18415 -3401 18737 -3400
rect 17992 -3748 18096 -3452
rect 17403 -3800 17725 -3799
rect 17403 -4120 17404 -3800
rect 17724 -4120 17725 -3800
rect 17403 -4121 17725 -4120
rect 16980 -4468 17084 -4172
rect 16391 -4520 16713 -4519
rect 16391 -4840 16392 -4520
rect 16712 -4840 16713 -4520
rect 16391 -4841 16713 -4840
rect 15968 -5188 16072 -4892
rect 15379 -5240 15701 -5239
rect 15379 -5560 15380 -5240
rect 15700 -5560 15701 -5240
rect 15379 -5561 15701 -5560
rect 14956 -5760 15060 -5612
rect 15488 -5760 15592 -5561
rect 15968 -5612 15988 -5188
rect 16052 -5612 16072 -5188
rect 16500 -5239 16604 -4841
rect 16980 -4892 17000 -4468
rect 17064 -4892 17084 -4468
rect 17512 -4519 17616 -4121
rect 17992 -4172 18012 -3748
rect 18076 -4172 18096 -3748
rect 18524 -3799 18628 -3401
rect 19004 -3452 19024 -3028
rect 19088 -3452 19108 -3028
rect 19536 -3079 19640 -2681
rect 20016 -2732 20036 -2308
rect 20100 -2732 20120 -2308
rect 20548 -2359 20652 -1961
rect 21028 -2012 21048 -1588
rect 21112 -2012 21132 -1588
rect 21560 -1639 21664 -1241
rect 22040 -1292 22060 -868
rect 22124 -1292 22144 -868
rect 22572 -919 22676 -521
rect 23052 -572 23072 -148
rect 23136 -572 23156 -148
rect 23584 -199 23688 199
rect 24064 148 24084 572
rect 24148 148 24168 572
rect 24596 521 24700 919
rect 25076 868 25096 1292
rect 25160 868 25180 1292
rect 25608 1241 25712 1639
rect 26088 1588 26108 2012
rect 26172 1588 26192 2012
rect 26620 1961 26724 2359
rect 27100 2308 27120 2732
rect 27184 2308 27204 2732
rect 27632 2681 27736 3079
rect 28112 3028 28132 3452
rect 28196 3028 28216 3452
rect 28644 3401 28748 3799
rect 29124 3748 29144 4172
rect 29208 3748 29228 4172
rect 29656 4121 29760 4519
rect 30136 4468 30156 4892
rect 30220 4468 30240 4892
rect 30668 4841 30772 5239
rect 31148 5188 31168 5612
rect 31232 5188 31252 5612
rect 31680 5561 31784 5760
rect 32160 5612 32264 5760
rect 31571 5560 31893 5561
rect 31571 5240 31572 5560
rect 31892 5240 31893 5560
rect 31571 5239 31893 5240
rect 31148 4892 31252 5188
rect 30559 4840 30881 4841
rect 30559 4520 30560 4840
rect 30880 4520 30881 4840
rect 30559 4519 30881 4520
rect 30136 4172 30240 4468
rect 29547 4120 29869 4121
rect 29547 3800 29548 4120
rect 29868 3800 29869 4120
rect 29547 3799 29869 3800
rect 29124 3452 29228 3748
rect 28535 3400 28857 3401
rect 28535 3080 28536 3400
rect 28856 3080 28857 3400
rect 28535 3079 28857 3080
rect 28112 2732 28216 3028
rect 27523 2680 27845 2681
rect 27523 2360 27524 2680
rect 27844 2360 27845 2680
rect 27523 2359 27845 2360
rect 27100 2012 27204 2308
rect 26511 1960 26833 1961
rect 26511 1640 26512 1960
rect 26832 1640 26833 1960
rect 26511 1639 26833 1640
rect 26088 1292 26192 1588
rect 25499 1240 25821 1241
rect 25499 920 25500 1240
rect 25820 920 25821 1240
rect 25499 919 25821 920
rect 25076 572 25180 868
rect 24487 520 24809 521
rect 24487 200 24488 520
rect 24808 200 24809 520
rect 24487 199 24809 200
rect 24064 -148 24168 148
rect 23475 -200 23797 -199
rect 23475 -520 23476 -200
rect 23796 -520 23797 -200
rect 23475 -521 23797 -520
rect 23052 -868 23156 -572
rect 22463 -920 22785 -919
rect 22463 -1240 22464 -920
rect 22784 -1240 22785 -920
rect 22463 -1241 22785 -1240
rect 22040 -1588 22144 -1292
rect 21451 -1640 21773 -1639
rect 21451 -1960 21452 -1640
rect 21772 -1960 21773 -1640
rect 21451 -1961 21773 -1960
rect 21028 -2308 21132 -2012
rect 20439 -2360 20761 -2359
rect 20439 -2680 20440 -2360
rect 20760 -2680 20761 -2360
rect 20439 -2681 20761 -2680
rect 20016 -3028 20120 -2732
rect 19427 -3080 19749 -3079
rect 19427 -3400 19428 -3080
rect 19748 -3400 19749 -3080
rect 19427 -3401 19749 -3400
rect 19004 -3748 19108 -3452
rect 18415 -3800 18737 -3799
rect 18415 -4120 18416 -3800
rect 18736 -4120 18737 -3800
rect 18415 -4121 18737 -4120
rect 17992 -4468 18096 -4172
rect 17403 -4520 17725 -4519
rect 17403 -4840 17404 -4520
rect 17724 -4840 17725 -4520
rect 17403 -4841 17725 -4840
rect 16980 -5188 17084 -4892
rect 16391 -5240 16713 -5239
rect 16391 -5560 16392 -5240
rect 16712 -5560 16713 -5240
rect 16391 -5561 16713 -5560
rect 15968 -5760 16072 -5612
rect 16500 -5760 16604 -5561
rect 16980 -5612 17000 -5188
rect 17064 -5612 17084 -5188
rect 17512 -5239 17616 -4841
rect 17992 -4892 18012 -4468
rect 18076 -4892 18096 -4468
rect 18524 -4519 18628 -4121
rect 19004 -4172 19024 -3748
rect 19088 -4172 19108 -3748
rect 19536 -3799 19640 -3401
rect 20016 -3452 20036 -3028
rect 20100 -3452 20120 -3028
rect 20548 -3079 20652 -2681
rect 21028 -2732 21048 -2308
rect 21112 -2732 21132 -2308
rect 21560 -2359 21664 -1961
rect 22040 -2012 22060 -1588
rect 22124 -2012 22144 -1588
rect 22572 -1639 22676 -1241
rect 23052 -1292 23072 -868
rect 23136 -1292 23156 -868
rect 23584 -919 23688 -521
rect 24064 -572 24084 -148
rect 24148 -572 24168 -148
rect 24596 -199 24700 199
rect 25076 148 25096 572
rect 25160 148 25180 572
rect 25608 521 25712 919
rect 26088 868 26108 1292
rect 26172 868 26192 1292
rect 26620 1241 26724 1639
rect 27100 1588 27120 2012
rect 27184 1588 27204 2012
rect 27632 1961 27736 2359
rect 28112 2308 28132 2732
rect 28196 2308 28216 2732
rect 28644 2681 28748 3079
rect 29124 3028 29144 3452
rect 29208 3028 29228 3452
rect 29656 3401 29760 3799
rect 30136 3748 30156 4172
rect 30220 3748 30240 4172
rect 30668 4121 30772 4519
rect 31148 4468 31168 4892
rect 31232 4468 31252 4892
rect 31680 4841 31784 5239
rect 32160 5188 32180 5612
rect 32244 5188 32264 5612
rect 32160 4892 32264 5188
rect 31571 4840 31893 4841
rect 31571 4520 31572 4840
rect 31892 4520 31893 4840
rect 31571 4519 31893 4520
rect 31148 4172 31252 4468
rect 30559 4120 30881 4121
rect 30559 3800 30560 4120
rect 30880 3800 30881 4120
rect 30559 3799 30881 3800
rect 30136 3452 30240 3748
rect 29547 3400 29869 3401
rect 29547 3080 29548 3400
rect 29868 3080 29869 3400
rect 29547 3079 29869 3080
rect 29124 2732 29228 3028
rect 28535 2680 28857 2681
rect 28535 2360 28536 2680
rect 28856 2360 28857 2680
rect 28535 2359 28857 2360
rect 28112 2012 28216 2308
rect 27523 1960 27845 1961
rect 27523 1640 27524 1960
rect 27844 1640 27845 1960
rect 27523 1639 27845 1640
rect 27100 1292 27204 1588
rect 26511 1240 26833 1241
rect 26511 920 26512 1240
rect 26832 920 26833 1240
rect 26511 919 26833 920
rect 26088 572 26192 868
rect 25499 520 25821 521
rect 25499 200 25500 520
rect 25820 200 25821 520
rect 25499 199 25821 200
rect 25076 -148 25180 148
rect 24487 -200 24809 -199
rect 24487 -520 24488 -200
rect 24808 -520 24809 -200
rect 24487 -521 24809 -520
rect 24064 -868 24168 -572
rect 23475 -920 23797 -919
rect 23475 -1240 23476 -920
rect 23796 -1240 23797 -920
rect 23475 -1241 23797 -1240
rect 23052 -1588 23156 -1292
rect 22463 -1640 22785 -1639
rect 22463 -1960 22464 -1640
rect 22784 -1960 22785 -1640
rect 22463 -1961 22785 -1960
rect 22040 -2308 22144 -2012
rect 21451 -2360 21773 -2359
rect 21451 -2680 21452 -2360
rect 21772 -2680 21773 -2360
rect 21451 -2681 21773 -2680
rect 21028 -3028 21132 -2732
rect 20439 -3080 20761 -3079
rect 20439 -3400 20440 -3080
rect 20760 -3400 20761 -3080
rect 20439 -3401 20761 -3400
rect 20016 -3748 20120 -3452
rect 19427 -3800 19749 -3799
rect 19427 -4120 19428 -3800
rect 19748 -4120 19749 -3800
rect 19427 -4121 19749 -4120
rect 19004 -4468 19108 -4172
rect 18415 -4520 18737 -4519
rect 18415 -4840 18416 -4520
rect 18736 -4840 18737 -4520
rect 18415 -4841 18737 -4840
rect 17992 -5188 18096 -4892
rect 17403 -5240 17725 -5239
rect 17403 -5560 17404 -5240
rect 17724 -5560 17725 -5240
rect 17403 -5561 17725 -5560
rect 16980 -5760 17084 -5612
rect 17512 -5760 17616 -5561
rect 17992 -5612 18012 -5188
rect 18076 -5612 18096 -5188
rect 18524 -5239 18628 -4841
rect 19004 -4892 19024 -4468
rect 19088 -4892 19108 -4468
rect 19536 -4519 19640 -4121
rect 20016 -4172 20036 -3748
rect 20100 -4172 20120 -3748
rect 20548 -3799 20652 -3401
rect 21028 -3452 21048 -3028
rect 21112 -3452 21132 -3028
rect 21560 -3079 21664 -2681
rect 22040 -2732 22060 -2308
rect 22124 -2732 22144 -2308
rect 22572 -2359 22676 -1961
rect 23052 -2012 23072 -1588
rect 23136 -2012 23156 -1588
rect 23584 -1639 23688 -1241
rect 24064 -1292 24084 -868
rect 24148 -1292 24168 -868
rect 24596 -919 24700 -521
rect 25076 -572 25096 -148
rect 25160 -572 25180 -148
rect 25608 -199 25712 199
rect 26088 148 26108 572
rect 26172 148 26192 572
rect 26620 521 26724 919
rect 27100 868 27120 1292
rect 27184 868 27204 1292
rect 27632 1241 27736 1639
rect 28112 1588 28132 2012
rect 28196 1588 28216 2012
rect 28644 1961 28748 2359
rect 29124 2308 29144 2732
rect 29208 2308 29228 2732
rect 29656 2681 29760 3079
rect 30136 3028 30156 3452
rect 30220 3028 30240 3452
rect 30668 3401 30772 3799
rect 31148 3748 31168 4172
rect 31232 3748 31252 4172
rect 31680 4121 31784 4519
rect 32160 4468 32180 4892
rect 32244 4468 32264 4892
rect 32160 4172 32264 4468
rect 31571 4120 31893 4121
rect 31571 3800 31572 4120
rect 31892 3800 31893 4120
rect 31571 3799 31893 3800
rect 31148 3452 31252 3748
rect 30559 3400 30881 3401
rect 30559 3080 30560 3400
rect 30880 3080 30881 3400
rect 30559 3079 30881 3080
rect 30136 2732 30240 3028
rect 29547 2680 29869 2681
rect 29547 2360 29548 2680
rect 29868 2360 29869 2680
rect 29547 2359 29869 2360
rect 29124 2012 29228 2308
rect 28535 1960 28857 1961
rect 28535 1640 28536 1960
rect 28856 1640 28857 1960
rect 28535 1639 28857 1640
rect 28112 1292 28216 1588
rect 27523 1240 27845 1241
rect 27523 920 27524 1240
rect 27844 920 27845 1240
rect 27523 919 27845 920
rect 27100 572 27204 868
rect 26511 520 26833 521
rect 26511 200 26512 520
rect 26832 200 26833 520
rect 26511 199 26833 200
rect 26088 -148 26192 148
rect 25499 -200 25821 -199
rect 25499 -520 25500 -200
rect 25820 -520 25821 -200
rect 25499 -521 25821 -520
rect 25076 -868 25180 -572
rect 24487 -920 24809 -919
rect 24487 -1240 24488 -920
rect 24808 -1240 24809 -920
rect 24487 -1241 24809 -1240
rect 24064 -1588 24168 -1292
rect 23475 -1640 23797 -1639
rect 23475 -1960 23476 -1640
rect 23796 -1960 23797 -1640
rect 23475 -1961 23797 -1960
rect 23052 -2308 23156 -2012
rect 22463 -2360 22785 -2359
rect 22463 -2680 22464 -2360
rect 22784 -2680 22785 -2360
rect 22463 -2681 22785 -2680
rect 22040 -3028 22144 -2732
rect 21451 -3080 21773 -3079
rect 21451 -3400 21452 -3080
rect 21772 -3400 21773 -3080
rect 21451 -3401 21773 -3400
rect 21028 -3748 21132 -3452
rect 20439 -3800 20761 -3799
rect 20439 -4120 20440 -3800
rect 20760 -4120 20761 -3800
rect 20439 -4121 20761 -4120
rect 20016 -4468 20120 -4172
rect 19427 -4520 19749 -4519
rect 19427 -4840 19428 -4520
rect 19748 -4840 19749 -4520
rect 19427 -4841 19749 -4840
rect 19004 -5188 19108 -4892
rect 18415 -5240 18737 -5239
rect 18415 -5560 18416 -5240
rect 18736 -5560 18737 -5240
rect 18415 -5561 18737 -5560
rect 17992 -5760 18096 -5612
rect 18524 -5760 18628 -5561
rect 19004 -5612 19024 -5188
rect 19088 -5612 19108 -5188
rect 19536 -5239 19640 -4841
rect 20016 -4892 20036 -4468
rect 20100 -4892 20120 -4468
rect 20548 -4519 20652 -4121
rect 21028 -4172 21048 -3748
rect 21112 -4172 21132 -3748
rect 21560 -3799 21664 -3401
rect 22040 -3452 22060 -3028
rect 22124 -3452 22144 -3028
rect 22572 -3079 22676 -2681
rect 23052 -2732 23072 -2308
rect 23136 -2732 23156 -2308
rect 23584 -2359 23688 -1961
rect 24064 -2012 24084 -1588
rect 24148 -2012 24168 -1588
rect 24596 -1639 24700 -1241
rect 25076 -1292 25096 -868
rect 25160 -1292 25180 -868
rect 25608 -919 25712 -521
rect 26088 -572 26108 -148
rect 26172 -572 26192 -148
rect 26620 -199 26724 199
rect 27100 148 27120 572
rect 27184 148 27204 572
rect 27632 521 27736 919
rect 28112 868 28132 1292
rect 28196 868 28216 1292
rect 28644 1241 28748 1639
rect 29124 1588 29144 2012
rect 29208 1588 29228 2012
rect 29656 1961 29760 2359
rect 30136 2308 30156 2732
rect 30220 2308 30240 2732
rect 30668 2681 30772 3079
rect 31148 3028 31168 3452
rect 31232 3028 31252 3452
rect 31680 3401 31784 3799
rect 32160 3748 32180 4172
rect 32244 3748 32264 4172
rect 32160 3452 32264 3748
rect 31571 3400 31893 3401
rect 31571 3080 31572 3400
rect 31892 3080 31893 3400
rect 31571 3079 31893 3080
rect 31148 2732 31252 3028
rect 30559 2680 30881 2681
rect 30559 2360 30560 2680
rect 30880 2360 30881 2680
rect 30559 2359 30881 2360
rect 30136 2012 30240 2308
rect 29547 1960 29869 1961
rect 29547 1640 29548 1960
rect 29868 1640 29869 1960
rect 29547 1639 29869 1640
rect 29124 1292 29228 1588
rect 28535 1240 28857 1241
rect 28535 920 28536 1240
rect 28856 920 28857 1240
rect 28535 919 28857 920
rect 28112 572 28216 868
rect 27523 520 27845 521
rect 27523 200 27524 520
rect 27844 200 27845 520
rect 27523 199 27845 200
rect 27100 -148 27204 148
rect 26511 -200 26833 -199
rect 26511 -520 26512 -200
rect 26832 -520 26833 -200
rect 26511 -521 26833 -520
rect 26088 -868 26192 -572
rect 25499 -920 25821 -919
rect 25499 -1240 25500 -920
rect 25820 -1240 25821 -920
rect 25499 -1241 25821 -1240
rect 25076 -1588 25180 -1292
rect 24487 -1640 24809 -1639
rect 24487 -1960 24488 -1640
rect 24808 -1960 24809 -1640
rect 24487 -1961 24809 -1960
rect 24064 -2308 24168 -2012
rect 23475 -2360 23797 -2359
rect 23475 -2680 23476 -2360
rect 23796 -2680 23797 -2360
rect 23475 -2681 23797 -2680
rect 23052 -3028 23156 -2732
rect 22463 -3080 22785 -3079
rect 22463 -3400 22464 -3080
rect 22784 -3400 22785 -3080
rect 22463 -3401 22785 -3400
rect 22040 -3748 22144 -3452
rect 21451 -3800 21773 -3799
rect 21451 -4120 21452 -3800
rect 21772 -4120 21773 -3800
rect 21451 -4121 21773 -4120
rect 21028 -4468 21132 -4172
rect 20439 -4520 20761 -4519
rect 20439 -4840 20440 -4520
rect 20760 -4840 20761 -4520
rect 20439 -4841 20761 -4840
rect 20016 -5188 20120 -4892
rect 19427 -5240 19749 -5239
rect 19427 -5560 19428 -5240
rect 19748 -5560 19749 -5240
rect 19427 -5561 19749 -5560
rect 19004 -5760 19108 -5612
rect 19536 -5760 19640 -5561
rect 20016 -5612 20036 -5188
rect 20100 -5612 20120 -5188
rect 20548 -5239 20652 -4841
rect 21028 -4892 21048 -4468
rect 21112 -4892 21132 -4468
rect 21560 -4519 21664 -4121
rect 22040 -4172 22060 -3748
rect 22124 -4172 22144 -3748
rect 22572 -3799 22676 -3401
rect 23052 -3452 23072 -3028
rect 23136 -3452 23156 -3028
rect 23584 -3079 23688 -2681
rect 24064 -2732 24084 -2308
rect 24148 -2732 24168 -2308
rect 24596 -2359 24700 -1961
rect 25076 -2012 25096 -1588
rect 25160 -2012 25180 -1588
rect 25608 -1639 25712 -1241
rect 26088 -1292 26108 -868
rect 26172 -1292 26192 -868
rect 26620 -919 26724 -521
rect 27100 -572 27120 -148
rect 27184 -572 27204 -148
rect 27632 -199 27736 199
rect 28112 148 28132 572
rect 28196 148 28216 572
rect 28644 521 28748 919
rect 29124 868 29144 1292
rect 29208 868 29228 1292
rect 29656 1241 29760 1639
rect 30136 1588 30156 2012
rect 30220 1588 30240 2012
rect 30668 1961 30772 2359
rect 31148 2308 31168 2732
rect 31232 2308 31252 2732
rect 31680 2681 31784 3079
rect 32160 3028 32180 3452
rect 32244 3028 32264 3452
rect 32160 2732 32264 3028
rect 31571 2680 31893 2681
rect 31571 2360 31572 2680
rect 31892 2360 31893 2680
rect 31571 2359 31893 2360
rect 31148 2012 31252 2308
rect 30559 1960 30881 1961
rect 30559 1640 30560 1960
rect 30880 1640 30881 1960
rect 30559 1639 30881 1640
rect 30136 1292 30240 1588
rect 29547 1240 29869 1241
rect 29547 920 29548 1240
rect 29868 920 29869 1240
rect 29547 919 29869 920
rect 29124 572 29228 868
rect 28535 520 28857 521
rect 28535 200 28536 520
rect 28856 200 28857 520
rect 28535 199 28857 200
rect 28112 -148 28216 148
rect 27523 -200 27845 -199
rect 27523 -520 27524 -200
rect 27844 -520 27845 -200
rect 27523 -521 27845 -520
rect 27100 -868 27204 -572
rect 26511 -920 26833 -919
rect 26511 -1240 26512 -920
rect 26832 -1240 26833 -920
rect 26511 -1241 26833 -1240
rect 26088 -1588 26192 -1292
rect 25499 -1640 25821 -1639
rect 25499 -1960 25500 -1640
rect 25820 -1960 25821 -1640
rect 25499 -1961 25821 -1960
rect 25076 -2308 25180 -2012
rect 24487 -2360 24809 -2359
rect 24487 -2680 24488 -2360
rect 24808 -2680 24809 -2360
rect 24487 -2681 24809 -2680
rect 24064 -3028 24168 -2732
rect 23475 -3080 23797 -3079
rect 23475 -3400 23476 -3080
rect 23796 -3400 23797 -3080
rect 23475 -3401 23797 -3400
rect 23052 -3748 23156 -3452
rect 22463 -3800 22785 -3799
rect 22463 -4120 22464 -3800
rect 22784 -4120 22785 -3800
rect 22463 -4121 22785 -4120
rect 22040 -4468 22144 -4172
rect 21451 -4520 21773 -4519
rect 21451 -4840 21452 -4520
rect 21772 -4840 21773 -4520
rect 21451 -4841 21773 -4840
rect 21028 -5188 21132 -4892
rect 20439 -5240 20761 -5239
rect 20439 -5560 20440 -5240
rect 20760 -5560 20761 -5240
rect 20439 -5561 20761 -5560
rect 20016 -5760 20120 -5612
rect 20548 -5760 20652 -5561
rect 21028 -5612 21048 -5188
rect 21112 -5612 21132 -5188
rect 21560 -5239 21664 -4841
rect 22040 -4892 22060 -4468
rect 22124 -4892 22144 -4468
rect 22572 -4519 22676 -4121
rect 23052 -4172 23072 -3748
rect 23136 -4172 23156 -3748
rect 23584 -3799 23688 -3401
rect 24064 -3452 24084 -3028
rect 24148 -3452 24168 -3028
rect 24596 -3079 24700 -2681
rect 25076 -2732 25096 -2308
rect 25160 -2732 25180 -2308
rect 25608 -2359 25712 -1961
rect 26088 -2012 26108 -1588
rect 26172 -2012 26192 -1588
rect 26620 -1639 26724 -1241
rect 27100 -1292 27120 -868
rect 27184 -1292 27204 -868
rect 27632 -919 27736 -521
rect 28112 -572 28132 -148
rect 28196 -572 28216 -148
rect 28644 -199 28748 199
rect 29124 148 29144 572
rect 29208 148 29228 572
rect 29656 521 29760 919
rect 30136 868 30156 1292
rect 30220 868 30240 1292
rect 30668 1241 30772 1639
rect 31148 1588 31168 2012
rect 31232 1588 31252 2012
rect 31680 1961 31784 2359
rect 32160 2308 32180 2732
rect 32244 2308 32264 2732
rect 32160 2012 32264 2308
rect 31571 1960 31893 1961
rect 31571 1640 31572 1960
rect 31892 1640 31893 1960
rect 31571 1639 31893 1640
rect 31148 1292 31252 1588
rect 30559 1240 30881 1241
rect 30559 920 30560 1240
rect 30880 920 30881 1240
rect 30559 919 30881 920
rect 30136 572 30240 868
rect 29547 520 29869 521
rect 29547 200 29548 520
rect 29868 200 29869 520
rect 29547 199 29869 200
rect 29124 -148 29228 148
rect 28535 -200 28857 -199
rect 28535 -520 28536 -200
rect 28856 -520 28857 -200
rect 28535 -521 28857 -520
rect 28112 -868 28216 -572
rect 27523 -920 27845 -919
rect 27523 -1240 27524 -920
rect 27844 -1240 27845 -920
rect 27523 -1241 27845 -1240
rect 27100 -1588 27204 -1292
rect 26511 -1640 26833 -1639
rect 26511 -1960 26512 -1640
rect 26832 -1960 26833 -1640
rect 26511 -1961 26833 -1960
rect 26088 -2308 26192 -2012
rect 25499 -2360 25821 -2359
rect 25499 -2680 25500 -2360
rect 25820 -2680 25821 -2360
rect 25499 -2681 25821 -2680
rect 25076 -3028 25180 -2732
rect 24487 -3080 24809 -3079
rect 24487 -3400 24488 -3080
rect 24808 -3400 24809 -3080
rect 24487 -3401 24809 -3400
rect 24064 -3748 24168 -3452
rect 23475 -3800 23797 -3799
rect 23475 -4120 23476 -3800
rect 23796 -4120 23797 -3800
rect 23475 -4121 23797 -4120
rect 23052 -4468 23156 -4172
rect 22463 -4520 22785 -4519
rect 22463 -4840 22464 -4520
rect 22784 -4840 22785 -4520
rect 22463 -4841 22785 -4840
rect 22040 -5188 22144 -4892
rect 21451 -5240 21773 -5239
rect 21451 -5560 21452 -5240
rect 21772 -5560 21773 -5240
rect 21451 -5561 21773 -5560
rect 21028 -5760 21132 -5612
rect 21560 -5760 21664 -5561
rect 22040 -5612 22060 -5188
rect 22124 -5612 22144 -5188
rect 22572 -5239 22676 -4841
rect 23052 -4892 23072 -4468
rect 23136 -4892 23156 -4468
rect 23584 -4519 23688 -4121
rect 24064 -4172 24084 -3748
rect 24148 -4172 24168 -3748
rect 24596 -3799 24700 -3401
rect 25076 -3452 25096 -3028
rect 25160 -3452 25180 -3028
rect 25608 -3079 25712 -2681
rect 26088 -2732 26108 -2308
rect 26172 -2732 26192 -2308
rect 26620 -2359 26724 -1961
rect 27100 -2012 27120 -1588
rect 27184 -2012 27204 -1588
rect 27632 -1639 27736 -1241
rect 28112 -1292 28132 -868
rect 28196 -1292 28216 -868
rect 28644 -919 28748 -521
rect 29124 -572 29144 -148
rect 29208 -572 29228 -148
rect 29656 -199 29760 199
rect 30136 148 30156 572
rect 30220 148 30240 572
rect 30668 521 30772 919
rect 31148 868 31168 1292
rect 31232 868 31252 1292
rect 31680 1241 31784 1639
rect 32160 1588 32180 2012
rect 32244 1588 32264 2012
rect 32160 1292 32264 1588
rect 31571 1240 31893 1241
rect 31571 920 31572 1240
rect 31892 920 31893 1240
rect 31571 919 31893 920
rect 31148 572 31252 868
rect 30559 520 30881 521
rect 30559 200 30560 520
rect 30880 200 30881 520
rect 30559 199 30881 200
rect 30136 -148 30240 148
rect 29547 -200 29869 -199
rect 29547 -520 29548 -200
rect 29868 -520 29869 -200
rect 29547 -521 29869 -520
rect 29124 -868 29228 -572
rect 28535 -920 28857 -919
rect 28535 -1240 28536 -920
rect 28856 -1240 28857 -920
rect 28535 -1241 28857 -1240
rect 28112 -1588 28216 -1292
rect 27523 -1640 27845 -1639
rect 27523 -1960 27524 -1640
rect 27844 -1960 27845 -1640
rect 27523 -1961 27845 -1960
rect 27100 -2308 27204 -2012
rect 26511 -2360 26833 -2359
rect 26511 -2680 26512 -2360
rect 26832 -2680 26833 -2360
rect 26511 -2681 26833 -2680
rect 26088 -3028 26192 -2732
rect 25499 -3080 25821 -3079
rect 25499 -3400 25500 -3080
rect 25820 -3400 25821 -3080
rect 25499 -3401 25821 -3400
rect 25076 -3748 25180 -3452
rect 24487 -3800 24809 -3799
rect 24487 -4120 24488 -3800
rect 24808 -4120 24809 -3800
rect 24487 -4121 24809 -4120
rect 24064 -4468 24168 -4172
rect 23475 -4520 23797 -4519
rect 23475 -4840 23476 -4520
rect 23796 -4840 23797 -4520
rect 23475 -4841 23797 -4840
rect 23052 -5188 23156 -4892
rect 22463 -5240 22785 -5239
rect 22463 -5560 22464 -5240
rect 22784 -5560 22785 -5240
rect 22463 -5561 22785 -5560
rect 22040 -5760 22144 -5612
rect 22572 -5760 22676 -5561
rect 23052 -5612 23072 -5188
rect 23136 -5612 23156 -5188
rect 23584 -5239 23688 -4841
rect 24064 -4892 24084 -4468
rect 24148 -4892 24168 -4468
rect 24596 -4519 24700 -4121
rect 25076 -4172 25096 -3748
rect 25160 -4172 25180 -3748
rect 25608 -3799 25712 -3401
rect 26088 -3452 26108 -3028
rect 26172 -3452 26192 -3028
rect 26620 -3079 26724 -2681
rect 27100 -2732 27120 -2308
rect 27184 -2732 27204 -2308
rect 27632 -2359 27736 -1961
rect 28112 -2012 28132 -1588
rect 28196 -2012 28216 -1588
rect 28644 -1639 28748 -1241
rect 29124 -1292 29144 -868
rect 29208 -1292 29228 -868
rect 29656 -919 29760 -521
rect 30136 -572 30156 -148
rect 30220 -572 30240 -148
rect 30668 -199 30772 199
rect 31148 148 31168 572
rect 31232 148 31252 572
rect 31680 521 31784 919
rect 32160 868 32180 1292
rect 32244 868 32264 1292
rect 32160 572 32264 868
rect 31571 520 31893 521
rect 31571 200 31572 520
rect 31892 200 31893 520
rect 31571 199 31893 200
rect 31148 -148 31252 148
rect 30559 -200 30881 -199
rect 30559 -520 30560 -200
rect 30880 -520 30881 -200
rect 30559 -521 30881 -520
rect 30136 -868 30240 -572
rect 29547 -920 29869 -919
rect 29547 -1240 29548 -920
rect 29868 -1240 29869 -920
rect 29547 -1241 29869 -1240
rect 29124 -1588 29228 -1292
rect 28535 -1640 28857 -1639
rect 28535 -1960 28536 -1640
rect 28856 -1960 28857 -1640
rect 28535 -1961 28857 -1960
rect 28112 -2308 28216 -2012
rect 27523 -2360 27845 -2359
rect 27523 -2680 27524 -2360
rect 27844 -2680 27845 -2360
rect 27523 -2681 27845 -2680
rect 27100 -3028 27204 -2732
rect 26511 -3080 26833 -3079
rect 26511 -3400 26512 -3080
rect 26832 -3400 26833 -3080
rect 26511 -3401 26833 -3400
rect 26088 -3748 26192 -3452
rect 25499 -3800 25821 -3799
rect 25499 -4120 25500 -3800
rect 25820 -4120 25821 -3800
rect 25499 -4121 25821 -4120
rect 25076 -4468 25180 -4172
rect 24487 -4520 24809 -4519
rect 24487 -4840 24488 -4520
rect 24808 -4840 24809 -4520
rect 24487 -4841 24809 -4840
rect 24064 -5188 24168 -4892
rect 23475 -5240 23797 -5239
rect 23475 -5560 23476 -5240
rect 23796 -5560 23797 -5240
rect 23475 -5561 23797 -5560
rect 23052 -5760 23156 -5612
rect 23584 -5760 23688 -5561
rect 24064 -5612 24084 -5188
rect 24148 -5612 24168 -5188
rect 24596 -5239 24700 -4841
rect 25076 -4892 25096 -4468
rect 25160 -4892 25180 -4468
rect 25608 -4519 25712 -4121
rect 26088 -4172 26108 -3748
rect 26172 -4172 26192 -3748
rect 26620 -3799 26724 -3401
rect 27100 -3452 27120 -3028
rect 27184 -3452 27204 -3028
rect 27632 -3079 27736 -2681
rect 28112 -2732 28132 -2308
rect 28196 -2732 28216 -2308
rect 28644 -2359 28748 -1961
rect 29124 -2012 29144 -1588
rect 29208 -2012 29228 -1588
rect 29656 -1639 29760 -1241
rect 30136 -1292 30156 -868
rect 30220 -1292 30240 -868
rect 30668 -919 30772 -521
rect 31148 -572 31168 -148
rect 31232 -572 31252 -148
rect 31680 -199 31784 199
rect 32160 148 32180 572
rect 32244 148 32264 572
rect 32160 -148 32264 148
rect 31571 -200 31893 -199
rect 31571 -520 31572 -200
rect 31892 -520 31893 -200
rect 31571 -521 31893 -520
rect 31148 -868 31252 -572
rect 30559 -920 30881 -919
rect 30559 -1240 30560 -920
rect 30880 -1240 30881 -920
rect 30559 -1241 30881 -1240
rect 30136 -1588 30240 -1292
rect 29547 -1640 29869 -1639
rect 29547 -1960 29548 -1640
rect 29868 -1960 29869 -1640
rect 29547 -1961 29869 -1960
rect 29124 -2308 29228 -2012
rect 28535 -2360 28857 -2359
rect 28535 -2680 28536 -2360
rect 28856 -2680 28857 -2360
rect 28535 -2681 28857 -2680
rect 28112 -3028 28216 -2732
rect 27523 -3080 27845 -3079
rect 27523 -3400 27524 -3080
rect 27844 -3400 27845 -3080
rect 27523 -3401 27845 -3400
rect 27100 -3748 27204 -3452
rect 26511 -3800 26833 -3799
rect 26511 -4120 26512 -3800
rect 26832 -4120 26833 -3800
rect 26511 -4121 26833 -4120
rect 26088 -4468 26192 -4172
rect 25499 -4520 25821 -4519
rect 25499 -4840 25500 -4520
rect 25820 -4840 25821 -4520
rect 25499 -4841 25821 -4840
rect 25076 -5188 25180 -4892
rect 24487 -5240 24809 -5239
rect 24487 -5560 24488 -5240
rect 24808 -5560 24809 -5240
rect 24487 -5561 24809 -5560
rect 24064 -5760 24168 -5612
rect 24596 -5760 24700 -5561
rect 25076 -5612 25096 -5188
rect 25160 -5612 25180 -5188
rect 25608 -5239 25712 -4841
rect 26088 -4892 26108 -4468
rect 26172 -4892 26192 -4468
rect 26620 -4519 26724 -4121
rect 27100 -4172 27120 -3748
rect 27184 -4172 27204 -3748
rect 27632 -3799 27736 -3401
rect 28112 -3452 28132 -3028
rect 28196 -3452 28216 -3028
rect 28644 -3079 28748 -2681
rect 29124 -2732 29144 -2308
rect 29208 -2732 29228 -2308
rect 29656 -2359 29760 -1961
rect 30136 -2012 30156 -1588
rect 30220 -2012 30240 -1588
rect 30668 -1639 30772 -1241
rect 31148 -1292 31168 -868
rect 31232 -1292 31252 -868
rect 31680 -919 31784 -521
rect 32160 -572 32180 -148
rect 32244 -572 32264 -148
rect 32160 -868 32264 -572
rect 31571 -920 31893 -919
rect 31571 -1240 31572 -920
rect 31892 -1240 31893 -920
rect 31571 -1241 31893 -1240
rect 31148 -1588 31252 -1292
rect 30559 -1640 30881 -1639
rect 30559 -1960 30560 -1640
rect 30880 -1960 30881 -1640
rect 30559 -1961 30881 -1960
rect 30136 -2308 30240 -2012
rect 29547 -2360 29869 -2359
rect 29547 -2680 29548 -2360
rect 29868 -2680 29869 -2360
rect 29547 -2681 29869 -2680
rect 29124 -3028 29228 -2732
rect 28535 -3080 28857 -3079
rect 28535 -3400 28536 -3080
rect 28856 -3400 28857 -3080
rect 28535 -3401 28857 -3400
rect 28112 -3748 28216 -3452
rect 27523 -3800 27845 -3799
rect 27523 -4120 27524 -3800
rect 27844 -4120 27845 -3800
rect 27523 -4121 27845 -4120
rect 27100 -4468 27204 -4172
rect 26511 -4520 26833 -4519
rect 26511 -4840 26512 -4520
rect 26832 -4840 26833 -4520
rect 26511 -4841 26833 -4840
rect 26088 -5188 26192 -4892
rect 25499 -5240 25821 -5239
rect 25499 -5560 25500 -5240
rect 25820 -5560 25821 -5240
rect 25499 -5561 25821 -5560
rect 25076 -5760 25180 -5612
rect 25608 -5760 25712 -5561
rect 26088 -5612 26108 -5188
rect 26172 -5612 26192 -5188
rect 26620 -5239 26724 -4841
rect 27100 -4892 27120 -4468
rect 27184 -4892 27204 -4468
rect 27632 -4519 27736 -4121
rect 28112 -4172 28132 -3748
rect 28196 -4172 28216 -3748
rect 28644 -3799 28748 -3401
rect 29124 -3452 29144 -3028
rect 29208 -3452 29228 -3028
rect 29656 -3079 29760 -2681
rect 30136 -2732 30156 -2308
rect 30220 -2732 30240 -2308
rect 30668 -2359 30772 -1961
rect 31148 -2012 31168 -1588
rect 31232 -2012 31252 -1588
rect 31680 -1639 31784 -1241
rect 32160 -1292 32180 -868
rect 32244 -1292 32264 -868
rect 32160 -1588 32264 -1292
rect 31571 -1640 31893 -1639
rect 31571 -1960 31572 -1640
rect 31892 -1960 31893 -1640
rect 31571 -1961 31893 -1960
rect 31148 -2308 31252 -2012
rect 30559 -2360 30881 -2359
rect 30559 -2680 30560 -2360
rect 30880 -2680 30881 -2360
rect 30559 -2681 30881 -2680
rect 30136 -3028 30240 -2732
rect 29547 -3080 29869 -3079
rect 29547 -3400 29548 -3080
rect 29868 -3400 29869 -3080
rect 29547 -3401 29869 -3400
rect 29124 -3748 29228 -3452
rect 28535 -3800 28857 -3799
rect 28535 -4120 28536 -3800
rect 28856 -4120 28857 -3800
rect 28535 -4121 28857 -4120
rect 28112 -4468 28216 -4172
rect 27523 -4520 27845 -4519
rect 27523 -4840 27524 -4520
rect 27844 -4840 27845 -4520
rect 27523 -4841 27845 -4840
rect 27100 -5188 27204 -4892
rect 26511 -5240 26833 -5239
rect 26511 -5560 26512 -5240
rect 26832 -5560 26833 -5240
rect 26511 -5561 26833 -5560
rect 26088 -5760 26192 -5612
rect 26620 -5760 26724 -5561
rect 27100 -5612 27120 -5188
rect 27184 -5612 27204 -5188
rect 27632 -5239 27736 -4841
rect 28112 -4892 28132 -4468
rect 28196 -4892 28216 -4468
rect 28644 -4519 28748 -4121
rect 29124 -4172 29144 -3748
rect 29208 -4172 29228 -3748
rect 29656 -3799 29760 -3401
rect 30136 -3452 30156 -3028
rect 30220 -3452 30240 -3028
rect 30668 -3079 30772 -2681
rect 31148 -2732 31168 -2308
rect 31232 -2732 31252 -2308
rect 31680 -2359 31784 -1961
rect 32160 -2012 32180 -1588
rect 32244 -2012 32264 -1588
rect 32160 -2308 32264 -2012
rect 31571 -2360 31893 -2359
rect 31571 -2680 31572 -2360
rect 31892 -2680 31893 -2360
rect 31571 -2681 31893 -2680
rect 31148 -3028 31252 -2732
rect 30559 -3080 30881 -3079
rect 30559 -3400 30560 -3080
rect 30880 -3400 30881 -3080
rect 30559 -3401 30881 -3400
rect 30136 -3748 30240 -3452
rect 29547 -3800 29869 -3799
rect 29547 -4120 29548 -3800
rect 29868 -4120 29869 -3800
rect 29547 -4121 29869 -4120
rect 29124 -4468 29228 -4172
rect 28535 -4520 28857 -4519
rect 28535 -4840 28536 -4520
rect 28856 -4840 28857 -4520
rect 28535 -4841 28857 -4840
rect 28112 -5188 28216 -4892
rect 27523 -5240 27845 -5239
rect 27523 -5560 27524 -5240
rect 27844 -5560 27845 -5240
rect 27523 -5561 27845 -5560
rect 27100 -5760 27204 -5612
rect 27632 -5760 27736 -5561
rect 28112 -5612 28132 -5188
rect 28196 -5612 28216 -5188
rect 28644 -5239 28748 -4841
rect 29124 -4892 29144 -4468
rect 29208 -4892 29228 -4468
rect 29656 -4519 29760 -4121
rect 30136 -4172 30156 -3748
rect 30220 -4172 30240 -3748
rect 30668 -3799 30772 -3401
rect 31148 -3452 31168 -3028
rect 31232 -3452 31252 -3028
rect 31680 -3079 31784 -2681
rect 32160 -2732 32180 -2308
rect 32244 -2732 32264 -2308
rect 32160 -3028 32264 -2732
rect 31571 -3080 31893 -3079
rect 31571 -3400 31572 -3080
rect 31892 -3400 31893 -3080
rect 31571 -3401 31893 -3400
rect 31148 -3748 31252 -3452
rect 30559 -3800 30881 -3799
rect 30559 -4120 30560 -3800
rect 30880 -4120 30881 -3800
rect 30559 -4121 30881 -4120
rect 30136 -4468 30240 -4172
rect 29547 -4520 29869 -4519
rect 29547 -4840 29548 -4520
rect 29868 -4840 29869 -4520
rect 29547 -4841 29869 -4840
rect 29124 -5188 29228 -4892
rect 28535 -5240 28857 -5239
rect 28535 -5560 28536 -5240
rect 28856 -5560 28857 -5240
rect 28535 -5561 28857 -5560
rect 28112 -5760 28216 -5612
rect 28644 -5760 28748 -5561
rect 29124 -5612 29144 -5188
rect 29208 -5612 29228 -5188
rect 29656 -5239 29760 -4841
rect 30136 -4892 30156 -4468
rect 30220 -4892 30240 -4468
rect 30668 -4519 30772 -4121
rect 31148 -4172 31168 -3748
rect 31232 -4172 31252 -3748
rect 31680 -3799 31784 -3401
rect 32160 -3452 32180 -3028
rect 32244 -3452 32264 -3028
rect 32160 -3748 32264 -3452
rect 31571 -3800 31893 -3799
rect 31571 -4120 31572 -3800
rect 31892 -4120 31893 -3800
rect 31571 -4121 31893 -4120
rect 31148 -4468 31252 -4172
rect 30559 -4520 30881 -4519
rect 30559 -4840 30560 -4520
rect 30880 -4840 30881 -4520
rect 30559 -4841 30881 -4840
rect 30136 -5188 30240 -4892
rect 29547 -5240 29869 -5239
rect 29547 -5560 29548 -5240
rect 29868 -5560 29869 -5240
rect 29547 -5561 29869 -5560
rect 29124 -5760 29228 -5612
rect 29656 -5760 29760 -5561
rect 30136 -5612 30156 -5188
rect 30220 -5612 30240 -5188
rect 30668 -5239 30772 -4841
rect 31148 -4892 31168 -4468
rect 31232 -4892 31252 -4468
rect 31680 -4519 31784 -4121
rect 32160 -4172 32180 -3748
rect 32244 -4172 32264 -3748
rect 32160 -4468 32264 -4172
rect 31571 -4520 31893 -4519
rect 31571 -4840 31572 -4520
rect 31892 -4840 31893 -4520
rect 31571 -4841 31893 -4840
rect 31148 -5188 31252 -4892
rect 30559 -5240 30881 -5239
rect 30559 -5560 30560 -5240
rect 30880 -5560 30881 -5240
rect 30559 -5561 30881 -5560
rect 30136 -5760 30240 -5612
rect 30668 -5760 30772 -5561
rect 31148 -5612 31168 -5188
rect 31232 -5612 31252 -5188
rect 31680 -5239 31784 -4841
rect 32160 -4892 32180 -4468
rect 32244 -4892 32264 -4468
rect 32160 -5188 32264 -4892
rect 31571 -5240 31893 -5239
rect 31571 -5560 31572 -5240
rect 31892 -5560 31893 -5240
rect 31571 -5561 31893 -5560
rect 31148 -5760 31252 -5612
rect 31680 -5760 31784 -5561
rect 32160 -5612 32180 -5188
rect 32244 -5612 32264 -5188
rect 32160 -5760 32264 -5612
<< properties >>
string FIXED_BBOX 31492 5160 31972 5640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 64 ny 16 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
