magic
tech sky130A
magscale 1 2
timestamp 1757893939
<< metal1 >>
rect 1421 2274 3012 2574
rect 4372 2264 4672 2564
rect -519 336 -269 360
rect -519 284 -355 336
rect -303 284 -269 336
rect -519 260 -269 284
rect -519 136 -69 160
rect -519 84 -155 136
rect -103 84 -69 136
rect -519 60 -69 84
rect 2978 -2538 4718 -2238
rect -519 -4466 -269 -4442
rect -519 -4518 -355 -4466
rect -303 -4518 -269 -4466
rect -519 -4542 -269 -4518
rect -519 -4666 -69 -4642
rect -519 -4718 -155 -4666
rect -103 -4718 -69 -4666
rect -519 -4742 -69 -4718
rect 1421 -7330 4718 -7030
rect -519 -9268 -273 -9244
rect -519 -9320 -359 -9268
rect -307 -9320 -273 -9268
rect -519 -9344 -273 -9320
rect -519 -9468 -69 -9444
rect -519 -9520 -155 -9468
rect -103 -9520 -69 -9468
rect -519 -9544 -69 -9520
rect 1421 -12132 3012 -11832
rect 4340 -12141 4640 -11841
rect -519 -14070 -269 -14046
rect -519 -14122 -355 -14070
rect -303 -14122 -269 -14070
rect -519 -14146 -269 -14122
rect -189 -14246 -69 -14245
rect -519 -14269 -69 -14246
rect -519 -14321 -155 -14269
rect -103 -14321 -69 -14269
rect -519 -14345 -69 -14321
rect -519 -14346 -79 -14345
rect 1421 -16934 3012 -16634
rect 4262 -16944 4562 -16644
rect -519 -18872 -269 -18848
rect -519 -18924 -355 -18872
rect -303 -18924 -269 -18872
rect -519 -18948 -269 -18924
rect -519 -19072 -69 -19048
rect -519 -19124 -155 -19072
rect -103 -19124 -69 -19072
rect -519 -19148 -69 -19124
rect 1631 -21736 3012 -21436
rect 4262 -21746 4562 -21446
rect -519 -23674 -269 -23650
rect -519 -23726 -355 -23674
rect -303 -23726 -269 -23674
rect -519 -23750 -269 -23726
rect -519 -23874 -69 -23850
rect -519 -23926 -155 -23874
rect -103 -23926 -69 -23874
rect -519 -23950 -69 -23926
rect 4214 -26548 4514 -26248
rect -519 -28453 -279 -28452
rect -519 -28477 -269 -28453
rect -519 -28529 -355 -28477
rect -303 -28529 -269 -28477
rect -519 -28552 -269 -28529
rect -389 -28553 -269 -28552
rect -519 -28676 -69 -28652
rect -519 -28728 -155 -28676
rect -103 -28728 -69 -28676
rect -519 -28752 -69 -28728
rect 1421 -31340 3012 -31040
rect 4218 -31350 4518 -31050
rect -519 -33278 -269 -33254
rect -519 -33330 -355 -33278
rect -303 -33330 -269 -33278
rect -519 -33354 -269 -33330
rect -519 -33478 -69 -33454
rect -519 -33530 -155 -33478
rect -103 -33530 -69 -33478
rect -519 -33554 -69 -33530
rect 2978 -36142 3012 -35842
rect 4232 -36152 4532 -35852
rect -519 -38080 -269 -38056
rect -519 -38132 -355 -38080
rect -303 -38132 -269 -38080
rect -519 -38156 -269 -38132
rect -519 -38280 -69 -38256
rect -519 -38332 -155 -38280
rect -103 -38332 -69 -38280
rect -519 -38356 -69 -38332
<< via1 >>
rect -355 284 -303 336
rect -155 84 -103 136
rect -355 -4518 -303 -4466
rect -155 -4718 -103 -4666
rect -359 -9320 -307 -9268
rect -155 -9520 -103 -9468
rect -355 -14122 -303 -14070
rect -155 -14321 -103 -14269
rect -355 -18924 -303 -18872
rect -155 -19124 -103 -19072
rect -355 -23726 -303 -23674
rect -155 -23926 -103 -23874
rect -355 -28529 -303 -28477
rect -155 -28728 -103 -28676
rect -355 -33330 -303 -33278
rect -155 -33530 -103 -33478
rect -355 -38132 -303 -38080
rect -155 -38332 -103 -38280
<< metal2 >>
rect -379 336 -279 370
rect -379 284 -355 336
rect -303 284 -279 336
rect -379 250 -279 284
rect -179 136 -79 170
rect -179 84 -155 136
rect -103 84 -79 136
rect -179 50 -79 84
rect -379 -4466 -279 -4432
rect -379 -4518 -355 -4466
rect -303 -4518 -279 -4466
rect -379 -4552 -279 -4518
rect -179 -4666 -79 -4632
rect -179 -4718 -155 -4666
rect -103 -4718 -79 -4666
rect -179 -4752 -79 -4718
rect -383 -9268 -283 -9234
rect -383 -9320 -359 -9268
rect -307 -9320 -283 -9268
rect -383 -9354 -283 -9320
rect -179 -9468 -79 -9434
rect -179 -9520 -155 -9468
rect -103 -9520 -79 -9468
rect -179 -9554 -79 -9520
rect -379 -14070 -279 -14036
rect -379 -14122 -355 -14070
rect -303 -14122 -279 -14070
rect -379 -14156 -279 -14122
rect -179 -14269 -79 -14235
rect -179 -14321 -155 -14269
rect -103 -14321 -79 -14269
rect -179 -14355 -79 -14321
rect -379 -18872 -279 -18835
rect -379 -18924 -355 -18872
rect -303 -18924 -279 -18872
rect -379 -18958 -279 -18924
rect -179 -19072 -79 -19038
rect -179 -19124 -155 -19072
rect -103 -19124 -79 -19072
rect -179 -19158 -79 -19124
rect -379 -23674 -279 -23640
rect -379 -23726 -355 -23674
rect -303 -23726 -279 -23674
rect -379 -23760 -279 -23726
rect -179 -23874 -79 -23840
rect -179 -23926 -155 -23874
rect -103 -23926 -79 -23874
rect -179 -23960 -79 -23926
rect -379 -28477 -279 -28443
rect -379 -28529 -355 -28477
rect -303 -28529 -279 -28477
rect -379 -28563 -279 -28529
rect -179 -28676 -79 -28642
rect -179 -28728 -155 -28676
rect -103 -28728 -79 -28676
rect -179 -28762 -79 -28728
rect -379 -33278 -279 -33244
rect -379 -33330 -355 -33278
rect -303 -33330 -279 -33278
rect -379 -33364 -279 -33330
rect -179 -33478 -79 -33444
rect -179 -33530 -155 -33478
rect -103 -33530 -79 -33478
rect -179 -33564 -79 -33530
rect -379 -38080 -279 -38046
rect -379 -38132 -355 -38080
rect -303 -38132 -279 -38080
rect -379 -38166 -279 -38132
rect -179 -38280 -79 -38246
rect 21 -38269 121 4462
rect 1021 -38269 1121 4728
rect 1221 -38269 1321 4634
rect -179 -38332 -155 -38280
rect -103 -38332 -79 -38280
rect -179 -38366 -79 -38332
use cdac_sw_3  cdac_sw_3_0
timestamp 1757893939
transform 1 0 1439 0 1 -6272
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_1
timestamp 1757893939
transform 1 0 1439 0 1 -1480
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_2
timestamp 1757893939
transform 1 0 1439 0 1 3322
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_3
timestamp 1757893939
transform 1 0 1439 0 1 -15886
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_4
timestamp 1757893939
transform 1 0 1439 0 1 -11083
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_5
timestamp 1757893939
transform 1 0 1439 0 1 -20688
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_6
timestamp 1757893939
transform 1 0 1439 0 1 -25490
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_7
timestamp 1757893939
transform 1 0 1439 0 1 -30292
box -1828 -3272 3610 1410
use cdac_sw_3  cdac_sw_3_8
timestamp 1757893939
transform 1 0 1439 0 1 -35094
box -1828 -3272 3610 1410
<< labels >>
flabel metal2 s 1052 4651 1092 4691 0 FreeSans 1000 0 0 0 VDD
port 1 nsew
flabel metal2 s 1249 4437 1289 4477 0 FreeSans 1000 0 0 0 VSS
port 2 nsew
flabel metal2 s 55 4351 95 4391 0 FreeSans 1000 0 0 0 VCM
port 3 nsew
flabel metal1 s -501 281 -461 321 0 FreeSans 1000 0 0 0 SW_IN[0]
port 4 nsew
flabel metal1 s -492 -4511 -452 -4471 0 FreeSans 1000 0 0 0 SW_IN[1]
port 5 nsew
flabel metal1 s -503 -9309 -463 -9269 0 FreeSans 1000 0 0 0 SW_IN[2]
port 6 nsew
flabel metal1 s -499 -14115 -459 -14075 0 FreeSans 1000 0 0 0 SW_IN[3]
port 7 nsew
flabel metal1 s -503 -18914 -463 -18874 0 FreeSans 1000 0 0 0 SW_IN[4]
port 8 nsew
flabel metal1 s -498 -23716 -458 -23676 0 FreeSans 1000 0 0 0 SW_IN[5]
port 9 nsew
flabel metal1 s -500 -28521 -460 -28481 0 FreeSans 1000 0 0 0 SW_IN[6]
port 10 nsew
flabel metal1 s -497 -33321 -457 -33281 0 FreeSans 1000 0 0 0 SW_IN[7]
port 11 nsew
flabel metal1 s -496 -38127 -456 -38087 0 FreeSans 1000 0 0 0 SW_IN[8]
port 12 nsew
flabel metal1 s -496 88 -456 128 0 FreeSans 1000 0 0 0 CF[0]
port 14 nsew
flabel metal1 s -497 -4710 -457 -4670 0 FreeSans 1000 0 0 0 CF[1]
port 15 nsew
flabel metal1 s -500 -9513 -460 -9473 0 FreeSans 1000 0 0 0 CF[2]
port 16 nsew
flabel metal1 s -490 -14319 -450 -14279 0 FreeSans 1000 0 0 0 CF[3]
port 17 nsew
flabel metal1 s -497 -19117 -457 -19077 0 FreeSans 1000 0 0 0 CF[4]
port 18 nsew
flabel metal1 s -495 -23917 -455 -23877 0 FreeSans 1000 0 0 0 CF[5]
port 19 nsew
flabel metal1 s -500 -28722 -460 -28682 0 FreeSans 1000 0 0 0 CF[6]
port 20 nsew
flabel metal1 s -497 -33525 -457 -33485 0 FreeSans 1000 0 0 0 CF[7]
port 21 nsew
flabel metal1 s -495 -38323 -455 -38283 0 FreeSans 1000 0 0 0 CF[8]
port 22 nsew
flabel metal1 4372 2264 4672 2564 0 FreeSans 1600 0 0 0 S[0]
port 24 nsew
flabel metal1 4320 -2538 4620 -2238 0 FreeSans 1600 0 0 0 S[1]
port 25 nsew
flabel metal1 4360 -7330 4660 -7030 0 FreeSans 1600 0 0 0 S[2]
port 26 nsew
flabel metal1 4340 -12141 4640 -11841 0 FreeSans 1600 0 0 0 S[3]
port 27 nsew
flabel metal1 4262 -16944 4562 -16644 0 FreeSans 1600 0 0 0 S[4]
port 28 nsew
flabel metal1 4262 -21746 4562 -21446 0 FreeSans 1600 0 0 0 S[5]
port 29 nsew
flabel metal1 4214 -26548 4514 -26248 0 FreeSans 1600 0 0 0 S[6]
port 30 nsew
flabel metal1 4218 -31350 4518 -31050 0 FreeSans 1600 0 0 0 S[7]
port 31 nsew
flabel metal1 4232 -36152 4532 -35852 0 FreeSans 1600 0 0 0 S[8]
port 32 nsew
<< end >>
