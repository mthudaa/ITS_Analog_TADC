magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< error_p >>
rect -29 441 29 447
rect -29 407 -17 441
rect -29 401 29 407
<< pwell >>
rect -201 -569 201 569
<< nmos >>
rect -15 -431 15 369
<< ndiff >>
rect -73 326 -15 369
rect -73 292 -61 326
rect -27 292 -15 326
rect -73 258 -15 292
rect -73 224 -61 258
rect -27 224 -15 258
rect -73 190 -15 224
rect -73 156 -61 190
rect -27 156 -15 190
rect -73 122 -15 156
rect -73 88 -61 122
rect -27 88 -15 122
rect -73 54 -15 88
rect -73 20 -61 54
rect -27 20 -15 54
rect -73 -14 -15 20
rect -73 -48 -61 -14
rect -27 -48 -15 -14
rect -73 -82 -15 -48
rect -73 -116 -61 -82
rect -27 -116 -15 -82
rect -73 -150 -15 -116
rect -73 -184 -61 -150
rect -27 -184 -15 -150
rect -73 -218 -15 -184
rect -73 -252 -61 -218
rect -27 -252 -15 -218
rect -73 -286 -15 -252
rect -73 -320 -61 -286
rect -27 -320 -15 -286
rect -73 -354 -15 -320
rect -73 -388 -61 -354
rect -27 -388 -15 -354
rect -73 -431 -15 -388
rect 15 326 73 369
rect 15 292 27 326
rect 61 292 73 326
rect 15 258 73 292
rect 15 224 27 258
rect 61 224 73 258
rect 15 190 73 224
rect 15 156 27 190
rect 61 156 73 190
rect 15 122 73 156
rect 15 88 27 122
rect 61 88 73 122
rect 15 54 73 88
rect 15 20 27 54
rect 61 20 73 54
rect 15 -14 73 20
rect 15 -48 27 -14
rect 61 -48 73 -14
rect 15 -82 73 -48
rect 15 -116 27 -82
rect 61 -116 73 -82
rect 15 -150 73 -116
rect 15 -184 27 -150
rect 61 -184 73 -150
rect 15 -218 73 -184
rect 15 -252 27 -218
rect 61 -252 73 -218
rect 15 -286 73 -252
rect 15 -320 27 -286
rect 61 -320 73 -286
rect 15 -354 73 -320
rect 15 -388 27 -354
rect 61 -388 73 -354
rect 15 -431 73 -388
<< ndiffc >>
rect -61 292 -27 326
rect -61 224 -27 258
rect -61 156 -27 190
rect -61 88 -27 122
rect -61 20 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -82
rect -61 -184 -27 -150
rect -61 -252 -27 -218
rect -61 -320 -27 -286
rect -61 -388 -27 -354
rect 27 292 61 326
rect 27 224 61 258
rect 27 156 61 190
rect 27 88 61 122
rect 27 20 61 54
rect 27 -48 61 -14
rect 27 -116 61 -82
rect 27 -184 61 -150
rect 27 -252 61 -218
rect 27 -320 61 -286
rect 27 -388 61 -354
<< psubdiff >>
rect -175 509 -51 543
rect -17 509 17 543
rect 51 509 175 543
rect -175 -509 -141 509
rect 141 425 175 509
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -509 175 -425
rect -175 -543 -51 -509
rect -17 -543 17 -509
rect 51 -543 175 -509
<< psubdiffcont >>
rect -51 509 -17 543
rect 17 509 51 543
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect -51 -543 -17 -509
rect 17 -543 51 -509
<< poly >>
rect -33 441 33 457
rect -33 407 -17 441
rect 17 407 33 441
rect -33 391 33 407
rect -15 369 15 391
rect -15 -457 15 -431
<< polycont >>
rect -17 407 17 441
<< locali >>
rect -175 509 -51 543
rect -17 509 17 543
rect 51 509 175 543
rect -175 -509 -141 509
rect -33 407 -17 441
rect 17 407 33 441
rect 141 425 175 509
rect -61 346 -27 373
rect -61 274 -27 292
rect -61 202 -27 224
rect -61 130 -27 156
rect -61 58 -27 88
rect -61 -14 -27 20
rect -61 -82 -27 -48
rect -61 -150 -27 -120
rect -61 -218 -27 -192
rect -61 -286 -27 -264
rect -61 -354 -27 -336
rect -61 -435 -27 -408
rect 27 346 61 373
rect 27 274 61 292
rect 27 202 61 224
rect 27 130 61 156
rect 27 58 61 88
rect 27 -14 61 20
rect 27 -82 61 -48
rect 27 -150 61 -120
rect 27 -218 61 -192
rect 27 -286 61 -264
rect 27 -354 61 -336
rect 27 -435 61 -408
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -509 175 -425
rect -175 -543 -51 -509
rect -17 -543 17 -509
rect 51 -543 175 -509
<< viali >>
rect -17 407 17 441
rect -61 326 -27 346
rect -61 312 -27 326
rect -61 258 -27 274
rect -61 240 -27 258
rect -61 190 -27 202
rect -61 168 -27 190
rect -61 122 -27 130
rect -61 96 -27 122
rect -61 54 -27 58
rect -61 24 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -86
rect -61 -120 -27 -116
rect -61 -184 -27 -158
rect -61 -192 -27 -184
rect -61 -252 -27 -230
rect -61 -264 -27 -252
rect -61 -320 -27 -302
rect -61 -336 -27 -320
rect -61 -388 -27 -374
rect -61 -408 -27 -388
rect 27 326 61 346
rect 27 312 61 326
rect 27 258 61 274
rect 27 240 61 258
rect 27 190 61 202
rect 27 168 61 190
rect 27 122 61 130
rect 27 96 61 122
rect 27 54 61 58
rect 27 24 61 54
rect 27 -48 61 -14
rect 27 -116 61 -86
rect 27 -120 61 -116
rect 27 -184 61 -158
rect 27 -192 61 -184
rect 27 -252 61 -230
rect 27 -264 61 -252
rect 27 -320 61 -302
rect 27 -336 61 -320
rect 27 -388 61 -374
rect 27 -408 61 -388
<< metal1 >>
rect -29 441 29 447
rect -29 407 -17 441
rect 17 407 29 441
rect -29 401 29 407
rect -67 346 -21 369
rect -67 312 -61 346
rect -27 312 -21 346
rect -67 274 -21 312
rect -67 240 -61 274
rect -27 240 -21 274
rect -67 202 -21 240
rect -67 168 -61 202
rect -27 168 -21 202
rect -67 130 -21 168
rect -67 96 -61 130
rect -27 96 -21 130
rect -67 58 -21 96
rect -67 24 -61 58
rect -27 24 -21 58
rect -67 -14 -21 24
rect -67 -48 -61 -14
rect -27 -48 -21 -14
rect -67 -86 -21 -48
rect -67 -120 -61 -86
rect -27 -120 -21 -86
rect -67 -158 -21 -120
rect -67 -192 -61 -158
rect -27 -192 -21 -158
rect -67 -230 -21 -192
rect -67 -264 -61 -230
rect -27 -264 -21 -230
rect -67 -302 -21 -264
rect -67 -336 -61 -302
rect -27 -336 -21 -302
rect -67 -374 -21 -336
rect -67 -408 -61 -374
rect -27 -408 -21 -374
rect -67 -431 -21 -408
rect 21 346 67 369
rect 21 312 27 346
rect 61 312 67 346
rect 21 274 67 312
rect 21 240 27 274
rect 61 240 67 274
rect 21 202 67 240
rect 21 168 27 202
rect 61 168 67 202
rect 21 130 67 168
rect 21 96 27 130
rect 61 96 67 130
rect 21 58 67 96
rect 21 24 27 58
rect 61 24 67 58
rect 21 -14 67 24
rect 21 -48 27 -14
rect 61 -48 67 -14
rect 21 -86 67 -48
rect 21 -120 27 -86
rect 61 -120 67 -86
rect 21 -158 67 -120
rect 21 -192 27 -158
rect 61 -192 67 -158
rect 21 -230 67 -192
rect 21 -264 27 -230
rect 61 -264 67 -230
rect 21 -302 67 -264
rect 21 -336 27 -302
rect 61 -336 67 -302
rect 21 -374 67 -336
rect 21 -408 27 -374
rect 61 -408 67 -374
rect 21 -431 67 -408
<< properties >>
string FIXED_BBOX -158 -526 158 526
<< end >>
