magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< pwell >>
rect -184 -126 184 126
<< nmos >>
rect -100 -100 100 100
<< ndiff >>
rect -158 85 -100 100
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -100 -100 -85
rect 100 85 158 100
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -100 158 -85
<< ndiffc >>
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
<< poly >>
rect -100 100 100 126
rect -100 -126 100 -100
<< locali >>
rect -146 85 -112 104
rect -146 17 -112 19
rect -146 -19 -112 -17
rect -146 -104 -112 -85
rect 112 85 146 104
rect 112 17 146 19
rect 112 -19 146 -17
rect 112 -104 146 -85
<< viali >>
rect -146 51 -112 53
rect -146 19 -112 51
rect -146 -51 -112 -19
rect -146 -53 -112 -51
rect 112 51 146 53
rect 112 19 146 51
rect 112 -51 146 -19
rect 112 -53 146 -51
<< metal1 >>
rect -152 53 -106 100
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -100 -106 -53
rect 106 53 152 100
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -100 152 -53
<< end >>
