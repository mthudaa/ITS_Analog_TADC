magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 9 403
rect 43 369 81 403
rect 115 369 153 403
rect 187 369 225 403
rect 259 369 297 403
rect 331 369 369 403
rect 403 369 441 403
rect 475 369 513 403
rect 547 369 585 403
rect 619 369 657 403
rect 691 369 729 403
rect 763 369 801 403
rect 835 369 873 403
rect 907 369 945 403
rect 979 369 1017 403
rect 1051 369 1077 403
rect 1149 -17 1173 17
rect 1207 -17 1245 17
rect 1279 -17 1317 17
rect 1351 -17 1389 17
rect 1423 -17 1461 17
rect 1495 -17 1533 17
rect 1567 -17 1605 17
rect 1639 -17 1677 17
rect 1711 -17 1749 17
rect 1783 -17 1807 17
<< viali >>
rect 9 369 43 403
rect 81 369 115 403
rect 153 369 187 403
rect 225 369 259 403
rect 297 369 331 403
rect 369 369 403 403
rect 441 369 475 403
rect 513 369 547 403
rect 585 369 619 403
rect 657 369 691 403
rect 729 369 763 403
rect 801 369 835 403
rect 873 369 907 403
rect 945 369 979 403
rect 1017 369 1051 403
rect 1173 -17 1207 17
rect 1245 -17 1279 17
rect 1317 -17 1351 17
rect 1389 -17 1423 17
rect 1461 -17 1495 17
rect 1533 -17 1567 17
rect 1605 -17 1639 17
rect 1677 -17 1711 17
rect 1749 -17 1783 17
<< metal1 >>
rect -53 403 1843 439
rect -53 369 9 403
rect 43 369 81 403
rect 115 369 153 403
rect 187 369 225 403
rect 259 369 297 403
rect 331 369 369 403
rect 403 369 441 403
rect 475 369 513 403
rect 547 369 585 403
rect 619 369 657 403
rect 691 369 729 403
rect 763 369 801 403
rect 835 369 873 403
rect 907 369 945 403
rect 979 369 1017 403
rect 1051 369 1843 403
rect -53 363 1843 369
rect -53 289 1633 323
rect -53 143 125 243
rect 1665 143 1843 243
rect 166 63 1843 97
rect -53 17 1843 23
rect -53 -17 1173 17
rect 1207 -17 1245 17
rect 1279 -17 1317 17
rect 1351 -17 1389 17
rect 1423 -17 1461 17
rect 1495 -17 1533 17
rect 1567 -17 1605 17
rect 1639 -17 1677 17
rect 1711 -17 1749 17
rect 1783 -17 1843 17
rect -53 -53 1843 -17
use sky130_fd_pr__pfet_01v8_SEQPU3  XM1
timestamp 1750100919
transform 0 1 530 -1 0 193
box -246 -583 246 583
use sky130_fd_pr__nfet_01v8_6AUVNX  XM2
timestamp 1750100919
transform 0 1 1478 -1 0 193
box -236 -355 236 355
<< labels >>
flabel metal1 s -41 397 -30 409 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -38 -26 -27 -14 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -46 303 -35 315 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -38 188 -27 200 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 1819 187 1830 199 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 1821 74 1832 86 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
