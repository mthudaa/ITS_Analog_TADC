magic
tech sky130A
magscale 1 2
timestamp 1757832914
<< error_p >>
rect -29 445 29 451
rect -29 411 -17 445
rect -29 405 29 411
<< nwell >>
rect -211 -584 211 584
<< pmos >>
rect -15 -436 15 364
<< pdiff >>
rect -73 321 -15 364
rect -73 287 -61 321
rect -27 287 -15 321
rect -73 253 -15 287
rect -73 219 -61 253
rect -27 219 -15 253
rect -73 185 -15 219
rect -73 151 -61 185
rect -27 151 -15 185
rect -73 117 -15 151
rect -73 83 -61 117
rect -27 83 -15 117
rect -73 49 -15 83
rect -73 15 -61 49
rect -27 15 -15 49
rect -73 -19 -15 15
rect -73 -53 -61 -19
rect -27 -53 -15 -19
rect -73 -87 -15 -53
rect -73 -121 -61 -87
rect -27 -121 -15 -87
rect -73 -155 -15 -121
rect -73 -189 -61 -155
rect -27 -189 -15 -155
rect -73 -223 -15 -189
rect -73 -257 -61 -223
rect -27 -257 -15 -223
rect -73 -291 -15 -257
rect -73 -325 -61 -291
rect -27 -325 -15 -291
rect -73 -359 -15 -325
rect -73 -393 -61 -359
rect -27 -393 -15 -359
rect -73 -436 -15 -393
rect 15 321 73 364
rect 15 287 27 321
rect 61 287 73 321
rect 15 253 73 287
rect 15 219 27 253
rect 61 219 73 253
rect 15 185 73 219
rect 15 151 27 185
rect 61 151 73 185
rect 15 117 73 151
rect 15 83 27 117
rect 61 83 73 117
rect 15 49 73 83
rect 15 15 27 49
rect 61 15 73 49
rect 15 -19 73 15
rect 15 -53 27 -19
rect 61 -53 73 -19
rect 15 -87 73 -53
rect 15 -121 27 -87
rect 61 -121 73 -87
rect 15 -155 73 -121
rect 15 -189 27 -155
rect 61 -189 73 -155
rect 15 -223 73 -189
rect 15 -257 27 -223
rect 61 -257 73 -223
rect 15 -291 73 -257
rect 15 -325 27 -291
rect 61 -325 73 -291
rect 15 -359 73 -325
rect 15 -393 27 -359
rect 61 -393 73 -359
rect 15 -436 73 -393
<< pdiffc >>
rect -61 287 -27 321
rect -61 219 -27 253
rect -61 151 -27 185
rect -61 83 -27 117
rect -61 15 -27 49
rect -61 -53 -27 -19
rect -61 -121 -27 -87
rect -61 -189 -27 -155
rect -61 -257 -27 -223
rect -61 -325 -27 -291
rect -61 -393 -27 -359
rect 27 287 61 321
rect 27 219 61 253
rect 27 151 61 185
rect 27 83 61 117
rect 27 15 61 49
rect 27 -53 61 -19
rect 27 -121 61 -87
rect 27 -189 61 -155
rect 27 -257 61 -223
rect 27 -325 61 -291
rect 27 -393 61 -359
<< nsubdiff >>
rect -175 514 -51 548
rect -17 514 17 548
rect 51 514 175 548
rect -175 425 -141 514
rect 141 425 175 514
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -514 -141 -425
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -514 175 -425
rect -175 -548 -51 -514
rect -17 -548 17 -514
rect 51 -548 175 -514
<< nsubdiffcont >>
rect -51 514 -17 548
rect 17 514 51 548
rect -175 391 -141 425
rect 141 391 175 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect -51 -548 -17 -514
rect 17 -548 51 -514
<< poly >>
rect -33 445 33 461
rect -33 411 -17 445
rect 17 411 33 445
rect -33 395 33 411
rect -15 364 15 395
rect -15 -462 15 -436
<< polycont >>
rect -17 411 17 445
<< locali >>
rect -175 514 -51 548
rect -17 514 17 548
rect 51 514 175 548
rect -175 425 -141 514
rect -33 411 -17 445
rect 17 411 33 445
rect 141 425 175 514
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -514 -141 -425
rect -61 341 -27 368
rect -61 269 -27 287
rect -61 197 -27 219
rect -61 125 -27 151
rect -61 53 -27 83
rect -61 -19 -27 15
rect -61 -87 -27 -53
rect -61 -155 -27 -125
rect -61 -223 -27 -197
rect -61 -291 -27 -269
rect -61 -359 -27 -341
rect -61 -440 -27 -413
rect 27 341 61 368
rect 27 269 61 287
rect 27 197 61 219
rect 27 125 61 151
rect 27 53 61 83
rect 27 -19 61 15
rect 27 -87 61 -53
rect 27 -155 61 -125
rect 27 -223 61 -197
rect 27 -291 61 -269
rect 27 -359 61 -341
rect 27 -440 61 -413
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -514 175 -425
rect -175 -548 -51 -514
rect -17 -548 17 -514
rect 51 -548 175 -514
<< viali >>
rect -17 411 17 445
rect -61 321 -27 341
rect -61 307 -27 321
rect -61 253 -27 269
rect -61 235 -27 253
rect -61 185 -27 197
rect -61 163 -27 185
rect -61 117 -27 125
rect -61 91 -27 117
rect -61 49 -27 53
rect -61 19 -27 49
rect -61 -53 -27 -19
rect -61 -121 -27 -91
rect -61 -125 -27 -121
rect -61 -189 -27 -163
rect -61 -197 -27 -189
rect -61 -257 -27 -235
rect -61 -269 -27 -257
rect -61 -325 -27 -307
rect -61 -341 -27 -325
rect -61 -393 -27 -379
rect -61 -413 -27 -393
rect 27 321 61 341
rect 27 307 61 321
rect 27 253 61 269
rect 27 235 61 253
rect 27 185 61 197
rect 27 163 61 185
rect 27 117 61 125
rect 27 91 61 117
rect 27 49 61 53
rect 27 19 61 49
rect 27 -53 61 -19
rect 27 -121 61 -91
rect 27 -125 61 -121
rect 27 -189 61 -163
rect 27 -197 61 -189
rect 27 -257 61 -235
rect 27 -269 61 -257
rect 27 -325 61 -307
rect 27 -341 61 -325
rect 27 -393 61 -379
rect 27 -413 61 -393
<< metal1 >>
rect -29 445 29 451
rect -29 411 -17 445
rect 17 411 29 445
rect -29 405 29 411
rect -67 341 -21 364
rect -67 307 -61 341
rect -27 307 -21 341
rect -67 269 -21 307
rect -67 235 -61 269
rect -27 235 -21 269
rect -67 197 -21 235
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -163 -21 -125
rect -67 -197 -61 -163
rect -27 -197 -21 -163
rect -67 -235 -21 -197
rect -67 -269 -61 -235
rect -27 -269 -21 -235
rect -67 -307 -21 -269
rect -67 -341 -61 -307
rect -27 -341 -21 -307
rect -67 -379 -21 -341
rect -67 -413 -61 -379
rect -27 -413 -21 -379
rect -67 -436 -21 -413
rect 21 341 67 364
rect 21 307 27 341
rect 61 307 67 341
rect 21 269 67 307
rect 21 235 27 269
rect 61 235 67 269
rect 21 197 67 235
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -163 67 -125
rect 21 -197 27 -163
rect 61 -197 67 -163
rect 21 -235 67 -197
rect 21 -269 27 -235
rect 61 -269 67 -235
rect 21 -307 67 -269
rect 21 -341 27 -307
rect 61 -341 67 -307
rect 21 -379 67 -341
rect 21 -413 27 -379
rect 61 -413 67 -379
rect 21 -436 67 -413
<< properties >>
string FIXED_BBOX -158 -531 158 531
<< end >>
