magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 1393 362 1433 365
rect 1393 328 1396 362
rect 1430 328 1433 362
rect 1393 325 1433 328
rect 967 277 1027 290
rect 805 261 865 274
rect 239 248 299 261
rect 77 245 117 248
rect 77 211 80 245
rect 114 211 117 245
rect 77 208 117 211
rect 239 214 252 248
rect 286 214 299 248
rect 239 201 299 214
rect 353 248 413 261
rect 353 214 366 248
rect 400 214 413 248
rect 353 201 413 214
rect 535 245 575 248
rect 535 211 538 245
rect 572 211 575 245
rect 805 227 818 261
rect 852 227 865 261
rect 967 243 980 277
rect 1014 243 1027 277
rect 967 230 1027 243
rect 805 214 865 227
rect 535 208 575 211
rect 241 150 281 153
rect 241 116 244 150
rect 278 116 281 150
rect 241 113 281 116
rect 529 71 569 74
rect 529 37 532 71
rect 566 37 569 71
rect 529 34 569 37
<< viali >>
rect 1396 328 1430 362
rect 80 211 114 245
rect 252 214 286 248
rect 366 214 400 248
rect 538 211 572 245
rect 818 227 852 261
rect 980 243 1014 277
rect 244 116 278 150
rect 532 37 566 71
<< metal1 >>
rect 38 568 1478 666
rect 0 507 875 511
rect 0 455 357 507
rect 409 455 809 507
rect 861 455 875 507
rect 0 451 875 455
rect 0 387 1037 391
rect 0 335 243 387
rect 295 335 971 387
rect 1023 335 1037 387
rect 0 331 1037 335
rect 1381 365 1445 371
rect 1381 362 1516 365
rect 1381 328 1396 362
rect 1430 328 1516 362
rect 1381 325 1516 328
rect 1381 319 1445 325
rect 955 286 1039 296
rect 793 270 877 280
rect 227 257 311 267
rect 65 245 129 254
rect 65 211 80 245
rect 114 211 129 245
rect 65 202 129 211
rect 227 205 243 257
rect 295 205 311 257
rect 77 74 117 202
rect 227 195 311 205
rect 341 257 425 267
rect 341 205 357 257
rect 409 205 425 257
rect 341 195 425 205
rect 523 245 587 254
rect 523 211 538 245
rect 572 211 587 245
rect 523 202 587 211
rect 793 218 809 270
rect 861 218 877 270
rect 955 234 971 286
rect 1023 234 1039 286
rect 955 224 1039 234
rect 793 208 877 218
rect 229 153 293 159
rect 535 153 575 202
rect 229 150 1516 153
rect 229 116 244 150
rect 278 116 1516 150
rect 229 113 1516 116
rect 229 107 293 113
rect 517 74 581 80
rect 77 71 1516 74
rect 77 37 532 71
rect 566 37 1516 71
rect 77 34 1516 37
rect 517 28 581 34
rect 38 -98 1478 0
<< via1 >>
rect 357 455 409 507
rect 809 455 861 507
rect 243 335 295 387
rect 971 335 1023 387
rect 243 248 295 257
rect 243 214 252 248
rect 252 214 286 248
rect 286 214 295 248
rect 243 205 295 214
rect 357 248 409 257
rect 357 214 366 248
rect 366 214 400 248
rect 400 214 409 248
rect 357 205 409 214
rect 809 261 861 270
rect 809 227 818 261
rect 818 227 852 261
rect 852 227 861 261
rect 809 218 861 227
rect 971 277 1023 286
rect 971 243 980 277
rect 980 243 1014 277
rect 1014 243 1023 277
rect 971 234 1023 243
<< metal2 >>
rect 353 507 413 521
rect 353 455 357 507
rect 409 455 413 507
rect 239 387 299 401
rect 239 335 243 387
rect 295 335 299 387
rect 239 257 299 335
rect 239 205 243 257
rect 295 205 299 257
rect 239 191 299 205
rect 353 257 413 455
rect 353 205 357 257
rect 409 205 413 257
rect 353 191 413 205
rect 805 507 865 521
rect 805 455 809 507
rect 861 455 865 507
rect 805 270 865 455
rect 805 218 809 270
rect 861 218 865 270
rect 967 387 1027 401
rect 967 335 971 387
rect 1023 335 1027 387
rect 967 286 1027 335
rect 967 234 971 286
rect 1023 234 1027 286
rect 967 220 1027 234
rect 805 204 865 218
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1750100919
transform 1 0 614 0 1 -49
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  x1
timestamp 1750100919
transform 1 0 38 0 1 -49
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  x2
timestamp 1750100919
transform 1 0 326 0 1 -49
box -38 -49 326 715
use sky130_fd_sc_hs__xor2_1  x3
timestamp 1750100919
transform 1 0 710 0 1 -49
box -38 -49 806 715
<< labels >>
flabel metal1 s 0 451 30 511 0 FreeSans 500 0 0 0 A
port 1 nsew
flabel metal1 s 0 331 30 391 0 FreeSans 500 0 0 0 B
port 2 nsew
flabel metal1 s 91 568 189 666 0 FreeSans 500 0 0 0 VDD
port 3 nsew
flabel metal1 s 95 -98 193 0 0 FreeSans 500 0 0 0 VSS
port 4 nsew
flabel metal1 s 1496 325 1516 365 0 FreeSans 500 0 0 0 RDY
port 5 nsew
flabel metal1 s 1476 113 1516 153 0 FreeSans 500 0 0 0 OUTP
port 6 nsew
flabel metal1 s 1476 34 1516 74 0 FreeSans 500 0 0 0 OUTN
port 7 nsew
<< end >>
