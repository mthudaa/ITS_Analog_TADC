magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect -246 -583 246 583
<< pmos >>
rect -50 64 50 364
rect -50 -364 50 -64
<< pdiff >>
rect -108 333 -50 364
rect -108 299 -96 333
rect -62 299 -50 333
rect -108 265 -50 299
rect -108 231 -96 265
rect -62 231 -50 265
rect -108 197 -50 231
rect -108 163 -96 197
rect -62 163 -50 197
rect -108 129 -50 163
rect -108 95 -96 129
rect -62 95 -50 129
rect -108 64 -50 95
rect 50 333 108 364
rect 50 299 62 333
rect 96 299 108 333
rect 50 265 108 299
rect 50 231 62 265
rect 96 231 108 265
rect 50 197 108 231
rect 50 163 62 197
rect 96 163 108 197
rect 50 129 108 163
rect 50 95 62 129
rect 96 95 108 129
rect 50 64 108 95
rect -108 -95 -50 -64
rect -108 -129 -96 -95
rect -62 -129 -50 -95
rect -108 -163 -50 -129
rect -108 -197 -96 -163
rect -62 -197 -50 -163
rect -108 -231 -50 -197
rect -108 -265 -96 -231
rect -62 -265 -50 -231
rect -108 -299 -50 -265
rect -108 -333 -96 -299
rect -62 -333 -50 -299
rect -108 -364 -50 -333
rect 50 -95 108 -64
rect 50 -129 62 -95
rect 96 -129 108 -95
rect 50 -163 108 -129
rect 50 -197 62 -163
rect 96 -197 108 -163
rect 50 -231 108 -197
rect 50 -265 62 -231
rect 96 -265 108 -231
rect 50 -299 108 -265
rect 50 -333 62 -299
rect 96 -333 108 -299
rect 50 -364 108 -333
<< pdiffc >>
rect -96 299 -62 333
rect -96 231 -62 265
rect -96 163 -62 197
rect -96 95 -62 129
rect 62 299 96 333
rect 62 231 96 265
rect 62 163 96 197
rect 62 95 96 129
rect -96 -129 -62 -95
rect -96 -197 -62 -163
rect -96 -265 -62 -231
rect -96 -333 -62 -299
rect 62 -129 96 -95
rect 62 -197 96 -163
rect 62 -265 96 -231
rect 62 -333 96 -299
<< nsubdiff >>
rect -210 513 -85 547
rect -51 513 -17 547
rect 17 513 51 547
rect 85 513 210 547
rect -210 425 -176 513
rect -210 357 -176 391
rect 176 425 210 513
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect -210 -513 -176 -425
rect 176 -391 210 -357
rect 176 -513 210 -425
rect -210 -547 -85 -513
rect -51 -547 -17 -513
rect 17 -547 51 -513
rect 85 -547 210 -513
<< nsubdiffcont >>
rect -85 513 -51 547
rect -17 513 17 547
rect 51 513 85 547
rect -210 391 -176 425
rect 176 391 210 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect -210 -425 -176 -391
rect 176 -425 210 -391
rect -85 -547 -51 -513
rect -17 -547 17 -513
rect 51 -547 85 -513
<< poly >>
rect -50 445 50 461
rect -50 411 -17 445
rect 17 411 50 445
rect -50 364 50 411
rect -50 17 50 64
rect -50 -17 -17 17
rect 17 -17 50 17
rect -50 -64 50 -17
rect -50 -411 50 -364
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect -50 -461 50 -445
<< polycont >>
rect -17 411 17 445
rect -17 -17 17 17
rect -17 -445 17 -411
<< locali >>
rect -210 513 -85 547
rect -51 513 -17 547
rect 17 513 51 547
rect 85 513 210 547
rect -210 425 -176 513
rect -50 411 -17 445
rect 17 411 50 445
rect 176 425 210 513
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -96 339 -62 368
rect -96 267 -62 299
rect -96 197 -62 231
rect -96 129 -62 161
rect -96 60 -62 89
rect 62 339 96 368
rect 62 267 96 299
rect 62 197 96 231
rect 62 129 96 161
rect 62 60 96 89
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect 176 17 210 51
rect -50 -17 -17 17
rect 17 -17 50 17
rect -210 -51 -176 -17
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -96 -89 -62 -60
rect -96 -161 -62 -129
rect -96 -231 -62 -197
rect -96 -299 -62 -267
rect -96 -368 -62 -339
rect 62 -89 96 -60
rect 62 -161 96 -129
rect 62 -231 96 -197
rect 62 -299 96 -267
rect 62 -368 96 -339
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect -210 -513 -176 -425
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect 176 -513 210 -425
rect -210 -547 -85 -513
rect -51 -547 -17 -513
rect 17 -547 51 -513
rect 85 -547 210 -513
<< viali >>
rect -17 411 17 445
rect -96 333 -62 339
rect -96 305 -62 333
rect -96 265 -62 267
rect -96 233 -62 265
rect -96 163 -62 195
rect -96 161 -62 163
rect -96 95 -62 123
rect -96 89 -62 95
rect 62 333 96 339
rect 62 305 96 333
rect 62 265 96 267
rect 62 233 96 265
rect 62 163 96 195
rect 62 161 96 163
rect 62 95 96 123
rect 62 89 96 95
rect -17 -17 17 17
rect -96 -95 -62 -89
rect -96 -123 -62 -95
rect -96 -163 -62 -161
rect -96 -195 -62 -163
rect -96 -265 -62 -233
rect -96 -267 -62 -265
rect -96 -333 -62 -305
rect -96 -339 -62 -333
rect 62 -95 96 -89
rect 62 -123 96 -95
rect 62 -163 96 -161
rect 62 -195 96 -163
rect 62 -265 96 -233
rect 62 -267 96 -265
rect 62 -333 96 -305
rect 62 -339 96 -333
rect -17 -445 17 -411
<< metal1 >>
rect -46 445 46 451
rect -46 411 -17 445
rect 17 411 46 445
rect -46 405 46 411
rect -102 339 -56 364
rect -102 305 -96 339
rect -62 305 -56 339
rect -102 267 -56 305
rect -102 233 -96 267
rect -62 233 -56 267
rect -102 195 -56 233
rect -102 161 -96 195
rect -62 161 -56 195
rect -102 123 -56 161
rect -102 89 -96 123
rect -62 89 -56 123
rect -102 64 -56 89
rect 56 339 102 364
rect 56 305 62 339
rect 96 305 102 339
rect 56 267 102 305
rect 56 233 62 267
rect 96 233 102 267
rect 56 195 102 233
rect 56 161 62 195
rect 96 161 102 195
rect 56 123 102 161
rect 56 89 62 123
rect 96 89 102 123
rect 56 64 102 89
rect -46 17 46 23
rect -46 -17 -17 17
rect 17 -17 46 17
rect -46 -23 46 -17
rect -102 -89 -56 -64
rect -102 -123 -96 -89
rect -62 -123 -56 -89
rect -102 -161 -56 -123
rect -102 -195 -96 -161
rect -62 -195 -56 -161
rect -102 -233 -56 -195
rect -102 -267 -96 -233
rect -62 -267 -56 -233
rect -102 -305 -56 -267
rect -102 -339 -96 -305
rect -62 -339 -56 -305
rect -102 -364 -56 -339
rect 56 -89 102 -64
rect 56 -123 62 -89
rect 96 -123 102 -89
rect 56 -161 102 -123
rect 56 -195 62 -161
rect 96 -195 102 -161
rect 56 -233 102 -195
rect 56 -267 62 -233
rect 96 -267 102 -233
rect 56 -305 102 -267
rect 56 -339 62 -305
rect 96 -339 102 -305
rect 56 -364 102 -339
rect -46 -411 46 -405
rect -46 -445 -17 -411
rect 17 -445 46 -411
rect -46 -451 46 -445
<< properties >>
string FIXED_BBOX -193 -530 193 530
<< end >>
