magic
tech sky130A
magscale 1 2
timestamp 1748343649
<< metal3 >>
rect -3410 2652 -2238 2680
rect -3410 1828 -2322 2652
rect -2258 1828 -2238 2652
rect -3410 1800 -2238 1828
rect -1998 2652 -826 2680
rect -1998 1828 -910 2652
rect -846 1828 -826 2652
rect -1998 1800 -826 1828
rect -586 2652 586 2680
rect -586 1828 502 2652
rect 566 1828 586 2652
rect -586 1800 586 1828
rect 826 2652 1998 2680
rect 826 1828 1914 2652
rect 1978 1828 1998 2652
rect 826 1800 1998 1828
rect 2238 2652 3410 2680
rect 2238 1828 3326 2652
rect 3390 1828 3410 2652
rect 2238 1800 3410 1828
rect -3410 1532 -2238 1560
rect -3410 708 -2322 1532
rect -2258 708 -2238 1532
rect -3410 680 -2238 708
rect -1998 1532 -826 1560
rect -1998 708 -910 1532
rect -846 708 -826 1532
rect -1998 680 -826 708
rect -586 1532 586 1560
rect -586 708 502 1532
rect 566 708 586 1532
rect -586 680 586 708
rect 826 1532 1998 1560
rect 826 708 1914 1532
rect 1978 708 1998 1532
rect 826 680 1998 708
rect 2238 1532 3410 1560
rect 2238 708 3326 1532
rect 3390 708 3410 1532
rect 2238 680 3410 708
rect -3410 412 -2238 440
rect -3410 -412 -2322 412
rect -2258 -412 -2238 412
rect -3410 -440 -2238 -412
rect -1998 412 -826 440
rect -1998 -412 -910 412
rect -846 -412 -826 412
rect -1998 -440 -826 -412
rect -586 412 586 440
rect -586 -412 502 412
rect 566 -412 586 412
rect -586 -440 586 -412
rect 826 412 1998 440
rect 826 -412 1914 412
rect 1978 -412 1998 412
rect 826 -440 1998 -412
rect 2238 412 3410 440
rect 2238 -412 3326 412
rect 3390 -412 3410 412
rect 2238 -440 3410 -412
rect -3410 -708 -2238 -680
rect -3410 -1532 -2322 -708
rect -2258 -1532 -2238 -708
rect -3410 -1560 -2238 -1532
rect -1998 -708 -826 -680
rect -1998 -1532 -910 -708
rect -846 -1532 -826 -708
rect -1998 -1560 -826 -1532
rect -586 -708 586 -680
rect -586 -1532 502 -708
rect 566 -1532 586 -708
rect -586 -1560 586 -1532
rect 826 -708 1998 -680
rect 826 -1532 1914 -708
rect 1978 -1532 1998 -708
rect 826 -1560 1998 -1532
rect 2238 -708 3410 -680
rect 2238 -1532 3326 -708
rect 3390 -1532 3410 -708
rect 2238 -1560 3410 -1532
rect -3410 -1828 -2238 -1800
rect -3410 -2652 -2322 -1828
rect -2258 -2652 -2238 -1828
rect -3410 -2680 -2238 -2652
rect -1998 -1828 -826 -1800
rect -1998 -2652 -910 -1828
rect -846 -2652 -826 -1828
rect -1998 -2680 -826 -2652
rect -586 -1828 586 -1800
rect -586 -2652 502 -1828
rect 566 -2652 586 -1828
rect -586 -2680 586 -2652
rect 826 -1828 1998 -1800
rect 826 -2652 1914 -1828
rect 1978 -2652 1998 -1828
rect 826 -2680 1998 -2652
rect 2238 -1828 3410 -1800
rect 2238 -2652 3326 -1828
rect 3390 -2652 3410 -1828
rect 2238 -2680 3410 -2652
<< via3 >>
rect -2322 1828 -2258 2652
rect -910 1828 -846 2652
rect 502 1828 566 2652
rect 1914 1828 1978 2652
rect 3326 1828 3390 2652
rect -2322 708 -2258 1532
rect -910 708 -846 1532
rect 502 708 566 1532
rect 1914 708 1978 1532
rect 3326 708 3390 1532
rect -2322 -412 -2258 412
rect -910 -412 -846 412
rect 502 -412 566 412
rect 1914 -412 1978 412
rect 3326 -412 3390 412
rect -2322 -1532 -2258 -708
rect -910 -1532 -846 -708
rect 502 -1532 566 -708
rect 1914 -1532 1978 -708
rect 3326 -1532 3390 -708
rect -2322 -2652 -2258 -1828
rect -910 -2652 -846 -1828
rect 502 -2652 566 -1828
rect 1914 -2652 1978 -1828
rect 3326 -2652 3390 -1828
<< mimcap >>
rect -3370 2600 -2570 2640
rect -3370 1880 -3330 2600
rect -2610 1880 -2570 2600
rect -3370 1840 -2570 1880
rect -1958 2600 -1158 2640
rect -1958 1880 -1918 2600
rect -1198 1880 -1158 2600
rect -1958 1840 -1158 1880
rect -546 2600 254 2640
rect -546 1880 -506 2600
rect 214 1880 254 2600
rect -546 1840 254 1880
rect 866 2600 1666 2640
rect 866 1880 906 2600
rect 1626 1880 1666 2600
rect 866 1840 1666 1880
rect 2278 2600 3078 2640
rect 2278 1880 2318 2600
rect 3038 1880 3078 2600
rect 2278 1840 3078 1880
rect -3370 1480 -2570 1520
rect -3370 760 -3330 1480
rect -2610 760 -2570 1480
rect -3370 720 -2570 760
rect -1958 1480 -1158 1520
rect -1958 760 -1918 1480
rect -1198 760 -1158 1480
rect -1958 720 -1158 760
rect -546 1480 254 1520
rect -546 760 -506 1480
rect 214 760 254 1480
rect -546 720 254 760
rect 866 1480 1666 1520
rect 866 760 906 1480
rect 1626 760 1666 1480
rect 866 720 1666 760
rect 2278 1480 3078 1520
rect 2278 760 2318 1480
rect 3038 760 3078 1480
rect 2278 720 3078 760
rect -3370 360 -2570 400
rect -3370 -360 -3330 360
rect -2610 -360 -2570 360
rect -3370 -400 -2570 -360
rect -1958 360 -1158 400
rect -1958 -360 -1918 360
rect -1198 -360 -1158 360
rect -1958 -400 -1158 -360
rect -546 360 254 400
rect -546 -360 -506 360
rect 214 -360 254 360
rect -546 -400 254 -360
rect 866 360 1666 400
rect 866 -360 906 360
rect 1626 -360 1666 360
rect 866 -400 1666 -360
rect 2278 360 3078 400
rect 2278 -360 2318 360
rect 3038 -360 3078 360
rect 2278 -400 3078 -360
rect -3370 -760 -2570 -720
rect -3370 -1480 -3330 -760
rect -2610 -1480 -2570 -760
rect -3370 -1520 -2570 -1480
rect -1958 -760 -1158 -720
rect -1958 -1480 -1918 -760
rect -1198 -1480 -1158 -760
rect -1958 -1520 -1158 -1480
rect -546 -760 254 -720
rect -546 -1480 -506 -760
rect 214 -1480 254 -760
rect -546 -1520 254 -1480
rect 866 -760 1666 -720
rect 866 -1480 906 -760
rect 1626 -1480 1666 -760
rect 866 -1520 1666 -1480
rect 2278 -760 3078 -720
rect 2278 -1480 2318 -760
rect 3038 -1480 3078 -760
rect 2278 -1520 3078 -1480
rect -3370 -1880 -2570 -1840
rect -3370 -2600 -3330 -1880
rect -2610 -2600 -2570 -1880
rect -3370 -2640 -2570 -2600
rect -1958 -1880 -1158 -1840
rect -1958 -2600 -1918 -1880
rect -1198 -2600 -1158 -1880
rect -1958 -2640 -1158 -2600
rect -546 -1880 254 -1840
rect -546 -2600 -506 -1880
rect 214 -2600 254 -1880
rect -546 -2640 254 -2600
rect 866 -1880 1666 -1840
rect 866 -2600 906 -1880
rect 1626 -2600 1666 -1880
rect 866 -2640 1666 -2600
rect 2278 -1880 3078 -1840
rect 2278 -2600 2318 -1880
rect 3038 -2600 3078 -1880
rect 2278 -2640 3078 -2600
<< mimcapcontact >>
rect -3330 1880 -2610 2600
rect -1918 1880 -1198 2600
rect -506 1880 214 2600
rect 906 1880 1626 2600
rect 2318 1880 3038 2600
rect -3330 760 -2610 1480
rect -1918 760 -1198 1480
rect -506 760 214 1480
rect 906 760 1626 1480
rect 2318 760 3038 1480
rect -3330 -360 -2610 360
rect -1918 -360 -1198 360
rect -506 -360 214 360
rect 906 -360 1626 360
rect 2318 -360 3038 360
rect -3330 -1480 -2610 -760
rect -1918 -1480 -1198 -760
rect -506 -1480 214 -760
rect 906 -1480 1626 -760
rect 2318 -1480 3038 -760
rect -3330 -2600 -2610 -1880
rect -1918 -2600 -1198 -1880
rect -506 -2600 214 -1880
rect 906 -2600 1626 -1880
rect 2318 -2600 3038 -1880
<< metal4 >>
rect -2338 2652 -2242 2668
rect -3331 2600 -2609 2601
rect -3331 1880 -3330 2600
rect -2610 1880 -2609 2600
rect -3331 1879 -2609 1880
rect -2338 1828 -2322 2652
rect -2258 1828 -2242 2652
rect -926 2652 -830 2668
rect -1919 2600 -1197 2601
rect -1919 1880 -1918 2600
rect -1198 1880 -1197 2600
rect -1919 1879 -1197 1880
rect -2338 1812 -2242 1828
rect -926 1828 -910 2652
rect -846 1828 -830 2652
rect 486 2652 582 2668
rect -507 2600 215 2601
rect -507 1880 -506 2600
rect 214 1880 215 2600
rect -507 1879 215 1880
rect -926 1812 -830 1828
rect 486 1828 502 2652
rect 566 1828 582 2652
rect 1898 2652 1994 2668
rect 905 2600 1627 2601
rect 905 1880 906 2600
rect 1626 1880 1627 2600
rect 905 1879 1627 1880
rect 486 1812 582 1828
rect 1898 1828 1914 2652
rect 1978 1828 1994 2652
rect 3310 2652 3406 2668
rect 2317 2600 3039 2601
rect 2317 1880 2318 2600
rect 3038 1880 3039 2600
rect 2317 1879 3039 1880
rect 1898 1812 1994 1828
rect 3310 1828 3326 2652
rect 3390 1828 3406 2652
rect 3310 1812 3406 1828
rect -2338 1532 -2242 1548
rect -3331 1480 -2609 1481
rect -3331 760 -3330 1480
rect -2610 760 -2609 1480
rect -3331 759 -2609 760
rect -2338 708 -2322 1532
rect -2258 708 -2242 1532
rect -926 1532 -830 1548
rect -1919 1480 -1197 1481
rect -1919 760 -1918 1480
rect -1198 760 -1197 1480
rect -1919 759 -1197 760
rect -2338 692 -2242 708
rect -926 708 -910 1532
rect -846 708 -830 1532
rect 486 1532 582 1548
rect -507 1480 215 1481
rect -507 760 -506 1480
rect 214 760 215 1480
rect -507 759 215 760
rect -926 692 -830 708
rect 486 708 502 1532
rect 566 708 582 1532
rect 1898 1532 1994 1548
rect 905 1480 1627 1481
rect 905 760 906 1480
rect 1626 760 1627 1480
rect 905 759 1627 760
rect 486 692 582 708
rect 1898 708 1914 1532
rect 1978 708 1994 1532
rect 3310 1532 3406 1548
rect 2317 1480 3039 1481
rect 2317 760 2318 1480
rect 3038 760 3039 1480
rect 2317 759 3039 760
rect 1898 692 1994 708
rect 3310 708 3326 1532
rect 3390 708 3406 1532
rect 3310 692 3406 708
rect -2338 412 -2242 428
rect -3331 360 -2609 361
rect -3331 -360 -3330 360
rect -2610 -360 -2609 360
rect -3331 -361 -2609 -360
rect -2338 -412 -2322 412
rect -2258 -412 -2242 412
rect -926 412 -830 428
rect -1919 360 -1197 361
rect -1919 -360 -1918 360
rect -1198 -360 -1197 360
rect -1919 -361 -1197 -360
rect -2338 -428 -2242 -412
rect -926 -412 -910 412
rect -846 -412 -830 412
rect 486 412 582 428
rect -507 360 215 361
rect -507 -360 -506 360
rect 214 -360 215 360
rect -507 -361 215 -360
rect -926 -428 -830 -412
rect 486 -412 502 412
rect 566 -412 582 412
rect 1898 412 1994 428
rect 905 360 1627 361
rect 905 -360 906 360
rect 1626 -360 1627 360
rect 905 -361 1627 -360
rect 486 -428 582 -412
rect 1898 -412 1914 412
rect 1978 -412 1994 412
rect 3310 412 3406 428
rect 2317 360 3039 361
rect 2317 -360 2318 360
rect 3038 -360 3039 360
rect 2317 -361 3039 -360
rect 1898 -428 1994 -412
rect 3310 -412 3326 412
rect 3390 -412 3406 412
rect 3310 -428 3406 -412
rect -2338 -708 -2242 -692
rect -3331 -760 -2609 -759
rect -3331 -1480 -3330 -760
rect -2610 -1480 -2609 -760
rect -3331 -1481 -2609 -1480
rect -2338 -1532 -2322 -708
rect -2258 -1532 -2242 -708
rect -926 -708 -830 -692
rect -1919 -760 -1197 -759
rect -1919 -1480 -1918 -760
rect -1198 -1480 -1197 -760
rect -1919 -1481 -1197 -1480
rect -2338 -1548 -2242 -1532
rect -926 -1532 -910 -708
rect -846 -1532 -830 -708
rect 486 -708 582 -692
rect -507 -760 215 -759
rect -507 -1480 -506 -760
rect 214 -1480 215 -760
rect -507 -1481 215 -1480
rect -926 -1548 -830 -1532
rect 486 -1532 502 -708
rect 566 -1532 582 -708
rect 1898 -708 1994 -692
rect 905 -760 1627 -759
rect 905 -1480 906 -760
rect 1626 -1480 1627 -760
rect 905 -1481 1627 -1480
rect 486 -1548 582 -1532
rect 1898 -1532 1914 -708
rect 1978 -1532 1994 -708
rect 3310 -708 3406 -692
rect 2317 -760 3039 -759
rect 2317 -1480 2318 -760
rect 3038 -1480 3039 -760
rect 2317 -1481 3039 -1480
rect 1898 -1548 1994 -1532
rect 3310 -1532 3326 -708
rect 3390 -1532 3406 -708
rect 3310 -1548 3406 -1532
rect -2338 -1828 -2242 -1812
rect -3331 -1880 -2609 -1879
rect -3331 -2600 -3330 -1880
rect -2610 -2600 -2609 -1880
rect -3331 -2601 -2609 -2600
rect -2338 -2652 -2322 -1828
rect -2258 -2652 -2242 -1828
rect -926 -1828 -830 -1812
rect -1919 -1880 -1197 -1879
rect -1919 -2600 -1918 -1880
rect -1198 -2600 -1197 -1880
rect -1919 -2601 -1197 -2600
rect -2338 -2668 -2242 -2652
rect -926 -2652 -910 -1828
rect -846 -2652 -830 -1828
rect 486 -1828 582 -1812
rect -507 -1880 215 -1879
rect -507 -2600 -506 -1880
rect 214 -2600 215 -1880
rect -507 -2601 215 -2600
rect -926 -2668 -830 -2652
rect 486 -2652 502 -1828
rect 566 -2652 582 -1828
rect 1898 -1828 1994 -1812
rect 905 -1880 1627 -1879
rect 905 -2600 906 -1880
rect 1626 -2600 1627 -1880
rect 905 -2601 1627 -2600
rect 486 -2668 582 -2652
rect 1898 -2652 1914 -1828
rect 1978 -2652 1994 -1828
rect 3310 -1828 3406 -1812
rect 2317 -1880 3039 -1879
rect 2317 -2600 2318 -1880
rect 3038 -2600 3039 -1880
rect 2317 -2601 3039 -2600
rect 1898 -2668 1994 -2652
rect 3310 -2652 3326 -1828
rect 3390 -2652 3406 -1828
rect 3310 -2668 3406 -2652
<< properties >>
string FIXED_BBOX 2238 1800 3118 2680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
